`timescale 1ns/1ns
import mAddAdd_package::*;

module mAddAdd(
  input logic clk,
  input logic reset,
  input Go_t \\QTree_Int_src_d ,
  output logic \\QTree_Int_src_r ,
  input QTree_Int_t dummy_write_QTree_Int_d,
  output logic dummy_write_QTree_Int_r,
  input Go_t sourceGo_d,
  output logic sourceGo_r,
  input Pointer_QTree_Int_t m1aen_0_d,
  output logic m1aen_0_r,
  input Pointer_QTree_Int_t m2aeo_1_d,
  output logic m2aeo_1_r,
  input Pointer_QTree_Int_t m3aep_2_d,
  output logic m3aep_2_r,
  output \Word16#_t  forkHP1_QTree_Int_snk_dout,
  input logic forkHP1_QTree_Int_snk_rout,
  output Pointer_QTree_Int_t dummy_write_QTree_Int_sink_dout,
  input logic dummy_write_QTree_Int_sink_rout,
  output Int_t \es_6_1I#_dout ,
  input logic \es_6_1I#_rout 
  );
  /* --define=INPUTS=((__05CQTree_Int_src, 0, 1, Go), (dummy_write_QTree_Int, 66, 73786976294838206464, QTree_Int), (sourceGo, 0, 1, Go), (m1aen_0, 16, 65536, Pointer_QTree_Int), (m2aeo_1, 16, 65536, Pointer_QTree_Int), (m3aep_2, 16, 65536, Pointer_QTree_Int)) */
  /* --define=TAPS=() */
  /* --define=OUTPUTS=((forkHP1_QTree_Int_snk, 16, 65536, Word16__023), (dummy_write_QTree_Int_sink, 16, 65536, Pointer_QTree_Int), (es_6_1I__023, 32, 4294967296, Int)) */
  /* TYPE_START
CT__024wnnz 16 3 (0,[0]) (1,[16p,16p,16p,16p]) (2,[32,16p,16p,16p]) (3,[32,32,16p,16p]) (4,[32,32,32,16p])
QTree_Int 16 2 (0,[0]) (1,[32]) (2,[16p,16p,16p,16p]) (3,[0])
CTf__027__027__027__027__027__027__027__027__027__027__027__027_f__027__027__027__027__027__027__027__027__027__027__027__027_Int 16 3 (0,[0]) (1,[16p,16p,16p,0,0,16p,16p,16p,16p]) (2,[16p,16p,16p,16p,0,0,16p,16p]) (3,[16p,16p,16p,16p,16p,0,0]) (4,[16p,16p,16p,16p])
CTf_f_Int 16 3 (0,[0]) (1,[16p,16p,16p,16p,0,0,16p,16p,16p,16p,16p,16p]) (2,[16p,16p,16p,16p,16p,0,0,16p,16p,16p]) (3,[16p,16p,16p,16p,16p,16p,0,0]) (4,[16p,16p,16p,16p])
TupGo___Pointer_QTree_Int 16 0 (0,[0,16p])
TupGo___Pointer_QTree_Int___Pointer_CT__024wnnz 16 0 (0,[0,16p,16p])
TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf__027__027__027__027__027__027__027__027__027__027__027__027_f__027__027__027__027__027__027__027__027__027__027__027__027_Int 16 0 (0,[0,16p,16p,0,0,16p])
TupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int 16 0 (0,[0,16p,16p,16p,0,0,16p])
TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int 16 0 (0,[0,16p,16p,0,0])
TupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int 16 0 (0,[0,16p,16p,16p,0,0])
TYPE_END */
  /*  */
  /*  */
  Go_t go_1_d;
  logic go_1_r;
  Go_t go_2_d;
  logic go_2_r;
  Go_t go_3_d;
  logic go_3_r;
  Go_t go_4_d;
  logic go_4_r;
  Go_t go__5_d;
  logic go__5_r;
  Go_t go__6_d;
  logic go__6_r;
  Go_t go__7_d;
  logic go__7_r;
  Go_t go__8_d;
  logic go__8_r;
  Go_t go__9_d;
  logic go__9_r;
  Go_t go__10_d;
  logic go__10_r;
  \Word16#_t  initHP_CT$wnnz_d;
  logic initHP_CT$wnnz_r;
  \Word16#_t  incrHP_CT$wnnz_d;
  logic incrHP_CT$wnnz_r;
  Go_t incrHP_mergeCT$wnnz_d;
  logic incrHP_mergeCT$wnnz_r;
  Go_t incrHP_CT$wnnz1_d;
  logic incrHP_CT$wnnz1_r;
  Go_t incrHP_CT$wnnz2_d;
  logic incrHP_CT$wnnz2_r;
  \Word16#_t  addHP_CT$wnnz_d;
  logic addHP_CT$wnnz_r;
  \Word16#_t  mergeHP_CT$wnnz_d;
  logic mergeHP_CT$wnnz_r;
  Go_t incrHP_mergeCT$wnnz_buf_d;
  logic incrHP_mergeCT$wnnz_buf_r;
  \Word16#_t  mergeHP_CT$wnnz_buf_d;
  logic mergeHP_CT$wnnz_buf_r;
  \Word16#_t  forkHP1_CT$wnnz_d;
  logic forkHP1_CT$wnnz_r;
  \Word16#_t  forkHP1_CT$wnn2_d;
  logic forkHP1_CT$wnn2_r;
  \Word16#_t  forkHP1_CT$wnn3_d;
  logic forkHP1_CT$wnn3_r;
  C2_t memMergeChoice_CT$wnnz_d;
  logic memMergeChoice_CT$wnnz_r;
  MemIn_CT$wnnz_t memMergeIn_CT$wnnz_d;
  logic memMergeIn_CT$wnnz_r;
  MemOut_CT$wnnz_t memOut_CT$wnnz_d;
  logic memOut_CT$wnnz_r;
  MemOut_CT$wnnz_t memReadOut_CT$wnnz_d;
  logic memReadOut_CT$wnnz_r;
  MemOut_CT$wnnz_t memWriteOut_CT$wnnz_d;
  logic memWriteOut_CT$wnnz_r;
  MemIn_CT$wnnz_t memMergeIn_CT$wnnz_dbuf_d;
  logic memMergeIn_CT$wnnz_dbuf_r;
  MemIn_CT$wnnz_t memMergeIn_CT$wnnz_rbuf_d;
  logic memMergeIn_CT$wnnz_rbuf_r;
  MemOut_CT$wnnz_t memOut_CT$wnnz_dbuf_d;
  logic memOut_CT$wnnz_dbuf_r;
  MemOut_CT$wnnz_t memOut_CT$wnnz_rbuf_d;
  logic memOut_CT$wnnz_rbuf_r;
  \Word16#_t  destructReadIn_CT$wnnz_d;
  logic destructReadIn_CT$wnnz_r;
  MemIn_CT$wnnz_t dconReadIn_CT$wnnz_d;
  logic dconReadIn_CT$wnnz_r;
  CT$wnnz_t readPointer_CT$wnnzscfarg_0_1_argbuf_d;
  logic readPointer_CT$wnnzscfarg_0_1_argbuf_r;
  C5_t writeMerge_choice_CT$wnnz_d;
  logic writeMerge_choice_CT$wnnz_r;
  CT$wnnz_t writeMerge_data_CT$wnnz_d;
  logic writeMerge_data_CT$wnnz_r;
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet0_1_argbuf_d;
  logic writeCT$wnnzlizzieLet0_1_argbuf_r;
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet59_1_argbuf_d;
  logic writeCT$wnnzlizzieLet59_1_argbuf_r;
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet5_1_argbuf_d;
  logic writeCT$wnnzlizzieLet5_1_argbuf_r;
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet60_1_argbuf_d;
  logic writeCT$wnnzlizzieLet60_1_argbuf_r;
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet61_1_argbuf_d;
  logic writeCT$wnnzlizzieLet61_1_argbuf_r;
  MemIn_CT$wnnz_t dconWriteIn_CT$wnnz_d;
  logic dconWriteIn_CT$wnnz_r;
  Pointer_CT$wnnz_t dconPtr_CT$wnnz_d;
  logic dconPtr_CT$wnnz_r;
  Pointer_CT$wnnz_t _259_d;
  logic _259_r;
  assign _259_r = 1'd1;
  Pointer_CT$wnnz_t demuxWriteResult_CT$wnnz_d;
  logic demuxWriteResult_CT$wnnz_r;
  \Word16#_t  initHP_QTree_Int_d;
  logic initHP_QTree_Int_r;
  \Word16#_t  incrHP_QTree_Int_d;
  logic incrHP_QTree_Int_r;
  Go_t incrHP_mergeQTree_Int_d;
  logic incrHP_mergeQTree_Int_r;
  Go_t incrHP_QTree_Int1_d;
  logic incrHP_QTree_Int1_r;
  Go_t incrHP_QTree_Int2_d;
  logic incrHP_QTree_Int2_r;
  \Word16#_t  addHP_QTree_Int_d;
  logic addHP_QTree_Int_r;
  \Word16#_t  mergeHP_QTree_Int_d;
  logic mergeHP_QTree_Int_r;
  Go_t incrHP_mergeQTree_Int_buf_d;
  logic incrHP_mergeQTree_Int_buf_r;
  \Word16#_t  mergeHP_QTree_Int_buf_d;
  logic mergeHP_QTree_Int_buf_r;
  Go_t go_1_dummy_write_QTree_Int_d;
  logic go_1_dummy_write_QTree_Int_r;
  Go_t go_2_dummy_write_QTree_Int_d;
  logic go_2_dummy_write_QTree_Int_r;
  \Word16#_t  forkHP1_QTree_Int_d;
  logic forkHP1_QTree_Int_r;
  \Word16#_t  forkHP1_QTree_Int_snk_d;
  logic forkHP1_QTree_Int_snk_r;
  \Word16#_t  forkHP1_QTree_In3_d;
  logic forkHP1_QTree_In3_r;
  \Word16#_t  forkHP1_QTree_In4_d;
  logic forkHP1_QTree_In4_r;
  C2_t memMergeChoice_QTree_Int_d;
  logic memMergeChoice_QTree_Int_r;
  MemIn_QTree_Int_t memMergeIn_QTree_Int_d;
  logic memMergeIn_QTree_Int_r;
  MemOut_QTree_Int_t memOut_QTree_Int_d;
  logic memOut_QTree_Int_r;
  MemOut_QTree_Int_t memReadOut_QTree_Int_d;
  logic memReadOut_QTree_Int_r;
  MemOut_QTree_Int_t memWriteOut_QTree_Int_d;
  logic memWriteOut_QTree_Int_r;
  MemIn_QTree_Int_t memMergeIn_QTree_Int_dbuf_d;
  logic memMergeIn_QTree_Int_dbuf_r;
  MemIn_QTree_Int_t memMergeIn_QTree_Int_rbuf_d;
  logic memMergeIn_QTree_Int_rbuf_r;
  MemOut_QTree_Int_t memOut_QTree_Int_dbuf_d;
  logic memOut_QTree_Int_dbuf_r;
  MemOut_QTree_Int_t memOut_QTree_Int_rbuf_d;
  logic memOut_QTree_Int_rbuf_r;
  C6_t readMerge_choice_QTree_Int_d;
  logic readMerge_choice_QTree_Int_r;
  Pointer_QTree_Int_t readMerge_data_QTree_Int_d;
  logic readMerge_data_QTree_Int_r;
  QTree_Int_t readPointer_QTree_Intm1aeq_1_argbuf_d;
  logic readPointer_QTree_Intm1aeq_1_argbuf_r;
  QTree_Int_t readPointer_QTree_Intm2aer_1_argbuf_d;
  logic readPointer_QTree_Intm2aer_1_argbuf_r;
  QTree_Int_t readPointer_QTree_Intm3aes_1_argbuf_d;
  logic readPointer_QTree_Intm3aes_1_argbuf_r;
  QTree_Int_t readPointer_QTree_Intq4afj_1_argbuf_d;
  logic readPointer_QTree_Intq4afj_1_argbuf_r;
  QTree_Int_t readPointer_QTree_Intt4afk_1_argbuf_d;
  logic readPointer_QTree_Intt4afk_1_argbuf_r;
  QTree_Int_t readPointer_QTree_Intwsmk_1_1_argbuf_d;
  logic readPointer_QTree_Intwsmk_1_1_argbuf_r;
  \Word16#_t  destructReadIn_QTree_Int_d;
  logic destructReadIn_QTree_Int_r;
  MemIn_QTree_Int_t dconReadIn_QTree_Int_d;
  logic dconReadIn_QTree_Int_r;
  QTree_Int_t destructReadOut_QTree_Int_d;
  logic destructReadOut_QTree_Int_r;
  C38_t writeMerge_choice_QTree_Int_d;
  logic writeMerge_choice_QTree_Int_r;
  QTree_Int_t writeMerge_data_QTree_Int_d;
  logic writeMerge_data_QTree_Int_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet10_1_argbuf_d;
  logic writeQTree_IntlizzieLet10_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet11_1_argbuf_d;
  logic writeQTree_IntlizzieLet11_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet13_1_argbuf_d;
  logic writeQTree_IntlizzieLet13_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet15_1_argbuf_d;
  logic writeQTree_IntlizzieLet15_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet16_1_argbuf_d;
  logic writeQTree_IntlizzieLet16_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet20_1_argbuf_d;
  logic writeQTree_IntlizzieLet20_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet21_1_argbuf_d;
  logic writeQTree_IntlizzieLet21_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet22_1_argbuf_d;
  logic writeQTree_IntlizzieLet22_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet23_1_argbuf_d;
  logic writeQTree_IntlizzieLet23_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet25_1_argbuf_d;
  logic writeQTree_IntlizzieLet25_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet26_1_argbuf_d;
  logic writeQTree_IntlizzieLet26_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet27_1_argbuf_d;
  logic writeQTree_IntlizzieLet27_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet28_1_argbuf_d;
  logic writeQTree_IntlizzieLet28_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet31_1_argbuf_d;
  logic writeQTree_IntlizzieLet31_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet32_1_argbuf_d;
  logic writeQTree_IntlizzieLet32_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet33_1_argbuf_d;
  logic writeQTree_IntlizzieLet33_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet34_1_argbuf_d;
  logic writeQTree_IntlizzieLet34_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet36_1_argbuf_d;
  logic writeQTree_IntlizzieLet36_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet37_2_1_argbuf_d;
  logic writeQTree_IntlizzieLet37_2_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet38_1_1_argbuf_d;
  logic writeQTree_IntlizzieLet38_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet39_1_1_argbuf_d;
  logic writeQTree_IntlizzieLet39_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet40_1_argbuf_d;
  logic writeQTree_IntlizzieLet40_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet41_1_argbuf_d;
  logic writeQTree_IntlizzieLet41_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet42_1_argbuf_d;
  logic writeQTree_IntlizzieLet42_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet45_1_argbuf_d;
  logic writeQTree_IntlizzieLet45_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet46_1_argbuf_d;
  logic writeQTree_IntlizzieLet46_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet47_1_argbuf_d;
  logic writeQTree_IntlizzieLet47_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet48_1_argbuf_d;
  logic writeQTree_IntlizzieLet48_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet50_1_argbuf_d;
  logic writeQTree_IntlizzieLet50_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet51_1_argbuf_d;
  logic writeQTree_IntlizzieLet51_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet53_1_argbuf_d;
  logic writeQTree_IntlizzieLet53_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet54_1_argbuf_d;
  logic writeQTree_IntlizzieLet54_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet55_1_argbuf_d;
  logic writeQTree_IntlizzieLet55_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet66_1_argbuf_d;
  logic writeQTree_IntlizzieLet66_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet71_1_argbuf_d;
  logic writeQTree_IntlizzieLet71_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet8_1_argbuf_d;
  logic writeQTree_IntlizzieLet8_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet9_1_argbuf_d;
  logic writeQTree_IntlizzieLet9_1_argbuf_r;
  Pointer_QTree_Int_t dummy_write_QTree_Int_sink_d;
  logic dummy_write_QTree_Int_sink_r;
  MemIn_QTree_Int_t dconWriteIn_QTree_Int_d;
  logic dconWriteIn_QTree_Int_r;
  Pointer_QTree_Int_t dconPtr_QTree_Int_d;
  logic dconPtr_QTree_Int_r;
  Pointer_QTree_Int_t _258_d;
  logic _258_r;
  assign _258_r = 1'd1;
  Pointer_QTree_Int_t demuxWriteResult_QTree_Int_d;
  logic demuxWriteResult_QTree_Int_r;
  \Word16#_t  \initHP_CTf''''''''''''_f''''''''''''_Int_d ;
  logic \initHP_CTf''''''''''''_f''''''''''''_Int_r ;
  \Word16#_t  \incrHP_CTf''''''''''''_f''''''''''''_Int_d ;
  logic \incrHP_CTf''''''''''''_f''''''''''''_Int_r ;
  Go_t \incrHP_mergeCTf''''''''''''_f''''''''''''_Int_d ;
  logic \incrHP_mergeCTf''''''''''''_f''''''''''''_Int_r ;
  Go_t \incrHP_CTf''''''''''''_f''''''''''''_Int1_d ;
  logic \incrHP_CTf''''''''''''_f''''''''''''_Int1_r ;
  Go_t \incrHP_CTf''''''''''''_f''''''''''''_Int2_d ;
  logic \incrHP_CTf''''''''''''_f''''''''''''_Int2_r ;
  \Word16#_t  \addHP_CTf''''''''''''_f''''''''''''_Int_d ;
  logic \addHP_CTf''''''''''''_f''''''''''''_Int_r ;
  \Word16#_t  \mergeHP_CTf''''''''''''_f''''''''''''_Int_d ;
  logic \mergeHP_CTf''''''''''''_f''''''''''''_Int_r ;
  Go_t \incrHP_mergeCTf''''''''''''_f''''''''''''_Int_buf_d ;
  logic \incrHP_mergeCTf''''''''''''_f''''''''''''_Int_buf_r ;
  \Word16#_t  \mergeHP_CTf''''''''''''_f''''''''''''_Int_buf_d ;
  logic \mergeHP_CTf''''''''''''_f''''''''''''_Int_buf_r ;
  \Word16#_t  \forkHP1_CTf''''''''''''_f''''''''''''_Int_d ;
  logic \forkHP1_CTf''''''''''''_f''''''''''''_Int_r ;
  \Word16#_t  \forkHP1_CTf''''''''''''_f''''''''''''_In2_d ;
  logic \forkHP1_CTf''''''''''''_f''''''''''''_In2_r ;
  \Word16#_t  \forkHP1_CTf''''''''''''_f''''''''''''_In3_d ;
  logic \forkHP1_CTf''''''''''''_f''''''''''''_In3_r ;
  C2_t \memMergeChoice_CTf''''''''''''_f''''''''''''_Int_d ;
  logic \memMergeChoice_CTf''''''''''''_f''''''''''''_Int_r ;
  \MemIn_CTf''''''''''''_f''''''''''''_Int_t  \memMergeIn_CTf''''''''''''_f''''''''''''_Int_d ;
  logic \memMergeIn_CTf''''''''''''_f''''''''''''_Int_r ;
  \MemOut_CTf''''''''''''_f''''''''''''_Int_t  \memOut_CTf''''''''''''_f''''''''''''_Int_d ;
  logic \memOut_CTf''''''''''''_f''''''''''''_Int_r ;
  \MemOut_CTf''''''''''''_f''''''''''''_Int_t  \memReadOut_CTf''''''''''''_f''''''''''''_Int_d ;
  logic \memReadOut_CTf''''''''''''_f''''''''''''_Int_r ;
  \MemOut_CTf''''''''''''_f''''''''''''_Int_t  \memWriteOut_CTf''''''''''''_f''''''''''''_Int_d ;
  logic \memWriteOut_CTf''''''''''''_f''''''''''''_Int_r ;
  \MemIn_CTf''''''''''''_f''''''''''''_Int_t  \memMergeIn_CTf''''''''''''_f''''''''''''_Int_dbuf_d ;
  logic \memMergeIn_CTf''''''''''''_f''''''''''''_Int_dbuf_r ;
  \MemIn_CTf''''''''''''_f''''''''''''_Int_t  \memMergeIn_CTf''''''''''''_f''''''''''''_Int_rbuf_d ;
  logic \memMergeIn_CTf''''''''''''_f''''''''''''_Int_rbuf_r ;
  \MemOut_CTf''''''''''''_f''''''''''''_Int_t  \memOut_CTf''''''''''''_f''''''''''''_Int_dbuf_d ;
  logic \memOut_CTf''''''''''''_f''''''''''''_Int_dbuf_r ;
  \MemOut_CTf''''''''''''_f''''''''''''_Int_t  \memOut_CTf''''''''''''_f''''''''''''_Int_rbuf_d ;
  logic \memOut_CTf''''''''''''_f''''''''''''_Int_rbuf_r ;
  \Word16#_t  \destructReadIn_CTf''''''''''''_f''''''''''''_Int_d ;
  logic \destructReadIn_CTf''''''''''''_f''''''''''''_Int_r ;
  \MemIn_CTf''''''''''''_f''''''''''''_Int_t  \dconReadIn_CTf''''''''''''_f''''''''''''_Int_d ;
  logic \dconReadIn_CTf''''''''''''_f''''''''''''_Int_r ;
  \CTf''''''''''''_f''''''''''''_Int_t  \readPointer_CTf''''''''''''_f''''''''''''_Intscfarg_0_1_1_argbuf_d ;
  logic \readPointer_CTf''''''''''''_f''''''''''''_Intscfarg_0_1_1_argbuf_r ;
  C5_t \writeMerge_choice_CTf''''''''''''_f''''''''''''_Int_d ;
  logic \writeMerge_choice_CTf''''''''''''_f''''''''''''_Int_r ;
  \CTf''''''''''''_f''''''''''''_Int_t  \writeMerge_data_CTf''''''''''''_f''''''''''''_Int_d ;
  logic \writeMerge_data_CTf''''''''''''_f''''''''''''_Int_r ;
  \Pointer_CTf''''''''''''_f''''''''''''_Int_t  \writeCTf''''''''''''_f''''''''''''_IntlizzieLet14_1_argbuf_d ;
  logic \writeCTf''''''''''''_f''''''''''''_IntlizzieLet14_1_argbuf_r ;
  \Pointer_CTf''''''''''''_f''''''''''''_Int_t  \writeCTf''''''''''''_f''''''''''''_IntlizzieLet56_1_argbuf_d ;
  logic \writeCTf''''''''''''_f''''''''''''_IntlizzieLet56_1_argbuf_r ;
  \Pointer_CTf''''''''''''_f''''''''''''_Int_t  \writeCTf''''''''''''_f''''''''''''_IntlizzieLet63_1_argbuf_d ;
  logic \writeCTf''''''''''''_f''''''''''''_IntlizzieLet63_1_argbuf_r ;
  \Pointer_CTf''''''''''''_f''''''''''''_Int_t  \writeCTf''''''''''''_f''''''''''''_IntlizzieLet64_1_argbuf_d ;
  logic \writeCTf''''''''''''_f''''''''''''_IntlizzieLet64_1_argbuf_r ;
  \Pointer_CTf''''''''''''_f''''''''''''_Int_t  \writeCTf''''''''''''_f''''''''''''_IntlizzieLet65_1_argbuf_d ;
  logic \writeCTf''''''''''''_f''''''''''''_IntlizzieLet65_1_argbuf_r ;
  \MemIn_CTf''''''''''''_f''''''''''''_Int_t  \dconWriteIn_CTf''''''''''''_f''''''''''''_Int_d ;
  logic \dconWriteIn_CTf''''''''''''_f''''''''''''_Int_r ;
  \Pointer_CTf''''''''''''_f''''''''''''_Int_t  \dconPtr_CTf''''''''''''_f''''''''''''_Int_d ;
  logic \dconPtr_CTf''''''''''''_f''''''''''''_Int_r ;
  \Pointer_CTf''''''''''''_f''''''''''''_Int_t  _257_d;
  logic _257_r;
  assign _257_r = 1'd1;
  \Pointer_CTf''''''''''''_f''''''''''''_Int_t  \demuxWriteResult_CTf''''''''''''_f''''''''''''_Int_d ;
  logic \demuxWriteResult_CTf''''''''''''_f''''''''''''_Int_r ;
  \Word16#_t  initHP_CTf_f_Int_d;
  logic initHP_CTf_f_Int_r;
  \Word16#_t  incrHP_CTf_f_Int_d;
  logic incrHP_CTf_f_Int_r;
  Go_t incrHP_mergeCTf_f_Int_d;
  logic incrHP_mergeCTf_f_Int_r;
  Go_t incrHP_CTf_f_Int1_d;
  logic incrHP_CTf_f_Int1_r;
  Go_t incrHP_CTf_f_Int2_d;
  logic incrHP_CTf_f_Int2_r;
  \Word16#_t  addHP_CTf_f_Int_d;
  logic addHP_CTf_f_Int_r;
  \Word16#_t  mergeHP_CTf_f_Int_d;
  logic mergeHP_CTf_f_Int_r;
  Go_t incrHP_mergeCTf_f_Int_buf_d;
  logic incrHP_mergeCTf_f_Int_buf_r;
  \Word16#_t  mergeHP_CTf_f_Int_buf_d;
  logic mergeHP_CTf_f_Int_buf_r;
  \Word16#_t  forkHP1_CTf_f_Int_d;
  logic forkHP1_CTf_f_Int_r;
  \Word16#_t  forkHP1_CTf_f_In2_d;
  logic forkHP1_CTf_f_In2_r;
  \Word16#_t  forkHP1_CTf_f_In3_d;
  logic forkHP1_CTf_f_In3_r;
  C2_t memMergeChoice_CTf_f_Int_d;
  logic memMergeChoice_CTf_f_Int_r;
  MemIn_CTf_f_Int_t memMergeIn_CTf_f_Int_d;
  logic memMergeIn_CTf_f_Int_r;
  MemOut_CTf_f_Int_t memOut_CTf_f_Int_d;
  logic memOut_CTf_f_Int_r;
  MemOut_CTf_f_Int_t memReadOut_CTf_f_Int_d;
  logic memReadOut_CTf_f_Int_r;
  MemOut_CTf_f_Int_t memWriteOut_CTf_f_Int_d;
  logic memWriteOut_CTf_f_Int_r;
  MemIn_CTf_f_Int_t memMergeIn_CTf_f_Int_dbuf_d;
  logic memMergeIn_CTf_f_Int_dbuf_r;
  MemIn_CTf_f_Int_t memMergeIn_CTf_f_Int_rbuf_d;
  logic memMergeIn_CTf_f_Int_rbuf_r;
  MemOut_CTf_f_Int_t memOut_CTf_f_Int_dbuf_d;
  logic memOut_CTf_f_Int_dbuf_r;
  MemOut_CTf_f_Int_t memOut_CTf_f_Int_rbuf_d;
  logic memOut_CTf_f_Int_rbuf_r;
  \Word16#_t  destructReadIn_CTf_f_Int_d;
  logic destructReadIn_CTf_f_Int_r;
  MemIn_CTf_f_Int_t dconReadIn_CTf_f_Int_d;
  logic dconReadIn_CTf_f_Int_r;
  CTf_f_Int_t readPointer_CTf_f_Intscfarg_0_2_1_argbuf_d;
  logic readPointer_CTf_f_Intscfarg_0_2_1_argbuf_r;
  C5_t writeMerge_choice_CTf_f_Int_d;
  logic writeMerge_choice_CTf_f_Int_r;
  CTf_f_Int_t writeMerge_data_CTf_f_Int_d;
  logic writeMerge_data_CTf_f_Int_r;
  Pointer_CTf_f_Int_t writeCTf_f_IntlizzieLet52_1_argbuf_d;
  logic writeCTf_f_IntlizzieLet52_1_argbuf_r;
  Pointer_CTf_f_Int_t writeCTf_f_IntlizzieLet57_1_argbuf_d;
  logic writeCTf_f_IntlizzieLet57_1_argbuf_r;
  Pointer_CTf_f_Int_t writeCTf_f_IntlizzieLet68_1_argbuf_d;
  logic writeCTf_f_IntlizzieLet68_1_argbuf_r;
  Pointer_CTf_f_Int_t writeCTf_f_IntlizzieLet69_1_argbuf_d;
  logic writeCTf_f_IntlizzieLet69_1_argbuf_r;
  Pointer_CTf_f_Int_t writeCTf_f_IntlizzieLet70_1_argbuf_d;
  logic writeCTf_f_IntlizzieLet70_1_argbuf_r;
  MemIn_CTf_f_Int_t dconWriteIn_CTf_f_Int_d;
  logic dconWriteIn_CTf_f_Int_r;
  Pointer_CTf_f_Int_t dconPtr_CTf_f_Int_d;
  logic dconPtr_CTf_f_Int_r;
  Pointer_CTf_f_Int_t _256_d;
  logic _256_r;
  assign _256_r = 1'd1;
  Pointer_CTf_f_Int_t demuxWriteResult_CTf_f_Int_d;
  logic demuxWriteResult_CTf_f_Int_r;
  Go_t \$wnnzTupGo___Pointer_QTree_Intgo_6_d ;
  logic \$wnnzTupGo___Pointer_QTree_Intgo_6_r ;
  Pointer_QTree_Int_t \$wnnzTupGo___Pointer_QTree_Intwsmk_d ;
  logic \$wnnzTupGo___Pointer_QTree_Intwsmk_r ;
  Go_t go_6_1_d;
  logic go_6_1_r;
  Go_t go_6_2_d;
  logic go_6_2_r;
  Pointer_QTree_Int_t wsmk_1_argbuf_d;
  logic wsmk_1_argbuf_r;
  Int_t \es_6_1I#_d ;
  logic \es_6_1I#_r ;
  C5_t applyfnInt_Bool_5_choice_d;
  logic applyfnInt_Bool_5_choice_r;
  TupGo___MyDTInt_Bool___Int_t applyfnInt_Bool_5_data_d;
  logic applyfnInt_Bool_5_data_r;
  MyDTInt_Bool_t arg0_1_d;
  logic arg0_1_r;
  MyDTInt_Bool_t arg0_2_d;
  logic arg0_2_r;
  MyDTInt_Bool_t arg0_3_d;
  logic arg0_3_r;
  MyBool_t applyfnInt_Bool_5_resbuf_d;
  logic applyfnInt_Bool_5_resbuf_r;
  MyBool_t applyfnInt_Bool_5_2_argbuf_d;
  logic applyfnInt_Bool_5_2_argbuf_r;
  MyBool_t es_2_1_d;
  logic es_2_1_r;
  MyBool_t es_2_2_d;
  logic es_2_2_r;
  MyBool_t es_2_3_d;
  logic es_2_3_r;
  MyBool_t es_2_4_d;
  logic es_2_4_r;
  MyBool_t es_2_5_d;
  logic es_2_5_r;
  MyBool_t applyfnInt_Bool_5_3_argbuf_d;
  logic applyfnInt_Bool_5_3_argbuf_r;
  MyBool_t es_10_1_d;
  logic es_10_1_r;
  MyBool_t es_10_2_d;
  logic es_10_2_r;
  MyBool_t es_10_3_d;
  logic es_10_3_r;
  MyBool_t es_10_4_d;
  logic es_10_4_r;
  MyBool_t es_10_5_d;
  logic es_10_5_r;
  MyBool_t applyfnInt_Bool_5_4_argbuf_d;
  logic applyfnInt_Bool_5_4_argbuf_r;
  MyBool_t es_14_1_d;
  logic es_14_1_r;
  MyBool_t es_14_2_d;
  logic es_14_2_r;
  MyBool_t es_14_3_d;
  logic es_14_3_r;
  MyBool_t es_14_4_d;
  logic es_14_4_r;
  MyBool_t es_14_5_d;
  logic es_14_5_r;
  MyBool_t es_14_6_d;
  logic es_14_6_r;
  MyBool_t es_14_7_d;
  logic es_14_7_r;
  MyBool_t es_14_8_d;
  logic es_14_8_r;
  MyBool_t applyfnInt_Bool_5_5_argbuf_d;
  logic applyfnInt_Bool_5_5_argbuf_r;
  MyBool_t es_21_1_d;
  logic es_21_1_r;
  MyBool_t es_21_2_d;
  logic es_21_2_r;
  MyBool_t es_21_3_d;
  logic es_21_3_r;
  MyBool_t es_21_4_d;
  logic es_21_4_r;
  MyBool_t es_21_5_d;
  logic es_21_5_r;
  MyBool_t es_21_6_d;
  logic es_21_6_r;
  MyBool_t applyfnInt_Bool_5_1_d;
  logic applyfnInt_Bool_5_1_r;
  MyBool_t applyfnInt_Bool_5_2_d;
  logic applyfnInt_Bool_5_2_r;
  MyBool_t applyfnInt_Bool_5_3_d;
  logic applyfnInt_Bool_5_3_r;
  MyBool_t applyfnInt_Bool_5_4_d;
  logic applyfnInt_Bool_5_4_r;
  MyBool_t applyfnInt_Bool_5_5_d;
  logic applyfnInt_Bool_5_5_r;
  Go_t applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intgo_7_d;
  logic applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intgo_7_r;
  MyDTInt_Bool_t applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_d;
  logic applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_r;
  Int_t applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg1_d;
  logic applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg1_r;
  MyBool_t es_2_1_1_d;
  logic es_2_1_1_r;
  MyBool_t es_2_1_2_d;
  logic es_2_1_2_r;
  MyBool_t es_2_1_3_d;
  logic es_2_1_3_r;
  MyBool_t es_2_1_4_d;
  logic es_2_1_4_r;
  MyBool_t es_2_1_5_d;
  logic es_2_1_5_r;
  C12_t applyfnInt_Int_Int_5_choice_d;
  logic applyfnInt_Int_Int_5_choice_r;
  TupMyDTInt_Int_Int___Int___Int_t applyfnInt_Int_Int_5_data_d;
  logic applyfnInt_Int_Int_5_data_r;
  MyDTInt_Int_Int_t arg0_2_1_d;
  logic arg0_2_1_r;
  MyDTInt_Int_Int_t arg0_2_2_d;
  logic arg0_2_2_r;
  MyDTInt_Int_Int_t arg0_2_3_d;
  logic arg0_2_3_r;
  Int_t applyfnInt_Int_Int_5_resbuf_d;
  logic applyfnInt_Int_Int_5_resbuf_r;
  Int_t applyfnInt_Int_Int_5_10_argbuf_d;
  logic applyfnInt_Int_Int_5_10_argbuf_r;
  Int_t es_17_1_argbuf_d;
  logic es_17_1_argbuf_r;
  Int_t applyfnInt_Int_Int_5_11_argbuf_d;
  logic applyfnInt_Int_Int_5_11_argbuf_r;
  Int_t es_24_1_argbuf_d;
  logic es_24_1_argbuf_r;
  Int_t applyfnInt_Int_Int_5_12_argbuf_d;
  logic applyfnInt_Int_Int_5_12_argbuf_r;
  QTree_Int_t es_22_1QVal_Int_d;
  logic es_22_1QVal_Int_r;
  Int_t applyfnInt_Int_Int_5_2_argbuf_d;
  logic applyfnInt_Int_Int_5_2_argbuf_r;
  QTree_Int_t es_3_1_1QVal_Int_d;
  logic es_3_1_1QVal_Int_r;
  Int_t applyfnInt_Int_Int_5_3_argbuf_d;
  logic applyfnInt_Int_Int_5_3_argbuf_r;
  Int_t es_1_1_argbuf_d;
  logic es_1_1_argbuf_r;
  Int_t applyfnInt_Int_Int_5_4_argbuf_d;
  logic applyfnInt_Int_Int_5_4_argbuf_r;
  QTree_Int_t es_3_1QVal_Int_d;
  logic es_3_1QVal_Int_r;
  Int_t applyfnInt_Int_Int_5_5_argbuf_d;
  logic applyfnInt_Int_Int_5_5_argbuf_r;
  Int_t es_9_1_argbuf_d;
  logic es_9_1_argbuf_r;
  Int_t applyfnInt_Int_Int_5_6_argbuf_d;
  logic applyfnInt_Int_Int_5_6_argbuf_r;
  QTree_Int_t es_11_1QVal_Int_d;
  logic es_11_1QVal_Int_r;
  Int_t applyfnInt_Int_Int_5_7_argbuf_d;
  logic applyfnInt_Int_Int_5_7_argbuf_r;
  Int_t es_13_1_argbuf_d;
  logic es_13_1_argbuf_r;
  Int_t applyfnInt_Int_Int_5_8_argbuf_d;
  logic applyfnInt_Int_Int_5_8_argbuf_r;
  QTree_Int_t es_15_1QVal_Int_d;
  logic es_15_1QVal_Int_r;
  Int_t applyfnInt_Int_Int_5_9_argbuf_d;
  logic applyfnInt_Int_Int_5_9_argbuf_r;
  Int_t es_19_1_argbuf_d;
  logic es_19_1_argbuf_r;
  Int_t applyfnInt_Int_Int_5_1_d;
  logic applyfnInt_Int_Int_5_1_r;
  Int_t applyfnInt_Int_Int_5_2_d;
  logic applyfnInt_Int_Int_5_2_r;
  Int_t applyfnInt_Int_Int_5_3_d;
  logic applyfnInt_Int_Int_5_3_r;
  Int_t applyfnInt_Int_Int_5_4_d;
  logic applyfnInt_Int_Int_5_4_r;
  Int_t applyfnInt_Int_Int_5_5_d;
  logic applyfnInt_Int_Int_5_5_r;
  Int_t applyfnInt_Int_Int_5_6_d;
  logic applyfnInt_Int_Int_5_6_r;
  Int_t applyfnInt_Int_Int_5_7_d;
  logic applyfnInt_Int_Int_5_7_r;
  Int_t applyfnInt_Int_Int_5_8_d;
  logic applyfnInt_Int_Int_5_8_r;
  Int_t applyfnInt_Int_Int_5_9_d;
  logic applyfnInt_Int_Int_5_9_r;
  Int_t applyfnInt_Int_Int_5_10_d;
  logic applyfnInt_Int_Int_5_10_r;
  Int_t applyfnInt_Int_Int_5_11_d;
  logic applyfnInt_Int_Int_5_11_r;
  Int_t applyfnInt_Int_Int_5_12_d;
  logic applyfnInt_Int_Int_5_12_r;
  MyDTInt_Int_Int_t applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_2_d;
  logic applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_2_r;
  Int_t applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg2_d;
  logic applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg2_r;
  Int_t applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg1_1_d;
  logic applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg1_1_r;
  Int_t es_1_1_1_argbuf_d;
  logic es_1_1_1_argbuf_r;
  Int_t arg0_1Dcon_isZ_d;
  logic arg0_1Dcon_isZ_r;
  Int_t arg0_1Dcon_isZ_1_d;
  logic arg0_1Dcon_isZ_1_r;
  Int_t arg0_1Dcon_isZ_2_d;
  logic arg0_1Dcon_isZ_2_r;
  Int_t arg0_1Dcon_isZ_3_d;
  logic arg0_1Dcon_isZ_3_r;
  Int_t arg0_1Dcon_isZ_4_d;
  logic arg0_1Dcon_isZ_4_r;
  \Int#_t  x1ajq_destruct_d;
  logic x1ajq_destruct_r;
  Int_t \arg0_1Dcon_isZ_1I#_d ;
  logic \arg0_1Dcon_isZ_1I#_r ;
  Go_t \arg0_1Dcon_isZ_3I#_d ;
  logic \arg0_1Dcon_isZ_3I#_r ;
  Go_t \arg0_1Dcon_isZ_3I#_1_d ;
  logic \arg0_1Dcon_isZ_3I#_1_r ;
  Go_t \arg0_1Dcon_isZ_3I#_2_d ;
  logic \arg0_1Dcon_isZ_3I#_2_r ;
  Go_t \arg0_1Dcon_isZ_3I#_3_d ;
  logic \arg0_1Dcon_isZ_3I#_3_r ;
  Go_t \arg0_1Dcon_isZ_3I#_1_argbuf_d ;
  logic \arg0_1Dcon_isZ_3I#_1_argbuf_r ;
  \Int#_t  \arg0_1Dcon_isZ_3I#_1_argbuf_0_d ;
  logic \arg0_1Dcon_isZ_3I#_1_argbuf_0_r ;
  Bool_t lizzieLet1_1wild1Xv_1_Eq_d;
  logic lizzieLet1_1wild1Xv_1_Eq_r;
  Go_t \arg0_1Dcon_isZ_3I#_2_argbuf_d ;
  logic \arg0_1Dcon_isZ_3I#_2_argbuf_r ;
  TupGo___Bool_t boolConvert_1TupGo___Bool_1_d;
  logic boolConvert_1TupGo___Bool_1_r;
  MyBool_t lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_d;
  logic lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_r;
  Go_t arg0_2Dcon_isZ_d;
  logic arg0_2Dcon_isZ_r;
  Int_t \arg0_2_1Dcon_$fNumInt_$c+_d ;
  logic \arg0_2_1Dcon_$fNumInt_$c+_r ;
  Int_t \arg0_2_2Dcon_$fNumInt_$c+_d ;
  logic \arg0_2_2Dcon_$fNumInt_$c+_r ;
  Int_t \arg0_2_2Dcon_$fNumInt_$c+_1_d ;
  logic \arg0_2_2Dcon_$fNumInt_$c+_1_r ;
  Int_t \arg0_2_2Dcon_$fNumInt_$c+_2_d ;
  logic \arg0_2_2Dcon_$fNumInt_$c+_2_r ;
  Int_t \arg0_2_2Dcon_$fNumInt_$c+_3_d ;
  logic \arg0_2_2Dcon_$fNumInt_$c+_3_r ;
  Int_t \arg0_2_2Dcon_$fNumInt_$c+_4_d ;
  logic \arg0_2_2Dcon_$fNumInt_$c+_4_r ;
  \Int#_t  xa1lV_destruct_d;
  logic xa1lV_destruct_r;
  Int_t \arg0_2_2Dcon_$fNumInt_$c+_1I#_d ;
  logic \arg0_2_2Dcon_$fNumInt_$c+_1I#_r ;
  Int_t \arg0_2_2Dcon_$fNumInt_$c+_3I#_d ;
  logic \arg0_2_2Dcon_$fNumInt_$c+_3I#_r ;
  Int_t \arg0_2_2Dcon_$fNumInt_$c+_3I#_1_d ;
  logic \arg0_2_2Dcon_$fNumInt_$c+_3I#_1_r ;
  Int_t \arg0_2_2Dcon_$fNumInt_$c+_3I#_2_d ;
  logic \arg0_2_2Dcon_$fNumInt_$c+_3I#_2_r ;
  Int_t \arg0_2_2Dcon_$fNumInt_$c+_3I#_3_d ;
  logic \arg0_2_2Dcon_$fNumInt_$c+_3I#_3_r ;
  Int_t \arg0_2_2Dcon_$fNumInt_$c+_3I#_4_d ;
  logic \arg0_2_2Dcon_$fNumInt_$c+_3I#_4_r ;
  \Int#_t  ya1lW_destruct_d;
  logic ya1lW_destruct_r;
  Int_t \arg0_2_2Dcon_$fNumInt_$c+_3I#_1I#_d ;
  logic \arg0_2_2Dcon_$fNumInt_$c+_3I#_1I#_r ;
  \Int#_t  \arg0_2_2Dcon_$fNumInt_$c+_3I#_3I#_d ;
  logic \arg0_2_2Dcon_$fNumInt_$c+_3I#_3I#_r ;
  \Int#_t  \arg0_2_2Dcon_$fNumInt_$c+_3I#_3I#_1ya1lW_1_Add32_d ;
  logic \arg0_2_2Dcon_$fNumInt_$c+_3I#_3I#_1ya1lW_1_Add32_r ;
  Int_t \es_0_1_1I#_d ;
  logic \es_0_1_1I#_r ;
  Int_t \es_0_1_1I#_mux_d ;
  logic \es_0_1_1I#_mux_r ;
  Int_t \es_0_1_1I#_mux_mux_d ;
  logic \es_0_1_1I#_mux_mux_r ;
  Int_t \es_0_1_1I#_mux_mux_mux_d ;
  logic \es_0_1_1I#_mux_mux_mux_r ;
  MyBool_t lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_d;
  logic lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_r;
  Go_t boolConvert_1TupGo___Boolgo_1_d;
  logic boolConvert_1TupGo___Boolgo_1_r;
  Bool_t boolConvert_1TupGo___Boolbool_d;
  logic boolConvert_1TupGo___Boolbool_r;
  Bool_t bool_1_d;
  logic bool_1_r;
  Bool_t bool_2_d;
  logic bool_2_r;
  MyBool_t lizzieLet3_1_d;
  logic lizzieLet3_1_r;
  MyBool_t lizzieLet3_2_d;
  logic lizzieLet3_2_r;
  Go_t bool_1False_d;
  logic bool_1False_r;
  Go_t bool_1True_d;
  logic bool_1True_r;
  MyBool_t bool_1False_1MyFalse_d;
  logic bool_1False_1MyFalse_r;
  MyBool_t boolConvert_1_resbuf_d;
  logic boolConvert_1_resbuf_r;
  MyBool_t bool_1True_1MyTrue_d;
  logic bool_1True_1MyTrue_r;
  MyBool_t bool_1False_1MyFalsebool_1True_1MyTrue_mux_d;
  logic bool_1False_1MyFalsebool_1True_1MyTrue_mux_r;
  Go_t call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnzgo_8_d;
  logic call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnzgo_8_r;
  Pointer_QTree_Int_t call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnzwsmk_1_d;
  logic call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnzwsmk_1_r;
  Pointer_CT$wnnz_t call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnzsc_0_d;
  logic call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnzsc_0_r;
  Go_t call_$wnnz_initBufi_d;
  logic call_$wnnz_initBufi_r;
  C5_t go_8_goMux_choice_d;
  logic go_8_goMux_choice_r;
  Go_t go_8_goMux_data_d;
  logic go_8_goMux_data_r;
  Go_t call_$wnnz_unlockFork1_d;
  logic call_$wnnz_unlockFork1_r;
  Go_t call_$wnnz_unlockFork2_d;
  logic call_$wnnz_unlockFork2_r;
  Go_t call_$wnnz_unlockFork3_d;
  logic call_$wnnz_unlockFork3_r;
  Go_t call_$wnnz_initBuf_d;
  logic call_$wnnz_initBuf_r;
  Go_t call_$wnnz_goMux1_d;
  logic call_$wnnz_goMux1_r;
  Pointer_QTree_Int_t call_$wnnz_goMux2_d;
  logic call_$wnnz_goMux2_r;
  Pointer_CT$wnnz_t call_$wnnz_goMux3_d;
  logic call_$wnnz_goMux3_r;
  Go_t \call_f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf''''''''''''_f''''''''''''_Intgo_9_d ;
  logic \call_f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf''''''''''''_f''''''''''''_Intgo_9_r ;
  Pointer_QTree_Int_t \call_f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf''''''''''''_f''''''''''''_Intq4afj_d ;
  logic \call_f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf''''''''''''_f''''''''''''_Intq4afj_r ;
  Pointer_QTree_Int_t \call_f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf''''''''''''_f''''''''''''_Intt4afk_d ;
  logic \call_f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf''''''''''''_f''''''''''''_Intt4afk_r ;
  MyDTInt_Bool_t \call_f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf''''''''''''_f''''''''''''_Intis_zafl_d ;
  logic \call_f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf''''''''''''_f''''''''''''_Intis_zafl_r ;
  MyDTInt_Int_Int_t \call_f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf''''''''''''_f''''''''''''_Intop_addafm_d ;
  logic \call_f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf''''''''''''_f''''''''''''_Intop_addafm_r ;
  \Pointer_CTf''''''''''''_f''''''''''''_Int_t  \call_f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf''''''''''''_f''''''''''''_Intsc_0_1_d ;
  logic \call_f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf''''''''''''_f''''''''''''_Intsc_0_1_r ;
  Go_t \call_f''''''''''''_f''''''''''''_Int_initBufi_d ;
  logic \call_f''''''''''''_f''''''''''''_Int_initBufi_r ;
  C5_t go_9_goMux_choice_d;
  logic go_9_goMux_choice_r;
  Go_t go_9_goMux_data_d;
  logic go_9_goMux_data_r;
  Go_t \call_f''''''''''''_f''''''''''''_Int_unlockFork1_d ;
  logic \call_f''''''''''''_f''''''''''''_Int_unlockFork1_r ;
  Go_t \call_f''''''''''''_f''''''''''''_Int_unlockFork2_d ;
  logic \call_f''''''''''''_f''''''''''''_Int_unlockFork2_r ;
  Go_t \call_f''''''''''''_f''''''''''''_Int_unlockFork3_d ;
  logic \call_f''''''''''''_f''''''''''''_Int_unlockFork3_r ;
  Go_t \call_f''''''''''''_f''''''''''''_Int_unlockFork4_d ;
  logic \call_f''''''''''''_f''''''''''''_Int_unlockFork4_r ;
  Go_t \call_f''''''''''''_f''''''''''''_Int_unlockFork5_d ;
  logic \call_f''''''''''''_f''''''''''''_Int_unlockFork5_r ;
  Go_t \call_f''''''''''''_f''''''''''''_Int_unlockFork6_d ;
  logic \call_f''''''''''''_f''''''''''''_Int_unlockFork6_r ;
  Go_t \call_f''''''''''''_f''''''''''''_Int_initBuf_d ;
  logic \call_f''''''''''''_f''''''''''''_Int_initBuf_r ;
  Go_t \call_f''''''''''''_f''''''''''''_Int_goMux1_d ;
  logic \call_f''''''''''''_f''''''''''''_Int_goMux1_r ;
  Pointer_QTree_Int_t \call_f''''''''''''_f''''''''''''_Int_goMux2_d ;
  logic \call_f''''''''''''_f''''''''''''_Int_goMux2_r ;
  Pointer_QTree_Int_t \call_f''''''''''''_f''''''''''''_Int_goMux3_d ;
  logic \call_f''''''''''''_f''''''''''''_Int_goMux3_r ;
  MyDTInt_Bool_t \call_f''''''''''''_f''''''''''''_Int_goMux4_d ;
  logic \call_f''''''''''''_f''''''''''''_Int_goMux4_r ;
  MyDTInt_Int_Int_t \call_f''''''''''''_f''''''''''''_Int_goMux5_d ;
  logic \call_f''''''''''''_f''''''''''''_Int_goMux5_r ;
  \Pointer_CTf''''''''''''_f''''''''''''_Int_t  \call_f''''''''''''_f''''''''''''_Int_goMux6_d ;
  logic \call_f''''''''''''_f''''''''''''_Int_goMux6_r ;
  Go_t call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intgo_10_d;
  logic call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intgo_10_r;
  Pointer_QTree_Int_t call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intm1aeq_d;
  logic call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intm1aeq_r;
  Pointer_QTree_Int_t call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intm2aer_d;
  logic call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intm2aer_r;
  Pointer_QTree_Int_t call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intm3aes_d;
  logic call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intm3aes_r;
  MyDTInt_Bool_t call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intis_zaet_d;
  logic call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intis_zaet_r;
  MyDTInt_Int_Int_t call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intop_addaeu_d;
  logic call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intop_addaeu_r;
  Pointer_CTf_f_Int_t call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intsc_0_2_d;
  logic call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intsc_0_2_r;
  Go_t call_f_f_Int_initBufi_d;
  logic call_f_f_Int_initBufi_r;
  C5_t go_10_goMux_choice_d;
  logic go_10_goMux_choice_r;
  Go_t go_10_goMux_data_d;
  logic go_10_goMux_data_r;
  Go_t call_f_f_Int_unlockFork1_d;
  logic call_f_f_Int_unlockFork1_r;
  Go_t call_f_f_Int_unlockFork2_d;
  logic call_f_f_Int_unlockFork2_r;
  Go_t call_f_f_Int_unlockFork3_d;
  logic call_f_f_Int_unlockFork3_r;
  Go_t call_f_f_Int_unlockFork4_d;
  logic call_f_f_Int_unlockFork4_r;
  Go_t call_f_f_Int_unlockFork5_d;
  logic call_f_f_Int_unlockFork5_r;
  Go_t call_f_f_Int_unlockFork6_d;
  logic call_f_f_Int_unlockFork6_r;
  Go_t call_f_f_Int_unlockFork7_d;
  logic call_f_f_Int_unlockFork7_r;
  Go_t call_f_f_Int_initBuf_d;
  logic call_f_f_Int_initBuf_r;
  Go_t call_f_f_Int_goMux1_d;
  logic call_f_f_Int_goMux1_r;
  Pointer_QTree_Int_t call_f_f_Int_goMux2_d;
  logic call_f_f_Int_goMux2_r;
  Pointer_QTree_Int_t call_f_f_Int_goMux3_d;
  logic call_f_f_Int_goMux3_r;
  Pointer_QTree_Int_t call_f_f_Int_goMux4_d;
  logic call_f_f_Int_goMux4_r;
  MyDTInt_Bool_t call_f_f_Int_goMux5_d;
  logic call_f_f_Int_goMux5_r;
  MyDTInt_Int_Int_t call_f_f_Int_goMux6_d;
  logic call_f_f_Int_goMux6_r;
  Pointer_CTf_f_Int_t call_f_f_Int_goMux7_d;
  logic call_f_f_Int_goMux7_r;
  Int_t es_10_1MyFalse_d;
  logic es_10_1MyFalse_r;
  Int_t _255_d;
  logic _255_r;
  assign _255_r = 1'd1;
  Int_t es_10_1MyFalse_1_argbuf_d;
  logic es_10_1MyFalse_1_argbuf_r;
  MyDTInt_Int_Int_t es_10_2MyFalse_d;
  logic es_10_2MyFalse_r;
  MyDTInt_Int_Int_t _254_d;
  logic _254_r;
  assign _254_r = 1'd1;
  MyDTInt_Int_Int_t es_10_2MyFalse_1_argbuf_d;
  logic es_10_2MyFalse_1_argbuf_r;
  TupMyDTInt_Int_Int___Int___Int_t applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int6_d;
  logic applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int6_r;
  Pointer_CTf_f_Int_t es_10_3MyFalse_d;
  logic es_10_3MyFalse_r;
  Pointer_CTf_f_Int_t es_10_3MyTrue_d;
  logic es_10_3MyTrue_r;
  Pointer_CTf_f_Int_t es_10_3MyFalse_1_argbuf_d;
  logic es_10_3MyFalse_1_argbuf_r;
  Pointer_CTf_f_Int_t es_10_3MyTrue_1_argbuf_d;
  logic es_10_3MyTrue_1_argbuf_r;
  Go_t es_10_4MyFalse_d;
  logic es_10_4MyFalse_r;
  Go_t es_10_4MyTrue_d;
  logic es_10_4MyTrue_r;
  Go_t es_10_4MyFalse_1_argbuf_d;
  logic es_10_4MyFalse_1_argbuf_r;
  Go_t es_10_4MyTrue_1_d;
  logic es_10_4MyTrue_1_r;
  Go_t es_10_4MyTrue_2_d;
  logic es_10_4MyTrue_2_r;
  QTree_Int_t es_10_4MyTrue_1QNone_Int_d;
  logic es_10_4MyTrue_1QNone_Int_r;
  QTree_Int_t lizzieLet32_1_argbuf_d;
  logic lizzieLet32_1_argbuf_r;
  Go_t es_10_4MyTrue_2_argbuf_d;
  logic es_10_4MyTrue_2_argbuf_r;
  Int_t es_10_5MyFalse_d;
  logic es_10_5MyFalse_r;
  Int_t _253_d;
  logic _253_r;
  assign _253_r = 1'd1;
  Int_t es_10_5MyFalse_1_argbuf_d;
  logic es_10_5MyFalse_1_argbuf_r;
  QTree_Int_t lizzieLet31_1_argbuf_d;
  logic lizzieLet31_1_argbuf_r;
  Int_t es_14_1MyFalse_d;
  logic es_14_1MyFalse_r;
  Int_t _252_d;
  logic _252_r;
  assign _252_r = 1'd1;
  MyDTInt_Int_Int_t es_14_2MyFalse_d;
  logic es_14_2MyFalse_r;
  MyDTInt_Int_Int_t _251_d;
  logic _251_r;
  assign _251_r = 1'd1;
  Pointer_CTf_f_Int_t es_14_3MyFalse_d;
  logic es_14_3MyFalse_r;
  Pointer_CTf_f_Int_t es_14_3MyTrue_d;
  logic es_14_3MyTrue_r;
  Pointer_CTf_f_Int_t es_14_3MyTrue_1_argbuf_d;
  logic es_14_3MyTrue_1_argbuf_r;
  Go_t es_14_4MyFalse_d;
  logic es_14_4MyFalse_r;
  Go_t es_14_4MyTrue_d;
  logic es_14_4MyTrue_r;
  Go_t es_14_4MyTrue_1_argbuf_d;
  logic es_14_4MyTrue_1_argbuf_r;
  MyDTInt_Bool_t es_14_5MyFalse_d;
  logic es_14_5MyFalse_r;
  MyDTInt_Bool_t _250_d;
  logic _250_r;
  assign _250_r = 1'd1;
  QTree_Int_t es_14_6MyFalse_d;
  logic es_14_6MyFalse_r;
  QTree_Int_t _249_d;
  logic _249_r;
  assign _249_r = 1'd1;
  QTree_Int_t es_14_6MyFalse_1_d;
  logic es_14_6MyFalse_1_r;
  QTree_Int_t es_14_6MyFalse_2_d;
  logic es_14_6MyFalse_2_r;
  QTree_Int_t es_14_6MyFalse_3_d;
  logic es_14_6MyFalse_3_r;
  QTree_Int_t es_14_6MyFalse_4_d;
  logic es_14_6MyFalse_4_r;
  QTree_Int_t es_14_6MyFalse_5_d;
  logic es_14_6MyFalse_5_r;
  QTree_Int_t es_14_6MyFalse_6_d;
  logic es_14_6MyFalse_6_r;
  QTree_Int_t es_14_6MyFalse_7_d;
  logic es_14_6MyFalse_7_r;
  QTree_Int_t es_14_6MyFalse_8_d;
  logic es_14_6MyFalse_8_r;
  Int_t \v'aeR_destruct_d ;
  logic \v'aeR_destruct_r ;
  QTree_Int_t _248_d;
  logic _248_r;
  assign _248_r = 1'd1;
  QTree_Int_t es_14_6MyFalse_1QVal_Int_d;
  logic es_14_6MyFalse_1QVal_Int_r;
  QTree_Int_t _247_d;
  logic _247_r;
  assign _247_r = 1'd1;
  QTree_Int_t _246_d;
  logic _246_r;
  assign _246_r = 1'd1;
  Int_t es_14_6MyFalse_3QNone_Int_d;
  logic es_14_6MyFalse_3QNone_Int_r;
  Int_t es_14_6MyFalse_3QVal_Int_d;
  logic es_14_6MyFalse_3QVal_Int_r;
  Int_t _245_d;
  logic _245_r;
  assign _245_r = 1'd1;
  Int_t _244_d;
  logic _244_r;
  assign _244_r = 1'd1;
  Int_t es_14_6MyFalse_3QNone_Int_1_argbuf_d;
  logic es_14_6MyFalse_3QNone_Int_1_argbuf_r;
  Int_t es_14_6MyFalse_3QVal_Int_1_d;
  logic es_14_6MyFalse_3QVal_Int_1_r;
  Int_t es_14_6MyFalse_3QVal_Int_2_d;
  logic es_14_6MyFalse_3QVal_Int_2_r;
  Int_t es_14_6MyFalse_3QVal_Int_1_argbuf_d;
  logic es_14_6MyFalse_3QVal_Int_1_argbuf_r;
  MyDTInt_Int_Int_t es_14_6MyFalse_4QNone_Int_d;
  logic es_14_6MyFalse_4QNone_Int_r;
  MyDTInt_Int_Int_t es_14_6MyFalse_4QVal_Int_d;
  logic es_14_6MyFalse_4QVal_Int_r;
  MyDTInt_Int_Int_t _243_d;
  logic _243_r;
  assign _243_r = 1'd1;
  MyDTInt_Int_Int_t _242_d;
  logic _242_r;
  assign _242_r = 1'd1;
  MyDTInt_Int_Int_t es_14_6MyFalse_4QNone_Int_1_argbuf_d;
  logic es_14_6MyFalse_4QNone_Int_1_argbuf_r;
  TupMyDTInt_Int_Int___Int___Int_t applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int8_d;
  logic applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int8_r;
  MyDTInt_Int_Int_t es_14_6MyFalse_4QVal_Int_1_d;
  logic es_14_6MyFalse_4QVal_Int_1_r;
  MyDTInt_Int_Int_t es_14_6MyFalse_4QVal_Int_2_d;
  logic es_14_6MyFalse_4QVal_Int_2_r;
  MyDTInt_Int_Int_t es_14_6MyFalse_4QVal_Int_3_d;
  logic es_14_6MyFalse_4QVal_Int_3_r;
  MyDTInt_Int_Int_t es_14_6MyFalse_4QVal_Int_1_argbuf_d;
  logic es_14_6MyFalse_4QVal_Int_1_argbuf_r;
  TupMyDTInt_Int_Int___Int___Int_t applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int9_d;
  logic applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int9_r;
  MyDTInt_Int_Int_t es_14_6MyFalse_4QVal_Int_2_argbuf_d;
  logic es_14_6MyFalse_4QVal_Int_2_argbuf_r;
  TupMyDTInt_Int_Int___Int___Int_t applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int10_d;
  logic applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int10_r;
  Pointer_CTf_f_Int_t es_14_6MyFalse_5QNone_Int_d;
  logic es_14_6MyFalse_5QNone_Int_r;
  Pointer_CTf_f_Int_t es_14_6MyFalse_5QVal_Int_d;
  logic es_14_6MyFalse_5QVal_Int_r;
  Pointer_CTf_f_Int_t es_14_6MyFalse_5QNode_Int_d;
  logic es_14_6MyFalse_5QNode_Int_r;
  Pointer_CTf_f_Int_t es_14_6MyFalse_5QError_Int_d;
  logic es_14_6MyFalse_5QError_Int_r;
  Pointer_CTf_f_Int_t es_14_6MyFalse_5QError_Int_1_argbuf_d;
  logic es_14_6MyFalse_5QError_Int_1_argbuf_r;
  Pointer_CTf_f_Int_t es_14_6MyFalse_5QNode_Int_1_argbuf_d;
  logic es_14_6MyFalse_5QNode_Int_1_argbuf_r;
  Pointer_CTf_f_Int_t es_14_6MyFalse_5QNone_Int_1_argbuf_d;
  logic es_14_6MyFalse_5QNone_Int_1_argbuf_r;
  Go_t es_14_6MyFalse_6QNone_Int_d;
  logic es_14_6MyFalse_6QNone_Int_r;
  Go_t es_14_6MyFalse_6QVal_Int_d;
  logic es_14_6MyFalse_6QVal_Int_r;
  Go_t es_14_6MyFalse_6QNode_Int_d;
  logic es_14_6MyFalse_6QNode_Int_r;
  Go_t es_14_6MyFalse_6QError_Int_d;
  logic es_14_6MyFalse_6QError_Int_r;
  Go_t es_14_6MyFalse_6QError_Int_1_d;
  logic es_14_6MyFalse_6QError_Int_1_r;
  Go_t es_14_6MyFalse_6QError_Int_2_d;
  logic es_14_6MyFalse_6QError_Int_2_r;
  QTree_Int_t es_14_6MyFalse_6QError_Int_1QError_Int_d;
  logic es_14_6MyFalse_6QError_Int_1QError_Int_r;
  QTree_Int_t lizzieLet40_1_argbuf_d;
  logic lizzieLet40_1_argbuf_r;
  Go_t es_14_6MyFalse_6QError_Int_2_argbuf_d;
  logic es_14_6MyFalse_6QError_Int_2_argbuf_r;
  Go_t es_14_6MyFalse_6QNode_Int_1_d;
  logic es_14_6MyFalse_6QNode_Int_1_r;
  Go_t es_14_6MyFalse_6QNode_Int_2_d;
  logic es_14_6MyFalse_6QNode_Int_2_r;
  QTree_Int_t es_14_6MyFalse_6QNode_Int_1QError_Int_d;
  logic es_14_6MyFalse_6QNode_Int_1QError_Int_r;
  QTree_Int_t lizzieLet39_1_1_argbuf_d;
  logic lizzieLet39_1_1_argbuf_r;
  Go_t es_14_6MyFalse_6QNode_Int_2_argbuf_d;
  logic es_14_6MyFalse_6QNode_Int_2_argbuf_r;
  Go_t es_14_6MyFalse_6QNone_Int_1_argbuf_d;
  logic es_14_6MyFalse_6QNone_Int_1_argbuf_r;
  Go_t es_14_6MyFalse_6QVal_Int_1_d;
  logic es_14_6MyFalse_6QVal_Int_1_r;
  Go_t es_14_6MyFalse_6QVal_Int_2_d;
  logic es_14_6MyFalse_6QVal_Int_2_r;
  Go_t es_14_6MyFalse_6QVal_Int_1_argbuf_d;
  logic es_14_6MyFalse_6QVal_Int_1_argbuf_r;
  TupGo___MyDTInt_Bool___Int_t applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int5_d;
  logic applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int5_r;
  MyDTInt_Bool_t _241_d;
  logic _241_r;
  assign _241_r = 1'd1;
  MyDTInt_Bool_t es_14_6MyFalse_7QVal_Int_d;
  logic es_14_6MyFalse_7QVal_Int_r;
  MyDTInt_Bool_t _240_d;
  logic _240_r;
  assign _240_r = 1'd1;
  MyDTInt_Bool_t _239_d;
  logic _239_r;
  assign _239_r = 1'd1;
  MyDTInt_Bool_t es_14_6MyFalse_7QVal_Int_1_argbuf_d;
  logic es_14_6MyFalse_7QVal_Int_1_argbuf_r;
  Int_t es_14_6MyFalse_8QNone_Int_d;
  logic es_14_6MyFalse_8QNone_Int_r;
  Int_t es_14_6MyFalse_8QVal_Int_d;
  logic es_14_6MyFalse_8QVal_Int_r;
  Int_t _238_d;
  logic _238_r;
  assign _238_r = 1'd1;
  Int_t _237_d;
  logic _237_r;
  assign _237_r = 1'd1;
  Int_t es_14_6MyFalse_8QNone_Int_1_argbuf_d;
  logic es_14_6MyFalse_8QNone_Int_1_argbuf_r;
  Int_t es_14_6MyFalse_8QVal_Int_1_d;
  logic es_14_6MyFalse_8QVal_Int_1_r;
  Int_t es_14_6MyFalse_8QVal_Int_2_d;
  logic es_14_6MyFalse_8QVal_Int_2_r;
  Int_t es_14_6MyFalse_8QVal_Int_1_argbuf_d;
  logic es_14_6MyFalse_8QVal_Int_1_argbuf_r;
  Pointer_QTree_Int_t _236_d;
  logic _236_r;
  assign _236_r = 1'd1;
  Pointer_QTree_Int_t es_14_7MyTrue_d;
  logic es_14_7MyTrue_r;
  Pointer_QTree_Int_t es_14_7MyTrue_1_argbuf_d;
  logic es_14_7MyTrue_1_argbuf_r;
  Int_t es_14_8MyFalse_d;
  logic es_14_8MyFalse_r;
  Int_t _235_d;
  logic _235_r;
  assign _235_r = 1'd1;
  QTree_Int_t lizzieLet36_1_argbuf_d;
  logic lizzieLet36_1_argbuf_r;
  Int_t es_21_1MyFalse_d;
  logic es_21_1MyFalse_r;
  Int_t _234_d;
  logic _234_r;
  assign _234_r = 1'd1;
  Int_t es_21_1MyFalse_1_argbuf_d;
  logic es_21_1MyFalse_1_argbuf_r;
  MyDTInt_Int_Int_t es_21_2MyFalse_d;
  logic es_21_2MyFalse_r;
  MyDTInt_Int_Int_t _233_d;
  logic _233_r;
  assign _233_r = 1'd1;
  MyDTInt_Int_Int_t es_21_2MyFalse_1_d;
  logic es_21_2MyFalse_1_r;
  MyDTInt_Int_Int_t es_21_2MyFalse_2_d;
  logic es_21_2MyFalse_2_r;
  MyDTInt_Int_Int_t es_21_2MyFalse_1_argbuf_d;
  logic es_21_2MyFalse_1_argbuf_r;
  TupMyDTInt_Int_Int___Int___Int_t applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int11_d;
  logic applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int11_r;
  MyDTInt_Int_Int_t es_21_2MyFalse_2_argbuf_d;
  logic es_21_2MyFalse_2_argbuf_r;
  TupMyDTInt_Int_Int___Int___Int_t applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int12_d;
  logic applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int12_r;
  Pointer_CTf_f_Int_t es_21_3MyFalse_d;
  logic es_21_3MyFalse_r;
  Pointer_CTf_f_Int_t es_21_3MyTrue_d;
  logic es_21_3MyTrue_r;
  Pointer_CTf_f_Int_t es_21_3MyFalse_1_argbuf_d;
  logic es_21_3MyFalse_1_argbuf_r;
  Pointer_CTf_f_Int_t es_21_3MyTrue_1_argbuf_d;
  logic es_21_3MyTrue_1_argbuf_r;
  Go_t es_21_4MyFalse_d;
  logic es_21_4MyFalse_r;
  Go_t es_21_4MyTrue_d;
  logic es_21_4MyTrue_r;
  Go_t es_21_4MyFalse_1_argbuf_d;
  logic es_21_4MyFalse_1_argbuf_r;
  Go_t es_21_4MyTrue_1_d;
  logic es_21_4MyTrue_1_r;
  Go_t es_21_4MyTrue_2_d;
  logic es_21_4MyTrue_2_r;
  QTree_Int_t es_21_4MyTrue_1QNone_Int_d;
  logic es_21_4MyTrue_1QNone_Int_r;
  QTree_Int_t lizzieLet38_1_1_argbuf_d;
  logic lizzieLet38_1_1_argbuf_r;
  Go_t es_21_4MyTrue_2_argbuf_d;
  logic es_21_4MyTrue_2_argbuf_r;
  Int_t es_21_5MyFalse_d;
  logic es_21_5MyFalse_r;
  Int_t _232_d;
  logic _232_r;
  assign _232_r = 1'd1;
  Int_t es_21_5MyFalse_1_argbuf_d;
  logic es_21_5MyFalse_1_argbuf_r;
  Int_t es_21_6MyFalse_d;
  logic es_21_6MyFalse_r;
  Int_t _231_d;
  logic _231_r;
  assign _231_r = 1'd1;
  Int_t es_21_6MyFalse_1_argbuf_d;
  logic es_21_6MyFalse_1_argbuf_r;
  QTree_Int_t lizzieLet37_2_1_argbuf_d;
  logic lizzieLet37_2_1_argbuf_r;
  QTree_Int_t lizzieLet46_1_argbuf_d;
  logic lizzieLet46_1_argbuf_r;
  Go_t es_2_1MyFalse_d;
  logic es_2_1MyFalse_r;
  Go_t es_2_1MyTrue_d;
  logic es_2_1MyTrue_r;
  Go_t es_2_1MyFalse_1_argbuf_d;
  logic es_2_1MyFalse_1_argbuf_r;
  Go_t es_2_1MyTrue_1_d;
  logic es_2_1MyTrue_1_r;
  Go_t es_2_1MyTrue_2_d;
  logic es_2_1MyTrue_2_r;
  QTree_Int_t es_2_1MyTrue_1QNone_Int_d;
  logic es_2_1MyTrue_1QNone_Int_r;
  QTree_Int_t lizzieLet9_1_argbuf_d;
  logic lizzieLet9_1_argbuf_r;
  Go_t es_2_1MyTrue_2_argbuf_d;
  logic es_2_1MyTrue_2_argbuf_r;
  MyDTInt_Int_Int_t es_2_1_1MyFalse_d;
  logic es_2_1_1MyFalse_r;
  MyDTInt_Int_Int_t _230_d;
  logic _230_r;
  assign _230_r = 1'd1;
  MyDTInt_Int_Int_t es_2_1_1MyFalse_1_argbuf_d;
  logic es_2_1_1MyFalse_1_argbuf_r;
  TupMyDTInt_Int_Int___Int___Int_t applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int2_d;
  logic applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int2_r;
  Pointer_CTf_f_Int_t es_2_1_2MyFalse_d;
  logic es_2_1_2MyFalse_r;
  Pointer_CTf_f_Int_t es_2_1_2MyTrue_d;
  logic es_2_1_2MyTrue_r;
  Pointer_CTf_f_Int_t es_2_1_2MyFalse_1_argbuf_d;
  logic es_2_1_2MyFalse_1_argbuf_r;
  Pointer_CTf_f_Int_t es_2_1_2MyTrue_1_argbuf_d;
  logic es_2_1_2MyTrue_1_argbuf_r;
  Go_t es_2_1_3MyFalse_d;
  logic es_2_1_3MyFalse_r;
  Go_t es_2_1_3MyTrue_d;
  logic es_2_1_3MyTrue_r;
  Go_t es_2_1_3MyFalse_1_argbuf_d;
  logic es_2_1_3MyFalse_1_argbuf_r;
  Go_t es_2_1_3MyTrue_1_d;
  logic es_2_1_3MyTrue_1_r;
  Go_t es_2_1_3MyTrue_2_d;
  logic es_2_1_3MyTrue_2_r;
  QTree_Int_t es_2_1_3MyTrue_1QNone_Int_d;
  logic es_2_1_3MyTrue_1QNone_Int_r;
  QTree_Int_t lizzieLet21_1_argbuf_d;
  logic lizzieLet21_1_argbuf_r;
  Go_t es_2_1_3MyTrue_2_argbuf_d;
  logic es_2_1_3MyTrue_2_argbuf_r;
  Int_t es_2_1_4MyFalse_d;
  logic es_2_1_4MyFalse_r;
  Int_t _229_d;
  logic _229_r;
  assign _229_r = 1'd1;
  Int_t es_2_1_4MyFalse_1_argbuf_d;
  logic es_2_1_4MyFalse_1_argbuf_r;
  Int_t es_2_1_5MyFalse_d;
  logic es_2_1_5MyFalse_r;
  Int_t _228_d;
  logic _228_r;
  assign _228_r = 1'd1;
  Int_t es_2_1_5MyFalse_1_argbuf_d;
  logic es_2_1_5MyFalse_1_argbuf_r;
  MyDTInt_Int_Int_t es_2_2MyFalse_d;
  logic es_2_2MyFalse_r;
  MyDTInt_Int_Int_t _227_d;
  logic _227_r;
  assign _227_r = 1'd1;
  MyDTInt_Int_Int_t es_2_2MyFalse_1_argbuf_d;
  logic es_2_2MyFalse_1_argbuf_r;
  TupMyDTInt_Int_Int___Int___Int_t applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int4_d;
  logic applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int4_r;
  \Pointer_CTf''''''''''''_f''''''''''''_Int_t  es_2_3MyFalse_d;
  logic es_2_3MyFalse_r;
  \Pointer_CTf''''''''''''_f''''''''''''_Int_t  es_2_3MyTrue_d;
  logic es_2_3MyTrue_r;
  \Pointer_CTf''''''''''''_f''''''''''''_Int_t  es_2_3MyFalse_1_argbuf_d;
  logic es_2_3MyFalse_1_argbuf_r;
  \Pointer_CTf''''''''''''_f''''''''''''_Int_t  es_2_3MyTrue_1_argbuf_d;
  logic es_2_3MyTrue_1_argbuf_r;
  Int_t es_2_4MyFalse_d;
  logic es_2_4MyFalse_r;
  Int_t _226_d;
  logic _226_r;
  assign _226_r = 1'd1;
  Int_t es_2_4MyFalse_1_argbuf_d;
  logic es_2_4MyFalse_1_argbuf_r;
  Int_t es_2_5MyFalse_d;
  logic es_2_5MyFalse_r;
  Int_t _225_d;
  logic _225_r;
  assign _225_r = 1'd1;
  Int_t es_2_5MyFalse_1_argbuf_d;
  logic es_2_5MyFalse_1_argbuf_r;
  QTree_Int_t lizzieLet50_1_argbuf_d;
  logic lizzieLet50_1_argbuf_r;
  QTree_Int_t lizzieLet8_1_argbuf_d;
  logic lizzieLet8_1_argbuf_r;
  QTree_Int_t lizzieLet20_1_argbuf_d;
  logic lizzieLet20_1_argbuf_r;
  QTree_Int_t lizzieLet26_1_argbuf_d;
  logic lizzieLet26_1_argbuf_r;
  \Int#_t  contRet_0_1_argbuf_d;
  logic contRet_0_1_argbuf_r;
  \Int#_t  es_4_2_1lizzieLet58_4Lcall_$wnnz0_1_Add32_d;
  logic es_4_2_1lizzieLet58_4Lcall_$wnnz0_1_Add32_r;
  C12_t \f''''''''''''_f''''''''''''_Int_choice_d ;
  logic \f''''''''''''_f''''''''''''_Int_choice_r ;
  TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_t \f''''''''''''_f''''''''''''_Int_data_d ;
  logic \f''''''''''''_f''''''''''''_Int_data_r ;
  Go_t go_11_1_d;
  logic go_11_1_r;
  Go_t go_11_2_d;
  logic go_11_2_r;
  MyDTInt_Bool_t is_zafl_1_1_argbuf_d;
  logic is_zafl_1_1_argbuf_r;
  MyDTInt_Int_Int_t op_addafm_1_1_argbuf_d;
  logic op_addafm_1_1_argbuf_r;
  Pointer_QTree_Int_t q4afj_1_1_argbuf_d;
  logic q4afj_1_1_argbuf_r;
  Pointer_QTree_Int_t t4afk_1_1_argbuf_d;
  logic t4afk_1_1_argbuf_r;
  Pointer_QTree_Int_t \f''''''''''''_f''''''''''''_Int_resbuf_d ;
  logic \f''''''''''''_f''''''''''''_Int_resbuf_r ;
  Pointer_QTree_Int_t \f''''''''''''_f''''''''''''_Int_10_argbuf_d ;
  logic \f''''''''''''_f''''''''''''_Int_10_argbuf_r ;
  Pointer_QTree_Int_t \f''''''''''''_f''''''''''''_Int_11_argbuf_d ;
  logic \f''''''''''''_f''''''''''''_Int_11_argbuf_r ;
  Pointer_QTree_Int_t \f''''''''''''_f''''''''''''_Int_12_argbuf_d ;
  logic \f''''''''''''_f''''''''''''_Int_12_argbuf_r ;
  QTree_Int_t es_30_1es_31_1es_32_1es_33_1QNode_Int_d;
  logic es_30_1es_31_1es_32_1es_33_1QNode_Int_r;
  Pointer_QTree_Int_t \f''''''''''''_f''''''''''''_Int_2_argbuf_d ;
  logic \f''''''''''''_f''''''''''''_Int_2_argbuf_r ;
  Pointer_QTree_Int_t \f''''''''''''_f''''''''''''_Int_3_argbuf_d ;
  logic \f''''''''''''_f''''''''''''_Int_3_argbuf_r ;
  Pointer_QTree_Int_t \f''''''''''''_f''''''''''''_Int_4_argbuf_d ;
  logic \f''''''''''''_f''''''''''''_Int_4_argbuf_r ;
  QTree_Int_t es_4_1_1es_5_1_1es_6_1_1es_7_1QNode_Int_d;
  logic es_4_1_1es_5_1_1es_6_1_1es_7_1QNode_Int_r;
  Pointer_QTree_Int_t \f''''''''''''_f''''''''''''_Int_5_argbuf_d ;
  logic \f''''''''''''_f''''''''''''_Int_5_argbuf_r ;
  Pointer_QTree_Int_t \f''''''''''''_f''''''''''''_Int_6_argbuf_d ;
  logic \f''''''''''''_f''''''''''''_Int_6_argbuf_r ;
  Pointer_QTree_Int_t \f''''''''''''_f''''''''''''_Int_7_argbuf_d ;
  logic \f''''''''''''_f''''''''''''_Int_7_argbuf_r ;
  Pointer_QTree_Int_t \f''''''''''''_f''''''''''''_Int_8_argbuf_d ;
  logic \f''''''''''''_f''''''''''''_Int_8_argbuf_r ;
  QTree_Int_t es_26_1es_27_1es_28_1es_29_1QNode_Int_d;
  logic es_26_1es_27_1es_28_1es_29_1QNode_Int_r;
  Pointer_QTree_Int_t \f''''''''''''_f''''''''''''_Int_9_argbuf_d ;
  logic \f''''''''''''_f''''''''''''_Int_9_argbuf_r ;
  Pointer_QTree_Int_t \f''''''''''''_f''''''''''''_Int_1_d ;
  logic \f''''''''''''_f''''''''''''_Int_1_r ;
  Pointer_QTree_Int_t \f''''''''''''_f''''''''''''_Int_2_d ;
  logic \f''''''''''''_f''''''''''''_Int_2_r ;
  Pointer_QTree_Int_t \f''''''''''''_f''''''''''''_Int_3_d ;
  logic \f''''''''''''_f''''''''''''_Int_3_r ;
  Pointer_QTree_Int_t \f''''''''''''_f''''''''''''_Int_4_d ;
  logic \f''''''''''''_f''''''''''''_Int_4_r ;
  Pointer_QTree_Int_t \f''''''''''''_f''''''''''''_Int_5_d ;
  logic \f''''''''''''_f''''''''''''_Int_5_r ;
  Pointer_QTree_Int_t \f''''''''''''_f''''''''''''_Int_6_d ;
  logic \f''''''''''''_f''''''''''''_Int_6_r ;
  Pointer_QTree_Int_t \f''''''''''''_f''''''''''''_Int_7_d ;
  logic \f''''''''''''_f''''''''''''_Int_7_r ;
  Pointer_QTree_Int_t \f''''''''''''_f''''''''''''_Int_8_d ;
  logic \f''''''''''''_f''''''''''''_Int_8_r ;
  Pointer_QTree_Int_t \f''''''''''''_f''''''''''''_Int_9_d ;
  logic \f''''''''''''_f''''''''''''_Int_9_r ;
  Pointer_QTree_Int_t \f''''''''''''_f''''''''''''_Int_10_d ;
  logic \f''''''''''''_f''''''''''''_Int_10_r ;
  Pointer_QTree_Int_t \f''''''''''''_f''''''''''''_Int_11_d ;
  logic \f''''''''''''_f''''''''''''_Int_11_r ;
  Pointer_QTree_Int_t \f''''''''''''_f''''''''''''_Int_12_d ;
  logic \f''''''''''''_f''''''''''''_Int_12_r ;
  Go_t \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intgo_11_d ;
  logic \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intgo_11_r ;
  Pointer_QTree_Int_t \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intq4afj_1_d ;
  logic \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intq4afj_1_r ;
  Pointer_QTree_Int_t \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intt4afk_1_d ;
  logic \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intt4afk_1_r ;
  MyDTInt_Bool_t \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zafl_1_d ;
  logic \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zafl_1_r ;
  MyDTInt_Int_Int_t \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addafm_1_d ;
  logic \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addafm_1_r ;
  Go_t f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intgo_12_d;
  logic f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intgo_12_r;
  Pointer_QTree_Int_t f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm1aeq_1_d;
  logic f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm1aeq_1_r;
  Pointer_QTree_Int_t f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm2aer_1_d;
  logic f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm2aer_1_r;
  Pointer_QTree_Int_t f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm3aes_1_d;
  logic f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm3aes_1_r;
  MyDTInt_Bool_t f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zaet_1_d;
  logic f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zaet_1_r;
  MyDTInt_Int_Int_t f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addaeu_1_d;
  logic f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addaeu_1_r;
  Go_t go_12_1_d;
  logic go_12_1_r;
  Go_t go_12_2_d;
  logic go_12_2_r;
  MyDTInt_Bool_t is_zaet_1_1_argbuf_d;
  logic is_zaet_1_1_argbuf_r;
  Pointer_QTree_Int_t m1aeq_1_1_argbuf_d;
  logic m1aeq_1_1_argbuf_r;
  Pointer_QTree_Int_t m2aer_1_1_argbuf_d;
  logic m2aer_1_1_argbuf_r;
  Pointer_QTree_Int_t m3aes_1_1_argbuf_d;
  logic m3aes_1_1_argbuf_r;
  MyDTInt_Int_Int_t op_addaeu_1_1_argbuf_d;
  logic op_addaeu_1_1_argbuf_r;
  Pointer_QTree_Int_t es_0_1_argbuf_d;
  logic es_0_1_argbuf_r;
  MyDTInt_Int_Int_t \go_1Dcon_$fNumInt_$c+_d ;
  logic \go_1Dcon_$fNumInt_$c+_r ;
  C5_t go_10_goMux_choice_1_d;
  logic go_10_goMux_choice_1_r;
  C5_t go_10_goMux_choice_2_d;
  logic go_10_goMux_choice_2_r;
  C5_t go_10_goMux_choice_3_d;
  logic go_10_goMux_choice_3_r;
  C5_t go_10_goMux_choice_4_d;
  logic go_10_goMux_choice_4_r;
  C5_t go_10_goMux_choice_5_d;
  logic go_10_goMux_choice_5_r;
  C5_t go_10_goMux_choice_6_d;
  logic go_10_goMux_choice_6_r;
  Pointer_QTree_Int_t m1aeq_goMux_mux_d;
  logic m1aeq_goMux_mux_r;
  Pointer_QTree_Int_t m2aer_goMux_mux_d;
  logic m2aer_goMux_mux_r;
  Pointer_QTree_Int_t m3aes_goMux_mux_d;
  logic m3aes_goMux_mux_r;
  MyDTInt_Bool_t is_zaet_goMux_mux_d;
  logic is_zaet_goMux_mux_r;
  MyDTInt_Int_Int_t op_addaeu_goMux_mux_d;
  logic op_addaeu_goMux_mux_r;
  Pointer_CTf_f_Int_t sc_0_2_goMux_mux_d;
  logic sc_0_2_goMux_mux_r;
  \CTf''''''''''''_f''''''''''''_Int_t  \go_11_1Lf''''''''''''_f''''''''''''_Intsbos_d ;
  logic \go_11_1Lf''''''''''''_f''''''''''''_Intsbos_r ;
  \CTf''''''''''''_f''''''''''''_Int_t  lizzieLet56_1_argbuf_d;
  logic lizzieLet56_1_argbuf_r;
  Go_t go_11_2_argbuf_d;
  logic go_11_2_argbuf_r;
  \TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf''''''''''''_f''''''''''''_Int_t  \call_f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf''''''''''''_f''''''''''''_Int_1_d ;
  logic \call_f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf''''''''''''_f''''''''''''_Int_1_r ;
  CTf_f_Int_t go_12_1Lf_f_Intsbos_d;
  logic go_12_1Lf_f_Intsbos_r;
  CTf_f_Int_t lizzieLet57_1_argbuf_d;
  logic lizzieLet57_1_argbuf_r;
  Go_t go_12_2_argbuf_d;
  logic go_12_2_argbuf_r;
  TupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_t call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_1_d;
  logic call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_1_r;
  C4_t go_13_goMux_choice_1_d;
  logic go_13_goMux_choice_1_r;
  C4_t go_13_goMux_choice_2_d;
  logic go_13_goMux_choice_2_r;
  \Int#_t  srtarg_0_goMux_mux_d;
  logic srtarg_0_goMux_mux_r;
  Pointer_CT$wnnz_t scfarg_0_goMux_mux_d;
  logic scfarg_0_goMux_mux_r;
  C11_t go_14_goMux_choice_1_d;
  logic go_14_goMux_choice_1_r;
  C11_t go_14_goMux_choice_2_d;
  logic go_14_goMux_choice_2_r;
  Pointer_QTree_Int_t srtarg_0_1_goMux_mux_d;
  logic srtarg_0_1_goMux_mux_r;
  \Pointer_CTf''''''''''''_f''''''''''''_Int_t  scfarg_0_1_goMux_mux_d;
  logic scfarg_0_1_goMux_mux_r;
  C35_t go_15_goMux_choice_1_d;
  logic go_15_goMux_choice_1_r;
  C35_t go_15_goMux_choice_2_d;
  logic go_15_goMux_choice_2_r;
  Pointer_QTree_Int_t srtarg_0_2_goMux_mux_d;
  logic srtarg_0_2_goMux_mux_r;
  Pointer_CTf_f_Int_t scfarg_0_2_goMux_mux_d;
  logic scfarg_0_2_goMux_mux_r;
  MyDTInt_Int_Int_t es_5_1_argbuf_d;
  logic es_5_1_argbuf_r;
  MyDTInt_Bool_t go_2Dcon_isZ_d;
  logic go_2Dcon_isZ_r;
  MyDTInt_Bool_t es_4_1_argbuf_d;
  logic es_4_1_argbuf_r;
  Go_t go_3_argbuf_d;
  logic go_3_argbuf_r;
  TupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_t f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_d;
  logic f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_r;
  Go_t go_4_argbuf_d;
  logic go_4_argbuf_r;
  TupGo___Pointer_QTree_Int_t \$wnnzTupGo___Pointer_QTree_Int_1_d ;
  logic \$wnnzTupGo___Pointer_QTree_Int_1_r ;
  CT$wnnz_t go_6_1L$wnnzsbos_d;
  logic go_6_1L$wnnzsbos_r;
  CT$wnnz_t lizzieLet0_1_argbuf_d;
  logic lizzieLet0_1_argbuf_r;
  Go_t go_6_2_argbuf_d;
  logic go_6_2_argbuf_r;
  TupGo___Pointer_QTree_Int___Pointer_CT$wnnz_t call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_1_d;
  logic call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_1_r;
  C5_t go_8_goMux_choice_1_d;
  logic go_8_goMux_choice_1_r;
  C5_t go_8_goMux_choice_2_d;
  logic go_8_goMux_choice_2_r;
  Pointer_QTree_Int_t wsmk_1_goMux_mux_d;
  logic wsmk_1_goMux_mux_r;
  Pointer_CT$wnnz_t sc_0_goMux_mux_d;
  logic sc_0_goMux_mux_r;
  C5_t go_9_goMux_choice_1_d;
  logic go_9_goMux_choice_1_r;
  C5_t go_9_goMux_choice_2_d;
  logic go_9_goMux_choice_2_r;
  C5_t go_9_goMux_choice_3_d;
  logic go_9_goMux_choice_3_r;
  C5_t go_9_goMux_choice_4_d;
  logic go_9_goMux_choice_4_r;
  C5_t go_9_goMux_choice_5_d;
  logic go_9_goMux_choice_5_r;
  Pointer_QTree_Int_t q4afj_goMux_mux_d;
  logic q4afj_goMux_mux_r;
  Pointer_QTree_Int_t t4afk_goMux_mux_d;
  logic t4afk_goMux_mux_r;
  MyDTInt_Bool_t is_zafl_goMux_mux_d;
  logic is_zafl_goMux_mux_r;
  MyDTInt_Int_Int_t op_addafm_goMux_mux_d;
  logic op_addafm_goMux_mux_r;
  \Pointer_CTf''''''''''''_f''''''''''''_Int_t  sc_0_1_goMux_mux_d;
  logic sc_0_1_goMux_mux_r;
  MyDTInt_Bool_t is_zaet_2_2_argbuf_d;
  logic is_zaet_2_2_argbuf_r;
  MyDTInt_Bool_t is_zaet_2_1_d;
  logic is_zaet_2_1_r;
  MyDTInt_Bool_t is_zaet_2_2_d;
  logic is_zaet_2_2_r;
  MyDTInt_Bool_t is_zaet_3_2_argbuf_d;
  logic is_zaet_3_2_argbuf_r;
  MyDTInt_Bool_t is_zaet_3_1_d;
  logic is_zaet_3_1_r;
  MyDTInt_Bool_t is_zaet_3_2_d;
  logic is_zaet_3_2_r;
  MyDTInt_Bool_t is_zaet_4_1_argbuf_d;
  logic is_zaet_4_1_argbuf_r;
  MyDTInt_Bool_t is_zafl_2_2_argbuf_d;
  logic is_zafl_2_2_argbuf_r;
  MyDTInt_Bool_t is_zafl_2_1_d;
  logic is_zafl_2_1_r;
  MyDTInt_Bool_t is_zafl_2_2_d;
  logic is_zafl_2_2_r;
  MyDTInt_Bool_t is_zafl_3_2_argbuf_d;
  logic is_zafl_3_2_argbuf_r;
  MyDTInt_Bool_t is_zafl_3_1_d;
  logic is_zafl_3_1_r;
  MyDTInt_Bool_t is_zafl_3_2_d;
  logic is_zafl_3_2_r;
  MyDTInt_Bool_t is_zafl_4_1_argbuf_d;
  logic is_zafl_4_1_argbuf_r;
  MyDTInt_Int_Int_t lizzieLet17_10QNone_Int_d;
  logic lizzieLet17_10QNone_Int_r;
  MyDTInt_Int_Int_t lizzieLet17_10QVal_Int_d;
  logic lizzieLet17_10QVal_Int_r;
  MyDTInt_Int_Int_t lizzieLet17_10QNode_Int_d;
  logic lizzieLet17_10QNode_Int_r;
  MyDTInt_Int_Int_t _224_d;
  logic _224_r;
  assign _224_r = 1'd1;
  Pointer_CTf_f_Int_t lizzieLet17_11QNone_Int_d;
  logic lizzieLet17_11QNone_Int_r;
  Pointer_CTf_f_Int_t lizzieLet17_11QVal_Int_d;
  logic lizzieLet17_11QVal_Int_r;
  Pointer_CTf_f_Int_t lizzieLet17_11QNode_Int_d;
  logic lizzieLet17_11QNode_Int_r;
  Pointer_CTf_f_Int_t lizzieLet17_11QError_Int_d;
  logic lizzieLet17_11QError_Int_r;
  Pointer_CTf_f_Int_t lizzieLet17_11QError_Int_1_argbuf_d;
  logic lizzieLet17_11QError_Int_1_argbuf_r;
  Pointer_QTree_Int_t q1af0_destruct_d;
  logic q1af0_destruct_r;
  Pointer_QTree_Int_t q2af1_destruct_d;
  logic q2af1_destruct_r;
  Pointer_QTree_Int_t q3af2_destruct_d;
  logic q3af2_destruct_r;
  Pointer_QTree_Int_t q4af3_destruct_d;
  logic q4af3_destruct_r;
  Int_t v1aeK_destruct_d;
  logic v1aeK_destruct_r;
  QTree_Int_t _223_d;
  logic _223_r;
  assign _223_r = 1'd1;
  QTree_Int_t lizzieLet17_1QVal_Int_d;
  logic lizzieLet17_1QVal_Int_r;
  QTree_Int_t lizzieLet17_1QNode_Int_d;
  logic lizzieLet17_1QNode_Int_r;
  QTree_Int_t _222_d;
  logic _222_r;
  assign _222_r = 1'd1;
  Go_t lizzieLet17_3QNone_Int_d;
  logic lizzieLet17_3QNone_Int_r;
  Go_t lizzieLet17_3QVal_Int_d;
  logic lizzieLet17_3QVal_Int_r;
  Go_t lizzieLet17_3QNode_Int_d;
  logic lizzieLet17_3QNode_Int_r;
  Go_t lizzieLet17_3QError_Int_d;
  logic lizzieLet17_3QError_Int_r;
  Go_t lizzieLet17_3QError_Int_1_d;
  logic lizzieLet17_3QError_Int_1_r;
  Go_t lizzieLet17_3QError_Int_2_d;
  logic lizzieLet17_3QError_Int_2_r;
  QTree_Int_t lizzieLet17_3QError_Int_1QError_Int_d;
  logic lizzieLet17_3QError_Int_1QError_Int_r;
  QTree_Int_t lizzieLet55_1_argbuf_d;
  logic lizzieLet55_1_argbuf_r;
  Go_t lizzieLet17_3QError_Int_2_argbuf_d;
  logic lizzieLet17_3QError_Int_2_argbuf_r;
  MyDTInt_Bool_t lizzieLet17_4QNone_Int_d;
  logic lizzieLet17_4QNone_Int_r;
  MyDTInt_Bool_t lizzieLet17_4QVal_Int_d;
  logic lizzieLet17_4QVal_Int_r;
  MyDTInt_Bool_t lizzieLet17_4QNode_Int_d;
  logic lizzieLet17_4QNode_Int_r;
  MyDTInt_Bool_t _221_d;
  logic _221_r;
  assign _221_r = 1'd1;
  QTree_Int_t lizzieLet17_5QNone_Int_d;
  logic lizzieLet17_5QNone_Int_r;
  QTree_Int_t lizzieLet17_5QVal_Int_d;
  logic lizzieLet17_5QVal_Int_r;
  QTree_Int_t lizzieLet17_5QNode_Int_d;
  logic lizzieLet17_5QNode_Int_r;
  QTree_Int_t _220_d;
  logic _220_r;
  assign _220_r = 1'd1;
  QTree_Int_t lizzieLet17_5QNode_Int_1_d;
  logic lizzieLet17_5QNode_Int_1_r;
  QTree_Int_t lizzieLet17_5QNode_Int_2_d;
  logic lizzieLet17_5QNode_Int_2_r;
  QTree_Int_t lizzieLet17_5QNode_Int_3_d;
  logic lizzieLet17_5QNode_Int_3_r;
  QTree_Int_t lizzieLet17_5QNode_Int_4_d;
  logic lizzieLet17_5QNode_Int_4_r;
  QTree_Int_t lizzieLet17_5QNode_Int_5_d;
  logic lizzieLet17_5QNode_Int_5_r;
  QTree_Int_t lizzieLet17_5QNode_Int_6_d;
  logic lizzieLet17_5QNode_Int_6_r;
  QTree_Int_t lizzieLet17_5QNode_Int_7_d;
  logic lizzieLet17_5QNode_Int_7_r;
  QTree_Int_t lizzieLet17_5QNode_Int_8_d;
  logic lizzieLet17_5QNode_Int_8_r;
  QTree_Int_t lizzieLet17_5QNode_Int_9_d;
  logic lizzieLet17_5QNode_Int_9_r;
  QTree_Int_t lizzieLet17_5QNode_Int_10_d;
  logic lizzieLet17_5QNode_Int_10_r;
  QTree_Int_t lizzieLet17_5QNode_Int_11_d;
  logic lizzieLet17_5QNode_Int_11_r;
  QTree_Int_t lizzieLet17_5QNode_Int_12_d;
  logic lizzieLet17_5QNode_Int_12_r;
  Pointer_QTree_Int_t lizzieLet17_5QNode_Int_10QNone_Int_d;
  logic lizzieLet17_5QNode_Int_10QNone_Int_r;
  Pointer_QTree_Int_t _219_d;
  logic _219_r;
  assign _219_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet17_5QNode_Int_10QNode_Int_d;
  logic lizzieLet17_5QNode_Int_10QNode_Int_r;
  Pointer_QTree_Int_t _218_d;
  logic _218_r;
  assign _218_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet17_5QNode_Int_11QNone_Int_d;
  logic lizzieLet17_5QNode_Int_11QNone_Int_r;
  Pointer_QTree_Int_t _217_d;
  logic _217_r;
  assign _217_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet17_5QNode_Int_11QNode_Int_d;
  logic lizzieLet17_5QNode_Int_11QNode_Int_r;
  Pointer_QTree_Int_t _216_d;
  logic _216_r;
  assign _216_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet17_5QNode_Int_12QNone_Int_d;
  logic lizzieLet17_5QNode_Int_12QNone_Int_r;
  Pointer_QTree_Int_t _215_d;
  logic _215_r;
  assign _215_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet17_5QNode_Int_12QNode_Int_d;
  logic lizzieLet17_5QNode_Int_12QNode_Int_r;
  Pointer_QTree_Int_t _214_d;
  logic _214_r;
  assign _214_r = 1'd1;
  Pointer_QTree_Int_t t1afa_destruct_d;
  logic t1afa_destruct_r;
  Pointer_QTree_Int_t t2afb_destruct_d;
  logic t2afb_destruct_r;
  Pointer_QTree_Int_t t3afc_destruct_d;
  logic t3afc_destruct_r;
  Pointer_QTree_Int_t t4afd_destruct_d;
  logic t4afd_destruct_r;
  QTree_Int_t _213_d;
  logic _213_r;
  assign _213_r = 1'd1;
  QTree_Int_t _212_d;
  logic _212_r;
  assign _212_r = 1'd1;
  QTree_Int_t lizzieLet17_5QNode_Int_1QNode_Int_d;
  logic lizzieLet17_5QNode_Int_1QNode_Int_r;
  QTree_Int_t _211_d;
  logic _211_r;
  assign _211_r = 1'd1;
  MyDTInt_Int_Int_t lizzieLet17_5QNode_Int_3QNone_Int_d;
  logic lizzieLet17_5QNode_Int_3QNone_Int_r;
  MyDTInt_Int_Int_t _210_d;
  logic _210_r;
  assign _210_r = 1'd1;
  MyDTInt_Int_Int_t lizzieLet17_5QNode_Int_3QNode_Int_d;
  logic lizzieLet17_5QNode_Int_3QNode_Int_r;
  MyDTInt_Int_Int_t _209_d;
  logic _209_r;
  assign _209_r = 1'd1;
  Pointer_CTf_f_Int_t lizzieLet17_5QNode_Int_4QNone_Int_d;
  logic lizzieLet17_5QNode_Int_4QNone_Int_r;
  Pointer_CTf_f_Int_t lizzieLet17_5QNode_Int_4QVal_Int_d;
  logic lizzieLet17_5QNode_Int_4QVal_Int_r;
  Pointer_CTf_f_Int_t lizzieLet17_5QNode_Int_4QNode_Int_d;
  logic lizzieLet17_5QNode_Int_4QNode_Int_r;
  Pointer_CTf_f_Int_t lizzieLet17_5QNode_Int_4QError_Int_d;
  logic lizzieLet17_5QNode_Int_4QError_Int_r;
  Pointer_CTf_f_Int_t lizzieLet17_5QNode_Int_4QError_Int_1_argbuf_d;
  logic lizzieLet17_5QNode_Int_4QError_Int_1_argbuf_r;
  Pointer_CTf_f_Int_t lizzieLet17_5QNode_Int_4QVal_Int_1_argbuf_d;
  logic lizzieLet17_5QNode_Int_4QVal_Int_1_argbuf_r;
  Go_t lizzieLet17_5QNode_Int_5QNone_Int_d;
  logic lizzieLet17_5QNode_Int_5QNone_Int_r;
  Go_t lizzieLet17_5QNode_Int_5QVal_Int_d;
  logic lizzieLet17_5QNode_Int_5QVal_Int_r;
  Go_t lizzieLet17_5QNode_Int_5QNode_Int_d;
  logic lizzieLet17_5QNode_Int_5QNode_Int_r;
  Go_t lizzieLet17_5QNode_Int_5QError_Int_d;
  logic lizzieLet17_5QNode_Int_5QError_Int_r;
  Go_t lizzieLet17_5QNode_Int_5QError_Int_1_d;
  logic lizzieLet17_5QNode_Int_5QError_Int_1_r;
  Go_t lizzieLet17_5QNode_Int_5QError_Int_2_d;
  logic lizzieLet17_5QNode_Int_5QError_Int_2_r;
  QTree_Int_t lizzieLet17_5QNode_Int_5QError_Int_1QError_Int_d;
  logic lizzieLet17_5QNode_Int_5QError_Int_1QError_Int_r;
  QTree_Int_t lizzieLet54_1_argbuf_d;
  logic lizzieLet54_1_argbuf_r;
  Go_t lizzieLet17_5QNode_Int_5QError_Int_2_argbuf_d;
  logic lizzieLet17_5QNode_Int_5QError_Int_2_argbuf_r;
  Go_t lizzieLet17_5QNode_Int_5QVal_Int_1_d;
  logic lizzieLet17_5QNode_Int_5QVal_Int_1_r;
  Go_t lizzieLet17_5QNode_Int_5QVal_Int_2_d;
  logic lizzieLet17_5QNode_Int_5QVal_Int_2_r;
  QTree_Int_t lizzieLet17_5QNode_Int_5QVal_Int_1QError_Int_d;
  logic lizzieLet17_5QNode_Int_5QVal_Int_1QError_Int_r;
  QTree_Int_t lizzieLet48_1_argbuf_d;
  logic lizzieLet48_1_argbuf_r;
  Go_t lizzieLet17_5QNode_Int_5QVal_Int_2_argbuf_d;
  logic lizzieLet17_5QNode_Int_5QVal_Int_2_argbuf_r;
  MyDTInt_Bool_t lizzieLet17_5QNode_Int_6QNone_Int_d;
  logic lizzieLet17_5QNode_Int_6QNone_Int_r;
  MyDTInt_Bool_t _208_d;
  logic _208_r;
  assign _208_r = 1'd1;
  MyDTInt_Bool_t lizzieLet17_5QNode_Int_6QNode_Int_d;
  logic lizzieLet17_5QNode_Int_6QNode_Int_r;
  MyDTInt_Bool_t _207_d;
  logic _207_r;
  assign _207_r = 1'd1;
  QTree_Int_t lizzieLet17_5QNode_Int_7QNone_Int_d;
  logic lizzieLet17_5QNode_Int_7QNone_Int_r;
  QTree_Int_t _206_d;
  logic _206_r;
  assign _206_r = 1'd1;
  QTree_Int_t lizzieLet17_5QNode_Int_7QNode_Int_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_r;
  QTree_Int_t _205_d;
  logic _205_r;
  assign _205_r = 1'd1;
  QTree_Int_t lizzieLet17_5QNode_Int_7QNode_Int_1_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_1_r;
  QTree_Int_t lizzieLet17_5QNode_Int_7QNode_Int_2_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_2_r;
  QTree_Int_t lizzieLet17_5QNode_Int_7QNode_Int_3_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_3_r;
  QTree_Int_t lizzieLet17_5QNode_Int_7QNode_Int_4_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_4_r;
  QTree_Int_t lizzieLet17_5QNode_Int_7QNode_Int_5_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_5_r;
  QTree_Int_t lizzieLet17_5QNode_Int_7QNode_Int_6_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_6_r;
  QTree_Int_t lizzieLet17_5QNode_Int_7QNode_Int_7_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_7_r;
  QTree_Int_t lizzieLet17_5QNode_Int_7QNode_Int_8_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_8_r;
  QTree_Int_t lizzieLet17_5QNode_Int_7QNode_Int_9_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_9_r;
  QTree_Int_t lizzieLet17_5QNode_Int_7QNode_Int_10_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_10_r;
  QTree_Int_t lizzieLet17_5QNode_Int_7QNode_Int_11_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_11_r;
  QTree_Int_t lizzieLet17_5QNode_Int_7QNode_Int_12_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_12_r;
  QTree_Int_t lizzieLet17_5QNode_Int_7QNode_Int_13_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_13_r;
  QTree_Int_t lizzieLet17_5QNode_Int_7QNode_Int_14_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_14_r;
  Pointer_QTree_Int_t lizzieLet17_5QNode_Int_7QNode_Int_10QNone_Int_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_10QNone_Int_r;
  Pointer_QTree_Int_t _204_d;
  logic _204_r;
  assign _204_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet17_5QNode_Int_7QNode_Int_10QNode_Int_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_10QNode_Int_r;
  Pointer_QTree_Int_t _203_d;
  logic _203_r;
  assign _203_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet17_5QNode_Int_7QNode_Int_10QNone_Int_1_argbuf_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_10QNone_Int_1_argbuf_r;
  Pointer_QTree_Int_t lizzieLet17_5QNode_Int_7QNode_Int_11QNone_Int_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_11QNone_Int_r;
  Pointer_QTree_Int_t _202_d;
  logic _202_r;
  assign _202_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet17_5QNode_Int_7QNode_Int_11QNode_Int_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_11QNode_Int_r;
  Pointer_QTree_Int_t _201_d;
  logic _201_r;
  assign _201_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet17_5QNode_Int_7QNode_Int_11QNone_Int_1_argbuf_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_11QNone_Int_1_argbuf_r;
  Pointer_QTree_Int_t lizzieLet17_5QNode_Int_7QNode_Int_12QNone_Int_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_12QNone_Int_r;
  Pointer_QTree_Int_t _200_d;
  logic _200_r;
  assign _200_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet17_5QNode_Int_7QNode_Int_12QNode_Int_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_12QNode_Int_r;
  Pointer_QTree_Int_t _199_d;
  logic _199_r;
  assign _199_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet17_5QNode_Int_7QNode_Int_12QNone_Int_1_argbuf_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_12QNone_Int_1_argbuf_r;
  Pointer_QTree_Int_t lizzieLet17_5QNode_Int_7QNode_Int_13QNone_Int_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_13QNone_Int_r;
  Pointer_QTree_Int_t _198_d;
  logic _198_r;
  assign _198_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet17_5QNode_Int_7QNode_Int_13QNode_Int_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_13QNode_Int_r;
  Pointer_QTree_Int_t _197_d;
  logic _197_r;
  assign _197_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet17_5QNode_Int_7QNode_Int_13QNone_Int_1_argbuf_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_13QNone_Int_1_argbuf_r;
  Pointer_QTree_Int_t lizzieLet17_5QNode_Int_7QNode_Int_14QNone_Int_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_14QNone_Int_r;
  Pointer_QTree_Int_t _196_d;
  logic _196_r;
  assign _196_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet17_5QNode_Int_7QNode_Int_14QNode_Int_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_14QNode_Int_r;
  Pointer_QTree_Int_t _195_d;
  logic _195_r;
  assign _195_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet17_5QNode_Int_7QNode_Int_14QNode_Int_1_argbuf_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_14QNode_Int_1_argbuf_r;
  Pointer_QTree_Int_t lizzieLet17_5QNode_Int_7QNode_Int_14QNone_Int_1_argbuf_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_14QNone_Int_1_argbuf_r;
  Pointer_QTree_Int_t \t1'aff_destruct_d ;
  logic \t1'aff_destruct_r ;
  Pointer_QTree_Int_t \t2'afg_destruct_d ;
  logic \t2'afg_destruct_r ;
  Pointer_QTree_Int_t \t3'afh_destruct_d ;
  logic \t3'afh_destruct_r ;
  Pointer_QTree_Int_t \t4'afi_destruct_d ;
  logic \t4'afi_destruct_r ;
  QTree_Int_t _194_d;
  logic _194_r;
  assign _194_r = 1'd1;
  QTree_Int_t _193_d;
  logic _193_r;
  assign _193_r = 1'd1;
  QTree_Int_t lizzieLet17_5QNode_Int_7QNode_Int_1QNode_Int_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_1QNode_Int_r;
  QTree_Int_t _192_d;
  logic _192_r;
  assign _192_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet17_5QNode_Int_7QNode_Int_3QNone_Int_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_3QNone_Int_r;
  Pointer_QTree_Int_t _191_d;
  logic _191_r;
  assign _191_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet17_5QNode_Int_7QNode_Int_3QNode_Int_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_3QNode_Int_r;
  Pointer_QTree_Int_t _190_d;
  logic _190_r;
  assign _190_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet17_5QNode_Int_7QNode_Int_3QNone_Int_1_argbuf_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_3QNone_Int_1_argbuf_r;
  Pointer_QTree_Int_t lizzieLet17_5QNode_Int_7QNode_Int_4QNone_Int_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_4QNone_Int_r;
  Pointer_QTree_Int_t _189_d;
  logic _189_r;
  assign _189_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet17_5QNode_Int_7QNode_Int_4QNode_Int_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_4QNode_Int_r;
  Pointer_QTree_Int_t _188_d;
  logic _188_r;
  assign _188_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet17_5QNode_Int_7QNode_Int_4QNone_Int_1_argbuf_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_4QNone_Int_1_argbuf_r;
  Pointer_QTree_Int_t lizzieLet17_5QNode_Int_7QNode_Int_5QNone_Int_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_5QNone_Int_r;
  Pointer_QTree_Int_t _187_d;
  logic _187_r;
  assign _187_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet17_5QNode_Int_7QNode_Int_5QNode_Int_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_5QNode_Int_r;
  Pointer_QTree_Int_t _186_d;
  logic _186_r;
  assign _186_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet17_5QNode_Int_7QNode_Int_5QNode_Int_1_argbuf_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_5QNode_Int_1_argbuf_r;
  Pointer_QTree_Int_t lizzieLet17_5QNode_Int_7QNode_Int_5QNone_Int_1_argbuf_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_5QNone_Int_1_argbuf_r;
  MyDTInt_Int_Int_t lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_r;
  MyDTInt_Int_Int_t _185_d;
  logic _185_r;
  assign _185_r = 1'd1;
  MyDTInt_Int_Int_t lizzieLet17_5QNode_Int_7QNode_Int_6QNode_Int_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_6QNode_Int_r;
  MyDTInt_Int_Int_t _184_d;
  logic _184_r;
  assign _184_r = 1'd1;
  MyDTInt_Int_Int_t lizzieLet17_5QNode_Int_7QNode_Int_6QNode_Int_1_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_6QNode_Int_1_r;
  MyDTInt_Int_Int_t lizzieLet17_5QNode_Int_7QNode_Int_6QNode_Int_2_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_6QNode_Int_2_r;
  MyDTInt_Int_Int_t lizzieLet17_5QNode_Int_7QNode_Int_6QNode_Int_2_argbuf_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_6QNode_Int_2_argbuf_r;
  MyDTInt_Int_Int_t lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_1_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_1_r;
  MyDTInt_Int_Int_t lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_2_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_2_r;
  MyDTInt_Int_Int_t lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_3_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_3_r;
  MyDTInt_Int_Int_t lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_4_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_4_r;
  MyDTInt_Int_Int_t lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_1_argbuf_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_1_argbuf_r;
  MyDTInt_Int_Int_t lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_2_argbuf_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_2_argbuf_r;
  MyDTInt_Int_Int_t lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_3_argbuf_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_3_argbuf_r;
  MyDTInt_Int_Int_t lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_4_argbuf_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_4_argbuf_r;
  Pointer_CTf_f_Int_t lizzieLet17_5QNode_Int_7QNode_Int_7QNone_Int_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_7QNone_Int_r;
  Pointer_CTf_f_Int_t lizzieLet17_5QNode_Int_7QNode_Int_7QVal_Int_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_7QVal_Int_r;
  Pointer_CTf_f_Int_t lizzieLet17_5QNode_Int_7QNode_Int_7QNode_Int_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_7QNode_Int_r;
  Pointer_CTf_f_Int_t lizzieLet17_5QNode_Int_7QNode_Int_7QError_Int_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_7QError_Int_r;
  Pointer_CTf_f_Int_t lizzieLet17_5QNode_Int_7QNode_Int_7QError_Int_1_argbuf_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_7QError_Int_1_argbuf_r;
  CTf_f_Int_t \lizzieLet17_5QNode_Int_7QNode_Int_7QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_10QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_11QNode_Int_1t1'aff_1lizzieLet17_5QNode_Int_7QNode_Int_9QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_6QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_3QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_12QNode_Int_1t2'afg_1lizzieLet17_5QNode_Int_7QNode_Int_4QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_13QNode_Int_1t3'afh_1Lcall_f_f_Int3_d ;
  logic \lizzieLet17_5QNode_Int_7QNode_Int_7QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_10QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_11QNode_Int_1t1'aff_1lizzieLet17_5QNode_Int_7QNode_Int_9QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_6QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_3QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_12QNode_Int_1t2'afg_1lizzieLet17_5QNode_Int_7QNode_Int_4QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_13QNode_Int_1t3'afh_1Lcall_f_f_Int3_r ;
  CTf_f_Int_t lizzieLet52_1_argbuf_d;
  logic lizzieLet52_1_argbuf_r;
  Pointer_CTf_f_Int_t lizzieLet17_5QNode_Int_7QNode_Int_7QNone_Int_1_argbuf_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_7QNone_Int_1_argbuf_r;
  Pointer_CTf_f_Int_t lizzieLet17_5QNode_Int_7QNode_Int_7QVal_Int_1_argbuf_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_7QVal_Int_1_argbuf_r;
  Go_t lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_r;
  Go_t lizzieLet17_5QNode_Int_7QNode_Int_8QVal_Int_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_8QVal_Int_r;
  Go_t lizzieLet17_5QNode_Int_7QNode_Int_8QNode_Int_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_8QNode_Int_r;
  Go_t lizzieLet17_5QNode_Int_7QNode_Int_8QError_Int_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_8QError_Int_r;
  Go_t lizzieLet17_5QNode_Int_7QNode_Int_8QError_Int_1_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_8QError_Int_1_r;
  Go_t lizzieLet17_5QNode_Int_7QNode_Int_8QError_Int_2_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_8QError_Int_2_r;
  QTree_Int_t lizzieLet17_5QNode_Int_7QNode_Int_8QError_Int_1QError_Int_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_8QError_Int_1QError_Int_r;
  QTree_Int_t lizzieLet53_1_argbuf_d;
  logic lizzieLet53_1_argbuf_r;
  Go_t lizzieLet17_5QNode_Int_7QNode_Int_8QError_Int_2_argbuf_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_8QError_Int_2_argbuf_r;
  Go_t lizzieLet17_5QNode_Int_7QNode_Int_8QNode_Int_1_argbuf_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_8QNode_Int_1_argbuf_r;
  Go_t lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_1_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_1_r;
  Go_t lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_2_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_2_r;
  Go_t lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_3_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_3_r;
  Go_t lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_4_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_4_r;
  Go_t lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_5_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_5_r;
  Go_t lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_1_argbuf_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_1_argbuf_r;
  TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_t \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int9_d ;
  logic \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int9_r ;
  Go_t lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_2_argbuf_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_2_argbuf_r;
  TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_t \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int10_d ;
  logic \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int10_r ;
  Go_t lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_3_argbuf_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_3_argbuf_r;
  TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_t \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int11_d ;
  logic \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int11_r ;
  Go_t lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_4_argbuf_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_4_argbuf_r;
  TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_t \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int12_d ;
  logic \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int12_r ;
  Go_t lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_5_argbuf_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_5_argbuf_r;
  Go_t lizzieLet17_5QNode_Int_7QNode_Int_8QVal_Int_1_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_8QVal_Int_1_r;
  Go_t lizzieLet17_5QNode_Int_7QNode_Int_8QVal_Int_2_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_8QVal_Int_2_r;
  QTree_Int_t lizzieLet17_5QNode_Int_7QNode_Int_8QVal_Int_1QError_Int_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_8QVal_Int_1QError_Int_r;
  QTree_Int_t lizzieLet51_1_argbuf_d;
  logic lizzieLet51_1_argbuf_r;
  Go_t lizzieLet17_5QNode_Int_7QNode_Int_8QVal_Int_2_argbuf_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_8QVal_Int_2_argbuf_r;
  MyDTInt_Bool_t lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_r;
  MyDTInt_Bool_t _183_d;
  logic _183_r;
  assign _183_r = 1'd1;
  MyDTInt_Bool_t lizzieLet17_5QNode_Int_7QNode_Int_9QNode_Int_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_9QNode_Int_r;
  MyDTInt_Bool_t _182_d;
  logic _182_r;
  assign _182_r = 1'd1;
  MyDTInt_Bool_t lizzieLet17_5QNode_Int_7QNode_Int_9QNode_Int_1_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_9QNode_Int_1_r;
  MyDTInt_Bool_t lizzieLet17_5QNode_Int_7QNode_Int_9QNode_Int_2_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_9QNode_Int_2_r;
  MyDTInt_Bool_t lizzieLet17_5QNode_Int_7QNode_Int_9QNode_Int_2_argbuf_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_9QNode_Int_2_argbuf_r;
  MyDTInt_Bool_t lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_1_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_1_r;
  MyDTInt_Bool_t lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_2_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_2_r;
  MyDTInt_Bool_t lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_3_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_3_r;
  MyDTInt_Bool_t lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_4_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_4_r;
  MyDTInt_Bool_t lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_1_argbuf_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_1_argbuf_r;
  MyDTInt_Bool_t lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_2_argbuf_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_2_argbuf_r;
  MyDTInt_Bool_t lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_3_argbuf_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_3_argbuf_r;
  MyDTInt_Bool_t lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_4_argbuf_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_4_argbuf_r;
  QTree_Int_t lizzieLet17_5QNode_Int_7QNone_Int_1_d;
  logic lizzieLet17_5QNode_Int_7QNone_Int_1_r;
  QTree_Int_t lizzieLet17_5QNode_Int_7QNone_Int_2_d;
  logic lizzieLet17_5QNode_Int_7QNone_Int_2_r;
  QTree_Int_t lizzieLet17_5QNode_Int_7QNone_Int_3_d;
  logic lizzieLet17_5QNode_Int_7QNone_Int_3_r;
  QTree_Int_t lizzieLet17_5QNode_Int_7QNone_Int_4_d;
  logic lizzieLet17_5QNode_Int_7QNone_Int_4_r;
  QTree_Int_t lizzieLet17_5QNode_Int_7QNone_Int_5_d;
  logic lizzieLet17_5QNode_Int_7QNone_Int_5_r;
  QTree_Int_t lizzieLet17_5QNode_Int_7QNone_Int_6_d;
  logic lizzieLet17_5QNode_Int_7QNone_Int_6_r;
  QTree_Int_t lizzieLet17_5QNode_Int_7QNone_Int_7_d;
  logic lizzieLet17_5QNode_Int_7QNone_Int_7_r;
  QTree_Int_t lizzieLet17_5QNode_Int_7QNone_Int_8_d;
  logic lizzieLet17_5QNode_Int_7QNone_Int_8_r;
  QTree_Int_t lizzieLet17_5QNode_Int_7QNone_Int_9_d;
  logic lizzieLet17_5QNode_Int_7QNone_Int_9_r;
  QTree_Int_t lizzieLet17_5QNode_Int_7QNone_Int_10_d;
  logic lizzieLet17_5QNode_Int_7QNone_Int_10_r;
  QTree_Int_t lizzieLet17_5QNode_Int_7QNone_Int_11_d;
  logic lizzieLet17_5QNode_Int_7QNone_Int_11_r;
  Pointer_QTree_Int_t lizzieLet17_5QNode_Int_7QNone_Int_10QNone_Int_d;
  logic lizzieLet17_5QNode_Int_7QNone_Int_10QNone_Int_r;
  Pointer_QTree_Int_t _181_d;
  logic _181_r;
  assign _181_r = 1'd1;
  Pointer_QTree_Int_t _180_d;
  logic _180_r;
  assign _180_r = 1'd1;
  Pointer_QTree_Int_t _179_d;
  logic _179_r;
  assign _179_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet17_5QNode_Int_7QNone_Int_10QNone_Int_1_argbuf_d;
  logic lizzieLet17_5QNode_Int_7QNone_Int_10QNone_Int_1_argbuf_r;
  Pointer_QTree_Int_t _178_d;
  logic _178_r;
  assign _178_r = 1'd1;
  Pointer_QTree_Int_t _177_d;
  logic _177_r;
  assign _177_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet17_5QNode_Int_7QNone_Int_11QNode_Int_d;
  logic lizzieLet17_5QNode_Int_7QNone_Int_11QNode_Int_r;
  Pointer_QTree_Int_t _176_d;
  logic _176_r;
  assign _176_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet17_5QNode_Int_7QNone_Int_11QNode_Int_1_argbuf_d;
  logic lizzieLet17_5QNode_Int_7QNone_Int_11QNode_Int_1_argbuf_r;
  Pointer_QTree_Int_t t1af5_destruct_d;
  logic t1af5_destruct_r;
  Pointer_QTree_Int_t t2af6_destruct_d;
  logic t2af6_destruct_r;
  Pointer_QTree_Int_t t3af7_destruct_d;
  logic t3af7_destruct_r;
  Pointer_QTree_Int_t t4af8_destruct_d;
  logic t4af8_destruct_r;
  QTree_Int_t _175_d;
  logic _175_r;
  assign _175_r = 1'd1;
  QTree_Int_t _174_d;
  logic _174_r;
  assign _174_r = 1'd1;
  QTree_Int_t lizzieLet17_5QNode_Int_7QNone_Int_1QNode_Int_d;
  logic lizzieLet17_5QNode_Int_7QNone_Int_1QNode_Int_r;
  QTree_Int_t _173_d;
  logic _173_r;
  assign _173_r = 1'd1;
  Pointer_QTree_Int_t _172_d;
  logic _172_r;
  assign _172_r = 1'd1;
  Pointer_QTree_Int_t _171_d;
  logic _171_r;
  assign _171_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet17_5QNode_Int_7QNone_Int_3QNode_Int_d;
  logic lizzieLet17_5QNode_Int_7QNone_Int_3QNode_Int_r;
  Pointer_QTree_Int_t _170_d;
  logic _170_r;
  assign _170_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet17_5QNode_Int_7QNone_Int_3QNode_Int_1_argbuf_d;
  logic lizzieLet17_5QNode_Int_7QNone_Int_3QNode_Int_1_argbuf_r;
  Pointer_QTree_Int_t _169_d;
  logic _169_r;
  assign _169_r = 1'd1;
  Pointer_QTree_Int_t _168_d;
  logic _168_r;
  assign _168_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet17_5QNode_Int_7QNone_Int_4QNode_Int_d;
  logic lizzieLet17_5QNode_Int_7QNone_Int_4QNode_Int_r;
  Pointer_QTree_Int_t _167_d;
  logic _167_r;
  assign _167_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet17_5QNode_Int_7QNone_Int_4QNode_Int_1_argbuf_d;
  logic lizzieLet17_5QNode_Int_7QNone_Int_4QNode_Int_1_argbuf_r;
  Pointer_QTree_Int_t _166_d;
  logic _166_r;
  assign _166_r = 1'd1;
  Pointer_QTree_Int_t _165_d;
  logic _165_r;
  assign _165_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet17_5QNode_Int_7QNone_Int_5QNode_Int_d;
  logic lizzieLet17_5QNode_Int_7QNone_Int_5QNode_Int_r;
  Pointer_QTree_Int_t _164_d;
  logic _164_r;
  assign _164_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet17_5QNode_Int_7QNone_Int_5QNode_Int_1_argbuf_d;
  logic lizzieLet17_5QNode_Int_7QNone_Int_5QNode_Int_1_argbuf_r;
  MyDTInt_Int_Int_t _163_d;
  logic _163_r;
  assign _163_r = 1'd1;
  MyDTInt_Int_Int_t _162_d;
  logic _162_r;
  assign _162_r = 1'd1;
  MyDTInt_Int_Int_t lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_d;
  logic lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_r;
  MyDTInt_Int_Int_t _161_d;
  logic _161_r;
  assign _161_r = 1'd1;
  MyDTInt_Int_Int_t lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_1_d;
  logic lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_1_r;
  MyDTInt_Int_Int_t lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_2_d;
  logic lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_2_r;
  MyDTInt_Int_Int_t lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_3_d;
  logic lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_3_r;
  MyDTInt_Int_Int_t lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_4_d;
  logic lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_4_r;
  MyDTInt_Int_Int_t lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_1_argbuf_d;
  logic lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_1_argbuf_r;
  MyDTInt_Int_Int_t lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_2_argbuf_d;
  logic lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_2_argbuf_r;
  MyDTInt_Int_Int_t lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_3_argbuf_d;
  logic lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_3_argbuf_r;
  MyDTInt_Int_Int_t lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_4_argbuf_d;
  logic lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_4_argbuf_r;
  Pointer_CTf_f_Int_t lizzieLet17_5QNode_Int_7QNone_Int_7QNone_Int_d;
  logic lizzieLet17_5QNode_Int_7QNone_Int_7QNone_Int_r;
  Pointer_CTf_f_Int_t lizzieLet17_5QNode_Int_7QNone_Int_7QVal_Int_d;
  logic lizzieLet17_5QNode_Int_7QNone_Int_7QVal_Int_r;
  Pointer_CTf_f_Int_t lizzieLet17_5QNode_Int_7QNone_Int_7QNode_Int_d;
  logic lizzieLet17_5QNode_Int_7QNone_Int_7QNode_Int_r;
  Pointer_CTf_f_Int_t lizzieLet17_5QNode_Int_7QNone_Int_7QError_Int_d;
  logic lizzieLet17_5QNode_Int_7QNone_Int_7QError_Int_r;
  Pointer_CTf_f_Int_t lizzieLet17_5QNode_Int_7QNone_Int_7QError_Int_1_argbuf_d;
  logic lizzieLet17_5QNode_Int_7QNone_Int_7QError_Int_1_argbuf_r;
  Pointer_CTf_f_Int_t lizzieLet17_5QNode_Int_7QNone_Int_7QNode_Int_1_argbuf_d;
  logic lizzieLet17_5QNode_Int_7QNone_Int_7QNode_Int_1_argbuf_r;
  Pointer_CTf_f_Int_t lizzieLet17_5QNode_Int_7QNone_Int_7QNone_Int_1_argbuf_d;
  logic lizzieLet17_5QNode_Int_7QNone_Int_7QNone_Int_1_argbuf_r;
  Pointer_CTf_f_Int_t lizzieLet17_5QNode_Int_7QNone_Int_7QVal_Int_1_argbuf_d;
  logic lizzieLet17_5QNode_Int_7QNone_Int_7QVal_Int_1_argbuf_r;
  Go_t lizzieLet17_5QNode_Int_7QNone_Int_8QNone_Int_d;
  logic lizzieLet17_5QNode_Int_7QNone_Int_8QNone_Int_r;
  Go_t lizzieLet17_5QNode_Int_7QNone_Int_8QVal_Int_d;
  logic lizzieLet17_5QNode_Int_7QNone_Int_8QVal_Int_r;
  Go_t lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_d;
  logic lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_r;
  Go_t lizzieLet17_5QNode_Int_7QNone_Int_8QError_Int_d;
  logic lizzieLet17_5QNode_Int_7QNone_Int_8QError_Int_r;
  Go_t lizzieLet17_5QNode_Int_7QNone_Int_8QError_Int_1_d;
  logic lizzieLet17_5QNode_Int_7QNone_Int_8QError_Int_1_r;
  Go_t lizzieLet17_5QNode_Int_7QNone_Int_8QError_Int_2_d;
  logic lizzieLet17_5QNode_Int_7QNone_Int_8QError_Int_2_r;
  QTree_Int_t lizzieLet17_5QNode_Int_7QNone_Int_8QError_Int_1QError_Int_d;
  logic lizzieLet17_5QNode_Int_7QNone_Int_8QError_Int_1QError_Int_r;
  QTree_Int_t lizzieLet47_1_argbuf_d;
  logic lizzieLet47_1_argbuf_r;
  Go_t lizzieLet17_5QNode_Int_7QNone_Int_8QError_Int_2_argbuf_d;
  logic lizzieLet17_5QNode_Int_7QNone_Int_8QError_Int_2_argbuf_r;
  Go_t lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_1_d;
  logic lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_1_r;
  Go_t lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_2_d;
  logic lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_2_r;
  Go_t lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_3_d;
  logic lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_3_r;
  Go_t lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_4_d;
  logic lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_4_r;
  Go_t lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_5_d;
  logic lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_5_r;
  Go_t lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_1_argbuf_d;
  logic lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_1_argbuf_r;
  TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_t \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int5_d ;
  logic \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int5_r ;
  Go_t lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_2_argbuf_d;
  logic lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_2_argbuf_r;
  TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_t \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int6_d ;
  logic \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int6_r ;
  Go_t lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_3_argbuf_d;
  logic lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_3_argbuf_r;
  TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_t \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int7_d ;
  logic \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int7_r ;
  Go_t lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_4_argbuf_d;
  logic lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_4_argbuf_r;
  TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_t \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int8_d ;
  logic \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int8_r ;
  Go_t lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_5_argbuf_d;
  logic lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_5_argbuf_r;
  Go_t lizzieLet17_5QNode_Int_7QNone_Int_8QNone_Int_1_argbuf_d;
  logic lizzieLet17_5QNode_Int_7QNone_Int_8QNone_Int_1_argbuf_r;
  Go_t lizzieLet17_5QNode_Int_7QNone_Int_8QVal_Int_1_d;
  logic lizzieLet17_5QNode_Int_7QNone_Int_8QVal_Int_1_r;
  Go_t lizzieLet17_5QNode_Int_7QNone_Int_8QVal_Int_2_d;
  logic lizzieLet17_5QNode_Int_7QNone_Int_8QVal_Int_2_r;
  QTree_Int_t lizzieLet17_5QNode_Int_7QNone_Int_8QVal_Int_1QError_Int_d;
  logic lizzieLet17_5QNode_Int_7QNone_Int_8QVal_Int_1QError_Int_r;
  QTree_Int_t lizzieLet45_1_argbuf_d;
  logic lizzieLet45_1_argbuf_r;
  Go_t lizzieLet17_5QNode_Int_7QNone_Int_8QVal_Int_2_argbuf_d;
  logic lizzieLet17_5QNode_Int_7QNone_Int_8QVal_Int_2_argbuf_r;
  MyDTInt_Bool_t _160_d;
  logic _160_r;
  assign _160_r = 1'd1;
  MyDTInt_Bool_t _159_d;
  logic _159_r;
  assign _159_r = 1'd1;
  MyDTInt_Bool_t lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_d;
  logic lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_r;
  MyDTInt_Bool_t _158_d;
  logic _158_r;
  assign _158_r = 1'd1;
  MyDTInt_Bool_t lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_1_d;
  logic lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_1_r;
  MyDTInt_Bool_t lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_2_d;
  logic lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_2_r;
  MyDTInt_Bool_t lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_3_d;
  logic lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_3_r;
  MyDTInt_Bool_t lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_4_d;
  logic lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_4_r;
  MyDTInt_Bool_t lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_1_argbuf_d;
  logic lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_1_argbuf_r;
  MyDTInt_Bool_t lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_2_argbuf_d;
  logic lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_2_argbuf_r;
  MyDTInt_Bool_t lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_3_argbuf_d;
  logic lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_3_argbuf_r;
  MyDTInt_Bool_t lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_4_argbuf_d;
  logic lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_4_argbuf_r;
  Pointer_QTree_Int_t lizzieLet17_5QNode_Int_8QNone_Int_d;
  logic lizzieLet17_5QNode_Int_8QNone_Int_r;
  Pointer_QTree_Int_t _157_d;
  logic _157_r;
  assign _157_r = 1'd1;
  Pointer_QTree_Int_t _156_d;
  logic _156_r;
  assign _156_r = 1'd1;
  Pointer_QTree_Int_t _155_d;
  logic _155_r;
  assign _155_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet17_5QNode_Int_9QNone_Int_d;
  logic lizzieLet17_5QNode_Int_9QNone_Int_r;
  Pointer_QTree_Int_t _154_d;
  logic _154_r;
  assign _154_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet17_5QNode_Int_9QNode_Int_d;
  logic lizzieLet17_5QNode_Int_9QNode_Int_r;
  Pointer_QTree_Int_t _153_d;
  logic _153_r;
  assign _153_r = 1'd1;
  QTree_Int_t lizzieLet17_5QNone_Int_1_d;
  logic lizzieLet17_5QNone_Int_1_r;
  QTree_Int_t lizzieLet17_5QNone_Int_2_d;
  logic lizzieLet17_5QNone_Int_2_r;
  QTree_Int_t lizzieLet17_5QNone_Int_3_d;
  logic lizzieLet17_5QNone_Int_3_r;
  QTree_Int_t lizzieLet17_5QNone_Int_4_d;
  logic lizzieLet17_5QNone_Int_4_r;
  QTree_Int_t lizzieLet17_5QNone_Int_5_d;
  logic lizzieLet17_5QNone_Int_5_r;
  QTree_Int_t lizzieLet17_5QNone_Int_6_d;
  logic lizzieLet17_5QNone_Int_6_r;
  QTree_Int_t lizzieLet17_5QNone_Int_7_d;
  logic lizzieLet17_5QNone_Int_7_r;
  QTree_Int_t lizzieLet17_5QNone_Int_8_d;
  logic lizzieLet17_5QNone_Int_8_r;
  QTree_Int_t lizzieLet17_5QNone_Int_9_d;
  logic lizzieLet17_5QNone_Int_9_r;
  Pointer_QTree_Int_t q1aeB_destruct_d;
  logic q1aeB_destruct_r;
  Pointer_QTree_Int_t q2aeC_destruct_d;
  logic q2aeC_destruct_r;
  Pointer_QTree_Int_t q3aeD_destruct_d;
  logic q3aeD_destruct_r;
  Pointer_QTree_Int_t q4aeE_destruct_d;
  logic q4aeE_destruct_r;
  Int_t v1aev_destruct_d;
  logic v1aev_destruct_r;
  QTree_Int_t _152_d;
  logic _152_r;
  assign _152_r = 1'd1;
  QTree_Int_t lizzieLet17_5QNone_Int_1QVal_Int_d;
  logic lizzieLet17_5QNone_Int_1QVal_Int_r;
  QTree_Int_t lizzieLet17_5QNone_Int_1QNode_Int_d;
  logic lizzieLet17_5QNone_Int_1QNode_Int_r;
  QTree_Int_t _151_d;
  logic _151_r;
  assign _151_r = 1'd1;
  MyDTInt_Int_Int_t _150_d;
  logic _150_r;
  assign _150_r = 1'd1;
  MyDTInt_Int_Int_t lizzieLet17_5QNone_Int_3QVal_Int_d;
  logic lizzieLet17_5QNone_Int_3QVal_Int_r;
  MyDTInt_Int_Int_t lizzieLet17_5QNone_Int_3QNode_Int_d;
  logic lizzieLet17_5QNone_Int_3QNode_Int_r;
  MyDTInt_Int_Int_t _149_d;
  logic _149_r;
  assign _149_r = 1'd1;
  Pointer_CTf_f_Int_t lizzieLet17_5QNone_Int_4QNone_Int_d;
  logic lizzieLet17_5QNone_Int_4QNone_Int_r;
  Pointer_CTf_f_Int_t lizzieLet17_5QNone_Int_4QVal_Int_d;
  logic lizzieLet17_5QNone_Int_4QVal_Int_r;
  Pointer_CTf_f_Int_t lizzieLet17_5QNone_Int_4QNode_Int_d;
  logic lizzieLet17_5QNone_Int_4QNode_Int_r;
  Pointer_CTf_f_Int_t lizzieLet17_5QNone_Int_4QError_Int_d;
  logic lizzieLet17_5QNone_Int_4QError_Int_r;
  Pointer_CTf_f_Int_t lizzieLet17_5QNone_Int_4QError_Int_1_argbuf_d;
  logic lizzieLet17_5QNone_Int_4QError_Int_1_argbuf_r;
  Pointer_CTf_f_Int_t lizzieLet17_5QNone_Int_4QNone_Int_1_argbuf_d;
  logic lizzieLet17_5QNone_Int_4QNone_Int_1_argbuf_r;
  Go_t lizzieLet17_5QNone_Int_5QNone_Int_d;
  logic lizzieLet17_5QNone_Int_5QNone_Int_r;
  Go_t lizzieLet17_5QNone_Int_5QVal_Int_d;
  logic lizzieLet17_5QNone_Int_5QVal_Int_r;
  Go_t lizzieLet17_5QNone_Int_5QNode_Int_d;
  logic lizzieLet17_5QNone_Int_5QNode_Int_r;
  Go_t lizzieLet17_5QNone_Int_5QError_Int_d;
  logic lizzieLet17_5QNone_Int_5QError_Int_r;
  Go_t lizzieLet17_5QNone_Int_5QError_Int_1_d;
  logic lizzieLet17_5QNone_Int_5QError_Int_1_r;
  Go_t lizzieLet17_5QNone_Int_5QError_Int_2_d;
  logic lizzieLet17_5QNone_Int_5QError_Int_2_r;
  QTree_Int_t lizzieLet17_5QNone_Int_5QError_Int_1QError_Int_d;
  logic lizzieLet17_5QNone_Int_5QError_Int_1QError_Int_r;
  QTree_Int_t lizzieLet28_1_argbuf_d;
  logic lizzieLet28_1_argbuf_r;
  Go_t lizzieLet17_5QNone_Int_5QError_Int_2_argbuf_d;
  logic lizzieLet17_5QNone_Int_5QError_Int_2_argbuf_r;
  Go_t lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_d;
  logic lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_r;
  C35_t go_15_goMux_choice_d;
  logic go_15_goMux_choice_r;
  Go_t go_15_goMux_data_d;
  logic go_15_goMux_data_r;
  MyDTInt_Bool_t _148_d;
  logic _148_r;
  assign _148_r = 1'd1;
  MyDTInt_Bool_t lizzieLet17_5QNone_Int_6QVal_Int_d;
  logic lizzieLet17_5QNone_Int_6QVal_Int_r;
  MyDTInt_Bool_t lizzieLet17_5QNone_Int_6QNode_Int_d;
  logic lizzieLet17_5QNone_Int_6QNode_Int_r;
  MyDTInt_Bool_t _147_d;
  logic _147_r;
  assign _147_r = 1'd1;
  QTree_Int_t _146_d;
  logic _146_r;
  assign _146_r = 1'd1;
  QTree_Int_t lizzieLet17_5QNone_Int_7QVal_Int_d;
  logic lizzieLet17_5QNone_Int_7QVal_Int_r;
  QTree_Int_t lizzieLet17_5QNone_Int_7QNode_Int_d;
  logic lizzieLet17_5QNone_Int_7QNode_Int_r;
  QTree_Int_t _145_d;
  logic _145_r;
  assign _145_r = 1'd1;
  QTree_Int_t lizzieLet17_5QNone_Int_7QNode_Int_1_d;
  logic lizzieLet17_5QNone_Int_7QNode_Int_1_r;
  QTree_Int_t lizzieLet17_5QNone_Int_7QNode_Int_2_d;
  logic lizzieLet17_5QNone_Int_7QNode_Int_2_r;
  QTree_Int_t lizzieLet17_5QNone_Int_7QNode_Int_3_d;
  logic lizzieLet17_5QNone_Int_7QNode_Int_3_r;
  QTree_Int_t lizzieLet17_5QNone_Int_7QNode_Int_4_d;
  logic lizzieLet17_5QNone_Int_7QNode_Int_4_r;
  QTree_Int_t lizzieLet17_5QNone_Int_7QNode_Int_5_d;
  logic lizzieLet17_5QNone_Int_7QNode_Int_5_r;
  QTree_Int_t lizzieLet17_5QNone_Int_7QNode_Int_6_d;
  logic lizzieLet17_5QNone_Int_7QNode_Int_6_r;
  QTree_Int_t lizzieLet17_5QNone_Int_7QNode_Int_7_d;
  logic lizzieLet17_5QNone_Int_7QNode_Int_7_r;
  QTree_Int_t lizzieLet17_5QNone_Int_7QNode_Int_8_d;
  logic lizzieLet17_5QNone_Int_7QNode_Int_8_r;
  QTree_Int_t lizzieLet17_5QNone_Int_7QNode_Int_9_d;
  logic lizzieLet17_5QNone_Int_7QNode_Int_9_r;
  QTree_Int_t lizzieLet17_5QNone_Int_7QNode_Int_10_d;
  logic lizzieLet17_5QNone_Int_7QNode_Int_10_r;
  QTree_Int_t lizzieLet17_5QNone_Int_7QNode_Int_11_d;
  logic lizzieLet17_5QNone_Int_7QNode_Int_11_r;
  Pointer_QTree_Int_t _144_d;
  logic _144_r;
  assign _144_r = 1'd1;
  Pointer_QTree_Int_t _143_d;
  logic _143_r;
  assign _143_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet17_5QNone_Int_7QNode_Int_10QNode_Int_d;
  logic lizzieLet17_5QNone_Int_7QNode_Int_10QNode_Int_r;
  Pointer_QTree_Int_t _142_d;
  logic _142_r;
  assign _142_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet17_5QNone_Int_7QNode_Int_10QNode_Int_1_argbuf_d;
  logic lizzieLet17_5QNone_Int_7QNode_Int_10QNode_Int_1_argbuf_r;
  Pointer_QTree_Int_t _141_d;
  logic _141_r;
  assign _141_r = 1'd1;
  Pointer_QTree_Int_t _140_d;
  logic _140_r;
  assign _140_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet17_5QNone_Int_7QNode_Int_11QNode_Int_d;
  logic lizzieLet17_5QNone_Int_7QNode_Int_11QNode_Int_r;
  Pointer_QTree_Int_t _139_d;
  logic _139_r;
  assign _139_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet17_5QNone_Int_7QNode_Int_11QNode_Int_1_argbuf_d;
  logic lizzieLet17_5QNone_Int_7QNode_Int_11QNode_Int_1_argbuf_r;
  Pointer_QTree_Int_t t1aeG_destruct_d;
  logic t1aeG_destruct_r;
  Pointer_QTree_Int_t t2aeH_destruct_d;
  logic t2aeH_destruct_r;
  Pointer_QTree_Int_t t3aeI_destruct_d;
  logic t3aeI_destruct_r;
  Pointer_QTree_Int_t t4aeJ_destruct_d;
  logic t4aeJ_destruct_r;
  QTree_Int_t _138_d;
  logic _138_r;
  assign _138_r = 1'd1;
  QTree_Int_t _137_d;
  logic _137_r;
  assign _137_r = 1'd1;
  QTree_Int_t lizzieLet17_5QNone_Int_7QNode_Int_1QNode_Int_d;
  logic lizzieLet17_5QNone_Int_7QNode_Int_1QNode_Int_r;
  QTree_Int_t _136_d;
  logic _136_r;
  assign _136_r = 1'd1;
  MyDTInt_Int_Int_t _135_d;
  logic _135_r;
  assign _135_r = 1'd1;
  MyDTInt_Int_Int_t _134_d;
  logic _134_r;
  assign _134_r = 1'd1;
  MyDTInt_Int_Int_t lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_d;
  logic lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_r;
  MyDTInt_Int_Int_t _133_d;
  logic _133_r;
  assign _133_r = 1'd1;
  MyDTInt_Int_Int_t lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_1_d;
  logic lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_1_r;
  MyDTInt_Int_Int_t lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_2_d;
  logic lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_2_r;
  MyDTInt_Int_Int_t lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_3_d;
  logic lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_3_r;
  MyDTInt_Int_Int_t lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_4_d;
  logic lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_4_r;
  MyDTInt_Int_Int_t lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_1_argbuf_d;
  logic lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_1_argbuf_r;
  MyDTInt_Int_Int_t lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_2_argbuf_d;
  logic lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_2_argbuf_r;
  MyDTInt_Int_Int_t lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_3_argbuf_d;
  logic lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_3_argbuf_r;
  MyDTInt_Int_Int_t lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_4_argbuf_d;
  logic lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_4_argbuf_r;
  Pointer_CTf_f_Int_t lizzieLet17_5QNone_Int_7QNode_Int_4QNone_Int_d;
  logic lizzieLet17_5QNone_Int_7QNode_Int_4QNone_Int_r;
  Pointer_CTf_f_Int_t lizzieLet17_5QNone_Int_7QNode_Int_4QVal_Int_d;
  logic lizzieLet17_5QNone_Int_7QNode_Int_4QVal_Int_r;
  Pointer_CTf_f_Int_t lizzieLet17_5QNone_Int_7QNode_Int_4QNode_Int_d;
  logic lizzieLet17_5QNone_Int_7QNode_Int_4QNode_Int_r;
  Pointer_CTf_f_Int_t lizzieLet17_5QNone_Int_7QNode_Int_4QError_Int_d;
  logic lizzieLet17_5QNone_Int_7QNode_Int_4QError_Int_r;
  Pointer_CTf_f_Int_t lizzieLet17_5QNone_Int_7QNode_Int_4QError_Int_1_argbuf_d;
  logic lizzieLet17_5QNone_Int_7QNode_Int_4QError_Int_1_argbuf_r;
  Pointer_CTf_f_Int_t lizzieLet17_5QNone_Int_7QNode_Int_4QNode_Int_1_argbuf_d;
  logic lizzieLet17_5QNone_Int_7QNode_Int_4QNode_Int_1_argbuf_r;
  Pointer_CTf_f_Int_t lizzieLet17_5QNone_Int_7QNode_Int_4QNone_Int_1_argbuf_d;
  logic lizzieLet17_5QNone_Int_7QNode_Int_4QNone_Int_1_argbuf_r;
  Pointer_CTf_f_Int_t lizzieLet17_5QNone_Int_7QNode_Int_4QVal_Int_1_argbuf_d;
  logic lizzieLet17_5QNone_Int_7QNode_Int_4QVal_Int_1_argbuf_r;
  Go_t lizzieLet17_5QNone_Int_7QNode_Int_5QNone_Int_d;
  logic lizzieLet17_5QNone_Int_7QNode_Int_5QNone_Int_r;
  Go_t lizzieLet17_5QNone_Int_7QNode_Int_5QVal_Int_d;
  logic lizzieLet17_5QNone_Int_7QNode_Int_5QVal_Int_r;
  Go_t lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_d;
  logic lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_r;
  Go_t lizzieLet17_5QNone_Int_7QNode_Int_5QError_Int_d;
  logic lizzieLet17_5QNone_Int_7QNode_Int_5QError_Int_r;
  Go_t lizzieLet17_5QNone_Int_7QNode_Int_5QError_Int_1_d;
  logic lizzieLet17_5QNone_Int_7QNode_Int_5QError_Int_1_r;
  Go_t lizzieLet17_5QNone_Int_7QNode_Int_5QError_Int_2_d;
  logic lizzieLet17_5QNone_Int_7QNode_Int_5QError_Int_2_r;
  QTree_Int_t lizzieLet17_5QNone_Int_7QNode_Int_5QError_Int_1QError_Int_d;
  logic lizzieLet17_5QNone_Int_7QNode_Int_5QError_Int_1QError_Int_r;
  QTree_Int_t lizzieLet27_1_argbuf_d;
  logic lizzieLet27_1_argbuf_r;
  Go_t lizzieLet17_5QNone_Int_7QNode_Int_5QError_Int_2_argbuf_d;
  logic lizzieLet17_5QNone_Int_7QNode_Int_5QError_Int_2_argbuf_r;
  Go_t lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_1_d;
  logic lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_1_r;
  Go_t lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_2_d;
  logic lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_2_r;
  Go_t lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_3_d;
  logic lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_3_r;
  Go_t lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_4_d;
  logic lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_4_r;
  Go_t lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_5_d;
  logic lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_5_r;
  Go_t lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_1_argbuf_d;
  logic lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_1_argbuf_r;
  TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_t \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_d ;
  logic \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_r ;
  Go_t lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_2_argbuf_d;
  logic lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_2_argbuf_r;
  TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_t \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int2_d ;
  logic \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int2_r ;
  Go_t lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_3_argbuf_d;
  logic lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_3_argbuf_r;
  TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_t \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int3_d ;
  logic \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int3_r ;
  Go_t lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_4_argbuf_d;
  logic lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_4_argbuf_r;
  TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_t \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int4_d ;
  logic \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int4_r ;
  Go_t lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_5_argbuf_d;
  logic lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_5_argbuf_r;
  Go_t lizzieLet17_5QNone_Int_7QNode_Int_5QNone_Int_1_argbuf_d;
  logic lizzieLet17_5QNone_Int_7QNode_Int_5QNone_Int_1_argbuf_r;
  Go_t lizzieLet17_5QNone_Int_7QNode_Int_5QVal_Int_1_d;
  logic lizzieLet17_5QNone_Int_7QNode_Int_5QVal_Int_1_r;
  Go_t lizzieLet17_5QNone_Int_7QNode_Int_5QVal_Int_2_d;
  logic lizzieLet17_5QNone_Int_7QNode_Int_5QVal_Int_2_r;
  QTree_Int_t lizzieLet17_5QNone_Int_7QNode_Int_5QVal_Int_1QError_Int_d;
  logic lizzieLet17_5QNone_Int_7QNode_Int_5QVal_Int_1QError_Int_r;
  QTree_Int_t lizzieLet25_1_argbuf_d;
  logic lizzieLet25_1_argbuf_r;
  Go_t lizzieLet17_5QNone_Int_7QNode_Int_5QVal_Int_2_argbuf_d;
  logic lizzieLet17_5QNone_Int_7QNode_Int_5QVal_Int_2_argbuf_r;
  MyDTInt_Bool_t _132_d;
  logic _132_r;
  assign _132_r = 1'd1;
  MyDTInt_Bool_t _131_d;
  logic _131_r;
  assign _131_r = 1'd1;
  MyDTInt_Bool_t lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_d;
  logic lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_r;
  MyDTInt_Bool_t _130_d;
  logic _130_r;
  assign _130_r = 1'd1;
  MyDTInt_Bool_t lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_1_d;
  logic lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_1_r;
  MyDTInt_Bool_t lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_2_d;
  logic lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_2_r;
  MyDTInt_Bool_t lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_3_d;
  logic lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_3_r;
  MyDTInt_Bool_t lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_4_d;
  logic lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_4_r;
  MyDTInt_Bool_t lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_1_argbuf_d;
  logic lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_1_argbuf_r;
  MyDTInt_Bool_t lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_2_argbuf_d;
  logic lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_2_argbuf_r;
  MyDTInt_Bool_t lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_3_argbuf_d;
  logic lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_3_argbuf_r;
  MyDTInt_Bool_t lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_4_argbuf_d;
  logic lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_4_argbuf_r;
  Pointer_QTree_Int_t lizzieLet17_5QNone_Int_7QNode_Int_7QNone_Int_d;
  logic lizzieLet17_5QNone_Int_7QNode_Int_7QNone_Int_r;
  Pointer_QTree_Int_t _129_d;
  logic _129_r;
  assign _129_r = 1'd1;
  Pointer_QTree_Int_t _128_d;
  logic _128_r;
  assign _128_r = 1'd1;
  Pointer_QTree_Int_t _127_d;
  logic _127_r;
  assign _127_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet17_5QNone_Int_7QNode_Int_7QNone_Int_1_argbuf_d;
  logic lizzieLet17_5QNone_Int_7QNode_Int_7QNone_Int_1_argbuf_r;
  Pointer_QTree_Int_t _126_d;
  logic _126_r;
  assign _126_r = 1'd1;
  Pointer_QTree_Int_t _125_d;
  logic _125_r;
  assign _125_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet17_5QNone_Int_7QNode_Int_8QNode_Int_d;
  logic lizzieLet17_5QNone_Int_7QNode_Int_8QNode_Int_r;
  Pointer_QTree_Int_t _124_d;
  logic _124_r;
  assign _124_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet17_5QNone_Int_7QNode_Int_8QNode_Int_1_argbuf_d;
  logic lizzieLet17_5QNone_Int_7QNode_Int_8QNode_Int_1_argbuf_r;
  Pointer_QTree_Int_t _123_d;
  logic _123_r;
  assign _123_r = 1'd1;
  Pointer_QTree_Int_t _122_d;
  logic _122_r;
  assign _122_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet17_5QNone_Int_7QNode_Int_9QNode_Int_d;
  logic lizzieLet17_5QNone_Int_7QNode_Int_9QNode_Int_r;
  Pointer_QTree_Int_t _121_d;
  logic _121_r;
  assign _121_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet17_5QNone_Int_7QNode_Int_9QNode_Int_1_argbuf_d;
  logic lizzieLet17_5QNone_Int_7QNode_Int_9QNode_Int_1_argbuf_r;
  QTree_Int_t lizzieLet17_5QNone_Int_7QVal_Int_1_d;
  logic lizzieLet17_5QNone_Int_7QVal_Int_1_r;
  QTree_Int_t lizzieLet17_5QNone_Int_7QVal_Int_2_d;
  logic lizzieLet17_5QNone_Int_7QVal_Int_2_r;
  QTree_Int_t lizzieLet17_5QNone_Int_7QVal_Int_3_d;
  logic lizzieLet17_5QNone_Int_7QVal_Int_3_r;
  QTree_Int_t lizzieLet17_5QNone_Int_7QVal_Int_4_d;
  logic lizzieLet17_5QNone_Int_7QVal_Int_4_r;
  QTree_Int_t lizzieLet17_5QNone_Int_7QVal_Int_5_d;
  logic lizzieLet17_5QNone_Int_7QVal_Int_5_r;
  QTree_Int_t lizzieLet17_5QNone_Int_7QVal_Int_6_d;
  logic lizzieLet17_5QNone_Int_7QVal_Int_6_r;
  QTree_Int_t lizzieLet17_5QNone_Int_7QVal_Int_7_d;
  logic lizzieLet17_5QNone_Int_7QVal_Int_7_r;
  QTree_Int_t lizzieLet17_5QNone_Int_7QVal_Int_8_d;
  logic lizzieLet17_5QNone_Int_7QVal_Int_8_r;
  Int_t vaew_destruct_d;
  logic vaew_destruct_r;
  QTree_Int_t _120_d;
  logic _120_r;
  assign _120_r = 1'd1;
  QTree_Int_t lizzieLet17_5QNone_Int_7QVal_Int_1QVal_Int_d;
  logic lizzieLet17_5QNone_Int_7QVal_Int_1QVal_Int_r;
  QTree_Int_t _119_d;
  logic _119_r;
  assign _119_r = 1'd1;
  QTree_Int_t _118_d;
  logic _118_r;
  assign _118_r = 1'd1;
  MyDTInt_Int_Int_t _117_d;
  logic _117_r;
  assign _117_r = 1'd1;
  MyDTInt_Int_Int_t lizzieLet17_5QNone_Int_7QVal_Int_3QVal_Int_d;
  logic lizzieLet17_5QNone_Int_7QVal_Int_3QVal_Int_r;
  MyDTInt_Int_Int_t _116_d;
  logic _116_r;
  assign _116_r = 1'd1;
  MyDTInt_Int_Int_t _115_d;
  logic _115_r;
  assign _115_r = 1'd1;
  MyDTInt_Int_Int_t lizzieLet17_5QNone_Int_7QVal_Int_3QVal_Int_1_d;
  logic lizzieLet17_5QNone_Int_7QVal_Int_3QVal_Int_1_r;
  MyDTInt_Int_Int_t lizzieLet17_5QNone_Int_7QVal_Int_3QVal_Int_2_d;
  logic lizzieLet17_5QNone_Int_7QVal_Int_3QVal_Int_2_r;
  MyDTInt_Int_Int_t lizzieLet17_5QNone_Int_7QVal_Int_3QVal_Int_1_argbuf_d;
  logic lizzieLet17_5QNone_Int_7QVal_Int_3QVal_Int_1_argbuf_r;
  TupMyDTInt_Int_Int___Int___Int_t applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_d;
  logic applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_r;
  Pointer_CTf_f_Int_t lizzieLet17_5QNone_Int_7QVal_Int_4QNone_Int_d;
  logic lizzieLet17_5QNone_Int_7QVal_Int_4QNone_Int_r;
  Pointer_CTf_f_Int_t lizzieLet17_5QNone_Int_7QVal_Int_4QVal_Int_d;
  logic lizzieLet17_5QNone_Int_7QVal_Int_4QVal_Int_r;
  Pointer_CTf_f_Int_t lizzieLet17_5QNone_Int_7QVal_Int_4QNode_Int_d;
  logic lizzieLet17_5QNone_Int_7QVal_Int_4QNode_Int_r;
  Pointer_CTf_f_Int_t lizzieLet17_5QNone_Int_7QVal_Int_4QError_Int_d;
  logic lizzieLet17_5QNone_Int_7QVal_Int_4QError_Int_r;
  Pointer_CTf_f_Int_t lizzieLet17_5QNone_Int_7QVal_Int_4QError_Int_1_argbuf_d;
  logic lizzieLet17_5QNone_Int_7QVal_Int_4QError_Int_1_argbuf_r;
  Pointer_CTf_f_Int_t lizzieLet17_5QNone_Int_7QVal_Int_4QNode_Int_1_argbuf_d;
  logic lizzieLet17_5QNone_Int_7QVal_Int_4QNode_Int_1_argbuf_r;
  Pointer_CTf_f_Int_t lizzieLet17_5QNone_Int_7QVal_Int_4QNone_Int_1_argbuf_d;
  logic lizzieLet17_5QNone_Int_7QVal_Int_4QNone_Int_1_argbuf_r;
  Go_t lizzieLet17_5QNone_Int_7QVal_Int_5QNone_Int_d;
  logic lizzieLet17_5QNone_Int_7QVal_Int_5QNone_Int_r;
  Go_t lizzieLet17_5QNone_Int_7QVal_Int_5QVal_Int_d;
  logic lizzieLet17_5QNone_Int_7QVal_Int_5QVal_Int_r;
  Go_t lizzieLet17_5QNone_Int_7QVal_Int_5QNode_Int_d;
  logic lizzieLet17_5QNone_Int_7QVal_Int_5QNode_Int_r;
  Go_t lizzieLet17_5QNone_Int_7QVal_Int_5QError_Int_d;
  logic lizzieLet17_5QNone_Int_7QVal_Int_5QError_Int_r;
  Go_t lizzieLet17_5QNone_Int_7QVal_Int_5QError_Int_1_d;
  logic lizzieLet17_5QNone_Int_7QVal_Int_5QError_Int_1_r;
  Go_t lizzieLet17_5QNone_Int_7QVal_Int_5QError_Int_2_d;
  logic lizzieLet17_5QNone_Int_7QVal_Int_5QError_Int_2_r;
  QTree_Int_t lizzieLet17_5QNone_Int_7QVal_Int_5QError_Int_1QError_Int_d;
  logic lizzieLet17_5QNone_Int_7QVal_Int_5QError_Int_1QError_Int_r;
  QTree_Int_t lizzieLet23_1_argbuf_d;
  logic lizzieLet23_1_argbuf_r;
  Go_t lizzieLet17_5QNone_Int_7QVal_Int_5QError_Int_2_argbuf_d;
  logic lizzieLet17_5QNone_Int_7QVal_Int_5QError_Int_2_argbuf_r;
  Go_t lizzieLet17_5QNone_Int_7QVal_Int_5QNode_Int_1_d;
  logic lizzieLet17_5QNone_Int_7QVal_Int_5QNode_Int_1_r;
  Go_t lizzieLet17_5QNone_Int_7QVal_Int_5QNode_Int_2_d;
  logic lizzieLet17_5QNone_Int_7QVal_Int_5QNode_Int_2_r;
  QTree_Int_t lizzieLet17_5QNone_Int_7QVal_Int_5QNode_Int_1QError_Int_d;
  logic lizzieLet17_5QNone_Int_7QVal_Int_5QNode_Int_1QError_Int_r;
  QTree_Int_t lizzieLet22_1_argbuf_d;
  logic lizzieLet22_1_argbuf_r;
  Go_t lizzieLet17_5QNone_Int_7QVal_Int_5QNode_Int_2_argbuf_d;
  logic lizzieLet17_5QNone_Int_7QVal_Int_5QNode_Int_2_argbuf_r;
  Go_t lizzieLet17_5QNone_Int_7QVal_Int_5QNone_Int_1_argbuf_d;
  logic lizzieLet17_5QNone_Int_7QVal_Int_5QNone_Int_1_argbuf_r;
  Go_t lizzieLet17_5QNone_Int_7QVal_Int_5QVal_Int_1_d;
  logic lizzieLet17_5QNone_Int_7QVal_Int_5QVal_Int_1_r;
  Go_t lizzieLet17_5QNone_Int_7QVal_Int_5QVal_Int_2_d;
  logic lizzieLet17_5QNone_Int_7QVal_Int_5QVal_Int_2_r;
  Go_t lizzieLet17_5QNone_Int_7QVal_Int_5QVal_Int_1_argbuf_d;
  logic lizzieLet17_5QNone_Int_7QVal_Int_5QVal_Int_1_argbuf_r;
  TupGo___MyDTInt_Bool___Int_t applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_d;
  logic applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_r;
  MyDTInt_Bool_t _114_d;
  logic _114_r;
  assign _114_r = 1'd1;
  MyDTInt_Bool_t lizzieLet17_5QNone_Int_7QVal_Int_6QVal_Int_d;
  logic lizzieLet17_5QNone_Int_7QVal_Int_6QVal_Int_r;
  MyDTInt_Bool_t _113_d;
  logic _113_r;
  assign _113_r = 1'd1;
  MyDTInt_Bool_t _112_d;
  logic _112_r;
  assign _112_r = 1'd1;
  MyDTInt_Bool_t lizzieLet17_5QNone_Int_7QVal_Int_6QVal_Int_1_argbuf_d;
  logic lizzieLet17_5QNone_Int_7QVal_Int_6QVal_Int_1_argbuf_r;
  Pointer_QTree_Int_t lizzieLet17_5QNone_Int_7QVal_Int_7QNone_Int_d;
  logic lizzieLet17_5QNone_Int_7QVal_Int_7QNone_Int_r;
  Pointer_QTree_Int_t _111_d;
  logic _111_r;
  assign _111_r = 1'd1;
  Pointer_QTree_Int_t _110_d;
  logic _110_r;
  assign _110_r = 1'd1;
  Pointer_QTree_Int_t _109_d;
  logic _109_r;
  assign _109_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet17_5QNone_Int_7QVal_Int_7QNone_Int_1_argbuf_d;
  logic lizzieLet17_5QNone_Int_7QVal_Int_7QNone_Int_1_argbuf_r;
  Int_t _108_d;
  logic _108_r;
  assign _108_r = 1'd1;
  Int_t lizzieLet17_5QNone_Int_7QVal_Int_8QVal_Int_d;
  logic lizzieLet17_5QNone_Int_7QVal_Int_8QVal_Int_r;
  Int_t _107_d;
  logic _107_r;
  assign _107_r = 1'd1;
  Int_t _106_d;
  logic _106_r;
  assign _106_r = 1'd1;
  Int_t lizzieLet17_5QNone_Int_7QVal_Int_8QVal_Int_1_d;
  logic lizzieLet17_5QNone_Int_7QVal_Int_8QVal_Int_1_r;
  Int_t lizzieLet17_5QNone_Int_7QVal_Int_8QVal_Int_2_d;
  logic lizzieLet17_5QNone_Int_7QVal_Int_8QVal_Int_2_r;
  Int_t lizzieLet17_5QNone_Int_7QVal_Int_8QVal_Int_1_argbuf_d;
  logic lizzieLet17_5QNone_Int_7QVal_Int_8QVal_Int_1_argbuf_r;
  Pointer_QTree_Int_t _105_d;
  logic _105_r;
  assign _105_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet17_5QNone_Int_8QVal_Int_d;
  logic lizzieLet17_5QNone_Int_8QVal_Int_r;
  Pointer_QTree_Int_t lizzieLet17_5QNone_Int_8QNode_Int_d;
  logic lizzieLet17_5QNone_Int_8QNode_Int_r;
  Pointer_QTree_Int_t _104_d;
  logic _104_r;
  assign _104_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet17_5QNone_Int_9QNone_Int_d;
  logic lizzieLet17_5QNone_Int_9QNone_Int_r;
  Pointer_QTree_Int_t _103_d;
  logic _103_r;
  assign _103_r = 1'd1;
  Pointer_QTree_Int_t _102_d;
  logic _102_r;
  assign _102_r = 1'd1;
  Pointer_QTree_Int_t _101_d;
  logic _101_r;
  assign _101_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet17_5QNone_Int_9QNone_Int_1_argbuf_d;
  logic lizzieLet17_5QNone_Int_9QNone_Int_1_argbuf_r;
  QTree_Int_t lizzieLet17_5QVal_Int_1_d;
  logic lizzieLet17_5QVal_Int_1_r;
  QTree_Int_t lizzieLet17_5QVal_Int_2_d;
  logic lizzieLet17_5QVal_Int_2_r;
  QTree_Int_t lizzieLet17_5QVal_Int_3_d;
  logic lizzieLet17_5QVal_Int_3_r;
  QTree_Int_t lizzieLet17_5QVal_Int_4_d;
  logic lizzieLet17_5QVal_Int_4_r;
  QTree_Int_t lizzieLet17_5QVal_Int_5_d;
  logic lizzieLet17_5QVal_Int_5_r;
  QTree_Int_t lizzieLet17_5QVal_Int_6_d;
  logic lizzieLet17_5QVal_Int_6_r;
  QTree_Int_t lizzieLet17_5QVal_Int_7_d;
  logic lizzieLet17_5QVal_Int_7_r;
  QTree_Int_t lizzieLet17_5QVal_Int_8_d;
  logic lizzieLet17_5QVal_Int_8_r;
  QTree_Int_t lizzieLet17_5QVal_Int_9_d;
  logic lizzieLet17_5QVal_Int_9_r;
  QTree_Int_t lizzieLet17_5QVal_Int_10_d;
  logic lizzieLet17_5QVal_Int_10_r;
  Int_t lizzieLet17_5QVal_Int_10QNone_Int_d;
  logic lizzieLet17_5QVal_Int_10QNone_Int_r;
  Int_t lizzieLet17_5QVal_Int_10QVal_Int_d;
  logic lizzieLet17_5QVal_Int_10QVal_Int_r;
  Int_t _100_d;
  logic _100_r;
  assign _100_r = 1'd1;
  Int_t _99_d;
  logic _99_r;
  assign _99_r = 1'd1;
  Int_t lizzieLet17_5QVal_Int_10QVal_Int_1_d;
  logic lizzieLet17_5QVal_Int_10QVal_Int_1_r;
  Int_t lizzieLet17_5QVal_Int_10QVal_Int_2_d;
  logic lizzieLet17_5QVal_Int_10QVal_Int_2_r;
  Int_t lizzieLet17_5QVal_Int_10QVal_Int_1_argbuf_d;
  logic lizzieLet17_5QVal_Int_10QVal_Int_1_argbuf_r;
  Int_t vaeQ_destruct_d;
  logic vaeQ_destruct_r;
  QTree_Int_t _98_d;
  logic _98_r;
  assign _98_r = 1'd1;
  QTree_Int_t lizzieLet17_5QVal_Int_1QVal_Int_d;
  logic lizzieLet17_5QVal_Int_1QVal_Int_r;
  QTree_Int_t _97_d;
  logic _97_r;
  assign _97_r = 1'd1;
  QTree_Int_t _96_d;
  logic _96_r;
  assign _96_r = 1'd1;
  MyDTInt_Int_Int_t lizzieLet17_5QVal_Int_3QNone_Int_d;
  logic lizzieLet17_5QVal_Int_3QNone_Int_r;
  MyDTInt_Int_Int_t lizzieLet17_5QVal_Int_3QVal_Int_d;
  logic lizzieLet17_5QVal_Int_3QVal_Int_r;
  MyDTInt_Int_Int_t _95_d;
  logic _95_r;
  assign _95_r = 1'd1;
  MyDTInt_Int_Int_t _94_d;
  logic _94_r;
  assign _94_r = 1'd1;
  MyDTInt_Int_Int_t lizzieLet17_5QVal_Int_3QVal_Int_1_d;
  logic lizzieLet17_5QVal_Int_3QVal_Int_1_r;
  MyDTInt_Int_Int_t lizzieLet17_5QVal_Int_3QVal_Int_2_d;
  logic lizzieLet17_5QVal_Int_3QVal_Int_2_r;
  MyDTInt_Int_Int_t lizzieLet17_5QVal_Int_3QVal_Int_1_argbuf_d;
  logic lizzieLet17_5QVal_Int_3QVal_Int_1_argbuf_r;
  TupMyDTInt_Int_Int___Int___Int_t applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int7_d;
  logic applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int7_r;
  Pointer_CTf_f_Int_t lizzieLet17_5QVal_Int_4QNone_Int_d;
  logic lizzieLet17_5QVal_Int_4QNone_Int_r;
  Pointer_CTf_f_Int_t lizzieLet17_5QVal_Int_4QVal_Int_d;
  logic lizzieLet17_5QVal_Int_4QVal_Int_r;
  Pointer_CTf_f_Int_t lizzieLet17_5QVal_Int_4QNode_Int_d;
  logic lizzieLet17_5QVal_Int_4QNode_Int_r;
  Pointer_CTf_f_Int_t lizzieLet17_5QVal_Int_4QError_Int_d;
  logic lizzieLet17_5QVal_Int_4QError_Int_r;
  Pointer_CTf_f_Int_t lizzieLet17_5QVal_Int_4QError_Int_1_argbuf_d;
  logic lizzieLet17_5QVal_Int_4QError_Int_1_argbuf_r;
  Pointer_CTf_f_Int_t lizzieLet17_5QVal_Int_4QNode_Int_1_argbuf_d;
  logic lizzieLet17_5QVal_Int_4QNode_Int_1_argbuf_r;
  Go_t lizzieLet17_5QVal_Int_5QNone_Int_d;
  logic lizzieLet17_5QVal_Int_5QNone_Int_r;
  Go_t lizzieLet17_5QVal_Int_5QVal_Int_d;
  logic lizzieLet17_5QVal_Int_5QVal_Int_r;
  Go_t lizzieLet17_5QVal_Int_5QNode_Int_d;
  logic lizzieLet17_5QVal_Int_5QNode_Int_r;
  Go_t lizzieLet17_5QVal_Int_5QError_Int_d;
  logic lizzieLet17_5QVal_Int_5QError_Int_r;
  Go_t lizzieLet17_5QVal_Int_5QError_Int_1_d;
  logic lizzieLet17_5QVal_Int_5QError_Int_1_r;
  Go_t lizzieLet17_5QVal_Int_5QError_Int_2_d;
  logic lizzieLet17_5QVal_Int_5QError_Int_2_r;
  QTree_Int_t lizzieLet17_5QVal_Int_5QError_Int_1QError_Int_d;
  logic lizzieLet17_5QVal_Int_5QError_Int_1QError_Int_r;
  QTree_Int_t lizzieLet42_1_argbuf_d;
  logic lizzieLet42_1_argbuf_r;
  Go_t lizzieLet17_5QVal_Int_5QError_Int_2_argbuf_d;
  logic lizzieLet17_5QVal_Int_5QError_Int_2_argbuf_r;
  Go_t lizzieLet17_5QVal_Int_5QNode_Int_1_d;
  logic lizzieLet17_5QVal_Int_5QNode_Int_1_r;
  Go_t lizzieLet17_5QVal_Int_5QNode_Int_2_d;
  logic lizzieLet17_5QVal_Int_5QNode_Int_2_r;
  QTree_Int_t lizzieLet17_5QVal_Int_5QNode_Int_1QError_Int_d;
  logic lizzieLet17_5QVal_Int_5QNode_Int_1QError_Int_r;
  QTree_Int_t lizzieLet41_1_argbuf_d;
  logic lizzieLet41_1_argbuf_r;
  Go_t lizzieLet17_5QVal_Int_5QNode_Int_2_argbuf_d;
  logic lizzieLet17_5QVal_Int_5QNode_Int_2_argbuf_r;
  Go_t lizzieLet17_5QVal_Int_5QVal_Int_1_d;
  logic lizzieLet17_5QVal_Int_5QVal_Int_1_r;
  Go_t lizzieLet17_5QVal_Int_5QVal_Int_2_d;
  logic lizzieLet17_5QVal_Int_5QVal_Int_2_r;
  Go_t lizzieLet17_5QVal_Int_5QVal_Int_1_argbuf_d;
  logic lizzieLet17_5QVal_Int_5QVal_Int_1_argbuf_r;
  TupGo___MyDTInt_Bool___Int_t applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int4_d;
  logic applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int4_r;
  MyDTInt_Bool_t lizzieLet17_5QVal_Int_6QNone_Int_d;
  logic lizzieLet17_5QVal_Int_6QNone_Int_r;
  MyDTInt_Bool_t lizzieLet17_5QVal_Int_6QVal_Int_d;
  logic lizzieLet17_5QVal_Int_6QVal_Int_r;
  MyDTInt_Bool_t _93_d;
  logic _93_r;
  assign _93_r = 1'd1;
  MyDTInt_Bool_t _92_d;
  logic _92_r;
  assign _92_r = 1'd1;
  MyDTInt_Bool_t lizzieLet17_5QVal_Int_6QVal_Int_1_d;
  logic lizzieLet17_5QVal_Int_6QVal_Int_1_r;
  MyDTInt_Bool_t lizzieLet17_5QVal_Int_6QVal_Int_2_d;
  logic lizzieLet17_5QVal_Int_6QVal_Int_2_r;
  MyDTInt_Bool_t lizzieLet17_5QVal_Int_6QVal_Int_1_argbuf_d;
  logic lizzieLet17_5QVal_Int_6QVal_Int_1_argbuf_r;
  QTree_Int_t lizzieLet17_5QVal_Int_7QNone_Int_d;
  logic lizzieLet17_5QVal_Int_7QNone_Int_r;
  QTree_Int_t lizzieLet17_5QVal_Int_7QVal_Int_d;
  logic lizzieLet17_5QVal_Int_7QVal_Int_r;
  QTree_Int_t _91_d;
  logic _91_r;
  assign _91_r = 1'd1;
  QTree_Int_t _90_d;
  logic _90_r;
  assign _90_r = 1'd1;
  QTree_Int_t lizzieLet17_5QVal_Int_7QNone_Int_1_d;
  logic lizzieLet17_5QVal_Int_7QNone_Int_1_r;
  QTree_Int_t lizzieLet17_5QVal_Int_7QNone_Int_2_d;
  logic lizzieLet17_5QVal_Int_7QNone_Int_2_r;
  QTree_Int_t lizzieLet17_5QVal_Int_7QNone_Int_3_d;
  logic lizzieLet17_5QVal_Int_7QNone_Int_3_r;
  QTree_Int_t lizzieLet17_5QVal_Int_7QNone_Int_4_d;
  logic lizzieLet17_5QVal_Int_7QNone_Int_4_r;
  QTree_Int_t lizzieLet17_5QVal_Int_7QNone_Int_5_d;
  logic lizzieLet17_5QVal_Int_7QNone_Int_5_r;
  QTree_Int_t lizzieLet17_5QVal_Int_7QNone_Int_6_d;
  logic lizzieLet17_5QVal_Int_7QNone_Int_6_r;
  QTree_Int_t lizzieLet17_5QVal_Int_7QNone_Int_7_d;
  logic lizzieLet17_5QVal_Int_7QNone_Int_7_r;
  QTree_Int_t lizzieLet17_5QVal_Int_7QNone_Int_8_d;
  logic lizzieLet17_5QVal_Int_7QNone_Int_8_r;
  Int_t vaeL_destruct_d;
  logic vaeL_destruct_r;
  QTree_Int_t _89_d;
  logic _89_r;
  assign _89_r = 1'd1;
  QTree_Int_t lizzieLet17_5QVal_Int_7QNone_Int_1QVal_Int_d;
  logic lizzieLet17_5QVal_Int_7QNone_Int_1QVal_Int_r;
  QTree_Int_t _88_d;
  logic _88_r;
  assign _88_r = 1'd1;
  QTree_Int_t _87_d;
  logic _87_r;
  assign _87_r = 1'd1;
  Int_t _86_d;
  logic _86_r;
  assign _86_r = 1'd1;
  Int_t lizzieLet17_5QVal_Int_7QNone_Int_3QVal_Int_d;
  logic lizzieLet17_5QVal_Int_7QNone_Int_3QVal_Int_r;
  Int_t _85_d;
  logic _85_r;
  assign _85_r = 1'd1;
  Int_t _84_d;
  logic _84_r;
  assign _84_r = 1'd1;
  Int_t lizzieLet17_5QVal_Int_7QNone_Int_3QVal_Int_1_d;
  logic lizzieLet17_5QVal_Int_7QNone_Int_3QVal_Int_1_r;
  Int_t lizzieLet17_5QVal_Int_7QNone_Int_3QVal_Int_2_d;
  logic lizzieLet17_5QVal_Int_7QNone_Int_3QVal_Int_2_r;
  Int_t lizzieLet17_5QVal_Int_7QNone_Int_3QVal_Int_1_argbuf_d;
  logic lizzieLet17_5QVal_Int_7QNone_Int_3QVal_Int_1_argbuf_r;
  MyDTInt_Int_Int_t _83_d;
  logic _83_r;
  assign _83_r = 1'd1;
  MyDTInt_Int_Int_t lizzieLet17_5QVal_Int_7QNone_Int_4QVal_Int_d;
  logic lizzieLet17_5QVal_Int_7QNone_Int_4QVal_Int_r;
  MyDTInt_Int_Int_t _82_d;
  logic _82_r;
  assign _82_r = 1'd1;
  MyDTInt_Int_Int_t _81_d;
  logic _81_r;
  assign _81_r = 1'd1;
  MyDTInt_Int_Int_t lizzieLet17_5QVal_Int_7QNone_Int_4QVal_Int_1_d;
  logic lizzieLet17_5QVal_Int_7QNone_Int_4QVal_Int_1_r;
  MyDTInt_Int_Int_t lizzieLet17_5QVal_Int_7QNone_Int_4QVal_Int_2_d;
  logic lizzieLet17_5QVal_Int_7QNone_Int_4QVal_Int_2_r;
  MyDTInt_Int_Int_t lizzieLet17_5QVal_Int_7QNone_Int_4QVal_Int_1_argbuf_d;
  logic lizzieLet17_5QVal_Int_7QNone_Int_4QVal_Int_1_argbuf_r;
  TupMyDTInt_Int_Int___Int___Int_t applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int5_d;
  logic applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int5_r;
  Pointer_CTf_f_Int_t lizzieLet17_5QVal_Int_7QNone_Int_5QNone_Int_d;
  logic lizzieLet17_5QVal_Int_7QNone_Int_5QNone_Int_r;
  Pointer_CTf_f_Int_t lizzieLet17_5QVal_Int_7QNone_Int_5QVal_Int_d;
  logic lizzieLet17_5QVal_Int_7QNone_Int_5QVal_Int_r;
  Pointer_CTf_f_Int_t lizzieLet17_5QVal_Int_7QNone_Int_5QNode_Int_d;
  logic lizzieLet17_5QVal_Int_7QNone_Int_5QNode_Int_r;
  Pointer_CTf_f_Int_t lizzieLet17_5QVal_Int_7QNone_Int_5QError_Int_d;
  logic lizzieLet17_5QVal_Int_7QNone_Int_5QError_Int_r;
  Pointer_CTf_f_Int_t lizzieLet17_5QVal_Int_7QNone_Int_5QError_Int_1_argbuf_d;
  logic lizzieLet17_5QVal_Int_7QNone_Int_5QError_Int_1_argbuf_r;
  Pointer_CTf_f_Int_t lizzieLet17_5QVal_Int_7QNone_Int_5QNode_Int_1_argbuf_d;
  logic lizzieLet17_5QVal_Int_7QNone_Int_5QNode_Int_1_argbuf_r;
  Pointer_CTf_f_Int_t lizzieLet17_5QVal_Int_7QNone_Int_5QNone_Int_1_argbuf_d;
  logic lizzieLet17_5QVal_Int_7QNone_Int_5QNone_Int_1_argbuf_r;
  Go_t lizzieLet17_5QVal_Int_7QNone_Int_6QNone_Int_d;
  logic lizzieLet17_5QVal_Int_7QNone_Int_6QNone_Int_r;
  Go_t lizzieLet17_5QVal_Int_7QNone_Int_6QVal_Int_d;
  logic lizzieLet17_5QVal_Int_7QNone_Int_6QVal_Int_r;
  Go_t lizzieLet17_5QVal_Int_7QNone_Int_6QNode_Int_d;
  logic lizzieLet17_5QVal_Int_7QNone_Int_6QNode_Int_r;
  Go_t lizzieLet17_5QVal_Int_7QNone_Int_6QError_Int_d;
  logic lizzieLet17_5QVal_Int_7QNone_Int_6QError_Int_r;
  Go_t lizzieLet17_5QVal_Int_7QNone_Int_6QError_Int_1_d;
  logic lizzieLet17_5QVal_Int_7QNone_Int_6QError_Int_1_r;
  Go_t lizzieLet17_5QVal_Int_7QNone_Int_6QError_Int_2_d;
  logic lizzieLet17_5QVal_Int_7QNone_Int_6QError_Int_2_r;
  QTree_Int_t lizzieLet17_5QVal_Int_7QNone_Int_6QError_Int_1QError_Int_d;
  logic lizzieLet17_5QVal_Int_7QNone_Int_6QError_Int_1QError_Int_r;
  QTree_Int_t lizzieLet34_1_argbuf_d;
  logic lizzieLet34_1_argbuf_r;
  Go_t lizzieLet17_5QVal_Int_7QNone_Int_6QError_Int_2_argbuf_d;
  logic lizzieLet17_5QVal_Int_7QNone_Int_6QError_Int_2_argbuf_r;
  Go_t lizzieLet17_5QVal_Int_7QNone_Int_6QNode_Int_1_d;
  logic lizzieLet17_5QVal_Int_7QNone_Int_6QNode_Int_1_r;
  Go_t lizzieLet17_5QVal_Int_7QNone_Int_6QNode_Int_2_d;
  logic lizzieLet17_5QVal_Int_7QNone_Int_6QNode_Int_2_r;
  QTree_Int_t lizzieLet17_5QVal_Int_7QNone_Int_6QNode_Int_1QError_Int_d;
  logic lizzieLet17_5QVal_Int_7QNone_Int_6QNode_Int_1QError_Int_r;
  QTree_Int_t lizzieLet33_1_argbuf_d;
  logic lizzieLet33_1_argbuf_r;
  Go_t lizzieLet17_5QVal_Int_7QNone_Int_6QNode_Int_2_argbuf_d;
  logic lizzieLet17_5QVal_Int_7QNone_Int_6QNode_Int_2_argbuf_r;
  Go_t lizzieLet17_5QVal_Int_7QNone_Int_6QNone_Int_1_argbuf_d;
  logic lizzieLet17_5QVal_Int_7QNone_Int_6QNone_Int_1_argbuf_r;
  Go_t lizzieLet17_5QVal_Int_7QNone_Int_6QVal_Int_1_d;
  logic lizzieLet17_5QVal_Int_7QNone_Int_6QVal_Int_1_r;
  Go_t lizzieLet17_5QVal_Int_7QNone_Int_6QVal_Int_2_d;
  logic lizzieLet17_5QVal_Int_7QNone_Int_6QVal_Int_2_r;
  Go_t lizzieLet17_5QVal_Int_7QNone_Int_6QVal_Int_1_argbuf_d;
  logic lizzieLet17_5QVal_Int_7QNone_Int_6QVal_Int_1_argbuf_r;
  TupGo___MyDTInt_Bool___Int_t applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int3_d;
  logic applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int3_r;
  MyDTInt_Bool_t _80_d;
  logic _80_r;
  assign _80_r = 1'd1;
  MyDTInt_Bool_t lizzieLet17_5QVal_Int_7QNone_Int_7QVal_Int_d;
  logic lizzieLet17_5QVal_Int_7QNone_Int_7QVal_Int_r;
  MyDTInt_Bool_t _79_d;
  logic _79_r;
  assign _79_r = 1'd1;
  MyDTInt_Bool_t _78_d;
  logic _78_r;
  assign _78_r = 1'd1;
  MyDTInt_Bool_t lizzieLet17_5QVal_Int_7QNone_Int_7QVal_Int_1_argbuf_d;
  logic lizzieLet17_5QVal_Int_7QNone_Int_7QVal_Int_1_argbuf_r;
  Pointer_QTree_Int_t lizzieLet17_5QVal_Int_7QNone_Int_8QNone_Int_d;
  logic lizzieLet17_5QVal_Int_7QNone_Int_8QNone_Int_r;
  Pointer_QTree_Int_t _77_d;
  logic _77_r;
  assign _77_r = 1'd1;
  Pointer_QTree_Int_t _76_d;
  logic _76_r;
  assign _76_r = 1'd1;
  Pointer_QTree_Int_t _75_d;
  logic _75_r;
  assign _75_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet17_5QVal_Int_7QNone_Int_8QNone_Int_1_argbuf_d;
  logic lizzieLet17_5QVal_Int_7QNone_Int_8QNone_Int_1_argbuf_r;
  Pointer_QTree_Int_t lizzieLet17_5QVal_Int_8QNone_Int_d;
  logic lizzieLet17_5QVal_Int_8QNone_Int_r;
  Pointer_QTree_Int_t _74_d;
  logic _74_r;
  assign _74_r = 1'd1;
  Pointer_QTree_Int_t _73_d;
  logic _73_r;
  assign _73_r = 1'd1;
  Pointer_QTree_Int_t _72_d;
  logic _72_r;
  assign _72_r = 1'd1;
  Pointer_QTree_Int_t _71_d;
  logic _71_r;
  assign _71_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet17_5QVal_Int_9QVal_Int_d;
  logic lizzieLet17_5QVal_Int_9QVal_Int_r;
  Pointer_QTree_Int_t _70_d;
  logic _70_r;
  assign _70_r = 1'd1;
  Pointer_QTree_Int_t _69_d;
  logic _69_r;
  assign _69_r = 1'd1;
  QTree_Int_t lizzieLet17_6QNone_Int_d;
  logic lizzieLet17_6QNone_Int_r;
  QTree_Int_t lizzieLet17_6QVal_Int_d;
  logic lizzieLet17_6QVal_Int_r;
  QTree_Int_t lizzieLet17_6QNode_Int_d;
  logic lizzieLet17_6QNode_Int_r;
  QTree_Int_t _68_d;
  logic _68_r;
  assign _68_r = 1'd1;
  Pointer_QTree_Int_t _67_d;
  logic _67_r;
  assign _67_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet17_7QVal_Int_d;
  logic lizzieLet17_7QVal_Int_r;
  Pointer_QTree_Int_t lizzieLet17_7QNode_Int_d;
  logic lizzieLet17_7QNode_Int_r;
  Pointer_QTree_Int_t _66_d;
  logic _66_r;
  assign _66_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet17_8QNone_Int_d;
  logic lizzieLet17_8QNone_Int_r;
  Pointer_QTree_Int_t _65_d;
  logic _65_r;
  assign _65_r = 1'd1;
  Pointer_QTree_Int_t _64_d;
  logic _64_r;
  assign _64_r = 1'd1;
  Pointer_QTree_Int_t _63_d;
  logic _63_r;
  assign _63_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet17_9QNone_Int_d;
  logic lizzieLet17_9QNone_Int_r;
  Pointer_QTree_Int_t lizzieLet17_9QVal_Int_d;
  logic lizzieLet17_9QVal_Int_r;
  Pointer_QTree_Int_t _62_d;
  logic _62_r;
  assign _62_r = 1'd1;
  Pointer_QTree_Int_t _61_d;
  logic _61_r;
  assign _61_r = 1'd1;
  Bool_t lizzieLet2_1_argbuf_d;
  logic lizzieLet2_1_argbuf_r;
  Go_t lizzieLet3_1MyFalse_d;
  logic lizzieLet3_1MyFalse_r;
  Go_t lizzieLet3_1MyTrue_d;
  logic lizzieLet3_1MyTrue_r;
  MyBool_t lizzieLet3_1MyFalse_1MyFalse_d;
  logic lizzieLet3_1MyFalse_1MyFalse_r;
  MyBool_t lizzieLet3_1MyTrue_1MyTrue_d;
  logic lizzieLet3_1MyTrue_1MyTrue_r;
  MyBool_t lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_d;
  logic lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_r;
  Pointer_QTree_Int_t q1a8r_destruct_d;
  logic q1a8r_destruct_r;
  Pointer_QTree_Int_t q2a8s_destruct_d;
  logic q2a8s_destruct_r;
  Pointer_QTree_Int_t q3a8t_destruct_d;
  logic q3a8t_destruct_r;
  Pointer_QTree_Int_t q4a8u_destruct_d;
  logic q4a8u_destruct_r;
  QTree_Int_t _60_d;
  logic _60_r;
  assign _60_r = 1'd1;
  QTree_Int_t _59_d;
  logic _59_r;
  assign _59_r = 1'd1;
  QTree_Int_t lizzieLet4_1QNode_Int_d;
  logic lizzieLet4_1QNode_Int_r;
  QTree_Int_t _58_d;
  logic _58_r;
  assign _58_r = 1'd1;
  Go_t lizzieLet4_3QNone_Int_d;
  logic lizzieLet4_3QNone_Int_r;
  Go_t lizzieLet4_3QVal_Int_d;
  logic lizzieLet4_3QVal_Int_r;
  Go_t lizzieLet4_3QNode_Int_d;
  logic lizzieLet4_3QNode_Int_r;
  Go_t lizzieLet4_3QError_Int_d;
  logic lizzieLet4_3QError_Int_r;
  Go_t lizzieLet4_3QError_Int_1_d;
  logic lizzieLet4_3QError_Int_1_r;
  Go_t lizzieLet4_3QError_Int_2_d;
  logic lizzieLet4_3QError_Int_2_r;
  Go_t lizzieLet4_3QError_Int_1_argbuf_d;
  logic lizzieLet4_3QError_Int_1_argbuf_r;
  \Int#_t  lizzieLet4_3QError_Int_1_argbuf_0_d;
  logic lizzieLet4_3QError_Int_1_argbuf_0_r;
  \Int#_t  lizzieLet37_1_1_argbuf_d;
  logic lizzieLet37_1_1_argbuf_r;
  Go_t lizzieLet4_3QError_Int_2_argbuf_d;
  logic lizzieLet4_3QError_Int_2_argbuf_r;
  Go_t lizzieLet4_3QNode_Int_1_argbuf_d;
  logic lizzieLet4_3QNode_Int_1_argbuf_r;
  Go_t lizzieLet4_3QNone_Int_1_d;
  logic lizzieLet4_3QNone_Int_1_r;
  Go_t lizzieLet4_3QNone_Int_2_d;
  logic lizzieLet4_3QNone_Int_2_r;
  Go_t lizzieLet4_3QNone_Int_1_argbuf_d;
  logic lizzieLet4_3QNone_Int_1_argbuf_r;
  \Int#_t  lizzieLet4_3QNone_Int_1_argbuf_0_d;
  logic lizzieLet4_3QNone_Int_1_argbuf_0_r;
  \Int#_t  lizzieLet37_1_argbuf_d;
  logic lizzieLet37_1_argbuf_r;
  Go_t lizzieLet4_3QNone_Int_2_argbuf_d;
  logic lizzieLet4_3QNone_Int_2_argbuf_r;
  C4_t go_13_goMux_choice_d;
  logic go_13_goMux_choice_r;
  Go_t go_13_goMux_data_d;
  logic go_13_goMux_data_r;
  Go_t lizzieLet4_3QVal_Int_1_d;
  logic lizzieLet4_3QVal_Int_1_r;
  Go_t lizzieLet4_3QVal_Int_2_d;
  logic lizzieLet4_3QVal_Int_2_r;
  Go_t lizzieLet4_3QVal_Int_1_argbuf_d;
  logic lizzieLet4_3QVal_Int_1_argbuf_r;
  \Int#_t  lizzieLet4_3QVal_Int_1_argbuf_1_d;
  logic lizzieLet4_3QVal_Int_1_argbuf_1_r;
  \Int#_t  lizzieLet38_1_argbuf_d;
  logic lizzieLet38_1_argbuf_r;
  Go_t lizzieLet4_3QVal_Int_2_argbuf_d;
  logic lizzieLet4_3QVal_Int_2_argbuf_r;
  Pointer_CT$wnnz_t lizzieLet4_4QNone_Int_d;
  logic lizzieLet4_4QNone_Int_r;
  Pointer_CT$wnnz_t lizzieLet4_4QVal_Int_d;
  logic lizzieLet4_4QVal_Int_r;
  Pointer_CT$wnnz_t lizzieLet4_4QNode_Int_d;
  logic lizzieLet4_4QNode_Int_r;
  Pointer_CT$wnnz_t lizzieLet4_4QError_Int_d;
  logic lizzieLet4_4QError_Int_r;
  Pointer_CT$wnnz_t lizzieLet4_4QError_Int_1_argbuf_d;
  logic lizzieLet4_4QError_Int_1_argbuf_r;
  CT$wnnz_t lizzieLet4_4QNode_Int_1q4a8u_1q3a8t_1q2a8s_1Lcall_$wnnz3_d;
  logic lizzieLet4_4QNode_Int_1q4a8u_1q3a8t_1q2a8s_1Lcall_$wnnz3_r;
  CT$wnnz_t lizzieLet5_1_argbuf_d;
  logic lizzieLet5_1_argbuf_r;
  Pointer_CT$wnnz_t lizzieLet4_4QNone_Int_1_argbuf_d;
  logic lizzieLet4_4QNone_Int_1_argbuf_r;
  Pointer_CT$wnnz_t lizzieLet4_4QVal_Int_1_argbuf_d;
  logic lizzieLet4_4QVal_Int_1_argbuf_r;
  \Int#_t  wwsmn_4_destruct_d;
  logic wwsmn_4_destruct_r;
  \Int#_t  ww1XmW_2_destruct_d;
  logic ww1XmW_2_destruct_r;
  \Int#_t  ww2XmZ_1_destruct_d;
  logic ww2XmZ_1_destruct_r;
  Pointer_CT$wnnz_t sc_0_6_destruct_d;
  logic sc_0_6_destruct_r;
  \Int#_t  wwsmn_3_destruct_d;
  logic wwsmn_3_destruct_r;
  \Int#_t  ww1XmW_1_destruct_d;
  logic ww1XmW_1_destruct_r;
  Pointer_CT$wnnz_t sc_0_5_destruct_d;
  logic sc_0_5_destruct_r;
  Pointer_QTree_Int_t q4a8u_3_destruct_d;
  logic q4a8u_3_destruct_r;
  \Int#_t  wwsmn_2_destruct_d;
  logic wwsmn_2_destruct_r;
  Pointer_CT$wnnz_t sc_0_4_destruct_d;
  logic sc_0_4_destruct_r;
  Pointer_QTree_Int_t q4a8u_2_destruct_d;
  logic q4a8u_2_destruct_r;
  Pointer_QTree_Int_t q3a8t_2_destruct_d;
  logic q3a8t_2_destruct_r;
  Pointer_CT$wnnz_t sc_0_3_destruct_d;
  logic sc_0_3_destruct_r;
  Pointer_QTree_Int_t q4a8u_1_destruct_d;
  logic q4a8u_1_destruct_r;
  Pointer_QTree_Int_t q3a8t_1_destruct_d;
  logic q3a8t_1_destruct_r;
  Pointer_QTree_Int_t q2a8s_1_destruct_d;
  logic q2a8s_1_destruct_r;
  CT$wnnz_t _57_d;
  logic _57_r;
  assign _57_r = 1'd1;
  CT$wnnz_t lizzieLet58_1Lcall_$wnnz3_d;
  logic lizzieLet58_1Lcall_$wnnz3_r;
  CT$wnnz_t lizzieLet58_1Lcall_$wnnz2_d;
  logic lizzieLet58_1Lcall_$wnnz2_r;
  CT$wnnz_t lizzieLet58_1Lcall_$wnnz1_d;
  logic lizzieLet58_1Lcall_$wnnz1_r;
  CT$wnnz_t lizzieLet58_1Lcall_$wnnz0_d;
  logic lizzieLet58_1Lcall_$wnnz0_r;
  Go_t _56_d;
  logic _56_r;
  assign _56_r = 1'd1;
  Go_t lizzieLet58_3Lcall_$wnnz3_d;
  logic lizzieLet58_3Lcall_$wnnz3_r;
  Go_t lizzieLet58_3Lcall_$wnnz2_d;
  logic lizzieLet58_3Lcall_$wnnz2_r;
  Go_t lizzieLet58_3Lcall_$wnnz1_d;
  logic lizzieLet58_3Lcall_$wnnz1_r;
  Go_t lizzieLet58_3Lcall_$wnnz0_d;
  logic lizzieLet58_3Lcall_$wnnz0_r;
  Go_t lizzieLet58_3Lcall_$wnnz0_1_argbuf_d;
  logic lizzieLet58_3Lcall_$wnnz0_1_argbuf_r;
  Go_t lizzieLet58_3Lcall_$wnnz1_1_argbuf_d;
  logic lizzieLet58_3Lcall_$wnnz1_1_argbuf_r;
  Go_t lizzieLet58_3Lcall_$wnnz2_1_argbuf_d;
  logic lizzieLet58_3Lcall_$wnnz2_1_argbuf_r;
  Go_t lizzieLet58_3Lcall_$wnnz3_1_argbuf_d;
  logic lizzieLet58_3Lcall_$wnnz3_1_argbuf_r;
  \Int#_t  lizzieLet58_4L$wnnzsbos_d;
  logic lizzieLet58_4L$wnnzsbos_r;
  \Int#_t  lizzieLet58_4Lcall_$wnnz3_d;
  logic lizzieLet58_4Lcall_$wnnz3_r;
  \Int#_t  lizzieLet58_4Lcall_$wnnz2_d;
  logic lizzieLet58_4Lcall_$wnnz2_r;
  \Int#_t  lizzieLet58_4Lcall_$wnnz1_d;
  logic lizzieLet58_4Lcall_$wnnz1_r;
  \Int#_t  lizzieLet58_4Lcall_$wnnz0_d;
  logic lizzieLet58_4Lcall_$wnnz0_r;
  \Int#_t  lizzieLet58_4L$wnnzsbos_1_merge_merge_fork_1_d;
  logic lizzieLet58_4L$wnnzsbos_1_merge_merge_fork_1_r;
  \Int#_t  lizzieLet58_4L$wnnzsbos_1_merge_merge_fork_2_d;
  logic lizzieLet58_4L$wnnzsbos_1_merge_merge_fork_2_r;
  Go_t call_$wnnz_goConst_d;
  logic call_$wnnz_goConst_r;
  \Int#_t  \$wnnz_resbuf_d ;
  logic \$wnnz_resbuf_r ;
  CT$wnnz_t lizzieLet58_4Lcall_$wnnz3_1sc_0_3_1q4a8u_1_1q3a8t_1_1Lcall_$wnnz2_d;
  logic lizzieLet58_4Lcall_$wnnz3_1sc_0_3_1q4a8u_1_1q3a8t_1_1Lcall_$wnnz2_r;
  CT$wnnz_t lizzieLet59_1_argbuf_d;
  logic lizzieLet59_1_argbuf_r;
  Pointer_QTree_Int_t es_5_2_destruct_d;
  logic es_5_2_destruct_r;
  Pointer_QTree_Int_t es_6_4_destruct_d;
  logic es_6_4_destruct_r;
  Pointer_QTree_Int_t es_7_3_destruct_d;
  logic es_7_3_destruct_r;
  \Pointer_CTf''''''''''''_f''''''''''''_Int_t  sc_0_10_destruct_d;
  logic sc_0_10_destruct_r;
  Pointer_QTree_Int_t es_6_3_destruct_d;
  logic es_6_3_destruct_r;
  Pointer_QTree_Int_t es_7_2_destruct_d;
  logic es_7_2_destruct_r;
  \Pointer_CTf''''''''''''_f''''''''''''_Int_t  sc_0_9_destruct_d;
  logic sc_0_9_destruct_r;
  Pointer_QTree_Int_t q1aft_3_destruct_d;
  logic q1aft_3_destruct_r;
  Pointer_QTree_Int_t t1afy_3_destruct_d;
  logic t1afy_3_destruct_r;
  MyDTInt_Bool_t is_zafl_4_destruct_d;
  logic is_zafl_4_destruct_r;
  MyDTInt_Int_Int_t op_addafm_4_destruct_d;
  logic op_addafm_4_destruct_r;
  Pointer_QTree_Int_t es_7_1_destruct_d;
  logic es_7_1_destruct_r;
  \Pointer_CTf''''''''''''_f''''''''''''_Int_t  sc_0_8_destruct_d;
  logic sc_0_8_destruct_r;
  Pointer_QTree_Int_t q1aft_2_destruct_d;
  logic q1aft_2_destruct_r;
  Pointer_QTree_Int_t t1afy_2_destruct_d;
  logic t1afy_2_destruct_r;
  MyDTInt_Bool_t is_zafl_3_destruct_d;
  logic is_zafl_3_destruct_r;
  MyDTInt_Int_Int_t op_addafm_3_destruct_d;
  logic op_addafm_3_destruct_r;
  Pointer_QTree_Int_t q2afu_2_destruct_d;
  logic q2afu_2_destruct_r;
  Pointer_QTree_Int_t t2afz_2_destruct_d;
  logic t2afz_2_destruct_r;
  \Pointer_CTf''''''''''''_f''''''''''''_Int_t  sc_0_7_destruct_d;
  logic sc_0_7_destruct_r;
  Pointer_QTree_Int_t q1aft_1_destruct_d;
  logic q1aft_1_destruct_r;
  Pointer_QTree_Int_t t1afy_1_destruct_d;
  logic t1afy_1_destruct_r;
  MyDTInt_Bool_t is_zafl_2_destruct_d;
  logic is_zafl_2_destruct_r;
  MyDTInt_Int_Int_t op_addafm_2_destruct_d;
  logic op_addafm_2_destruct_r;
  Pointer_QTree_Int_t q2afu_1_destruct_d;
  logic q2afu_1_destruct_r;
  Pointer_QTree_Int_t t2afz_1_destruct_d;
  logic t2afz_1_destruct_r;
  Pointer_QTree_Int_t q3afv_1_destruct_d;
  logic q3afv_1_destruct_r;
  Pointer_QTree_Int_t t3afA_1_destruct_d;
  logic t3afA_1_destruct_r;
  \CTf''''''''''''_f''''''''''''_Int_t  _55_d;
  logic _55_r;
  assign _55_r = 1'd1;
  \CTf''''''''''''_f''''''''''''_Int_t  \lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int3_d ;
  logic \lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int3_r ;
  \CTf''''''''''''_f''''''''''''_Int_t  \lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int2_d ;
  logic \lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int2_r ;
  \CTf''''''''''''_f''''''''''''_Int_t  \lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int1_d ;
  logic \lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int1_r ;
  \CTf''''''''''''_f''''''''''''_Int_t  \lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int0_d ;
  logic \lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int0_r ;
  Go_t _54_d;
  logic _54_r;
  assign _54_r = 1'd1;
  Go_t \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int3_d ;
  logic \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int3_r ;
  Go_t \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int2_d ;
  logic \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int2_r ;
  Go_t \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int1_d ;
  logic \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int1_r ;
  Go_t \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int0_d ;
  logic \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int0_r ;
  Go_t \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int0_1_argbuf_d ;
  logic \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int0_1_argbuf_r ;
  Go_t \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int1_1_argbuf_d ;
  logic \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int1_1_argbuf_r ;
  Go_t \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int2_1_argbuf_d ;
  logic \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int2_1_argbuf_r ;
  Go_t \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int3_1_argbuf_d ;
  logic \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int3_1_argbuf_r ;
  Pointer_QTree_Int_t \lizzieLet62_4Lf''''''''''''_f''''''''''''_Intsbos_d ;
  logic \lizzieLet62_4Lf''''''''''''_f''''''''''''_Intsbos_r ;
  Pointer_QTree_Int_t \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int3_d ;
  logic \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int3_r ;
  Pointer_QTree_Int_t \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int2_d ;
  logic \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int2_r ;
  Pointer_QTree_Int_t \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int1_d ;
  logic \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int1_r ;
  Pointer_QTree_Int_t \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int0_d ;
  logic \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int0_r ;
  QTree_Int_t \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int0_1es_5_2_1es_6_4_1es_7_3_1QNode_Int_d ;
  logic \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int0_1es_5_2_1es_6_4_1es_7_3_1QNode_Int_r ;
  QTree_Int_t lizzieLet66_1_argbuf_d;
  logic lizzieLet66_1_argbuf_r;
  \CTf''''''''''''_f''''''''''''_Int_t  \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int1_1es_6_3_1es_7_2_1sc_0_9_1Lcall_f''''''''''''_f''''''''''''_Int0_d ;
  logic \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int1_1es_6_3_1es_7_2_1sc_0_9_1Lcall_f''''''''''''_f''''''''''''_Int0_r ;
  \CTf''''''''''''_f''''''''''''_Int_t  lizzieLet65_1_argbuf_d;
  logic lizzieLet65_1_argbuf_r;
  \CTf''''''''''''_f''''''''''''_Int_t  \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int2_1es_7_1_1sc_0_8_1q1aft_2_1t1afy_2_1is_zafl_3_1op_addafm_3_1Lcall_f''''''''''''_f''''''''''''_Int1_d ;
  logic \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int2_1es_7_1_1sc_0_8_1q1aft_2_1t1afy_2_1is_zafl_3_1op_addafm_3_1Lcall_f''''''''''''_f''''''''''''_Int1_r ;
  \CTf''''''''''''_f''''''''''''_Int_t  lizzieLet64_1_argbuf_d;
  logic lizzieLet64_1_argbuf_r;
  \CTf''''''''''''_f''''''''''''_Int_t  \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int3_1sc_0_7_1q1aft_1_1t1afy_1_1is_zafl_2_1op_addafm_2_1q2afu_1_1t2afz_1_1Lcall_f''''''''''''_f''''''''''''_Int2_d ;
  logic \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int3_1sc_0_7_1q1aft_1_1t1afy_1_1is_zafl_2_1op_addafm_2_1q2afu_1_1t2afz_1_1Lcall_f''''''''''''_f''''''''''''_Int2_r ;
  \CTf''''''''''''_f''''''''''''_Int_t  lizzieLet63_1_argbuf_d;
  logic lizzieLet63_1_argbuf_r;
  Pointer_QTree_Int_t \lizzieLet62_4Lf''''''''''''_f''''''''''''_Intsbos_1_merge_merge_fork_1_d ;
  logic \lizzieLet62_4Lf''''''''''''_f''''''''''''_Intsbos_1_merge_merge_fork_1_r ;
  Pointer_QTree_Int_t \lizzieLet62_4Lf''''''''''''_f''''''''''''_Intsbos_1_merge_merge_fork_2_d ;
  logic \lizzieLet62_4Lf''''''''''''_f''''''''''''_Intsbos_1_merge_merge_fork_2_r ;
  Go_t \call_f''''''''''''_f''''''''''''_Int_goConst_d ;
  logic \call_f''''''''''''_f''''''''''''_Int_goConst_r ;
  Pointer_QTree_Int_t es_35_destruct_d;
  logic es_35_destruct_r;
  Pointer_QTree_Int_t es_36_1_destruct_d;
  logic es_36_1_destruct_r;
  Pointer_QTree_Int_t es_37_2_destruct_d;
  logic es_37_2_destruct_r;
  Pointer_CTf_f_Int_t sc_0_14_destruct_d;
  logic sc_0_14_destruct_r;
  Pointer_QTree_Int_t es_36_destruct_d;
  logic es_36_destruct_r;
  Pointer_QTree_Int_t es_37_1_destruct_d;
  logic es_37_1_destruct_r;
  Pointer_CTf_f_Int_t sc_0_13_destruct_d;
  logic sc_0_13_destruct_r;
  Pointer_QTree_Int_t q1af0_3_destruct_d;
  logic q1af0_3_destruct_r;
  Pointer_QTree_Int_t t1afa_3_destruct_d;
  logic t1afa_3_destruct_r;
  Pointer_QTree_Int_t \t1'aff_3_destruct_d ;
  logic \t1'aff_3_destruct_r ;
  MyDTInt_Bool_t is_zaet_4_destruct_d;
  logic is_zaet_4_destruct_r;
  MyDTInt_Int_Int_t op_addaeu_4_destruct_d;
  logic op_addaeu_4_destruct_r;
  Pointer_QTree_Int_t es_37_destruct_d;
  logic es_37_destruct_r;
  Pointer_CTf_f_Int_t sc_0_12_destruct_d;
  logic sc_0_12_destruct_r;
  Pointer_QTree_Int_t q1af0_2_destruct_d;
  logic q1af0_2_destruct_r;
  Pointer_QTree_Int_t t1afa_2_destruct_d;
  logic t1afa_2_destruct_r;
  Pointer_QTree_Int_t \t1'aff_2_destruct_d ;
  logic \t1'aff_2_destruct_r ;
  MyDTInt_Bool_t is_zaet_3_destruct_d;
  logic is_zaet_3_destruct_r;
  MyDTInt_Int_Int_t op_addaeu_3_destruct_d;
  logic op_addaeu_3_destruct_r;
  Pointer_QTree_Int_t q2af1_2_destruct_d;
  logic q2af1_2_destruct_r;
  Pointer_QTree_Int_t t2afb_2_destruct_d;
  logic t2afb_2_destruct_r;
  Pointer_QTree_Int_t \t2'afg_2_destruct_d ;
  logic \t2'afg_2_destruct_r ;
  Pointer_CTf_f_Int_t sc_0_11_destruct_d;
  logic sc_0_11_destruct_r;
  Pointer_QTree_Int_t q1af0_1_destruct_d;
  logic q1af0_1_destruct_r;
  Pointer_QTree_Int_t t1afa_1_destruct_d;
  logic t1afa_1_destruct_r;
  Pointer_QTree_Int_t \t1'aff_1_destruct_d ;
  logic \t1'aff_1_destruct_r ;
  MyDTInt_Bool_t is_zaet_2_destruct_d;
  logic is_zaet_2_destruct_r;
  MyDTInt_Int_Int_t op_addaeu_2_destruct_d;
  logic op_addaeu_2_destruct_r;
  Pointer_QTree_Int_t q2af1_1_destruct_d;
  logic q2af1_1_destruct_r;
  Pointer_QTree_Int_t t2afb_1_destruct_d;
  logic t2afb_1_destruct_r;
  Pointer_QTree_Int_t \t2'afg_1_destruct_d ;
  logic \t2'afg_1_destruct_r ;
  Pointer_QTree_Int_t q3af2_1_destruct_d;
  logic q3af2_1_destruct_r;
  Pointer_QTree_Int_t t3afc_1_destruct_d;
  logic t3afc_1_destruct_r;
  Pointer_QTree_Int_t \t3'afh_1_destruct_d ;
  logic \t3'afh_1_destruct_r ;
  CTf_f_Int_t _53_d;
  logic _53_r;
  assign _53_r = 1'd1;
  CTf_f_Int_t lizzieLet67_1Lcall_f_f_Int3_d;
  logic lizzieLet67_1Lcall_f_f_Int3_r;
  CTf_f_Int_t lizzieLet67_1Lcall_f_f_Int2_d;
  logic lizzieLet67_1Lcall_f_f_Int2_r;
  CTf_f_Int_t lizzieLet67_1Lcall_f_f_Int1_d;
  logic lizzieLet67_1Lcall_f_f_Int1_r;
  CTf_f_Int_t lizzieLet67_1Lcall_f_f_Int0_d;
  logic lizzieLet67_1Lcall_f_f_Int0_r;
  Go_t _52_d;
  logic _52_r;
  assign _52_r = 1'd1;
  Go_t lizzieLet67_3Lcall_f_f_Int3_d;
  logic lizzieLet67_3Lcall_f_f_Int3_r;
  Go_t lizzieLet67_3Lcall_f_f_Int2_d;
  logic lizzieLet67_3Lcall_f_f_Int2_r;
  Go_t lizzieLet67_3Lcall_f_f_Int1_d;
  logic lizzieLet67_3Lcall_f_f_Int1_r;
  Go_t lizzieLet67_3Lcall_f_f_Int0_d;
  logic lizzieLet67_3Lcall_f_f_Int0_r;
  Go_t lizzieLet67_3Lcall_f_f_Int0_1_argbuf_d;
  logic lizzieLet67_3Lcall_f_f_Int0_1_argbuf_r;
  Go_t lizzieLet67_3Lcall_f_f_Int1_1_argbuf_d;
  logic lizzieLet67_3Lcall_f_f_Int1_1_argbuf_r;
  Go_t lizzieLet67_3Lcall_f_f_Int2_1_argbuf_d;
  logic lizzieLet67_3Lcall_f_f_Int2_1_argbuf_r;
  Go_t lizzieLet67_3Lcall_f_f_Int3_1_argbuf_d;
  logic lizzieLet67_3Lcall_f_f_Int3_1_argbuf_r;
  Pointer_QTree_Int_t lizzieLet67_4Lf_f_Intsbos_d;
  logic lizzieLet67_4Lf_f_Intsbos_r;
  Pointer_QTree_Int_t lizzieLet67_4Lcall_f_f_Int3_d;
  logic lizzieLet67_4Lcall_f_f_Int3_r;
  Pointer_QTree_Int_t lizzieLet67_4Lcall_f_f_Int2_d;
  logic lizzieLet67_4Lcall_f_f_Int2_r;
  Pointer_QTree_Int_t lizzieLet67_4Lcall_f_f_Int1_d;
  logic lizzieLet67_4Lcall_f_f_Int1_r;
  Pointer_QTree_Int_t lizzieLet67_4Lcall_f_f_Int0_d;
  logic lizzieLet67_4Lcall_f_f_Int0_r;
  QTree_Int_t lizzieLet67_4Lcall_f_f_Int0_1es_35_1es_36_1_1es_37_2_1QNode_Int_d;
  logic lizzieLet67_4Lcall_f_f_Int0_1es_35_1es_36_1_1es_37_2_1QNode_Int_r;
  QTree_Int_t lizzieLet71_1_argbuf_d;
  logic lizzieLet71_1_argbuf_r;
  CTf_f_Int_t lizzieLet67_4Lcall_f_f_Int1_1es_36_1es_37_1_1sc_0_13_1Lcall_f_f_Int0_d;
  logic lizzieLet67_4Lcall_f_f_Int1_1es_36_1es_37_1_1sc_0_13_1Lcall_f_f_Int0_r;
  CTf_f_Int_t lizzieLet70_1_argbuf_d;
  logic lizzieLet70_1_argbuf_r;
  CTf_f_Int_t \lizzieLet67_4Lcall_f_f_Int2_1es_37_1sc_0_12_1q1af0_2_1t1afa_2_1t1'aff_2_1is_zaet_3_1op_addaeu_3_1Lcall_f_f_Int1_d ;
  logic \lizzieLet67_4Lcall_f_f_Int2_1es_37_1sc_0_12_1q1af0_2_1t1afa_2_1t1'aff_2_1is_zaet_3_1op_addaeu_3_1Lcall_f_f_Int1_r ;
  CTf_f_Int_t lizzieLet69_1_argbuf_d;
  logic lizzieLet69_1_argbuf_r;
  CTf_f_Int_t \lizzieLet67_4Lcall_f_f_Int3_1sc_0_11_1q1af0_1_1t1afa_1_1t1'aff_1_1is_zaet_2_1op_addaeu_2_1q2af1_1_1t2afb_1_1t2'afg_1_1Lcall_f_f_Int2_d ;
  logic \lizzieLet67_4Lcall_f_f_Int3_1sc_0_11_1q1af0_1_1t1afa_1_1t1'aff_1_1is_zaet_2_1op_addaeu_2_1q2af1_1_1t2afb_1_1t2'afg_1_1Lcall_f_f_Int2_r ;
  CTf_f_Int_t lizzieLet68_1_argbuf_d;
  logic lizzieLet68_1_argbuf_r;
  Pointer_QTree_Int_t lizzieLet67_4Lf_f_Intsbos_1_merge_merge_merge_fork_1_d;
  logic lizzieLet67_4Lf_f_Intsbos_1_merge_merge_merge_fork_1_r;
  Pointer_QTree_Int_t lizzieLet67_4Lf_f_Intsbos_1_merge_merge_merge_fork_2_d;
  logic lizzieLet67_4Lf_f_Intsbos_1_merge_merge_merge_fork_2_r;
  Go_t call_f_f_Int_goConst_d;
  logic call_f_f_Int_goConst_r;
  Pointer_QTree_Int_t f_f_Int_resbuf_d;
  logic f_f_Int_resbuf_r;
  Pointer_QTree_Int_t q1aft_destruct_d;
  logic q1aft_destruct_r;
  Pointer_QTree_Int_t q2afu_destruct_d;
  logic q2afu_destruct_r;
  Pointer_QTree_Int_t q3afv_destruct_d;
  logic q3afv_destruct_r;
  Pointer_QTree_Int_t q5afw_destruct_d;
  logic q5afw_destruct_r;
  Int_t v1afn_destruct_d;
  logic v1afn_destruct_r;
  QTree_Int_t _51_d;
  logic _51_r;
  assign _51_r = 1'd1;
  QTree_Int_t lizzieLet6_1QVal_Int_d;
  logic lizzieLet6_1QVal_Int_r;
  QTree_Int_t lizzieLet6_1QNode_Int_d;
  logic lizzieLet6_1QNode_Int_r;
  QTree_Int_t _50_d;
  logic _50_r;
  assign _50_r = 1'd1;
  Go_t lizzieLet6_3QNone_Int_d;
  logic lizzieLet6_3QNone_Int_r;
  Go_t lizzieLet6_3QVal_Int_d;
  logic lizzieLet6_3QVal_Int_r;
  Go_t lizzieLet6_3QNode_Int_d;
  logic lizzieLet6_3QNode_Int_r;
  Go_t lizzieLet6_3QError_Int_d;
  logic lizzieLet6_3QError_Int_r;
  Go_t lizzieLet6_3QError_Int_1_d;
  logic lizzieLet6_3QError_Int_1_r;
  Go_t lizzieLet6_3QError_Int_2_d;
  logic lizzieLet6_3QError_Int_2_r;
  QTree_Int_t lizzieLet6_3QError_Int_1QError_Int_d;
  logic lizzieLet6_3QError_Int_1QError_Int_r;
  QTree_Int_t lizzieLet16_1_argbuf_d;
  logic lizzieLet16_1_argbuf_r;
  Go_t lizzieLet6_3QError_Int_2_argbuf_d;
  logic lizzieLet6_3QError_Int_2_argbuf_r;
  Go_t lizzieLet6_3QNone_Int_1_argbuf_d;
  logic lizzieLet6_3QNone_Int_1_argbuf_r;
  C11_t go_14_goMux_choice_d;
  logic go_14_goMux_choice_r;
  Go_t go_14_goMux_data_d;
  logic go_14_goMux_data_r;
  MyDTInt_Bool_t _49_d;
  logic _49_r;
  assign _49_r = 1'd1;
  MyDTInt_Bool_t lizzieLet6_4QVal_Int_d;
  logic lizzieLet6_4QVal_Int_r;
  MyDTInt_Bool_t lizzieLet6_4QNode_Int_d;
  logic lizzieLet6_4QNode_Int_r;
  MyDTInt_Bool_t _48_d;
  logic _48_r;
  assign _48_r = 1'd1;
  QTree_Int_t _47_d;
  logic _47_r;
  assign _47_r = 1'd1;
  QTree_Int_t lizzieLet6_5QVal_Int_d;
  logic lizzieLet6_5QVal_Int_r;
  QTree_Int_t lizzieLet6_5QNode_Int_d;
  logic lizzieLet6_5QNode_Int_r;
  QTree_Int_t _46_d;
  logic _46_r;
  assign _46_r = 1'd1;
  QTree_Int_t lizzieLet6_5QNode_Int_1_d;
  logic lizzieLet6_5QNode_Int_1_r;
  QTree_Int_t lizzieLet6_5QNode_Int_2_d;
  logic lizzieLet6_5QNode_Int_2_r;
  QTree_Int_t lizzieLet6_5QNode_Int_3_d;
  logic lizzieLet6_5QNode_Int_3_r;
  QTree_Int_t lizzieLet6_5QNode_Int_4_d;
  logic lizzieLet6_5QNode_Int_4_r;
  QTree_Int_t lizzieLet6_5QNode_Int_5_d;
  logic lizzieLet6_5QNode_Int_5_r;
  QTree_Int_t lizzieLet6_5QNode_Int_6_d;
  logic lizzieLet6_5QNode_Int_6_r;
  QTree_Int_t lizzieLet6_5QNode_Int_7_d;
  logic lizzieLet6_5QNode_Int_7_r;
  QTree_Int_t lizzieLet6_5QNode_Int_8_d;
  logic lizzieLet6_5QNode_Int_8_r;
  QTree_Int_t lizzieLet6_5QNode_Int_9_d;
  logic lizzieLet6_5QNode_Int_9_r;
  QTree_Int_t lizzieLet6_5QNode_Int_10_d;
  logic lizzieLet6_5QNode_Int_10_r;
  QTree_Int_t lizzieLet6_5QNode_Int_11_d;
  logic lizzieLet6_5QNode_Int_11_r;
  Pointer_QTree_Int_t _45_d;
  logic _45_r;
  assign _45_r = 1'd1;
  Pointer_QTree_Int_t _44_d;
  logic _44_r;
  assign _44_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet6_5QNode_Int_10QNode_Int_d;
  logic lizzieLet6_5QNode_Int_10QNode_Int_r;
  Pointer_QTree_Int_t _43_d;
  logic _43_r;
  assign _43_r = 1'd1;
  Pointer_QTree_Int_t _42_d;
  logic _42_r;
  assign _42_r = 1'd1;
  Pointer_QTree_Int_t _41_d;
  logic _41_r;
  assign _41_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet6_5QNode_Int_11QNode_Int_d;
  logic lizzieLet6_5QNode_Int_11QNode_Int_r;
  Pointer_QTree_Int_t _40_d;
  logic _40_r;
  assign _40_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet6_5QNode_Int_11QNode_Int_1_argbuf_d;
  logic lizzieLet6_5QNode_Int_11QNode_Int_1_argbuf_r;
  Pointer_QTree_Int_t t1afy_destruct_d;
  logic t1afy_destruct_r;
  Pointer_QTree_Int_t t2afz_destruct_d;
  logic t2afz_destruct_r;
  Pointer_QTree_Int_t t3afA_destruct_d;
  logic t3afA_destruct_r;
  Pointer_QTree_Int_t t5afB_destruct_d;
  logic t5afB_destruct_r;
  QTree_Int_t _39_d;
  logic _39_r;
  assign _39_r = 1'd1;
  QTree_Int_t _38_d;
  logic _38_r;
  assign _38_r = 1'd1;
  QTree_Int_t lizzieLet6_5QNode_Int_1QNode_Int_d;
  logic lizzieLet6_5QNode_Int_1QNode_Int_r;
  QTree_Int_t _37_d;
  logic _37_r;
  assign _37_r = 1'd1;
  Go_t lizzieLet6_5QNode_Int_3QNone_Int_d;
  logic lizzieLet6_5QNode_Int_3QNone_Int_r;
  Go_t lizzieLet6_5QNode_Int_3QVal_Int_d;
  logic lizzieLet6_5QNode_Int_3QVal_Int_r;
  Go_t lizzieLet6_5QNode_Int_3QNode_Int_d;
  logic lizzieLet6_5QNode_Int_3QNode_Int_r;
  Go_t lizzieLet6_5QNode_Int_3QError_Int_d;
  logic lizzieLet6_5QNode_Int_3QError_Int_r;
  Go_t lizzieLet6_5QNode_Int_3QError_Int_1_d;
  logic lizzieLet6_5QNode_Int_3QError_Int_1_r;
  Go_t lizzieLet6_5QNode_Int_3QError_Int_2_d;
  logic lizzieLet6_5QNode_Int_3QError_Int_2_r;
  QTree_Int_t lizzieLet6_5QNode_Int_3QError_Int_1QError_Int_d;
  logic lizzieLet6_5QNode_Int_3QError_Int_1QError_Int_r;
  QTree_Int_t lizzieLet15_1_argbuf_d;
  logic lizzieLet15_1_argbuf_r;
  Go_t lizzieLet6_5QNode_Int_3QError_Int_2_argbuf_d;
  logic lizzieLet6_5QNode_Int_3QError_Int_2_argbuf_r;
  Go_t lizzieLet6_5QNode_Int_3QNode_Int_1_argbuf_d;
  logic lizzieLet6_5QNode_Int_3QNode_Int_1_argbuf_r;
  Go_t lizzieLet6_5QNode_Int_3QNone_Int_1_argbuf_d;
  logic lizzieLet6_5QNode_Int_3QNone_Int_1_argbuf_r;
  Go_t lizzieLet6_5QNode_Int_3QVal_Int_1_d;
  logic lizzieLet6_5QNode_Int_3QVal_Int_1_r;
  Go_t lizzieLet6_5QNode_Int_3QVal_Int_2_d;
  logic lizzieLet6_5QNode_Int_3QVal_Int_2_r;
  QTree_Int_t lizzieLet6_5QNode_Int_3QVal_Int_1QError_Int_d;
  logic lizzieLet6_5QNode_Int_3QVal_Int_1QError_Int_r;
  QTree_Int_t lizzieLet13_1_argbuf_d;
  logic lizzieLet13_1_argbuf_r;
  Go_t lizzieLet6_5QNode_Int_3QVal_Int_2_argbuf_d;
  logic lizzieLet6_5QNode_Int_3QVal_Int_2_argbuf_r;
  MyDTInt_Bool_t _36_d;
  logic _36_r;
  assign _36_r = 1'd1;
  MyDTInt_Bool_t _35_d;
  logic _35_r;
  assign _35_r = 1'd1;
  MyDTInt_Bool_t lizzieLet6_5QNode_Int_4QNode_Int_d;
  logic lizzieLet6_5QNode_Int_4QNode_Int_r;
  MyDTInt_Bool_t _34_d;
  logic _34_r;
  assign _34_r = 1'd1;
  MyDTInt_Bool_t lizzieLet6_5QNode_Int_4QNode_Int_1_d;
  logic lizzieLet6_5QNode_Int_4QNode_Int_1_r;
  MyDTInt_Bool_t lizzieLet6_5QNode_Int_4QNode_Int_2_d;
  logic lizzieLet6_5QNode_Int_4QNode_Int_2_r;
  MyDTInt_Bool_t lizzieLet6_5QNode_Int_4QNode_Int_2_argbuf_d;
  logic lizzieLet6_5QNode_Int_4QNode_Int_2_argbuf_r;
  MyDTInt_Int_Int_t _33_d;
  logic _33_r;
  assign _33_r = 1'd1;
  MyDTInt_Int_Int_t _32_d;
  logic _32_r;
  assign _32_r = 1'd1;
  MyDTInt_Int_Int_t lizzieLet6_5QNode_Int_5QNode_Int_d;
  logic lizzieLet6_5QNode_Int_5QNode_Int_r;
  MyDTInt_Int_Int_t _31_d;
  logic _31_r;
  assign _31_r = 1'd1;
  MyDTInt_Int_Int_t lizzieLet6_5QNode_Int_5QNode_Int_1_d;
  logic lizzieLet6_5QNode_Int_5QNode_Int_1_r;
  MyDTInt_Int_Int_t lizzieLet6_5QNode_Int_5QNode_Int_2_d;
  logic lizzieLet6_5QNode_Int_5QNode_Int_2_r;
  MyDTInt_Int_Int_t lizzieLet6_5QNode_Int_5QNode_Int_2_argbuf_d;
  logic lizzieLet6_5QNode_Int_5QNode_Int_2_argbuf_r;
  Pointer_QTree_Int_t lizzieLet6_5QNode_Int_6QNone_Int_d;
  logic lizzieLet6_5QNode_Int_6QNone_Int_r;
  Pointer_QTree_Int_t _30_d;
  logic _30_r;
  assign _30_r = 1'd1;
  Pointer_QTree_Int_t _29_d;
  logic _29_r;
  assign _29_r = 1'd1;
  Pointer_QTree_Int_t _28_d;
  logic _28_r;
  assign _28_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet6_5QNode_Int_6QNone_Int_1_argbuf_d;
  logic lizzieLet6_5QNode_Int_6QNone_Int_1_argbuf_r;
  \Pointer_CTf''''''''''''_f''''''''''''_Int_t  lizzieLet6_5QNode_Int_7QNone_Int_d;
  logic lizzieLet6_5QNode_Int_7QNone_Int_r;
  \Pointer_CTf''''''''''''_f''''''''''''_Int_t  lizzieLet6_5QNode_Int_7QVal_Int_d;
  logic lizzieLet6_5QNode_Int_7QVal_Int_r;
  \Pointer_CTf''''''''''''_f''''''''''''_Int_t  lizzieLet6_5QNode_Int_7QNode_Int_d;
  logic lizzieLet6_5QNode_Int_7QNode_Int_r;
  \Pointer_CTf''''''''''''_f''''''''''''_Int_t  lizzieLet6_5QNode_Int_7QError_Int_d;
  logic lizzieLet6_5QNode_Int_7QError_Int_r;
  \Pointer_CTf''''''''''''_f''''''''''''_Int_t  lizzieLet6_5QNode_Int_7QError_Int_1_argbuf_d;
  logic lizzieLet6_5QNode_Int_7QError_Int_1_argbuf_r;
  \CTf''''''''''''_f''''''''''''_Int_t  \lizzieLet6_5QNode_Int_7QNode_Int_1lizzieLet6_5QNode_Int_8QNode_Int_1t1afy_1lizzieLet6_5QNode_Int_4QNode_Int_1lizzieLet6_5QNode_Int_5QNode_Int_1lizzieLet6_5QNode_Int_9QNode_Int_1t2afz_1lizzieLet6_5QNode_Int_10QNode_Int_1t3afA_1Lcall_f''''''''''''_f''''''''''''_Int3_d ;
  logic \lizzieLet6_5QNode_Int_7QNode_Int_1lizzieLet6_5QNode_Int_8QNode_Int_1t1afy_1lizzieLet6_5QNode_Int_4QNode_Int_1lizzieLet6_5QNode_Int_5QNode_Int_1lizzieLet6_5QNode_Int_9QNode_Int_1t2afz_1lizzieLet6_5QNode_Int_10QNode_Int_1t3afA_1Lcall_f''''''''''''_f''''''''''''_Int3_r ;
  \CTf''''''''''''_f''''''''''''_Int_t  lizzieLet14_1_argbuf_d;
  logic lizzieLet14_1_argbuf_r;
  \Pointer_CTf''''''''''''_f''''''''''''_Int_t  lizzieLet6_5QNode_Int_7QNone_Int_1_argbuf_d;
  logic lizzieLet6_5QNode_Int_7QNone_Int_1_argbuf_r;
  \Pointer_CTf''''''''''''_f''''''''''''_Int_t  lizzieLet6_5QNode_Int_7QVal_Int_1_argbuf_d;
  logic lizzieLet6_5QNode_Int_7QVal_Int_1_argbuf_r;
  Pointer_QTree_Int_t _27_d;
  logic _27_r;
  assign _27_r = 1'd1;
  Pointer_QTree_Int_t _26_d;
  logic _26_r;
  assign _26_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet6_5QNode_Int_8QNode_Int_d;
  logic lizzieLet6_5QNode_Int_8QNode_Int_r;
  Pointer_QTree_Int_t _25_d;
  logic _25_r;
  assign _25_r = 1'd1;
  Pointer_QTree_Int_t _24_d;
  logic _24_r;
  assign _24_r = 1'd1;
  Pointer_QTree_Int_t _23_d;
  logic _23_r;
  assign _23_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet6_5QNode_Int_9QNode_Int_d;
  logic lizzieLet6_5QNode_Int_9QNode_Int_r;
  Pointer_QTree_Int_t _22_d;
  logic _22_r;
  assign _22_r = 1'd1;
  QTree_Int_t lizzieLet6_5QVal_Int_1_d;
  logic lizzieLet6_5QVal_Int_1_r;
  QTree_Int_t lizzieLet6_5QVal_Int_2_d;
  logic lizzieLet6_5QVal_Int_2_r;
  QTree_Int_t lizzieLet6_5QVal_Int_3_d;
  logic lizzieLet6_5QVal_Int_3_r;
  QTree_Int_t lizzieLet6_5QVal_Int_4_d;
  logic lizzieLet6_5QVal_Int_4_r;
  QTree_Int_t lizzieLet6_5QVal_Int_5_d;
  logic lizzieLet6_5QVal_Int_5_r;
  QTree_Int_t lizzieLet6_5QVal_Int_6_d;
  logic lizzieLet6_5QVal_Int_6_r;
  QTree_Int_t lizzieLet6_5QVal_Int_7_d;
  logic lizzieLet6_5QVal_Int_7_r;
  QTree_Int_t lizzieLet6_5QVal_Int_8_d;
  logic lizzieLet6_5QVal_Int_8_r;
  Int_t vafo_destruct_d;
  logic vafo_destruct_r;
  QTree_Int_t _21_d;
  logic _21_r;
  assign _21_r = 1'd1;
  QTree_Int_t lizzieLet6_5QVal_Int_1QVal_Int_d;
  logic lizzieLet6_5QVal_Int_1QVal_Int_r;
  QTree_Int_t _20_d;
  logic _20_r;
  assign _20_r = 1'd1;
  QTree_Int_t _19_d;
  logic _19_r;
  assign _19_r = 1'd1;
  Go_t lizzieLet6_5QVal_Int_3QNone_Int_d;
  logic lizzieLet6_5QVal_Int_3QNone_Int_r;
  Go_t lizzieLet6_5QVal_Int_3QVal_Int_d;
  logic lizzieLet6_5QVal_Int_3QVal_Int_r;
  Go_t lizzieLet6_5QVal_Int_3QNode_Int_d;
  logic lizzieLet6_5QVal_Int_3QNode_Int_r;
  Go_t lizzieLet6_5QVal_Int_3QError_Int_d;
  logic lizzieLet6_5QVal_Int_3QError_Int_r;
  Go_t lizzieLet6_5QVal_Int_3QError_Int_1_d;
  logic lizzieLet6_5QVal_Int_3QError_Int_1_r;
  Go_t lizzieLet6_5QVal_Int_3QError_Int_2_d;
  logic lizzieLet6_5QVal_Int_3QError_Int_2_r;
  QTree_Int_t lizzieLet6_5QVal_Int_3QError_Int_1QError_Int_d;
  logic lizzieLet6_5QVal_Int_3QError_Int_1QError_Int_r;
  QTree_Int_t lizzieLet11_1_argbuf_d;
  logic lizzieLet11_1_argbuf_r;
  Go_t lizzieLet6_5QVal_Int_3QError_Int_2_argbuf_d;
  logic lizzieLet6_5QVal_Int_3QError_Int_2_argbuf_r;
  Go_t lizzieLet6_5QVal_Int_3QNode_Int_1_d;
  logic lizzieLet6_5QVal_Int_3QNode_Int_1_r;
  Go_t lizzieLet6_5QVal_Int_3QNode_Int_2_d;
  logic lizzieLet6_5QVal_Int_3QNode_Int_2_r;
  QTree_Int_t lizzieLet6_5QVal_Int_3QNode_Int_1QError_Int_d;
  logic lizzieLet6_5QVal_Int_3QNode_Int_1QError_Int_r;
  QTree_Int_t lizzieLet10_1_argbuf_d;
  logic lizzieLet10_1_argbuf_r;
  Go_t lizzieLet6_5QVal_Int_3QNode_Int_2_argbuf_d;
  logic lizzieLet6_5QVal_Int_3QNode_Int_2_argbuf_r;
  Go_t lizzieLet6_5QVal_Int_3QNone_Int_1_argbuf_d;
  logic lizzieLet6_5QVal_Int_3QNone_Int_1_argbuf_r;
  Go_t lizzieLet6_5QVal_Int_3QVal_Int_1_d;
  logic lizzieLet6_5QVal_Int_3QVal_Int_1_r;
  Go_t lizzieLet6_5QVal_Int_3QVal_Int_2_d;
  logic lizzieLet6_5QVal_Int_3QVal_Int_2_r;
  Go_t lizzieLet6_5QVal_Int_3QVal_Int_1_argbuf_d;
  logic lizzieLet6_5QVal_Int_3QVal_Int_1_argbuf_r;
  TupGo___MyDTInt_Bool___Int_t applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int2_d;
  logic applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int2_r;
  MyDTInt_Bool_t _18_d;
  logic _18_r;
  assign _18_r = 1'd1;
  MyDTInt_Bool_t lizzieLet6_5QVal_Int_4QVal_Int_d;
  logic lizzieLet6_5QVal_Int_4QVal_Int_r;
  MyDTInt_Bool_t _17_d;
  logic _17_r;
  assign _17_r = 1'd1;
  MyDTInt_Bool_t _16_d;
  logic _16_r;
  assign _16_r = 1'd1;
  MyDTInt_Bool_t lizzieLet6_5QVal_Int_4QVal_Int_1_argbuf_d;
  logic lizzieLet6_5QVal_Int_4QVal_Int_1_argbuf_r;
  MyDTInt_Int_Int_t _15_d;
  logic _15_r;
  assign _15_r = 1'd1;
  MyDTInt_Int_Int_t lizzieLet6_5QVal_Int_5QVal_Int_d;
  logic lizzieLet6_5QVal_Int_5QVal_Int_r;
  MyDTInt_Int_Int_t _14_d;
  logic _14_r;
  assign _14_r = 1'd1;
  MyDTInt_Int_Int_t _13_d;
  logic _13_r;
  assign _13_r = 1'd1;
  MyDTInt_Int_Int_t lizzieLet6_5QVal_Int_5QVal_Int_1_d;
  logic lizzieLet6_5QVal_Int_5QVal_Int_1_r;
  MyDTInt_Int_Int_t lizzieLet6_5QVal_Int_5QVal_Int_2_d;
  logic lizzieLet6_5QVal_Int_5QVal_Int_2_r;
  MyDTInt_Int_Int_t lizzieLet6_5QVal_Int_5QVal_Int_1_argbuf_d;
  logic lizzieLet6_5QVal_Int_5QVal_Int_1_argbuf_r;
  TupMyDTInt_Int_Int___Int___Int_t applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int3_d;
  logic applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int3_r;
  Pointer_QTree_Int_t lizzieLet6_5QVal_Int_6QNone_Int_d;
  logic lizzieLet6_5QVal_Int_6QNone_Int_r;
  Pointer_QTree_Int_t _12_d;
  logic _12_r;
  assign _12_r = 1'd1;
  Pointer_QTree_Int_t _11_d;
  logic _11_r;
  assign _11_r = 1'd1;
  Pointer_QTree_Int_t _10_d;
  logic _10_r;
  assign _10_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet6_5QVal_Int_6QNone_Int_1_argbuf_d;
  logic lizzieLet6_5QVal_Int_6QNone_Int_1_argbuf_r;
  \Pointer_CTf''''''''''''_f''''''''''''_Int_t  lizzieLet6_5QVal_Int_7QNone_Int_d;
  logic lizzieLet6_5QVal_Int_7QNone_Int_r;
  \Pointer_CTf''''''''''''_f''''''''''''_Int_t  lizzieLet6_5QVal_Int_7QVal_Int_d;
  logic lizzieLet6_5QVal_Int_7QVal_Int_r;
  \Pointer_CTf''''''''''''_f''''''''''''_Int_t  lizzieLet6_5QVal_Int_7QNode_Int_d;
  logic lizzieLet6_5QVal_Int_7QNode_Int_r;
  \Pointer_CTf''''''''''''_f''''''''''''_Int_t  lizzieLet6_5QVal_Int_7QError_Int_d;
  logic lizzieLet6_5QVal_Int_7QError_Int_r;
  \Pointer_CTf''''''''''''_f''''''''''''_Int_t  lizzieLet6_5QVal_Int_7QError_Int_1_argbuf_d;
  logic lizzieLet6_5QVal_Int_7QError_Int_1_argbuf_r;
  \Pointer_CTf''''''''''''_f''''''''''''_Int_t  lizzieLet6_5QVal_Int_7QNode_Int_1_argbuf_d;
  logic lizzieLet6_5QVal_Int_7QNode_Int_1_argbuf_r;
  \Pointer_CTf''''''''''''_f''''''''''''_Int_t  lizzieLet6_5QVal_Int_7QNone_Int_1_argbuf_d;
  logic lizzieLet6_5QVal_Int_7QNone_Int_1_argbuf_r;
  Int_t _9_d;
  logic _9_r;
  assign _9_r = 1'd1;
  Int_t lizzieLet6_5QVal_Int_8QVal_Int_d;
  logic lizzieLet6_5QVal_Int_8QVal_Int_r;
  Int_t _8_d;
  logic _8_r;
  assign _8_r = 1'd1;
  Int_t _7_d;
  logic _7_r;
  assign _7_r = 1'd1;
  Int_t lizzieLet6_5QVal_Int_8QVal_Int_1_d;
  logic lizzieLet6_5QVal_Int_8QVal_Int_1_r;
  Int_t lizzieLet6_5QVal_Int_8QVal_Int_2_d;
  logic lizzieLet6_5QVal_Int_8QVal_Int_2_r;
  Int_t lizzieLet6_5QVal_Int_8QVal_Int_1_argbuf_d;
  logic lizzieLet6_5QVal_Int_8QVal_Int_1_argbuf_r;
  MyDTInt_Int_Int_t _6_d;
  logic _6_r;
  assign _6_r = 1'd1;
  MyDTInt_Int_Int_t lizzieLet6_6QVal_Int_d;
  logic lizzieLet6_6QVal_Int_r;
  MyDTInt_Int_Int_t lizzieLet6_6QNode_Int_d;
  logic lizzieLet6_6QNode_Int_r;
  MyDTInt_Int_Int_t _5_d;
  logic _5_r;
  assign _5_r = 1'd1;
  Pointer_QTree_Int_t _4_d;
  logic _4_r;
  assign _4_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet6_7QVal_Int_d;
  logic lizzieLet6_7QVal_Int_r;
  Pointer_QTree_Int_t lizzieLet6_7QNode_Int_d;
  logic lizzieLet6_7QNode_Int_r;
  Pointer_QTree_Int_t _3_d;
  logic _3_r;
  assign _3_r = 1'd1;
  \Pointer_CTf''''''''''''_f''''''''''''_Int_t  lizzieLet6_8QNone_Int_d;
  logic lizzieLet6_8QNone_Int_r;
  \Pointer_CTf''''''''''''_f''''''''''''_Int_t  lizzieLet6_8QVal_Int_d;
  logic lizzieLet6_8QVal_Int_r;
  \Pointer_CTf''''''''''''_f''''''''''''_Int_t  lizzieLet6_8QNode_Int_d;
  logic lizzieLet6_8QNode_Int_r;
  \Pointer_CTf''''''''''''_f''''''''''''_Int_t  lizzieLet6_8QError_Int_d;
  logic lizzieLet6_8QError_Int_r;
  \Pointer_CTf''''''''''''_f''''''''''''_Int_t  lizzieLet6_8QError_Int_1_argbuf_d;
  logic lizzieLet6_8QError_Int_1_argbuf_r;
  \Pointer_CTf''''''''''''_f''''''''''''_Int_t  lizzieLet6_8QNone_Int_1_argbuf_d;
  logic lizzieLet6_8QNone_Int_1_argbuf_r;
  Pointer_QTree_Int_t lizzieLet6_9QNone_Int_d;
  logic lizzieLet6_9QNone_Int_r;
  Pointer_QTree_Int_t _2_d;
  logic _2_r;
  assign _2_r = 1'd1;
  Pointer_QTree_Int_t _1_d;
  logic _1_r;
  assign _1_r = 1'd1;
  Pointer_QTree_Int_t _0_d;
  logic _0_r;
  assign _0_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet6_9QNone_Int_1_argbuf_d;
  logic lizzieLet6_9QNone_Int_1_argbuf_r;
  Pointer_QTree_Int_t m1aeq_1_argbuf_d;
  logic m1aeq_1_argbuf_r;
  Pointer_QTree_Int_t m1aeq_1_d;
  logic m1aeq_1_r;
  Pointer_QTree_Int_t m1aeq_2_d;
  logic m1aeq_2_r;
  Pointer_QTree_Int_t m2aer_1_argbuf_d;
  logic m2aer_1_argbuf_r;
  Pointer_QTree_Int_t m2aer_1_d;
  logic m2aer_1_r;
  Pointer_QTree_Int_t m2aer_2_d;
  logic m2aer_2_r;
  Pointer_QTree_Int_t m3aes_1_argbuf_d;
  logic m3aes_1_argbuf_r;
  Pointer_QTree_Int_t m3aes_1_d;
  logic m3aes_1_r;
  Pointer_QTree_Int_t m3aes_2_d;
  logic m3aes_2_r;
  MyDTInt_Int_Int_t op_addaeu_2_2_argbuf_d;
  logic op_addaeu_2_2_argbuf_r;
  MyDTInt_Int_Int_t op_addaeu_2_1_d;
  logic op_addaeu_2_1_r;
  MyDTInt_Int_Int_t op_addaeu_2_2_d;
  logic op_addaeu_2_2_r;
  MyDTInt_Int_Int_t op_addaeu_3_2_argbuf_d;
  logic op_addaeu_3_2_argbuf_r;
  MyDTInt_Int_Int_t op_addaeu_3_1_d;
  logic op_addaeu_3_1_r;
  MyDTInt_Int_Int_t op_addaeu_3_2_d;
  logic op_addaeu_3_2_r;
  MyDTInt_Int_Int_t op_addaeu_4_1_argbuf_d;
  logic op_addaeu_4_1_argbuf_r;
  MyDTInt_Int_Int_t op_addafm_2_2_argbuf_d;
  logic op_addafm_2_2_argbuf_r;
  MyDTInt_Int_Int_t op_addafm_2_1_d;
  logic op_addafm_2_1_r;
  MyDTInt_Int_Int_t op_addafm_2_2_d;
  logic op_addafm_2_2_r;
  MyDTInt_Int_Int_t op_addafm_3_2_argbuf_d;
  logic op_addafm_3_2_argbuf_r;
  MyDTInt_Int_Int_t op_addafm_3_1_d;
  logic op_addafm_3_1_r;
  MyDTInt_Int_Int_t op_addafm_3_2_d;
  logic op_addafm_3_2_r;
  MyDTInt_Int_Int_t op_addafm_4_1_argbuf_d;
  logic op_addafm_4_1_argbuf_r;
  Pointer_QTree_Int_t q1a8r_1_argbuf_d;
  logic q1a8r_1_argbuf_r;
  Pointer_QTree_Int_t q1af0_3_1_argbuf_d;
  logic q1af0_3_1_argbuf_r;
  Pointer_QTree_Int_t q1aft_3_1_argbuf_d;
  logic q1aft_3_1_argbuf_r;
  Pointer_QTree_Int_t q2a8s_1_1_argbuf_d;
  logic q2a8s_1_1_argbuf_r;
  Pointer_QTree_Int_t q2af1_2_1_argbuf_d;
  logic q2af1_2_1_argbuf_r;
  Pointer_QTree_Int_t q2afu_2_1_argbuf_d;
  logic q2afu_2_1_argbuf_r;
  Pointer_QTree_Int_t q3a8t_2_1_argbuf_d;
  logic q3a8t_2_1_argbuf_r;
  Pointer_QTree_Int_t q3af2_1_1_argbuf_d;
  logic q3af2_1_1_argbuf_r;
  Pointer_QTree_Int_t q3afv_1_1_argbuf_d;
  logic q3afv_1_1_argbuf_r;
  Pointer_QTree_Int_t q4a8u_3_1_argbuf_d;
  logic q4a8u_3_1_argbuf_r;
  Pointer_QTree_Int_t q4afj_1_argbuf_d;
  logic q4afj_1_argbuf_r;
  Pointer_QTree_Int_t q4afj_1_d;
  logic q4afj_1_r;
  Pointer_QTree_Int_t q4afj_2_d;
  logic q4afj_2_r;
  CT$wnnz_t readPointer_CT$wnnzscfarg_0_1_argbuf_rwb_d;
  logic readPointer_CT$wnnzscfarg_0_1_argbuf_rwb_r;
  CT$wnnz_t lizzieLet58_1_d;
  logic lizzieLet58_1_r;
  CT$wnnz_t lizzieLet58_2_d;
  logic lizzieLet58_2_r;
  CT$wnnz_t lizzieLet58_3_d;
  logic lizzieLet58_3_r;
  CT$wnnz_t lizzieLet58_4_d;
  logic lizzieLet58_4_r;
  \CTf''''''''''''_f''''''''''''_Int_t  \readPointer_CTf''''''''''''_f''''''''''''_Intscfarg_0_1_1_argbuf_rwb_d ;
  logic \readPointer_CTf''''''''''''_f''''''''''''_Intscfarg_0_1_1_argbuf_rwb_r ;
  \CTf''''''''''''_f''''''''''''_Int_t  lizzieLet62_1_d;
  logic lizzieLet62_1_r;
  \CTf''''''''''''_f''''''''''''_Int_t  lizzieLet62_2_d;
  logic lizzieLet62_2_r;
  \CTf''''''''''''_f''''''''''''_Int_t  lizzieLet62_3_d;
  logic lizzieLet62_3_r;
  \CTf''''''''''''_f''''''''''''_Int_t  lizzieLet62_4_d;
  logic lizzieLet62_4_r;
  CTf_f_Int_t readPointer_CTf_f_Intscfarg_0_2_1_argbuf_rwb_d;
  logic readPointer_CTf_f_Intscfarg_0_2_1_argbuf_rwb_r;
  CTf_f_Int_t lizzieLet67_1_d;
  logic lizzieLet67_1_r;
  CTf_f_Int_t lizzieLet67_2_d;
  logic lizzieLet67_2_r;
  CTf_f_Int_t lizzieLet67_3_d;
  logic lizzieLet67_3_r;
  CTf_f_Int_t lizzieLet67_4_d;
  logic lizzieLet67_4_r;
  QTree_Int_t readPointer_QTree_Intm1aeq_1_argbuf_rwb_d;
  logic readPointer_QTree_Intm1aeq_1_argbuf_rwb_r;
  QTree_Int_t lizzieLet17_1_d;
  logic lizzieLet17_1_r;
  QTree_Int_t lizzieLet17_2_d;
  logic lizzieLet17_2_r;
  QTree_Int_t lizzieLet17_3_d;
  logic lizzieLet17_3_r;
  QTree_Int_t lizzieLet17_4_d;
  logic lizzieLet17_4_r;
  QTree_Int_t lizzieLet17_5_d;
  logic lizzieLet17_5_r;
  QTree_Int_t lizzieLet17_6_d;
  logic lizzieLet17_6_r;
  QTree_Int_t lizzieLet17_7_d;
  logic lizzieLet17_7_r;
  QTree_Int_t lizzieLet17_8_d;
  logic lizzieLet17_8_r;
  QTree_Int_t lizzieLet17_9_d;
  logic lizzieLet17_9_r;
  QTree_Int_t lizzieLet17_10_d;
  logic lizzieLet17_10_r;
  QTree_Int_t lizzieLet17_11_d;
  logic lizzieLet17_11_r;
  QTree_Int_t readPointer_QTree_Intm2aer_1_argbuf_rwb_d;
  logic readPointer_QTree_Intm2aer_1_argbuf_rwb_r;
  QTree_Int_t readPointer_QTree_Intm3aes_1_argbuf_rwb_d;
  logic readPointer_QTree_Intm3aes_1_argbuf_rwb_r;
  QTree_Int_t readPointer_QTree_Intq4afj_1_argbuf_rwb_d;
  logic readPointer_QTree_Intq4afj_1_argbuf_rwb_r;
  QTree_Int_t lizzieLet6_1_d;
  logic lizzieLet6_1_r;
  QTree_Int_t lizzieLet6_2_d;
  logic lizzieLet6_2_r;
  QTree_Int_t lizzieLet6_3_d;
  logic lizzieLet6_3_r;
  QTree_Int_t lizzieLet6_4_d;
  logic lizzieLet6_4_r;
  QTree_Int_t lizzieLet6_5_d;
  logic lizzieLet6_5_r;
  QTree_Int_t lizzieLet6_6_d;
  logic lizzieLet6_6_r;
  QTree_Int_t lizzieLet6_7_d;
  logic lizzieLet6_7_r;
  QTree_Int_t lizzieLet6_8_d;
  logic lizzieLet6_8_r;
  QTree_Int_t lizzieLet6_9_d;
  logic lizzieLet6_9_r;
  QTree_Int_t readPointer_QTree_Intt4afk_1_argbuf_rwb_d;
  logic readPointer_QTree_Intt4afk_1_argbuf_rwb_r;
  QTree_Int_t readPointer_QTree_Intwsmk_1_1_argbuf_rwb_d;
  logic readPointer_QTree_Intwsmk_1_1_argbuf_rwb_r;
  QTree_Int_t lizzieLet4_1_d;
  logic lizzieLet4_1_r;
  QTree_Int_t lizzieLet4_2_d;
  logic lizzieLet4_2_r;
  QTree_Int_t lizzieLet4_3_d;
  logic lizzieLet4_3_r;
  QTree_Int_t lizzieLet4_4_d;
  logic lizzieLet4_4_r;
  \Pointer_CTf''''''''''''_f''''''''''''_Int_t  sc_0_10_1_argbuf_d;
  logic sc_0_10_1_argbuf_r;
  Pointer_CTf_f_Int_t sc_0_14_1_argbuf_d;
  logic sc_0_14_1_argbuf_r;
  Pointer_CT$wnnz_t sc_0_6_1_argbuf_d;
  logic sc_0_6_1_argbuf_r;
  \Pointer_CTf''''''''''''_f''''''''''''_Int_t  scfarg_0_1_1_argbuf_d;
  logic scfarg_0_1_1_argbuf_r;
  Pointer_CTf_f_Int_t scfarg_0_2_1_argbuf_d;
  logic scfarg_0_2_1_argbuf_r;
  Pointer_CT$wnnz_t scfarg_0_1_argbuf_d;
  logic scfarg_0_1_argbuf_r;
  Pointer_QTree_Int_t \t1'aff_3_1_argbuf_d ;
  logic \t1'aff_3_1_argbuf_r ;
  Pointer_QTree_Int_t t1aeG_1_argbuf_d;
  logic t1aeG_1_argbuf_r;
  Pointer_QTree_Int_t t1af5_1_argbuf_d;
  logic t1af5_1_argbuf_r;
  Pointer_QTree_Int_t t1afa_3_1_argbuf_d;
  logic t1afa_3_1_argbuf_r;
  Pointer_QTree_Int_t t1afy_3_1_argbuf_d;
  logic t1afy_3_1_argbuf_r;
  Pointer_QTree_Int_t \t2'afg_2_1_argbuf_d ;
  logic \t2'afg_2_1_argbuf_r ;
  Pointer_QTree_Int_t t2aeH_1_argbuf_d;
  logic t2aeH_1_argbuf_r;
  Pointer_QTree_Int_t t2af6_1_argbuf_d;
  logic t2af6_1_argbuf_r;
  Pointer_QTree_Int_t t2afb_2_1_argbuf_d;
  logic t2afb_2_1_argbuf_r;
  Pointer_QTree_Int_t t2afz_2_1_argbuf_d;
  logic t2afz_2_1_argbuf_r;
  Pointer_QTree_Int_t \t3'afh_1_1_argbuf_d ;
  logic \t3'afh_1_1_argbuf_r ;
  Pointer_QTree_Int_t t3aeI_1_argbuf_d;
  logic t3aeI_1_argbuf_r;
  Pointer_QTree_Int_t t3af7_1_argbuf_d;
  logic t3af7_1_argbuf_r;
  Pointer_QTree_Int_t t3afA_1_1_argbuf_d;
  logic t3afA_1_1_argbuf_r;
  Pointer_QTree_Int_t t3afc_1_1_argbuf_d;
  logic t3afc_1_1_argbuf_r;
  Pointer_QTree_Int_t \t4'afi_1_argbuf_d ;
  logic \t4'afi_1_argbuf_r ;
  Pointer_QTree_Int_t t4aeJ_1_argbuf_d;
  logic t4aeJ_1_argbuf_r;
  Pointer_QTree_Int_t t4af8_1_argbuf_d;
  logic t4af8_1_argbuf_r;
  Pointer_QTree_Int_t t4afk_1_argbuf_d;
  logic t4afk_1_argbuf_r;
  Pointer_QTree_Int_t t4afk_1_d;
  logic t4afk_1_r;
  Pointer_QTree_Int_t t4afk_2_d;
  logic t4afk_2_r;
  Pointer_QTree_Int_t t5afB_1_argbuf_d;
  logic t5afB_1_argbuf_r;
  Int_t \v'aeR_1_argbuf_d ;
  logic \v'aeR_1_argbuf_r ;
  Int_t \v'aeR_1_d ;
  logic \v'aeR_1_r ;
  Int_t \v'aeR_2_d ;
  logic \v'aeR_2_r ;
  Int_t vaeL_1_argbuf_d;
  logic vaeL_1_argbuf_r;
  Int_t vaeL_1_d;
  logic vaeL_1_r;
  Int_t vaeL_2_d;
  logic vaeL_2_r;
  Int_t vaeQ_1_argbuf_d;
  logic vaeQ_1_argbuf_r;
  Int_t vaeQ_1_d;
  logic vaeQ_1_r;
  Int_t vaeQ_2_d;
  logic vaeQ_2_r;
  Int_t vaew_1_argbuf_d;
  logic vaew_1_argbuf_r;
  Int_t vaew_1_d;
  logic vaew_1_r;
  Int_t vaew_2_d;
  logic vaew_2_r;
  Int_t vafo_1_argbuf_d;
  logic vafo_1_argbuf_r;
  Int_t vafo_1_d;
  logic vafo_1_r;
  Int_t vafo_2_d;
  logic vafo_2_r;
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet0_1_argbuf_rwb_d;
  logic writeCT$wnnzlizzieLet0_1_argbuf_rwb_r;
  Pointer_CT$wnnz_t lizzieLet39_1_argbuf_d;
  logic lizzieLet39_1_argbuf_r;
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet59_1_argbuf_rwb_d;
  logic writeCT$wnnzlizzieLet59_1_argbuf_rwb_r;
  Pointer_CT$wnnz_t sca2_1_argbuf_d;
  logic sca2_1_argbuf_r;
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet5_1_argbuf_rwb_d;
  logic writeCT$wnnzlizzieLet5_1_argbuf_rwb_r;
  Pointer_CT$wnnz_t sca3_1_argbuf_d;
  logic sca3_1_argbuf_r;
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet60_1_argbuf_rwb_d;
  logic writeCT$wnnzlizzieLet60_1_argbuf_rwb_r;
  Pointer_CT$wnnz_t sca1_1_argbuf_d;
  logic sca1_1_argbuf_r;
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet61_1_argbuf_rwb_d;
  logic writeCT$wnnzlizzieLet61_1_argbuf_rwb_r;
  Pointer_CT$wnnz_t sca0_1_argbuf_d;
  logic sca0_1_argbuf_r;
  \Pointer_CTf''''''''''''_f''''''''''''_Int_t  \writeCTf''''''''''''_f''''''''''''_IntlizzieLet14_1_argbuf_rwb_d ;
  logic \writeCTf''''''''''''_f''''''''''''_IntlizzieLet14_1_argbuf_rwb_r ;
  \Pointer_CTf''''''''''''_f''''''''''''_Int_t  sca3_1_1_argbuf_d;
  logic sca3_1_1_argbuf_r;
  \Pointer_CTf''''''''''''_f''''''''''''_Int_t  \writeCTf''''''''''''_f''''''''''''_IntlizzieLet56_1_argbuf_rwb_d ;
  logic \writeCTf''''''''''''_f''''''''''''_IntlizzieLet56_1_argbuf_rwb_r ;
  \Pointer_CTf''''''''''''_f''''''''''''_Int_t  lizzieLet7_1_1_argbuf_d;
  logic lizzieLet7_1_1_argbuf_r;
  \Pointer_CTf''''''''''''_f''''''''''''_Int_t  \writeCTf''''''''''''_f''''''''''''_IntlizzieLet63_1_argbuf_rwb_d ;
  logic \writeCTf''''''''''''_f''''''''''''_IntlizzieLet63_1_argbuf_rwb_r ;
  \Pointer_CTf''''''''''''_f''''''''''''_Int_t  sca2_1_1_argbuf_d;
  logic sca2_1_1_argbuf_r;
  \Pointer_CTf''''''''''''_f''''''''''''_Int_t  \writeCTf''''''''''''_f''''''''''''_IntlizzieLet64_1_argbuf_rwb_d ;
  logic \writeCTf''''''''''''_f''''''''''''_IntlizzieLet64_1_argbuf_rwb_r ;
  \Pointer_CTf''''''''''''_f''''''''''''_Int_t  sca1_1_1_argbuf_d;
  logic sca1_1_1_argbuf_r;
  \Pointer_CTf''''''''''''_f''''''''''''_Int_t  \writeCTf''''''''''''_f''''''''''''_IntlizzieLet65_1_argbuf_rwb_d ;
  logic \writeCTf''''''''''''_f''''''''''''_IntlizzieLet65_1_argbuf_rwb_r ;
  \Pointer_CTf''''''''''''_f''''''''''''_Int_t  sca0_1_1_argbuf_d;
  logic sca0_1_1_argbuf_r;
  Pointer_CTf_f_Int_t writeCTf_f_IntlizzieLet52_1_argbuf_rwb_d;
  logic writeCTf_f_IntlizzieLet52_1_argbuf_rwb_r;
  Pointer_CTf_f_Int_t sca3_2_1_argbuf_d;
  logic sca3_2_1_argbuf_r;
  Pointer_CTf_f_Int_t writeCTf_f_IntlizzieLet57_1_argbuf_rwb_d;
  logic writeCTf_f_IntlizzieLet57_1_argbuf_rwb_r;
  Pointer_CTf_f_Int_t lizzieLet36_1_1_argbuf_d;
  logic lizzieLet36_1_1_argbuf_r;
  Pointer_CTf_f_Int_t writeCTf_f_IntlizzieLet68_1_argbuf_rwb_d;
  logic writeCTf_f_IntlizzieLet68_1_argbuf_rwb_r;
  Pointer_CTf_f_Int_t sca2_2_1_argbuf_d;
  logic sca2_2_1_argbuf_r;
  Pointer_CTf_f_Int_t writeCTf_f_IntlizzieLet69_1_argbuf_rwb_d;
  logic writeCTf_f_IntlizzieLet69_1_argbuf_rwb_r;
  Pointer_CTf_f_Int_t sca1_2_1_argbuf_d;
  logic sca1_2_1_argbuf_r;
  Pointer_CTf_f_Int_t writeCTf_f_IntlizzieLet70_1_argbuf_rwb_d;
  logic writeCTf_f_IntlizzieLet70_1_argbuf_rwb_r;
  Pointer_CTf_f_Int_t sca0_2_1_argbuf_d;
  logic sca0_2_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet10_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet10_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet2_1_1_argbuf_d;
  logic lizzieLet2_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet11_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet11_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet3_1_1_argbuf_d;
  logic lizzieLet3_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet13_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet13_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet4_1_1_argbuf_d;
  logic lizzieLet4_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet15_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet15_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet5_1_1_argbuf_d;
  logic lizzieLet5_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet16_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet16_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet6_1_1_argbuf_d;
  logic lizzieLet6_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet20_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet20_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet8_1_1_argbuf_d;
  logic lizzieLet8_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet21_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet21_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet9_1_1_argbuf_d;
  logic lizzieLet9_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet22_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet22_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet10_1_1_argbuf_d;
  logic lizzieLet10_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet23_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet23_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet11_1_1_argbuf_d;
  logic lizzieLet11_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet25_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet25_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet12_1_argbuf_d;
  logic lizzieLet12_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet26_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet26_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet13_1_1_argbuf_d;
  logic lizzieLet13_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet27_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet27_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet14_1_1_argbuf_d;
  logic lizzieLet14_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet28_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet28_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet15_1_1_argbuf_d;
  logic lizzieLet15_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet31_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet31_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet16_1_1_argbuf_d;
  logic lizzieLet16_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet32_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet32_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet17_1_1_argbuf_d;
  logic lizzieLet17_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet33_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet33_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet18_1_1_argbuf_d;
  logic lizzieLet18_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet34_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet34_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet19_1_1_argbuf_d;
  logic lizzieLet19_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet36_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet36_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet20_1_1_argbuf_d;
  logic lizzieLet20_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet37_2_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet37_2_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet21_1_1_argbuf_d;
  logic lizzieLet21_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet38_1_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet38_1_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet22_1_1_argbuf_d;
  logic lizzieLet22_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet39_1_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet39_1_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet23_1_1_argbuf_d;
  logic lizzieLet23_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet40_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet40_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet24_1_argbuf_d;
  logic lizzieLet24_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet41_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet41_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet25_1_1_argbuf_d;
  logic lizzieLet25_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet42_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet42_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet26_1_1_argbuf_d;
  logic lizzieLet26_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet45_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet45_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet27_1_1_argbuf_d;
  logic lizzieLet27_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet46_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet46_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet28_1_1_argbuf_d;
  logic lizzieLet28_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet47_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet47_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet29_1_argbuf_d;
  logic lizzieLet29_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet48_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet48_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet30_1_argbuf_d;
  logic lizzieLet30_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet50_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet50_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet31_1_1_argbuf_d;
  logic lizzieLet31_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet51_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet51_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet32_1_1_argbuf_d;
  logic lizzieLet32_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet53_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet53_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet33_1_1_argbuf_d;
  logic lizzieLet33_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet54_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet54_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet34_1_1_argbuf_d;
  logic lizzieLet34_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet55_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet55_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet35_1_argbuf_d;
  logic lizzieLet35_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet66_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet66_1_argbuf_rwb_r;
  Pointer_QTree_Int_t contRet_0_1_1_argbuf_d;
  logic contRet_0_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet71_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet71_1_argbuf_rwb_r;
  Pointer_QTree_Int_t contRet_0_2_1_argbuf_d;
  logic contRet_0_2_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet8_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet8_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet0_1_1_argbuf_d;
  logic lizzieLet0_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet9_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet9_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet1_1_1_argbuf_d;
  logic lizzieLet1_1_1_argbuf_r;
  Pointer_QTree_Int_t wsmk_1_1_argbuf_d;
  logic wsmk_1_1_argbuf_r;
  CT$wnnz_t lizzieLet60_1_argbuf_d;
  logic lizzieLet60_1_argbuf_r;
  CT$wnnz_t wwsmn_2_1lizzieLet58_4Lcall_$wnnz2_1sc_0_4_1q4a8u_2_1Lcall_$wnnz1_d;
  logic wwsmn_2_1lizzieLet58_4Lcall_$wnnz2_1sc_0_4_1q4a8u_2_1Lcall_$wnnz1_r;
  CT$wnnz_t lizzieLet61_1_argbuf_d;
  logic lizzieLet61_1_argbuf_r;
  CT$wnnz_t wwsmn_3_1ww1XmW_1_1lizzieLet58_4Lcall_$wnnz1_1sc_0_5_1Lcall_$wnnz0_d;
  logic wwsmn_3_1ww1XmW_1_1lizzieLet58_4Lcall_$wnnz1_1sc_0_5_1Lcall_$wnnz0_r;
  \Int#_t  es_6_2_1ww2XmZ_1_1_Add32_d;
  logic es_6_2_1ww2XmZ_1_1_Add32_r;
  \Int#_t  wwsmn_4_1ww1XmW_2_1_Add32_d;
  logic wwsmn_4_1ww1XmW_2_1_Add32_r;
  
  /* fork (Ty Go) : (sourceGo,Go) > [(go_1,Go),
                                (go_2,Go),
                                (go_3,Go),
                                (go_4,Go),
                                (go__5,Go),
                                (go__6,Go),
                                (go__7,Go),
                                (go__8,Go),
                                (go__9,Go),
                                (go__10,Go)] */
  logic [9:0] sourceGo_emitted;
  logic [9:0] sourceGo_done;
  assign go_1_d = (sourceGo_d[0] && (! sourceGo_emitted[0]));
  assign go_2_d = (sourceGo_d[0] && (! sourceGo_emitted[1]));
  assign go_3_d = (sourceGo_d[0] && (! sourceGo_emitted[2]));
  assign go_4_d = (sourceGo_d[0] && (! sourceGo_emitted[3]));
  assign go__5_d = (sourceGo_d[0] && (! sourceGo_emitted[4]));
  assign go__6_d = (sourceGo_d[0] && (! sourceGo_emitted[5]));
  assign go__7_d = (sourceGo_d[0] && (! sourceGo_emitted[6]));
  assign go__8_d = (sourceGo_d[0] && (! sourceGo_emitted[7]));
  assign go__9_d = (sourceGo_d[0] && (! sourceGo_emitted[8]));
  assign go__10_d = (sourceGo_d[0] && (! sourceGo_emitted[9]));
  assign sourceGo_done = (sourceGo_emitted | ({go__10_d[0],
                                               go__9_d[0],
                                               go__8_d[0],
                                               go__7_d[0],
                                               go__6_d[0],
                                               go__5_d[0],
                                               go_4_d[0],
                                               go_3_d[0],
                                               go_2_d[0],
                                               go_1_d[0]} & {go__10_r,
                                                             go__9_r,
                                                             go__8_r,
                                                             go__7_r,
                                                             go__6_r,
                                                             go__5_r,
                                                             go_4_r,
                                                             go_3_r,
                                                             go_2_r,
                                                             go_1_r}));
  assign sourceGo_r = (& sourceGo_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) sourceGo_emitted <= 10'd0;
    else
      sourceGo_emitted <= (sourceGo_r ? 10'd0 :
                           sourceGo_done);
  
  /* const (Ty Word16#,Lit 0) : (go__5,Go) > (initHP_CT$wnnz,Word16#) */
  assign initHP_CT$wnnz_d = {16'd0, go__5_d[0]};
  assign go__5_r = initHP_CT$wnnz_r;
  
  /* const (Ty Word16#,
       Lit 1) : (incrHP_CT$wnnz1,Go) > (incrHP_CT$wnnz,Word16#) */
  assign incrHP_CT$wnnz_d = {16'd1, incrHP_CT$wnnz1_d[0]};
  assign incrHP_CT$wnnz1_r = incrHP_CT$wnnz_r;
  
  /* merge (Ty Go) : [(go__6,Go),
                 (incrHP_CT$wnnz2,Go)] > (incrHP_mergeCT$wnnz,Go) */
  logic [1:0] incrHP_mergeCT$wnnz_selected;
  logic [1:0] incrHP_mergeCT$wnnz_select;
  always_comb
    begin
      incrHP_mergeCT$wnnz_selected = 2'd0;
      if ((| incrHP_mergeCT$wnnz_select))
        incrHP_mergeCT$wnnz_selected = incrHP_mergeCT$wnnz_select;
      else
        if (go__6_d[0]) incrHP_mergeCT$wnnz_selected[0] = 1'd1;
        else if (incrHP_CT$wnnz2_d[0])
          incrHP_mergeCT$wnnz_selected[1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeCT$wnnz_select <= 2'd0;
    else
      incrHP_mergeCT$wnnz_select <= (incrHP_mergeCT$wnnz_r ? 2'd0 :
                                     incrHP_mergeCT$wnnz_selected);
  always_comb
    if (incrHP_mergeCT$wnnz_selected[0])
      incrHP_mergeCT$wnnz_d = go__6_d;
    else if (incrHP_mergeCT$wnnz_selected[1])
      incrHP_mergeCT$wnnz_d = incrHP_CT$wnnz2_d;
    else incrHP_mergeCT$wnnz_d = 1'd0;
  assign {incrHP_CT$wnnz2_r,
          go__6_r} = (incrHP_mergeCT$wnnz_r ? incrHP_mergeCT$wnnz_selected :
                      2'd0);
  
  /* fork (Ty Go) : (incrHP_mergeCT$wnnz_buf,Go) > [(incrHP_CT$wnnz1,Go),
                                               (incrHP_CT$wnnz2,Go)] */
  logic [1:0] incrHP_mergeCT$wnnz_buf_emitted;
  logic [1:0] incrHP_mergeCT$wnnz_buf_done;
  assign incrHP_CT$wnnz1_d = (incrHP_mergeCT$wnnz_buf_d[0] && (! incrHP_mergeCT$wnnz_buf_emitted[0]));
  assign incrHP_CT$wnnz2_d = (incrHP_mergeCT$wnnz_buf_d[0] && (! incrHP_mergeCT$wnnz_buf_emitted[1]));
  assign incrHP_mergeCT$wnnz_buf_done = (incrHP_mergeCT$wnnz_buf_emitted | ({incrHP_CT$wnnz2_d[0],
                                                                             incrHP_CT$wnnz1_d[0]} & {incrHP_CT$wnnz2_r,
                                                                                                      incrHP_CT$wnnz1_r}));
  assign incrHP_mergeCT$wnnz_buf_r = (& incrHP_mergeCT$wnnz_buf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeCT$wnnz_buf_emitted <= 2'd0;
    else
      incrHP_mergeCT$wnnz_buf_emitted <= (incrHP_mergeCT$wnnz_buf_r ? 2'd0 :
                                          incrHP_mergeCT$wnnz_buf_done);
  
  /* op_add (Ty Word16#) : (incrHP_CT$wnnz,Word16#) (forkHP1_CT$wnnz,Word16#) > (addHP_CT$wnnz,Word16#) */
  assign addHP_CT$wnnz_d = {(incrHP_CT$wnnz_d[16:1] + forkHP1_CT$wnnz_d[16:1]),
                            (incrHP_CT$wnnz_d[0] && forkHP1_CT$wnnz_d[0])};
  assign {incrHP_CT$wnnz_r,
          forkHP1_CT$wnnz_r} = {2 {(addHP_CT$wnnz_r && addHP_CT$wnnz_d[0])}};
  
  /* merge (Ty Word16#) : [(initHP_CT$wnnz,Word16#),
                      (addHP_CT$wnnz,Word16#)] > (mergeHP_CT$wnnz,Word16#) */
  logic [1:0] mergeHP_CT$wnnz_selected;
  logic [1:0] mergeHP_CT$wnnz_select;
  always_comb
    begin
      mergeHP_CT$wnnz_selected = 2'd0;
      if ((| mergeHP_CT$wnnz_select))
        mergeHP_CT$wnnz_selected = mergeHP_CT$wnnz_select;
      else
        if (initHP_CT$wnnz_d[0]) mergeHP_CT$wnnz_selected[0] = 1'd1;
        else if (addHP_CT$wnnz_d[0]) mergeHP_CT$wnnz_selected[1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_CT$wnnz_select <= 2'd0;
    else
      mergeHP_CT$wnnz_select <= (mergeHP_CT$wnnz_r ? 2'd0 :
                                 mergeHP_CT$wnnz_selected);
  always_comb
    if (mergeHP_CT$wnnz_selected[0])
      mergeHP_CT$wnnz_d = initHP_CT$wnnz_d;
    else if (mergeHP_CT$wnnz_selected[1])
      mergeHP_CT$wnnz_d = addHP_CT$wnnz_d;
    else mergeHP_CT$wnnz_d = {16'd0, 1'd0};
  assign {addHP_CT$wnnz_r,
          initHP_CT$wnnz_r} = (mergeHP_CT$wnnz_r ? mergeHP_CT$wnnz_selected :
                               2'd0);
  
  /* buf (Ty Go) : (incrHP_mergeCT$wnnz,Go) > (incrHP_mergeCT$wnnz_buf,Go) */
  Go_t incrHP_mergeCT$wnnz_bufchan_d;
  logic incrHP_mergeCT$wnnz_bufchan_r;
  assign incrHP_mergeCT$wnnz_r = ((! incrHP_mergeCT$wnnz_bufchan_d[0]) || incrHP_mergeCT$wnnz_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeCT$wnnz_bufchan_d <= 1'd0;
    else
      if (incrHP_mergeCT$wnnz_r)
        incrHP_mergeCT$wnnz_bufchan_d <= incrHP_mergeCT$wnnz_d;
  Go_t incrHP_mergeCT$wnnz_bufchan_buf;
  assign incrHP_mergeCT$wnnz_bufchan_r = (! incrHP_mergeCT$wnnz_bufchan_buf[0]);
  assign incrHP_mergeCT$wnnz_buf_d = (incrHP_mergeCT$wnnz_bufchan_buf[0] ? incrHP_mergeCT$wnnz_bufchan_buf :
                                      incrHP_mergeCT$wnnz_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeCT$wnnz_bufchan_buf <= 1'd0;
    else
      if ((incrHP_mergeCT$wnnz_buf_r && incrHP_mergeCT$wnnz_bufchan_buf[0]))
        incrHP_mergeCT$wnnz_bufchan_buf <= 1'd0;
      else if (((! incrHP_mergeCT$wnnz_buf_r) && (! incrHP_mergeCT$wnnz_bufchan_buf[0])))
        incrHP_mergeCT$wnnz_bufchan_buf <= incrHP_mergeCT$wnnz_bufchan_d;
  
  /* buf (Ty Word16#) : (mergeHP_CT$wnnz,Word16#) > (mergeHP_CT$wnnz_buf,Word16#) */
  \Word16#_t  mergeHP_CT$wnnz_bufchan_d;
  logic mergeHP_CT$wnnz_bufchan_r;
  assign mergeHP_CT$wnnz_r = ((! mergeHP_CT$wnnz_bufchan_d[0]) || mergeHP_CT$wnnz_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_CT$wnnz_bufchan_d <= {16'd0, 1'd0};
    else
      if (mergeHP_CT$wnnz_r)
        mergeHP_CT$wnnz_bufchan_d <= mergeHP_CT$wnnz_d;
  \Word16#_t  mergeHP_CT$wnnz_bufchan_buf;
  assign mergeHP_CT$wnnz_bufchan_r = (! mergeHP_CT$wnnz_bufchan_buf[0]);
  assign mergeHP_CT$wnnz_buf_d = (mergeHP_CT$wnnz_bufchan_buf[0] ? mergeHP_CT$wnnz_bufchan_buf :
                                  mergeHP_CT$wnnz_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_CT$wnnz_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((mergeHP_CT$wnnz_buf_r && mergeHP_CT$wnnz_bufchan_buf[0]))
        mergeHP_CT$wnnz_bufchan_buf <= {16'd0, 1'd0};
      else if (((! mergeHP_CT$wnnz_buf_r) && (! mergeHP_CT$wnnz_bufchan_buf[0])))
        mergeHP_CT$wnnz_bufchan_buf <= mergeHP_CT$wnnz_bufchan_d;
  
  /* fork (Ty Word16#) : (mergeHP_CT$wnnz_buf,Word16#) > [(forkHP1_CT$wnnz,Word16#),
                                                     (forkHP1_CT$wnn2,Word16#),
                                                     (forkHP1_CT$wnn3,Word16#)] */
  logic [2:0] mergeHP_CT$wnnz_buf_emitted;
  logic [2:0] mergeHP_CT$wnnz_buf_done;
  assign forkHP1_CT$wnnz_d = {mergeHP_CT$wnnz_buf_d[16:1],
                              (mergeHP_CT$wnnz_buf_d[0] && (! mergeHP_CT$wnnz_buf_emitted[0]))};
  assign forkHP1_CT$wnn2_d = {mergeHP_CT$wnnz_buf_d[16:1],
                              (mergeHP_CT$wnnz_buf_d[0] && (! mergeHP_CT$wnnz_buf_emitted[1]))};
  assign forkHP1_CT$wnn3_d = {mergeHP_CT$wnnz_buf_d[16:1],
                              (mergeHP_CT$wnnz_buf_d[0] && (! mergeHP_CT$wnnz_buf_emitted[2]))};
  assign mergeHP_CT$wnnz_buf_done = (mergeHP_CT$wnnz_buf_emitted | ({forkHP1_CT$wnn3_d[0],
                                                                     forkHP1_CT$wnn2_d[0],
                                                                     forkHP1_CT$wnnz_d[0]} & {forkHP1_CT$wnn3_r,
                                                                                              forkHP1_CT$wnn2_r,
                                                                                              forkHP1_CT$wnnz_r}));
  assign mergeHP_CT$wnnz_buf_r = (& mergeHP_CT$wnnz_buf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_CT$wnnz_buf_emitted <= 3'd0;
    else
      mergeHP_CT$wnnz_buf_emitted <= (mergeHP_CT$wnnz_buf_r ? 3'd0 :
                                      mergeHP_CT$wnnz_buf_done);
  
  /* mergectrl (Ty C2,
           Ty MemIn_CT$wnnz) : [(dconReadIn_CT$wnnz,MemIn_CT$wnnz),
                                (dconWriteIn_CT$wnnz,MemIn_CT$wnnz)] > (memMergeChoice_CT$wnnz,C2) (memMergeIn_CT$wnnz,MemIn_CT$wnnz) */
  logic [1:0] dconReadIn_CT$wnnz_select_d;
  assign dconReadIn_CT$wnnz_select_d = ((| dconReadIn_CT$wnnz_select_q) ? dconReadIn_CT$wnnz_select_q :
                                        (dconReadIn_CT$wnnz_d[0] ? 2'd1 :
                                         (dconWriteIn_CT$wnnz_d[0] ? 2'd2 :
                                          2'd0)));
  logic [1:0] dconReadIn_CT$wnnz_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) dconReadIn_CT$wnnz_select_q <= 2'd0;
    else
      dconReadIn_CT$wnnz_select_q <= (dconReadIn_CT$wnnz_done ? 2'd0 :
                                      dconReadIn_CT$wnnz_select_d);
  logic [1:0] dconReadIn_CT$wnnz_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) dconReadIn_CT$wnnz_emit_q <= 2'd0;
    else
      dconReadIn_CT$wnnz_emit_q <= (dconReadIn_CT$wnnz_done ? 2'd0 :
                                    dconReadIn_CT$wnnz_emit_d);
  logic [1:0] dconReadIn_CT$wnnz_emit_d;
  assign dconReadIn_CT$wnnz_emit_d = (dconReadIn_CT$wnnz_emit_q | ({memMergeChoice_CT$wnnz_d[0],
                                                                    memMergeIn_CT$wnnz_d[0]} & {memMergeChoice_CT$wnnz_r,
                                                                                                memMergeIn_CT$wnnz_r}));
  logic dconReadIn_CT$wnnz_done;
  assign dconReadIn_CT$wnnz_done = (& dconReadIn_CT$wnnz_emit_d);
  assign {dconWriteIn_CT$wnnz_r,
          dconReadIn_CT$wnnz_r} = (dconReadIn_CT$wnnz_done ? dconReadIn_CT$wnnz_select_d :
                                   2'd0);
  assign memMergeIn_CT$wnnz_d = ((dconReadIn_CT$wnnz_select_d[0] && (! dconReadIn_CT$wnnz_emit_q[0])) ? dconReadIn_CT$wnnz_d :
                                 ((dconReadIn_CT$wnnz_select_d[1] && (! dconReadIn_CT$wnnz_emit_q[0])) ? dconWriteIn_CT$wnnz_d :
                                  {132'd0, 1'd0}));
  assign memMergeChoice_CT$wnnz_d = ((dconReadIn_CT$wnnz_select_d[0] && (! dconReadIn_CT$wnnz_emit_q[1])) ? C1_2_dc(1'd1) :
                                     ((dconReadIn_CT$wnnz_select_d[1] && (! dconReadIn_CT$wnnz_emit_q[1])) ? C2_2_dc(1'd1) :
                                      {1'd0, 1'd0}));
  
  /* bram (Ty MemIn_CT$wnnz,
      Ty MemOut_CT$wnnz) : (memMergeIn_CT$wnnz_dbuf,MemIn_CT$wnnz) > (memOut_CT$wnnz,MemOut_CT$wnnz) */
  logic [114:0] memMergeIn_CT$wnnz_dbuf_mem[65535:0];
  logic [15:0] memMergeIn_CT$wnnz_dbuf_address;
  logic [114:0] memMergeIn_CT$wnnz_dbuf_din;
  logic [114:0] memOut_CT$wnnz_q;
  logic memOut_CT$wnnz_valid;
  logic memMergeIn_CT$wnnz_dbuf_we;
  logic memOut_CT$wnnz_we;
  assign memMergeIn_CT$wnnz_dbuf_din = memMergeIn_CT$wnnz_dbuf_d[132:18];
  assign memMergeIn_CT$wnnz_dbuf_address = memMergeIn_CT$wnnz_dbuf_d[17:2];
  assign memMergeIn_CT$wnnz_dbuf_we = (memMergeIn_CT$wnnz_dbuf_d[1:1] && memMergeIn_CT$wnnz_dbuf_d[0]);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        memOut_CT$wnnz_we <= 1'd0;
        memOut_CT$wnnz_valid <= 1'd0;
      end
    else
      begin
        memOut_CT$wnnz_we <= memMergeIn_CT$wnnz_dbuf_we;
        memOut_CT$wnnz_valid <= memMergeIn_CT$wnnz_dbuf_d[0];
        if (memMergeIn_CT$wnnz_dbuf_we)
          begin
            memMergeIn_CT$wnnz_dbuf_mem[memMergeIn_CT$wnnz_dbuf_address] <= memMergeIn_CT$wnnz_dbuf_din;
            memOut_CT$wnnz_q <= memMergeIn_CT$wnnz_dbuf_din;
          end
        else
          memOut_CT$wnnz_q <= memMergeIn_CT$wnnz_dbuf_mem[memMergeIn_CT$wnnz_dbuf_address];
      end
  assign memOut_CT$wnnz_d = {memOut_CT$wnnz_q,
                             memOut_CT$wnnz_we,
                             memOut_CT$wnnz_valid};
  assign memMergeIn_CT$wnnz_dbuf_r = ((! memOut_CT$wnnz_valid) || memOut_CT$wnnz_r);
  logic [31:0] profiling_MemIn_CT$wnnz_read;
  logic [31:0] profiling_MemIn_CT$wnnz_write;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        profiling_MemIn_CT$wnnz_write <= 0;
        profiling_MemIn_CT$wnnz_read <= 0;
      end
    else
      if ((memMergeIn_CT$wnnz_dbuf_we == 1'd1))
        profiling_MemIn_CT$wnnz_write <= (profiling_MemIn_CT$wnnz_write + 1);
      else
        if ((memOut_CT$wnnz_valid == 1'd1))
          profiling_MemIn_CT$wnnz_read <= (profiling_MemIn_CT$wnnz_read + 1);
  
  /* demux (Ty C2,
       Ty MemOut_CT$wnnz) : (memMergeChoice_CT$wnnz,C2) (memOut_CT$wnnz_dbuf,MemOut_CT$wnnz) > [(memReadOut_CT$wnnz,MemOut_CT$wnnz),
                                                                                                (memWriteOut_CT$wnnz,MemOut_CT$wnnz)] */
  logic [1:0] memOut_CT$wnnz_dbuf_onehotd;
  always_comb
    if ((memMergeChoice_CT$wnnz_d[0] && memOut_CT$wnnz_dbuf_d[0]))
      unique case (memMergeChoice_CT$wnnz_d[1:1])
        1'd0: memOut_CT$wnnz_dbuf_onehotd = 2'd1;
        1'd1: memOut_CT$wnnz_dbuf_onehotd = 2'd2;
        default: memOut_CT$wnnz_dbuf_onehotd = 2'd0;
      endcase
    else memOut_CT$wnnz_dbuf_onehotd = 2'd0;
  assign memReadOut_CT$wnnz_d = {memOut_CT$wnnz_dbuf_d[116:1],
                                 memOut_CT$wnnz_dbuf_onehotd[0]};
  assign memWriteOut_CT$wnnz_d = {memOut_CT$wnnz_dbuf_d[116:1],
                                  memOut_CT$wnnz_dbuf_onehotd[1]};
  assign memOut_CT$wnnz_dbuf_r = (| (memOut_CT$wnnz_dbuf_onehotd & {memWriteOut_CT$wnnz_r,
                                                                    memReadOut_CT$wnnz_r}));
  assign memMergeChoice_CT$wnnz_r = memOut_CT$wnnz_dbuf_r;
  
  /* dbuf (Ty MemIn_CT$wnnz) : (memMergeIn_CT$wnnz_rbuf,MemIn_CT$wnnz) > (memMergeIn_CT$wnnz_dbuf,MemIn_CT$wnnz) */
  assign memMergeIn_CT$wnnz_rbuf_r = ((! memMergeIn_CT$wnnz_dbuf_d[0]) || memMergeIn_CT$wnnz_dbuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memMergeIn_CT$wnnz_dbuf_d <= {132'd0, 1'd0};
    else
      if (memMergeIn_CT$wnnz_rbuf_r)
        memMergeIn_CT$wnnz_dbuf_d <= memMergeIn_CT$wnnz_rbuf_d;
  
  /* rbuf (Ty MemIn_CT$wnnz) : (memMergeIn_CT$wnnz,MemIn_CT$wnnz) > (memMergeIn_CT$wnnz_rbuf,MemIn_CT$wnnz) */
  MemIn_CT$wnnz_t memMergeIn_CT$wnnz_buf;
  assign memMergeIn_CT$wnnz_r = (! memMergeIn_CT$wnnz_buf[0]);
  assign memMergeIn_CT$wnnz_rbuf_d = (memMergeIn_CT$wnnz_buf[0] ? memMergeIn_CT$wnnz_buf :
                                      memMergeIn_CT$wnnz_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memMergeIn_CT$wnnz_buf <= {132'd0, 1'd0};
    else
      if ((memMergeIn_CT$wnnz_rbuf_r && memMergeIn_CT$wnnz_buf[0]))
        memMergeIn_CT$wnnz_buf <= {132'd0, 1'd0};
      else if (((! memMergeIn_CT$wnnz_rbuf_r) && (! memMergeIn_CT$wnnz_buf[0])))
        memMergeIn_CT$wnnz_buf <= memMergeIn_CT$wnnz_d;
  
  /* dbuf (Ty MemOut_CT$wnnz) : (memOut_CT$wnnz_rbuf,MemOut_CT$wnnz) > (memOut_CT$wnnz_dbuf,MemOut_CT$wnnz) */
  assign memOut_CT$wnnz_rbuf_r = ((! memOut_CT$wnnz_dbuf_d[0]) || memOut_CT$wnnz_dbuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memOut_CT$wnnz_dbuf_d <= {116'd0, 1'd0};
    else
      if (memOut_CT$wnnz_rbuf_r)
        memOut_CT$wnnz_dbuf_d <= memOut_CT$wnnz_rbuf_d;
  
  /* rbuf (Ty MemOut_CT$wnnz) : (memOut_CT$wnnz,MemOut_CT$wnnz) > (memOut_CT$wnnz_rbuf,MemOut_CT$wnnz) */
  MemOut_CT$wnnz_t memOut_CT$wnnz_buf;
  assign memOut_CT$wnnz_r = (! memOut_CT$wnnz_buf[0]);
  assign memOut_CT$wnnz_rbuf_d = (memOut_CT$wnnz_buf[0] ? memOut_CT$wnnz_buf :
                                  memOut_CT$wnnz_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memOut_CT$wnnz_buf <= {116'd0, 1'd0};
    else
      if ((memOut_CT$wnnz_rbuf_r && memOut_CT$wnnz_buf[0]))
        memOut_CT$wnnz_buf <= {116'd0, 1'd0};
      else if (((! memOut_CT$wnnz_rbuf_r) && (! memOut_CT$wnnz_buf[0])))
        memOut_CT$wnnz_buf <= memOut_CT$wnnz_d;
  
  /* destruct (Ty Pointer_CT$wnnz,
          Dcon Pointer_CT$wnnz) : (scfarg_0_1_argbuf,Pointer_CT$wnnz) > [(destructReadIn_CT$wnnz,Word16#)] */
  assign destructReadIn_CT$wnnz_d = {scfarg_0_1_argbuf_d[16:1],
                                     scfarg_0_1_argbuf_d[0]};
  assign scfarg_0_1_argbuf_r = destructReadIn_CT$wnnz_r;
  
  /* dcon (Ty MemIn_CT$wnnz,
      Dcon ReadIn_CT$wnnz) : [(destructReadIn_CT$wnnz,Word16#)] > (dconReadIn_CT$wnnz,MemIn_CT$wnnz) */
  assign dconReadIn_CT$wnnz_d = ReadIn_CT$wnnz_dc((& {destructReadIn_CT$wnnz_d[0]}), destructReadIn_CT$wnnz_d);
  assign {destructReadIn_CT$wnnz_r} = {1 {(dconReadIn_CT$wnnz_r && dconReadIn_CT$wnnz_d[0])}};
  
  /* destruct (Ty MemOut_CT$wnnz,
          Dcon ReadOut_CT$wnnz) : (memReadOut_CT$wnnz,MemOut_CT$wnnz) > [(readPointer_CT$wnnzscfarg_0_1_argbuf,CT$wnnz)] */
  assign readPointer_CT$wnnzscfarg_0_1_argbuf_d = {memReadOut_CT$wnnz_d[116:2],
                                                   memReadOut_CT$wnnz_d[0]};
  assign memReadOut_CT$wnnz_r = readPointer_CT$wnnzscfarg_0_1_argbuf_r;
  
  /* mergectrl (Ty C5,Ty CT$wnnz) : [(lizzieLet0_1_argbuf,CT$wnnz),
                                (lizzieLet59_1_argbuf,CT$wnnz),
                                (lizzieLet5_1_argbuf,CT$wnnz),
                                (lizzieLet60_1_argbuf,CT$wnnz),
                                (lizzieLet61_1_argbuf,CT$wnnz)] > (writeMerge_choice_CT$wnnz,C5) (writeMerge_data_CT$wnnz,CT$wnnz) */
  logic [4:0] lizzieLet0_1_argbuf_select_d;
  assign lizzieLet0_1_argbuf_select_d = ((| lizzieLet0_1_argbuf_select_q) ? lizzieLet0_1_argbuf_select_q :
                                         (lizzieLet0_1_argbuf_d[0] ? 5'd1 :
                                          (lizzieLet59_1_argbuf_d[0] ? 5'd2 :
                                           (lizzieLet5_1_argbuf_d[0] ? 5'd4 :
                                            (lizzieLet60_1_argbuf_d[0] ? 5'd8 :
                                             (lizzieLet61_1_argbuf_d[0] ? 5'd16 :
                                              5'd0))))));
  logic [4:0] lizzieLet0_1_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet0_1_argbuf_select_q <= 5'd0;
    else
      lizzieLet0_1_argbuf_select_q <= (lizzieLet0_1_argbuf_done ? 5'd0 :
                                       lizzieLet0_1_argbuf_select_d);
  logic [1:0] lizzieLet0_1_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet0_1_argbuf_emit_q <= 2'd0;
    else
      lizzieLet0_1_argbuf_emit_q <= (lizzieLet0_1_argbuf_done ? 2'd0 :
                                     lizzieLet0_1_argbuf_emit_d);
  logic [1:0] lizzieLet0_1_argbuf_emit_d;
  assign lizzieLet0_1_argbuf_emit_d = (lizzieLet0_1_argbuf_emit_q | ({writeMerge_choice_CT$wnnz_d[0],
                                                                      writeMerge_data_CT$wnnz_d[0]} & {writeMerge_choice_CT$wnnz_r,
                                                                                                       writeMerge_data_CT$wnnz_r}));
  logic lizzieLet0_1_argbuf_done;
  assign lizzieLet0_1_argbuf_done = (& lizzieLet0_1_argbuf_emit_d);
  assign {lizzieLet61_1_argbuf_r,
          lizzieLet60_1_argbuf_r,
          lizzieLet5_1_argbuf_r,
          lizzieLet59_1_argbuf_r,
          lizzieLet0_1_argbuf_r} = (lizzieLet0_1_argbuf_done ? lizzieLet0_1_argbuf_select_d :
                                    5'd0);
  assign writeMerge_data_CT$wnnz_d = ((lizzieLet0_1_argbuf_select_d[0] && (! lizzieLet0_1_argbuf_emit_q[0])) ? lizzieLet0_1_argbuf_d :
                                      ((lizzieLet0_1_argbuf_select_d[1] && (! lizzieLet0_1_argbuf_emit_q[0])) ? lizzieLet59_1_argbuf_d :
                                       ((lizzieLet0_1_argbuf_select_d[2] && (! lizzieLet0_1_argbuf_emit_q[0])) ? lizzieLet5_1_argbuf_d :
                                        ((lizzieLet0_1_argbuf_select_d[3] && (! lizzieLet0_1_argbuf_emit_q[0])) ? lizzieLet60_1_argbuf_d :
                                         ((lizzieLet0_1_argbuf_select_d[4] && (! lizzieLet0_1_argbuf_emit_q[0])) ? lizzieLet61_1_argbuf_d :
                                          {115'd0, 1'd0})))));
  assign writeMerge_choice_CT$wnnz_d = ((lizzieLet0_1_argbuf_select_d[0] && (! lizzieLet0_1_argbuf_emit_q[1])) ? C1_5_dc(1'd1) :
                                        ((lizzieLet0_1_argbuf_select_d[1] && (! lizzieLet0_1_argbuf_emit_q[1])) ? C2_5_dc(1'd1) :
                                         ((lizzieLet0_1_argbuf_select_d[2] && (! lizzieLet0_1_argbuf_emit_q[1])) ? C3_5_dc(1'd1) :
                                          ((lizzieLet0_1_argbuf_select_d[3] && (! lizzieLet0_1_argbuf_emit_q[1])) ? C4_5_dc(1'd1) :
                                           ((lizzieLet0_1_argbuf_select_d[4] && (! lizzieLet0_1_argbuf_emit_q[1])) ? C5_5_dc(1'd1) :
                                            {3'd0, 1'd0})))));
  
  /* demux (Ty C5,
       Ty Pointer_CT$wnnz) : (writeMerge_choice_CT$wnnz,C5) (demuxWriteResult_CT$wnnz,Pointer_CT$wnnz) > [(writeCT$wnnzlizzieLet0_1_argbuf,Pointer_CT$wnnz),
                                                                                                          (writeCT$wnnzlizzieLet59_1_argbuf,Pointer_CT$wnnz),
                                                                                                          (writeCT$wnnzlizzieLet5_1_argbuf,Pointer_CT$wnnz),
                                                                                                          (writeCT$wnnzlizzieLet60_1_argbuf,Pointer_CT$wnnz),
                                                                                                          (writeCT$wnnzlizzieLet61_1_argbuf,Pointer_CT$wnnz)] */
  logic [4:0] demuxWriteResult_CT$wnnz_onehotd;
  always_comb
    if ((writeMerge_choice_CT$wnnz_d[0] && demuxWriteResult_CT$wnnz_d[0]))
      unique case (writeMerge_choice_CT$wnnz_d[3:1])
        3'd0: demuxWriteResult_CT$wnnz_onehotd = 5'd1;
        3'd1: demuxWriteResult_CT$wnnz_onehotd = 5'd2;
        3'd2: demuxWriteResult_CT$wnnz_onehotd = 5'd4;
        3'd3: demuxWriteResult_CT$wnnz_onehotd = 5'd8;
        3'd4: demuxWriteResult_CT$wnnz_onehotd = 5'd16;
        default: demuxWriteResult_CT$wnnz_onehotd = 5'd0;
      endcase
    else demuxWriteResult_CT$wnnz_onehotd = 5'd0;
  assign writeCT$wnnzlizzieLet0_1_argbuf_d = {demuxWriteResult_CT$wnnz_d[16:1],
                                              demuxWriteResult_CT$wnnz_onehotd[0]};
  assign writeCT$wnnzlizzieLet59_1_argbuf_d = {demuxWriteResult_CT$wnnz_d[16:1],
                                               demuxWriteResult_CT$wnnz_onehotd[1]};
  assign writeCT$wnnzlizzieLet5_1_argbuf_d = {demuxWriteResult_CT$wnnz_d[16:1],
                                              demuxWriteResult_CT$wnnz_onehotd[2]};
  assign writeCT$wnnzlizzieLet60_1_argbuf_d = {demuxWriteResult_CT$wnnz_d[16:1],
                                               demuxWriteResult_CT$wnnz_onehotd[3]};
  assign writeCT$wnnzlizzieLet61_1_argbuf_d = {demuxWriteResult_CT$wnnz_d[16:1],
                                               demuxWriteResult_CT$wnnz_onehotd[4]};
  assign demuxWriteResult_CT$wnnz_r = (| (demuxWriteResult_CT$wnnz_onehotd & {writeCT$wnnzlizzieLet61_1_argbuf_r,
                                                                              writeCT$wnnzlizzieLet60_1_argbuf_r,
                                                                              writeCT$wnnzlizzieLet5_1_argbuf_r,
                                                                              writeCT$wnnzlizzieLet59_1_argbuf_r,
                                                                              writeCT$wnnzlizzieLet0_1_argbuf_r}));
  assign writeMerge_choice_CT$wnnz_r = demuxWriteResult_CT$wnnz_r;
  
  /* dcon (Ty MemIn_CT$wnnz,
      Dcon WriteIn_CT$wnnz) : [(forkHP1_CT$wnn2,Word16#),
                               (writeMerge_data_CT$wnnz,CT$wnnz)] > (dconWriteIn_CT$wnnz,MemIn_CT$wnnz) */
  assign dconWriteIn_CT$wnnz_d = WriteIn_CT$wnnz_dc((& {forkHP1_CT$wnn2_d[0],
                                                        writeMerge_data_CT$wnnz_d[0]}), forkHP1_CT$wnn2_d, writeMerge_data_CT$wnnz_d);
  assign {forkHP1_CT$wnn2_r,
          writeMerge_data_CT$wnnz_r} = {2 {(dconWriteIn_CT$wnnz_r && dconWriteIn_CT$wnnz_d[0])}};
  
  /* dcon (Ty Pointer_CT$wnnz,
      Dcon Pointer_CT$wnnz) : [(forkHP1_CT$wnn3,Word16#)] > (dconPtr_CT$wnnz,Pointer_CT$wnnz) */
  assign dconPtr_CT$wnnz_d = Pointer_CT$wnnz_dc((& {forkHP1_CT$wnn3_d[0]}), forkHP1_CT$wnn3_d);
  assign {forkHP1_CT$wnn3_r} = {1 {(dconPtr_CT$wnnz_r && dconPtr_CT$wnnz_d[0])}};
  
  /* demux (Ty MemOut_CT$wnnz,
       Ty Pointer_CT$wnnz) : (memWriteOut_CT$wnnz,MemOut_CT$wnnz) (dconPtr_CT$wnnz,Pointer_CT$wnnz) > [(_259,Pointer_CT$wnnz),
                                                                                                       (demuxWriteResult_CT$wnnz,Pointer_CT$wnnz)] */
  logic [1:0] dconPtr_CT$wnnz_onehotd;
  always_comb
    if ((memWriteOut_CT$wnnz_d[0] && dconPtr_CT$wnnz_d[0]))
      unique case (memWriteOut_CT$wnnz_d[1:1])
        1'd0: dconPtr_CT$wnnz_onehotd = 2'd1;
        1'd1: dconPtr_CT$wnnz_onehotd = 2'd2;
        default: dconPtr_CT$wnnz_onehotd = 2'd0;
      endcase
    else dconPtr_CT$wnnz_onehotd = 2'd0;
  assign _259_d = {dconPtr_CT$wnnz_d[16:1],
                   dconPtr_CT$wnnz_onehotd[0]};
  assign demuxWriteResult_CT$wnnz_d = {dconPtr_CT$wnnz_d[16:1],
                                       dconPtr_CT$wnnz_onehotd[1]};
  assign dconPtr_CT$wnnz_r = (| (dconPtr_CT$wnnz_onehotd & {demuxWriteResult_CT$wnnz_r,
                                                            _259_r}));
  assign memWriteOut_CT$wnnz_r = dconPtr_CT$wnnz_r;
  
  /* const (Ty Word16#,
       Lit 0) : (go_1_dummy_write_QTree_Int,Go) > (initHP_QTree_Int,Word16#) */
  assign initHP_QTree_Int_d = {16'd0,
                               go_1_dummy_write_QTree_Int_d[0]};
  assign go_1_dummy_write_QTree_Int_r = initHP_QTree_Int_r;
  
  /* const (Ty Word16#,
       Lit 1) : (incrHP_QTree_Int1,Go) > (incrHP_QTree_Int,Word16#) */
  assign incrHP_QTree_Int_d = {16'd1, incrHP_QTree_Int1_d[0]};
  assign incrHP_QTree_Int1_r = incrHP_QTree_Int_r;
  
  /* merge (Ty Go) : [(go_2_dummy_write_QTree_Int,Go),
                 (incrHP_QTree_Int2,Go)] > (incrHP_mergeQTree_Int,Go) */
  logic [1:0] incrHP_mergeQTree_Int_selected;
  logic [1:0] incrHP_mergeQTree_Int_select;
  always_comb
    begin
      incrHP_mergeQTree_Int_selected = 2'd0;
      if ((| incrHP_mergeQTree_Int_select))
        incrHP_mergeQTree_Int_selected = incrHP_mergeQTree_Int_select;
      else
        if (go_2_dummy_write_QTree_Int_d[0])
          incrHP_mergeQTree_Int_selected[0] = 1'd1;
        else if (incrHP_QTree_Int2_d[0])
          incrHP_mergeQTree_Int_selected[1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeQTree_Int_select <= 2'd0;
    else
      incrHP_mergeQTree_Int_select <= (incrHP_mergeQTree_Int_r ? 2'd0 :
                                       incrHP_mergeQTree_Int_selected);
  always_comb
    if (incrHP_mergeQTree_Int_selected[0])
      incrHP_mergeQTree_Int_d = go_2_dummy_write_QTree_Int_d;
    else if (incrHP_mergeQTree_Int_selected[1])
      incrHP_mergeQTree_Int_d = incrHP_QTree_Int2_d;
    else incrHP_mergeQTree_Int_d = 1'd0;
  assign {incrHP_QTree_Int2_r,
          go_2_dummy_write_QTree_Int_r} = (incrHP_mergeQTree_Int_r ? incrHP_mergeQTree_Int_selected :
                                           2'd0);
  
  /* fork (Ty Go) : (incrHP_mergeQTree_Int_buf,Go) > [(incrHP_QTree_Int1,Go),
                                                 (incrHP_QTree_Int2,Go)] */
  logic [1:0] incrHP_mergeQTree_Int_buf_emitted;
  logic [1:0] incrHP_mergeQTree_Int_buf_done;
  assign incrHP_QTree_Int1_d = (incrHP_mergeQTree_Int_buf_d[0] && (! incrHP_mergeQTree_Int_buf_emitted[0]));
  assign incrHP_QTree_Int2_d = (incrHP_mergeQTree_Int_buf_d[0] && (! incrHP_mergeQTree_Int_buf_emitted[1]));
  assign incrHP_mergeQTree_Int_buf_done = (incrHP_mergeQTree_Int_buf_emitted | ({incrHP_QTree_Int2_d[0],
                                                                                 incrHP_QTree_Int1_d[0]} & {incrHP_QTree_Int2_r,
                                                                                                            incrHP_QTree_Int1_r}));
  assign incrHP_mergeQTree_Int_buf_r = (& incrHP_mergeQTree_Int_buf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeQTree_Int_buf_emitted <= 2'd0;
    else
      incrHP_mergeQTree_Int_buf_emitted <= (incrHP_mergeQTree_Int_buf_r ? 2'd0 :
                                            incrHP_mergeQTree_Int_buf_done);
  
  /* op_add (Ty Word16#) : (incrHP_QTree_Int,Word16#) (forkHP1_QTree_Int,Word16#) > (addHP_QTree_Int,Word16#) */
  assign addHP_QTree_Int_d = {(incrHP_QTree_Int_d[16:1] + forkHP1_QTree_Int_d[16:1]),
                              (incrHP_QTree_Int_d[0] && forkHP1_QTree_Int_d[0])};
  assign {incrHP_QTree_Int_r,
          forkHP1_QTree_Int_r} = {2 {(addHP_QTree_Int_r && addHP_QTree_Int_d[0])}};
  
  /* merge (Ty Word16#) : [(initHP_QTree_Int,Word16#),
                      (addHP_QTree_Int,Word16#)] > (mergeHP_QTree_Int,Word16#) */
  logic [1:0] mergeHP_QTree_Int_selected;
  logic [1:0] mergeHP_QTree_Int_select;
  always_comb
    begin
      mergeHP_QTree_Int_selected = 2'd0;
      if ((| mergeHP_QTree_Int_select))
        mergeHP_QTree_Int_selected = mergeHP_QTree_Int_select;
      else
        if (initHP_QTree_Int_d[0]) mergeHP_QTree_Int_selected[0] = 1'd1;
        else if (addHP_QTree_Int_d[0])
          mergeHP_QTree_Int_selected[1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_QTree_Int_select <= 2'd0;
    else
      mergeHP_QTree_Int_select <= (mergeHP_QTree_Int_r ? 2'd0 :
                                   mergeHP_QTree_Int_selected);
  always_comb
    if (mergeHP_QTree_Int_selected[0])
      mergeHP_QTree_Int_d = initHP_QTree_Int_d;
    else if (mergeHP_QTree_Int_selected[1])
      mergeHP_QTree_Int_d = addHP_QTree_Int_d;
    else mergeHP_QTree_Int_d = {16'd0, 1'd0};
  assign {addHP_QTree_Int_r,
          initHP_QTree_Int_r} = (mergeHP_QTree_Int_r ? mergeHP_QTree_Int_selected :
                                 2'd0);
  
  /* buf (Ty Go) : (incrHP_mergeQTree_Int,Go) > (incrHP_mergeQTree_Int_buf,Go) */
  Go_t incrHP_mergeQTree_Int_bufchan_d;
  logic incrHP_mergeQTree_Int_bufchan_r;
  assign incrHP_mergeQTree_Int_r = ((! incrHP_mergeQTree_Int_bufchan_d[0]) || incrHP_mergeQTree_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeQTree_Int_bufchan_d <= 1'd0;
    else
      if (incrHP_mergeQTree_Int_r)
        incrHP_mergeQTree_Int_bufchan_d <= incrHP_mergeQTree_Int_d;
  Go_t incrHP_mergeQTree_Int_bufchan_buf;
  assign incrHP_mergeQTree_Int_bufchan_r = (! incrHP_mergeQTree_Int_bufchan_buf[0]);
  assign incrHP_mergeQTree_Int_buf_d = (incrHP_mergeQTree_Int_bufchan_buf[0] ? incrHP_mergeQTree_Int_bufchan_buf :
                                        incrHP_mergeQTree_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeQTree_Int_bufchan_buf <= 1'd0;
    else
      if ((incrHP_mergeQTree_Int_buf_r && incrHP_mergeQTree_Int_bufchan_buf[0]))
        incrHP_mergeQTree_Int_bufchan_buf <= 1'd0;
      else if (((! incrHP_mergeQTree_Int_buf_r) && (! incrHP_mergeQTree_Int_bufchan_buf[0])))
        incrHP_mergeQTree_Int_bufchan_buf <= incrHP_mergeQTree_Int_bufchan_d;
  
  /* buf (Ty Word16#) : (mergeHP_QTree_Int,Word16#) > (mergeHP_QTree_Int_buf,Word16#) */
  \Word16#_t  mergeHP_QTree_Int_bufchan_d;
  logic mergeHP_QTree_Int_bufchan_r;
  assign mergeHP_QTree_Int_r = ((! mergeHP_QTree_Int_bufchan_d[0]) || mergeHP_QTree_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_QTree_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (mergeHP_QTree_Int_r)
        mergeHP_QTree_Int_bufchan_d <= mergeHP_QTree_Int_d;
  \Word16#_t  mergeHP_QTree_Int_bufchan_buf;
  assign mergeHP_QTree_Int_bufchan_r = (! mergeHP_QTree_Int_bufchan_buf[0]);
  assign mergeHP_QTree_Int_buf_d = (mergeHP_QTree_Int_bufchan_buf[0] ? mergeHP_QTree_Int_bufchan_buf :
                                    mergeHP_QTree_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      mergeHP_QTree_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((mergeHP_QTree_Int_buf_r && mergeHP_QTree_Int_bufchan_buf[0]))
        mergeHP_QTree_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! mergeHP_QTree_Int_buf_r) && (! mergeHP_QTree_Int_bufchan_buf[0])))
        mergeHP_QTree_Int_bufchan_buf <= mergeHP_QTree_Int_bufchan_d;
  
  /* sink (Ty Word16#) : (forkHP1_QTree_Int_snk,Word16#) > */
  assign {forkHP1_QTree_Int_snk_r,
          forkHP1_QTree_Int_snk_dout} = {forkHP1_QTree_Int_snk_rout,
                                         forkHP1_QTree_Int_snk_d};
  
  /* source (Ty Go) : > (\QTree_Int_src,Go) */
  
  /* fork (Ty Go) : (\QTree_Int_src,Go) > [(go_1_dummy_write_QTree_Int,Go),
                                      (go_2_dummy_write_QTree_Int,Go)] */
  logic [1:0] \\QTree_Int_src_emitted ;
  logic [1:0] \\QTree_Int_src_done ;
  assign go_1_dummy_write_QTree_Int_d = (\\QTree_Int_src_d [0] && (! \\QTree_Int_src_emitted [0]));
  assign go_2_dummy_write_QTree_Int_d = (\\QTree_Int_src_d [0] && (! \\QTree_Int_src_emitted [1]));
  assign \\QTree_Int_src_done  = (\\QTree_Int_src_emitted  | ({go_2_dummy_write_QTree_Int_d[0],
                                                               go_1_dummy_write_QTree_Int_d[0]} & {go_2_dummy_write_QTree_Int_r,
                                                                                                   go_1_dummy_write_QTree_Int_r}));
  assign \\QTree_Int_src_r  = (& \\QTree_Int_src_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \\QTree_Int_src_emitted  <= 2'd0;
    else
      \\QTree_Int_src_emitted  <= (\\QTree_Int_src_r  ? 2'd0 :
                                   \\QTree_Int_src_done );
  
  /* source (Ty QTree_Int) : > (dummy_write_QTree_Int,QTree_Int) */
  
  /* sink (Ty Pointer_QTree_Int) : (dummy_write_QTree_Int_sink,Pointer_QTree_Int) > */
  assign {dummy_write_QTree_Int_sink_r,
          dummy_write_QTree_Int_sink_dout} = {dummy_write_QTree_Int_sink_rout,
                                              dummy_write_QTree_Int_sink_d};
  
  /* fork (Ty Word16#) : (mergeHP_QTree_Int_buf,Word16#) > [(forkHP1_QTree_Int,Word16#),
                                                       (forkHP1_QTree_Int_snk,Word16#),
                                                       (forkHP1_QTree_In3,Word16#),
                                                       (forkHP1_QTree_In4,Word16#)] */
  logic [3:0] mergeHP_QTree_Int_buf_emitted;
  logic [3:0] mergeHP_QTree_Int_buf_done;
  assign forkHP1_QTree_Int_d = {mergeHP_QTree_Int_buf_d[16:1],
                                (mergeHP_QTree_Int_buf_d[0] && (! mergeHP_QTree_Int_buf_emitted[0]))};
  assign forkHP1_QTree_Int_snk_d = {mergeHP_QTree_Int_buf_d[16:1],
                                    (mergeHP_QTree_Int_buf_d[0] && (! mergeHP_QTree_Int_buf_emitted[1]))};
  assign forkHP1_QTree_In3_d = {mergeHP_QTree_Int_buf_d[16:1],
                                (mergeHP_QTree_Int_buf_d[0] && (! mergeHP_QTree_Int_buf_emitted[2]))};
  assign forkHP1_QTree_In4_d = {mergeHP_QTree_Int_buf_d[16:1],
                                (mergeHP_QTree_Int_buf_d[0] && (! mergeHP_QTree_Int_buf_emitted[3]))};
  assign mergeHP_QTree_Int_buf_done = (mergeHP_QTree_Int_buf_emitted | ({forkHP1_QTree_In4_d[0],
                                                                         forkHP1_QTree_In3_d[0],
                                                                         forkHP1_QTree_Int_snk_d[0],
                                                                         forkHP1_QTree_Int_d[0]} & {forkHP1_QTree_In4_r,
                                                                                                    forkHP1_QTree_In3_r,
                                                                                                    forkHP1_QTree_Int_snk_r,
                                                                                                    forkHP1_QTree_Int_r}));
  assign mergeHP_QTree_Int_buf_r = (& mergeHP_QTree_Int_buf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_QTree_Int_buf_emitted <= 4'd0;
    else
      mergeHP_QTree_Int_buf_emitted <= (mergeHP_QTree_Int_buf_r ? 4'd0 :
                                        mergeHP_QTree_Int_buf_done);
  
  /* mergectrl (Ty C2,
           Ty MemIn_QTree_Int) : [(dconReadIn_QTree_Int,MemIn_QTree_Int),
                                  (dconWriteIn_QTree_Int,MemIn_QTree_Int)] > (memMergeChoice_QTree_Int,C2) (memMergeIn_QTree_Int,MemIn_QTree_Int) */
  logic [1:0] dconReadIn_QTree_Int_select_d;
  assign dconReadIn_QTree_Int_select_d = ((| dconReadIn_QTree_Int_select_q) ? dconReadIn_QTree_Int_select_q :
                                          (dconReadIn_QTree_Int_d[0] ? 2'd1 :
                                           (dconWriteIn_QTree_Int_d[0] ? 2'd2 :
                                            2'd0)));
  logic [1:0] dconReadIn_QTree_Int_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) dconReadIn_QTree_Int_select_q <= 2'd0;
    else
      dconReadIn_QTree_Int_select_q <= (dconReadIn_QTree_Int_done ? 2'd0 :
                                        dconReadIn_QTree_Int_select_d);
  logic [1:0] dconReadIn_QTree_Int_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) dconReadIn_QTree_Int_emit_q <= 2'd0;
    else
      dconReadIn_QTree_Int_emit_q <= (dconReadIn_QTree_Int_done ? 2'd0 :
                                      dconReadIn_QTree_Int_emit_d);
  logic [1:0] dconReadIn_QTree_Int_emit_d;
  assign dconReadIn_QTree_Int_emit_d = (dconReadIn_QTree_Int_emit_q | ({memMergeChoice_QTree_Int_d[0],
                                                                        memMergeIn_QTree_Int_d[0]} & {memMergeChoice_QTree_Int_r,
                                                                                                      memMergeIn_QTree_Int_r}));
  logic dconReadIn_QTree_Int_done;
  assign dconReadIn_QTree_Int_done = (& dconReadIn_QTree_Int_emit_d);
  assign {dconWriteIn_QTree_Int_r,
          dconReadIn_QTree_Int_r} = (dconReadIn_QTree_Int_done ? dconReadIn_QTree_Int_select_d :
                                     2'd0);
  assign memMergeIn_QTree_Int_d = ((dconReadIn_QTree_Int_select_d[0] && (! dconReadIn_QTree_Int_emit_q[0])) ? dconReadIn_QTree_Int_d :
                                   ((dconReadIn_QTree_Int_select_d[1] && (! dconReadIn_QTree_Int_emit_q[0])) ? dconWriteIn_QTree_Int_d :
                                    {83'd0, 1'd0}));
  assign memMergeChoice_QTree_Int_d = ((dconReadIn_QTree_Int_select_d[0] && (! dconReadIn_QTree_Int_emit_q[1])) ? C1_2_dc(1'd1) :
                                       ((dconReadIn_QTree_Int_select_d[1] && (! dconReadIn_QTree_Int_emit_q[1])) ? C2_2_dc(1'd1) :
                                        {1'd0, 1'd0}));
  
  /* bram (Ty MemIn_QTree_Int,
      Ty MemOut_QTree_Int) : (memMergeIn_QTree_Int_dbuf,MemIn_QTree_Int) > (memOut_QTree_Int,MemOut_QTree_Int) */
  logic [65:0] memMergeIn_QTree_Int_dbuf_mem[65535:0];
  logic [15:0] memMergeIn_QTree_Int_dbuf_address;
  logic [65:0] memMergeIn_QTree_Int_dbuf_din;
  logic [65:0] memOut_QTree_Int_q;
  logic memOut_QTree_Int_valid;
  logic memMergeIn_QTree_Int_dbuf_we;
  logic memOut_QTree_Int_we;
  assign memMergeIn_QTree_Int_dbuf_din = memMergeIn_QTree_Int_dbuf_d[83:18];
  assign memMergeIn_QTree_Int_dbuf_address = memMergeIn_QTree_Int_dbuf_d[17:2];
  assign memMergeIn_QTree_Int_dbuf_we = (memMergeIn_QTree_Int_dbuf_d[1:1] && memMergeIn_QTree_Int_dbuf_d[0]);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        memOut_QTree_Int_we <= 1'd0;
        memOut_QTree_Int_valid <= 1'd0;
      end
    else
      begin
        memOut_QTree_Int_we <= memMergeIn_QTree_Int_dbuf_we;
        memOut_QTree_Int_valid <= memMergeIn_QTree_Int_dbuf_d[0];
        if (memMergeIn_QTree_Int_dbuf_we)
          begin
            memMergeIn_QTree_Int_dbuf_mem[memMergeIn_QTree_Int_dbuf_address] <= memMergeIn_QTree_Int_dbuf_din;
            memOut_QTree_Int_q <= memMergeIn_QTree_Int_dbuf_din;
          end
        else
          memOut_QTree_Int_q <= memMergeIn_QTree_Int_dbuf_mem[memMergeIn_QTree_Int_dbuf_address];
      end
  assign memOut_QTree_Int_d = {memOut_QTree_Int_q,
                               memOut_QTree_Int_we,
                               memOut_QTree_Int_valid};
  assign memMergeIn_QTree_Int_dbuf_r = ((! memOut_QTree_Int_valid) || memOut_QTree_Int_r);
  logic [31:0] profiling_MemIn_QTree_Int_read;
  logic [31:0] profiling_MemIn_QTree_Int_write;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        profiling_MemIn_QTree_Int_write <= 0;
        profiling_MemIn_QTree_Int_read <= 0;
      end
    else
      if ((memMergeIn_QTree_Int_dbuf_we == 1'd1))
        profiling_MemIn_QTree_Int_write <= (profiling_MemIn_QTree_Int_write + 1);
      else
        if ((memOut_QTree_Int_valid == 1'd1))
          profiling_MemIn_QTree_Int_read <= (profiling_MemIn_QTree_Int_read + 1);
  
  /* demux (Ty C2,
       Ty MemOut_QTree_Int) : (memMergeChoice_QTree_Int,C2) (memOut_QTree_Int_dbuf,MemOut_QTree_Int) > [(memReadOut_QTree_Int,MemOut_QTree_Int),
                                                                                                        (memWriteOut_QTree_Int,MemOut_QTree_Int)] */
  logic [1:0] memOut_QTree_Int_dbuf_onehotd;
  always_comb
    if ((memMergeChoice_QTree_Int_d[0] && memOut_QTree_Int_dbuf_d[0]))
      unique case (memMergeChoice_QTree_Int_d[1:1])
        1'd0: memOut_QTree_Int_dbuf_onehotd = 2'd1;
        1'd1: memOut_QTree_Int_dbuf_onehotd = 2'd2;
        default: memOut_QTree_Int_dbuf_onehotd = 2'd0;
      endcase
    else memOut_QTree_Int_dbuf_onehotd = 2'd0;
  assign memReadOut_QTree_Int_d = {memOut_QTree_Int_dbuf_d[67:1],
                                   memOut_QTree_Int_dbuf_onehotd[0]};
  assign memWriteOut_QTree_Int_d = {memOut_QTree_Int_dbuf_d[67:1],
                                    memOut_QTree_Int_dbuf_onehotd[1]};
  assign memOut_QTree_Int_dbuf_r = (| (memOut_QTree_Int_dbuf_onehotd & {memWriteOut_QTree_Int_r,
                                                                        memReadOut_QTree_Int_r}));
  assign memMergeChoice_QTree_Int_r = memOut_QTree_Int_dbuf_r;
  
  /* dbuf (Ty MemIn_QTree_Int) : (memMergeIn_QTree_Int_rbuf,MemIn_QTree_Int) > (memMergeIn_QTree_Int_dbuf,MemIn_QTree_Int) */
  assign memMergeIn_QTree_Int_rbuf_r = ((! memMergeIn_QTree_Int_dbuf_d[0]) || memMergeIn_QTree_Int_dbuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memMergeIn_QTree_Int_dbuf_d <= {83'd0, 1'd0};
    else
      if (memMergeIn_QTree_Int_rbuf_r)
        memMergeIn_QTree_Int_dbuf_d <= memMergeIn_QTree_Int_rbuf_d;
  
  /* rbuf (Ty MemIn_QTree_Int) : (memMergeIn_QTree_Int,MemIn_QTree_Int) > (memMergeIn_QTree_Int_rbuf,MemIn_QTree_Int) */
  MemIn_QTree_Int_t memMergeIn_QTree_Int_buf;
  assign memMergeIn_QTree_Int_r = (! memMergeIn_QTree_Int_buf[0]);
  assign memMergeIn_QTree_Int_rbuf_d = (memMergeIn_QTree_Int_buf[0] ? memMergeIn_QTree_Int_buf :
                                        memMergeIn_QTree_Int_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memMergeIn_QTree_Int_buf <= {83'd0, 1'd0};
    else
      if ((memMergeIn_QTree_Int_rbuf_r && memMergeIn_QTree_Int_buf[0]))
        memMergeIn_QTree_Int_buf <= {83'd0, 1'd0};
      else if (((! memMergeIn_QTree_Int_rbuf_r) && (! memMergeIn_QTree_Int_buf[0])))
        memMergeIn_QTree_Int_buf <= memMergeIn_QTree_Int_d;
  
  /* dbuf (Ty MemOut_QTree_Int) : (memOut_QTree_Int_rbuf,MemOut_QTree_Int) > (memOut_QTree_Int_dbuf,MemOut_QTree_Int) */
  assign memOut_QTree_Int_rbuf_r = ((! memOut_QTree_Int_dbuf_d[0]) || memOut_QTree_Int_dbuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memOut_QTree_Int_dbuf_d <= {67'd0, 1'd0};
    else
      if (memOut_QTree_Int_rbuf_r)
        memOut_QTree_Int_dbuf_d <= memOut_QTree_Int_rbuf_d;
  
  /* rbuf (Ty MemOut_QTree_Int) : (memOut_QTree_Int,MemOut_QTree_Int) > (memOut_QTree_Int_rbuf,MemOut_QTree_Int) */
  MemOut_QTree_Int_t memOut_QTree_Int_buf;
  assign memOut_QTree_Int_r = (! memOut_QTree_Int_buf[0]);
  assign memOut_QTree_Int_rbuf_d = (memOut_QTree_Int_buf[0] ? memOut_QTree_Int_buf :
                                    memOut_QTree_Int_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memOut_QTree_Int_buf <= {67'd0, 1'd0};
    else
      if ((memOut_QTree_Int_rbuf_r && memOut_QTree_Int_buf[0]))
        memOut_QTree_Int_buf <= {67'd0, 1'd0};
      else if (((! memOut_QTree_Int_rbuf_r) && (! memOut_QTree_Int_buf[0])))
        memOut_QTree_Int_buf <= memOut_QTree_Int_d;
  
  /* mergectrl (Ty C6,
           Ty Pointer_QTree_Int) : [(m1aeq_1_argbuf,Pointer_QTree_Int),
                                    (m2aer_1_argbuf,Pointer_QTree_Int),
                                    (m3aes_1_argbuf,Pointer_QTree_Int),
                                    (q4afj_1_argbuf,Pointer_QTree_Int),
                                    (t4afk_1_argbuf,Pointer_QTree_Int),
                                    (wsmk_1_1_argbuf,Pointer_QTree_Int)] > (readMerge_choice_QTree_Int,C6) (readMerge_data_QTree_Int,Pointer_QTree_Int) */
  logic [5:0] m1aeq_1_argbuf_select_d;
  assign m1aeq_1_argbuf_select_d = ((| m1aeq_1_argbuf_select_q) ? m1aeq_1_argbuf_select_q :
                                    (m1aeq_1_argbuf_d[0] ? 6'd1 :
                                     (m2aer_1_argbuf_d[0] ? 6'd2 :
                                      (m3aes_1_argbuf_d[0] ? 6'd4 :
                                       (q4afj_1_argbuf_d[0] ? 6'd8 :
                                        (t4afk_1_argbuf_d[0] ? 6'd16 :
                                         (wsmk_1_1_argbuf_d[0] ? 6'd32 :
                                          6'd0)))))));
  logic [5:0] m1aeq_1_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m1aeq_1_argbuf_select_q <= 6'd0;
    else
      m1aeq_1_argbuf_select_q <= (m1aeq_1_argbuf_done ? 6'd0 :
                                  m1aeq_1_argbuf_select_d);
  logic [1:0] m1aeq_1_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m1aeq_1_argbuf_emit_q <= 2'd0;
    else
      m1aeq_1_argbuf_emit_q <= (m1aeq_1_argbuf_done ? 2'd0 :
                                m1aeq_1_argbuf_emit_d);
  logic [1:0] m1aeq_1_argbuf_emit_d;
  assign m1aeq_1_argbuf_emit_d = (m1aeq_1_argbuf_emit_q | ({readMerge_choice_QTree_Int_d[0],
                                                            readMerge_data_QTree_Int_d[0]} & {readMerge_choice_QTree_Int_r,
                                                                                              readMerge_data_QTree_Int_r}));
  logic m1aeq_1_argbuf_done;
  assign m1aeq_1_argbuf_done = (& m1aeq_1_argbuf_emit_d);
  assign {wsmk_1_1_argbuf_r,
          t4afk_1_argbuf_r,
          q4afj_1_argbuf_r,
          m3aes_1_argbuf_r,
          m2aer_1_argbuf_r,
          m1aeq_1_argbuf_r} = (m1aeq_1_argbuf_done ? m1aeq_1_argbuf_select_d :
                               6'd0);
  assign readMerge_data_QTree_Int_d = ((m1aeq_1_argbuf_select_d[0] && (! m1aeq_1_argbuf_emit_q[0])) ? m1aeq_1_argbuf_d :
                                       ((m1aeq_1_argbuf_select_d[1] && (! m1aeq_1_argbuf_emit_q[0])) ? m2aer_1_argbuf_d :
                                        ((m1aeq_1_argbuf_select_d[2] && (! m1aeq_1_argbuf_emit_q[0])) ? m3aes_1_argbuf_d :
                                         ((m1aeq_1_argbuf_select_d[3] && (! m1aeq_1_argbuf_emit_q[0])) ? q4afj_1_argbuf_d :
                                          ((m1aeq_1_argbuf_select_d[4] && (! m1aeq_1_argbuf_emit_q[0])) ? t4afk_1_argbuf_d :
                                           ((m1aeq_1_argbuf_select_d[5] && (! m1aeq_1_argbuf_emit_q[0])) ? wsmk_1_1_argbuf_d :
                                            {16'd0, 1'd0}))))));
  assign readMerge_choice_QTree_Int_d = ((m1aeq_1_argbuf_select_d[0] && (! m1aeq_1_argbuf_emit_q[1])) ? C1_6_dc(1'd1) :
                                         ((m1aeq_1_argbuf_select_d[1] && (! m1aeq_1_argbuf_emit_q[1])) ? C2_6_dc(1'd1) :
                                          ((m1aeq_1_argbuf_select_d[2] && (! m1aeq_1_argbuf_emit_q[1])) ? C3_6_dc(1'd1) :
                                           ((m1aeq_1_argbuf_select_d[3] && (! m1aeq_1_argbuf_emit_q[1])) ? C4_6_dc(1'd1) :
                                            ((m1aeq_1_argbuf_select_d[4] && (! m1aeq_1_argbuf_emit_q[1])) ? C5_6_dc(1'd1) :
                                             ((m1aeq_1_argbuf_select_d[5] && (! m1aeq_1_argbuf_emit_q[1])) ? C6_6_dc(1'd1) :
                                              {3'd0, 1'd0}))))));
  
  /* demux (Ty C6,
       Ty QTree_Int) : (readMerge_choice_QTree_Int,C6) (destructReadOut_QTree_Int,QTree_Int) > [(readPointer_QTree_Intm1aeq_1_argbuf,QTree_Int),
                                                                                                (readPointer_QTree_Intm2aer_1_argbuf,QTree_Int),
                                                                                                (readPointer_QTree_Intm3aes_1_argbuf,QTree_Int),
                                                                                                (readPointer_QTree_Intq4afj_1_argbuf,QTree_Int),
                                                                                                (readPointer_QTree_Intt4afk_1_argbuf,QTree_Int),
                                                                                                (readPointer_QTree_Intwsmk_1_1_argbuf,QTree_Int)] */
  logic [5:0] destructReadOut_QTree_Int_onehotd;
  always_comb
    if ((readMerge_choice_QTree_Int_d[0] && destructReadOut_QTree_Int_d[0]))
      unique case (readMerge_choice_QTree_Int_d[3:1])
        3'd0: destructReadOut_QTree_Int_onehotd = 6'd1;
        3'd1: destructReadOut_QTree_Int_onehotd = 6'd2;
        3'd2: destructReadOut_QTree_Int_onehotd = 6'd4;
        3'd3: destructReadOut_QTree_Int_onehotd = 6'd8;
        3'd4: destructReadOut_QTree_Int_onehotd = 6'd16;
        3'd5: destructReadOut_QTree_Int_onehotd = 6'd32;
        default: destructReadOut_QTree_Int_onehotd = 6'd0;
      endcase
    else destructReadOut_QTree_Int_onehotd = 6'd0;
  assign readPointer_QTree_Intm1aeq_1_argbuf_d = {destructReadOut_QTree_Int_d[66:1],
                                                  destructReadOut_QTree_Int_onehotd[0]};
  assign readPointer_QTree_Intm2aer_1_argbuf_d = {destructReadOut_QTree_Int_d[66:1],
                                                  destructReadOut_QTree_Int_onehotd[1]};
  assign readPointer_QTree_Intm3aes_1_argbuf_d = {destructReadOut_QTree_Int_d[66:1],
                                                  destructReadOut_QTree_Int_onehotd[2]};
  assign readPointer_QTree_Intq4afj_1_argbuf_d = {destructReadOut_QTree_Int_d[66:1],
                                                  destructReadOut_QTree_Int_onehotd[3]};
  assign readPointer_QTree_Intt4afk_1_argbuf_d = {destructReadOut_QTree_Int_d[66:1],
                                                  destructReadOut_QTree_Int_onehotd[4]};
  assign readPointer_QTree_Intwsmk_1_1_argbuf_d = {destructReadOut_QTree_Int_d[66:1],
                                                   destructReadOut_QTree_Int_onehotd[5]};
  assign destructReadOut_QTree_Int_r = (| (destructReadOut_QTree_Int_onehotd & {readPointer_QTree_Intwsmk_1_1_argbuf_r,
                                                                                readPointer_QTree_Intt4afk_1_argbuf_r,
                                                                                readPointer_QTree_Intq4afj_1_argbuf_r,
                                                                                readPointer_QTree_Intm3aes_1_argbuf_r,
                                                                                readPointer_QTree_Intm2aer_1_argbuf_r,
                                                                                readPointer_QTree_Intm1aeq_1_argbuf_r}));
  assign readMerge_choice_QTree_Int_r = destructReadOut_QTree_Int_r;
  
  /* destruct (Ty Pointer_QTree_Int,
          Dcon Pointer_QTree_Int) : (readMerge_data_QTree_Int,Pointer_QTree_Int) > [(destructReadIn_QTree_Int,Word16#)] */
  assign destructReadIn_QTree_Int_d = {readMerge_data_QTree_Int_d[16:1],
                                       readMerge_data_QTree_Int_d[0]};
  assign readMerge_data_QTree_Int_r = destructReadIn_QTree_Int_r;
  
  /* dcon (Ty MemIn_QTree_Int,
      Dcon ReadIn_QTree_Int) : [(destructReadIn_QTree_Int,Word16#)] > (dconReadIn_QTree_Int,MemIn_QTree_Int) */
  assign dconReadIn_QTree_Int_d = ReadIn_QTree_Int_dc((& {destructReadIn_QTree_Int_d[0]}), destructReadIn_QTree_Int_d);
  assign {destructReadIn_QTree_Int_r} = {1 {(dconReadIn_QTree_Int_r && dconReadIn_QTree_Int_d[0])}};
  
  /* destruct (Ty MemOut_QTree_Int,
          Dcon ReadOut_QTree_Int) : (memReadOut_QTree_Int,MemOut_QTree_Int) > [(destructReadOut_QTree_Int,QTree_Int)] */
  assign destructReadOut_QTree_Int_d = {memReadOut_QTree_Int_d[67:2],
                                        memReadOut_QTree_Int_d[0]};
  assign memReadOut_QTree_Int_r = destructReadOut_QTree_Int_r;
  
  /* mergectrl (Ty C38,
           Ty QTree_Int) : [(lizzieLet10_1_argbuf,QTree_Int),
                            (lizzieLet11_1_argbuf,QTree_Int),
                            (lizzieLet13_1_argbuf,QTree_Int),
                            (lizzieLet15_1_argbuf,QTree_Int),
                            (lizzieLet16_1_argbuf,QTree_Int),
                            (lizzieLet20_1_argbuf,QTree_Int),
                            (lizzieLet21_1_argbuf,QTree_Int),
                            (lizzieLet22_1_argbuf,QTree_Int),
                            (lizzieLet23_1_argbuf,QTree_Int),
                            (lizzieLet25_1_argbuf,QTree_Int),
                            (lizzieLet26_1_argbuf,QTree_Int),
                            (lizzieLet27_1_argbuf,QTree_Int),
                            (lizzieLet28_1_argbuf,QTree_Int),
                            (lizzieLet31_1_argbuf,QTree_Int),
                            (lizzieLet32_1_argbuf,QTree_Int),
                            (lizzieLet33_1_argbuf,QTree_Int),
                            (lizzieLet34_1_argbuf,QTree_Int),
                            (lizzieLet36_1_argbuf,QTree_Int),
                            (lizzieLet37_2_1_argbuf,QTree_Int),
                            (lizzieLet38_1_1_argbuf,QTree_Int),
                            (lizzieLet39_1_1_argbuf,QTree_Int),
                            (lizzieLet40_1_argbuf,QTree_Int),
                            (lizzieLet41_1_argbuf,QTree_Int),
                            (lizzieLet42_1_argbuf,QTree_Int),
                            (lizzieLet45_1_argbuf,QTree_Int),
                            (lizzieLet46_1_argbuf,QTree_Int),
                            (lizzieLet47_1_argbuf,QTree_Int),
                            (lizzieLet48_1_argbuf,QTree_Int),
                            (lizzieLet50_1_argbuf,QTree_Int),
                            (lizzieLet51_1_argbuf,QTree_Int),
                            (lizzieLet53_1_argbuf,QTree_Int),
                            (lizzieLet54_1_argbuf,QTree_Int),
                            (lizzieLet55_1_argbuf,QTree_Int),
                            (lizzieLet66_1_argbuf,QTree_Int),
                            (lizzieLet71_1_argbuf,QTree_Int),
                            (lizzieLet8_1_argbuf,QTree_Int),
                            (lizzieLet9_1_argbuf,QTree_Int),
                            (dummy_write_QTree_Int,QTree_Int)] > (writeMerge_choice_QTree_Int,C38) (writeMerge_data_QTree_Int,QTree_Int) */
  logic [37:0] lizzieLet10_1_argbuf_select_d;
  assign lizzieLet10_1_argbuf_select_d = ((| lizzieLet10_1_argbuf_select_q) ? lizzieLet10_1_argbuf_select_q :
                                          (lizzieLet10_1_argbuf_d[0] ? 38'd1 :
                                           (lizzieLet11_1_argbuf_d[0] ? 38'd2 :
                                            (lizzieLet13_1_argbuf_d[0] ? 38'd4 :
                                             (lizzieLet15_1_argbuf_d[0] ? 38'd8 :
                                              (lizzieLet16_1_argbuf_d[0] ? 38'd16 :
                                               (lizzieLet20_1_argbuf_d[0] ? 38'd32 :
                                                (lizzieLet21_1_argbuf_d[0] ? 38'd64 :
                                                 (lizzieLet22_1_argbuf_d[0] ? 38'd128 :
                                                  (lizzieLet23_1_argbuf_d[0] ? 38'd256 :
                                                   (lizzieLet25_1_argbuf_d[0] ? 38'd512 :
                                                    (lizzieLet26_1_argbuf_d[0] ? 38'd1024 :
                                                     (lizzieLet27_1_argbuf_d[0] ? 38'd2048 :
                                                      (lizzieLet28_1_argbuf_d[0] ? 38'd4096 :
                                                       (lizzieLet31_1_argbuf_d[0] ? 38'd8192 :
                                                        (lizzieLet32_1_argbuf_d[0] ? 38'd16384 :
                                                         (lizzieLet33_1_argbuf_d[0] ? 38'd32768 :
                                                          (lizzieLet34_1_argbuf_d[0] ? 38'd65536 :
                                                           (lizzieLet36_1_argbuf_d[0] ? 38'd131072 :
                                                            (lizzieLet37_2_1_argbuf_d[0] ? 38'd262144 :
                                                             (lizzieLet38_1_1_argbuf_d[0] ? 38'd524288 :
                                                              (lizzieLet39_1_1_argbuf_d[0] ? 38'd1048576 :
                                                               (lizzieLet40_1_argbuf_d[0] ? 38'd2097152 :
                                                                (lizzieLet41_1_argbuf_d[0] ? 38'd4194304 :
                                                                 (lizzieLet42_1_argbuf_d[0] ? 38'd8388608 :
                                                                  (lizzieLet45_1_argbuf_d[0] ? 38'd16777216 :
                                                                   (lizzieLet46_1_argbuf_d[0] ? 38'd33554432 :
                                                                    (lizzieLet47_1_argbuf_d[0] ? 38'd67108864 :
                                                                     (lizzieLet48_1_argbuf_d[0] ? 38'd134217728 :
                                                                      (lizzieLet50_1_argbuf_d[0] ? 38'd268435456 :
                                                                       (lizzieLet51_1_argbuf_d[0] ? 38'd536870912 :
                                                                        (lizzieLet53_1_argbuf_d[0] ? 38'd1073741824 :
                                                                         (lizzieLet54_1_argbuf_d[0] ? 38'd2147483648 :
                                                                          (lizzieLet55_1_argbuf_d[0] ? 38'd4294967296 :
                                                                           (lizzieLet66_1_argbuf_d[0] ? 38'd8589934592 :
                                                                            (lizzieLet71_1_argbuf_d[0] ? 38'd17179869184 :
                                                                             (lizzieLet8_1_argbuf_d[0] ? 38'd34359738368 :
                                                                              (lizzieLet9_1_argbuf_d[0] ? 38'd68719476736 :
                                                                               (dummy_write_QTree_Int_d[0] ? 38'd137438953472 :
                                                                                38'd0)))))))))))))))))))))))))))))))))))))));
  logic [37:0] lizzieLet10_1_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet10_1_argbuf_select_q <= 38'd0;
    else
      lizzieLet10_1_argbuf_select_q <= (lizzieLet10_1_argbuf_done ? 38'd0 :
                                        lizzieLet10_1_argbuf_select_d);
  logic [1:0] lizzieLet10_1_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet10_1_argbuf_emit_q <= 2'd0;
    else
      lizzieLet10_1_argbuf_emit_q <= (lizzieLet10_1_argbuf_done ? 2'd0 :
                                      lizzieLet10_1_argbuf_emit_d);
  logic [1:0] lizzieLet10_1_argbuf_emit_d;
  assign lizzieLet10_1_argbuf_emit_d = (lizzieLet10_1_argbuf_emit_q | ({writeMerge_choice_QTree_Int_d[0],
                                                                        writeMerge_data_QTree_Int_d[0]} & {writeMerge_choice_QTree_Int_r,
                                                                                                           writeMerge_data_QTree_Int_r}));
  logic lizzieLet10_1_argbuf_done;
  assign lizzieLet10_1_argbuf_done = (& lizzieLet10_1_argbuf_emit_d);
  assign {dummy_write_QTree_Int_r,
          lizzieLet9_1_argbuf_r,
          lizzieLet8_1_argbuf_r,
          lizzieLet71_1_argbuf_r,
          lizzieLet66_1_argbuf_r,
          lizzieLet55_1_argbuf_r,
          lizzieLet54_1_argbuf_r,
          lizzieLet53_1_argbuf_r,
          lizzieLet51_1_argbuf_r,
          lizzieLet50_1_argbuf_r,
          lizzieLet48_1_argbuf_r,
          lizzieLet47_1_argbuf_r,
          lizzieLet46_1_argbuf_r,
          lizzieLet45_1_argbuf_r,
          lizzieLet42_1_argbuf_r,
          lizzieLet41_1_argbuf_r,
          lizzieLet40_1_argbuf_r,
          lizzieLet39_1_1_argbuf_r,
          lizzieLet38_1_1_argbuf_r,
          lizzieLet37_2_1_argbuf_r,
          lizzieLet36_1_argbuf_r,
          lizzieLet34_1_argbuf_r,
          lizzieLet33_1_argbuf_r,
          lizzieLet32_1_argbuf_r,
          lizzieLet31_1_argbuf_r,
          lizzieLet28_1_argbuf_r,
          lizzieLet27_1_argbuf_r,
          lizzieLet26_1_argbuf_r,
          lizzieLet25_1_argbuf_r,
          lizzieLet23_1_argbuf_r,
          lizzieLet22_1_argbuf_r,
          lizzieLet21_1_argbuf_r,
          lizzieLet20_1_argbuf_r,
          lizzieLet16_1_argbuf_r,
          lizzieLet15_1_argbuf_r,
          lizzieLet13_1_argbuf_r,
          lizzieLet11_1_argbuf_r,
          lizzieLet10_1_argbuf_r} = (lizzieLet10_1_argbuf_done ? lizzieLet10_1_argbuf_select_d :
                                     38'd0);
  assign writeMerge_data_QTree_Int_d = ((lizzieLet10_1_argbuf_select_d[0] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet10_1_argbuf_d :
                                        ((lizzieLet10_1_argbuf_select_d[1] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet11_1_argbuf_d :
                                         ((lizzieLet10_1_argbuf_select_d[2] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet13_1_argbuf_d :
                                          ((lizzieLet10_1_argbuf_select_d[3] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet15_1_argbuf_d :
                                           ((lizzieLet10_1_argbuf_select_d[4] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet16_1_argbuf_d :
                                            ((lizzieLet10_1_argbuf_select_d[5] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet20_1_argbuf_d :
                                             ((lizzieLet10_1_argbuf_select_d[6] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet21_1_argbuf_d :
                                              ((lizzieLet10_1_argbuf_select_d[7] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet22_1_argbuf_d :
                                               ((lizzieLet10_1_argbuf_select_d[8] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet23_1_argbuf_d :
                                                ((lizzieLet10_1_argbuf_select_d[9] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet25_1_argbuf_d :
                                                 ((lizzieLet10_1_argbuf_select_d[10] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet26_1_argbuf_d :
                                                  ((lizzieLet10_1_argbuf_select_d[11] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet27_1_argbuf_d :
                                                   ((lizzieLet10_1_argbuf_select_d[12] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet28_1_argbuf_d :
                                                    ((lizzieLet10_1_argbuf_select_d[13] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet31_1_argbuf_d :
                                                     ((lizzieLet10_1_argbuf_select_d[14] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet32_1_argbuf_d :
                                                      ((lizzieLet10_1_argbuf_select_d[15] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet33_1_argbuf_d :
                                                       ((lizzieLet10_1_argbuf_select_d[16] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet34_1_argbuf_d :
                                                        ((lizzieLet10_1_argbuf_select_d[17] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet36_1_argbuf_d :
                                                         ((lizzieLet10_1_argbuf_select_d[18] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet37_2_1_argbuf_d :
                                                          ((lizzieLet10_1_argbuf_select_d[19] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet38_1_1_argbuf_d :
                                                           ((lizzieLet10_1_argbuf_select_d[20] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet39_1_1_argbuf_d :
                                                            ((lizzieLet10_1_argbuf_select_d[21] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet40_1_argbuf_d :
                                                             ((lizzieLet10_1_argbuf_select_d[22] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet41_1_argbuf_d :
                                                              ((lizzieLet10_1_argbuf_select_d[23] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet42_1_argbuf_d :
                                                               ((lizzieLet10_1_argbuf_select_d[24] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet45_1_argbuf_d :
                                                                ((lizzieLet10_1_argbuf_select_d[25] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet46_1_argbuf_d :
                                                                 ((lizzieLet10_1_argbuf_select_d[26] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet47_1_argbuf_d :
                                                                  ((lizzieLet10_1_argbuf_select_d[27] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet48_1_argbuf_d :
                                                                   ((lizzieLet10_1_argbuf_select_d[28] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet50_1_argbuf_d :
                                                                    ((lizzieLet10_1_argbuf_select_d[29] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet51_1_argbuf_d :
                                                                     ((lizzieLet10_1_argbuf_select_d[30] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet53_1_argbuf_d :
                                                                      ((lizzieLet10_1_argbuf_select_d[31] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet54_1_argbuf_d :
                                                                       ((lizzieLet10_1_argbuf_select_d[32] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet55_1_argbuf_d :
                                                                        ((lizzieLet10_1_argbuf_select_d[33] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet66_1_argbuf_d :
                                                                         ((lizzieLet10_1_argbuf_select_d[34] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet71_1_argbuf_d :
                                                                          ((lizzieLet10_1_argbuf_select_d[35] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet8_1_argbuf_d :
                                                                           ((lizzieLet10_1_argbuf_select_d[36] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet9_1_argbuf_d :
                                                                            ((lizzieLet10_1_argbuf_select_d[37] && (! lizzieLet10_1_argbuf_emit_q[0])) ? dummy_write_QTree_Int_d :
                                                                             {66'd0,
                                                                              1'd0}))))))))))))))))))))))))))))))))))))));
  assign writeMerge_choice_QTree_Int_d = ((lizzieLet10_1_argbuf_select_d[0] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C1_38_dc(1'd1) :
                                          ((lizzieLet10_1_argbuf_select_d[1] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C2_38_dc(1'd1) :
                                           ((lizzieLet10_1_argbuf_select_d[2] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C3_38_dc(1'd1) :
                                            ((lizzieLet10_1_argbuf_select_d[3] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C4_38_dc(1'd1) :
                                             ((lizzieLet10_1_argbuf_select_d[4] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C5_38_dc(1'd1) :
                                              ((lizzieLet10_1_argbuf_select_d[5] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C6_38_dc(1'd1) :
                                               ((lizzieLet10_1_argbuf_select_d[6] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C7_38_dc(1'd1) :
                                                ((lizzieLet10_1_argbuf_select_d[7] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C8_38_dc(1'd1) :
                                                 ((lizzieLet10_1_argbuf_select_d[8] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C9_38_dc(1'd1) :
                                                  ((lizzieLet10_1_argbuf_select_d[9] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C10_38_dc(1'd1) :
                                                   ((lizzieLet10_1_argbuf_select_d[10] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C11_38_dc(1'd1) :
                                                    ((lizzieLet10_1_argbuf_select_d[11] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C12_38_dc(1'd1) :
                                                     ((lizzieLet10_1_argbuf_select_d[12] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C13_38_dc(1'd1) :
                                                      ((lizzieLet10_1_argbuf_select_d[13] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C14_38_dc(1'd1) :
                                                       ((lizzieLet10_1_argbuf_select_d[14] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C15_38_dc(1'd1) :
                                                        ((lizzieLet10_1_argbuf_select_d[15] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C16_38_dc(1'd1) :
                                                         ((lizzieLet10_1_argbuf_select_d[16] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C17_38_dc(1'd1) :
                                                          ((lizzieLet10_1_argbuf_select_d[17] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C18_38_dc(1'd1) :
                                                           ((lizzieLet10_1_argbuf_select_d[18] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C19_38_dc(1'd1) :
                                                            ((lizzieLet10_1_argbuf_select_d[19] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C20_38_dc(1'd1) :
                                                             ((lizzieLet10_1_argbuf_select_d[20] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C21_38_dc(1'd1) :
                                                              ((lizzieLet10_1_argbuf_select_d[21] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C22_38_dc(1'd1) :
                                                               ((lizzieLet10_1_argbuf_select_d[22] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C23_38_dc(1'd1) :
                                                                ((lizzieLet10_1_argbuf_select_d[23] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C24_38_dc(1'd1) :
                                                                 ((lizzieLet10_1_argbuf_select_d[24] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C25_38_dc(1'd1) :
                                                                  ((lizzieLet10_1_argbuf_select_d[25] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C26_38_dc(1'd1) :
                                                                   ((lizzieLet10_1_argbuf_select_d[26] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C27_38_dc(1'd1) :
                                                                    ((lizzieLet10_1_argbuf_select_d[27] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C28_38_dc(1'd1) :
                                                                     ((lizzieLet10_1_argbuf_select_d[28] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C29_38_dc(1'd1) :
                                                                      ((lizzieLet10_1_argbuf_select_d[29] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C30_38_dc(1'd1) :
                                                                       ((lizzieLet10_1_argbuf_select_d[30] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C31_38_dc(1'd1) :
                                                                        ((lizzieLet10_1_argbuf_select_d[31] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C32_38_dc(1'd1) :
                                                                         ((lizzieLet10_1_argbuf_select_d[32] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C33_38_dc(1'd1) :
                                                                          ((lizzieLet10_1_argbuf_select_d[33] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C34_38_dc(1'd1) :
                                                                           ((lizzieLet10_1_argbuf_select_d[34] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C35_38_dc(1'd1) :
                                                                            ((lizzieLet10_1_argbuf_select_d[35] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C36_38_dc(1'd1) :
                                                                             ((lizzieLet10_1_argbuf_select_d[36] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C37_38_dc(1'd1) :
                                                                              ((lizzieLet10_1_argbuf_select_d[37] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C38_38_dc(1'd1) :
                                                                               {6'd0,
                                                                                1'd0}))))))))))))))))))))))))))))))))))))));
  
  /* demux (Ty C38,
       Ty Pointer_QTree_Int) : (writeMerge_choice_QTree_Int,C38) (demuxWriteResult_QTree_Int,Pointer_QTree_Int) > [(writeQTree_IntlizzieLet10_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet11_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet13_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet15_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet16_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet20_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet21_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet22_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet23_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet25_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet26_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet27_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet28_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet31_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet32_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet33_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet34_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet36_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet37_2_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet38_1_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet39_1_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet40_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet41_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet42_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet45_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet46_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet47_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet48_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet50_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet51_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet53_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet54_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet55_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet66_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet71_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet8_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet9_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (dummy_write_QTree_Int_sink,Pointer_QTree_Int)] */
  logic [37:0] demuxWriteResult_QTree_Int_onehotd;
  always_comb
    if ((writeMerge_choice_QTree_Int_d[0] && demuxWriteResult_QTree_Int_d[0]))
      unique case (writeMerge_choice_QTree_Int_d[6:1])
        6'd0: demuxWriteResult_QTree_Int_onehotd = 38'd1;
        6'd1: demuxWriteResult_QTree_Int_onehotd = 38'd2;
        6'd2: demuxWriteResult_QTree_Int_onehotd = 38'd4;
        6'd3: demuxWriteResult_QTree_Int_onehotd = 38'd8;
        6'd4: demuxWriteResult_QTree_Int_onehotd = 38'd16;
        6'd5: demuxWriteResult_QTree_Int_onehotd = 38'd32;
        6'd6: demuxWriteResult_QTree_Int_onehotd = 38'd64;
        6'd7: demuxWriteResult_QTree_Int_onehotd = 38'd128;
        6'd8: demuxWriteResult_QTree_Int_onehotd = 38'd256;
        6'd9: demuxWriteResult_QTree_Int_onehotd = 38'd512;
        6'd10: demuxWriteResult_QTree_Int_onehotd = 38'd1024;
        6'd11: demuxWriteResult_QTree_Int_onehotd = 38'd2048;
        6'd12: demuxWriteResult_QTree_Int_onehotd = 38'd4096;
        6'd13: demuxWriteResult_QTree_Int_onehotd = 38'd8192;
        6'd14: demuxWriteResult_QTree_Int_onehotd = 38'd16384;
        6'd15: demuxWriteResult_QTree_Int_onehotd = 38'd32768;
        6'd16: demuxWriteResult_QTree_Int_onehotd = 38'd65536;
        6'd17: demuxWriteResult_QTree_Int_onehotd = 38'd131072;
        6'd18: demuxWriteResult_QTree_Int_onehotd = 38'd262144;
        6'd19: demuxWriteResult_QTree_Int_onehotd = 38'd524288;
        6'd20: demuxWriteResult_QTree_Int_onehotd = 38'd1048576;
        6'd21: demuxWriteResult_QTree_Int_onehotd = 38'd2097152;
        6'd22: demuxWriteResult_QTree_Int_onehotd = 38'd4194304;
        6'd23: demuxWriteResult_QTree_Int_onehotd = 38'd8388608;
        6'd24: demuxWriteResult_QTree_Int_onehotd = 38'd16777216;
        6'd25: demuxWriteResult_QTree_Int_onehotd = 38'd33554432;
        6'd26: demuxWriteResult_QTree_Int_onehotd = 38'd67108864;
        6'd27: demuxWriteResult_QTree_Int_onehotd = 38'd134217728;
        6'd28: demuxWriteResult_QTree_Int_onehotd = 38'd268435456;
        6'd29: demuxWriteResult_QTree_Int_onehotd = 38'd536870912;
        6'd30: demuxWriteResult_QTree_Int_onehotd = 38'd1073741824;
        6'd31: demuxWriteResult_QTree_Int_onehotd = 38'd2147483648;
        6'd32: demuxWriteResult_QTree_Int_onehotd = 38'd4294967296;
        6'd33: demuxWriteResult_QTree_Int_onehotd = 38'd8589934592;
        6'd34: demuxWriteResult_QTree_Int_onehotd = 38'd17179869184;
        6'd35: demuxWriteResult_QTree_Int_onehotd = 38'd34359738368;
        6'd36: demuxWriteResult_QTree_Int_onehotd = 38'd68719476736;
        6'd37: demuxWriteResult_QTree_Int_onehotd = 38'd137438953472;
        default: demuxWriteResult_QTree_Int_onehotd = 38'd0;
      endcase
    else demuxWriteResult_QTree_Int_onehotd = 38'd0;
  assign writeQTree_IntlizzieLet10_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                 demuxWriteResult_QTree_Int_onehotd[0]};
  assign writeQTree_IntlizzieLet11_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                 demuxWriteResult_QTree_Int_onehotd[1]};
  assign writeQTree_IntlizzieLet13_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                 demuxWriteResult_QTree_Int_onehotd[2]};
  assign writeQTree_IntlizzieLet15_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                 demuxWriteResult_QTree_Int_onehotd[3]};
  assign writeQTree_IntlizzieLet16_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                 demuxWriteResult_QTree_Int_onehotd[4]};
  assign writeQTree_IntlizzieLet20_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                 demuxWriteResult_QTree_Int_onehotd[5]};
  assign writeQTree_IntlizzieLet21_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                 demuxWriteResult_QTree_Int_onehotd[6]};
  assign writeQTree_IntlizzieLet22_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                 demuxWriteResult_QTree_Int_onehotd[7]};
  assign writeQTree_IntlizzieLet23_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                 demuxWriteResult_QTree_Int_onehotd[8]};
  assign writeQTree_IntlizzieLet25_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                 demuxWriteResult_QTree_Int_onehotd[9]};
  assign writeQTree_IntlizzieLet26_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                 demuxWriteResult_QTree_Int_onehotd[10]};
  assign writeQTree_IntlizzieLet27_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                 demuxWriteResult_QTree_Int_onehotd[11]};
  assign writeQTree_IntlizzieLet28_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                 demuxWriteResult_QTree_Int_onehotd[12]};
  assign writeQTree_IntlizzieLet31_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                 demuxWriteResult_QTree_Int_onehotd[13]};
  assign writeQTree_IntlizzieLet32_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                 demuxWriteResult_QTree_Int_onehotd[14]};
  assign writeQTree_IntlizzieLet33_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                 demuxWriteResult_QTree_Int_onehotd[15]};
  assign writeQTree_IntlizzieLet34_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                 demuxWriteResult_QTree_Int_onehotd[16]};
  assign writeQTree_IntlizzieLet36_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                 demuxWriteResult_QTree_Int_onehotd[17]};
  assign writeQTree_IntlizzieLet37_2_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                   demuxWriteResult_QTree_Int_onehotd[18]};
  assign writeQTree_IntlizzieLet38_1_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                   demuxWriteResult_QTree_Int_onehotd[19]};
  assign writeQTree_IntlizzieLet39_1_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                   demuxWriteResult_QTree_Int_onehotd[20]};
  assign writeQTree_IntlizzieLet40_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                 demuxWriteResult_QTree_Int_onehotd[21]};
  assign writeQTree_IntlizzieLet41_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                 demuxWriteResult_QTree_Int_onehotd[22]};
  assign writeQTree_IntlizzieLet42_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                 demuxWriteResult_QTree_Int_onehotd[23]};
  assign writeQTree_IntlizzieLet45_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                 demuxWriteResult_QTree_Int_onehotd[24]};
  assign writeQTree_IntlizzieLet46_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                 demuxWriteResult_QTree_Int_onehotd[25]};
  assign writeQTree_IntlizzieLet47_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                 demuxWriteResult_QTree_Int_onehotd[26]};
  assign writeQTree_IntlizzieLet48_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                 demuxWriteResult_QTree_Int_onehotd[27]};
  assign writeQTree_IntlizzieLet50_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                 demuxWriteResult_QTree_Int_onehotd[28]};
  assign writeQTree_IntlizzieLet51_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                 demuxWriteResult_QTree_Int_onehotd[29]};
  assign writeQTree_IntlizzieLet53_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                 demuxWriteResult_QTree_Int_onehotd[30]};
  assign writeQTree_IntlizzieLet54_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                 demuxWriteResult_QTree_Int_onehotd[31]};
  assign writeQTree_IntlizzieLet55_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                 demuxWriteResult_QTree_Int_onehotd[32]};
  assign writeQTree_IntlizzieLet66_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                 demuxWriteResult_QTree_Int_onehotd[33]};
  assign writeQTree_IntlizzieLet71_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                 demuxWriteResult_QTree_Int_onehotd[34]};
  assign writeQTree_IntlizzieLet8_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                demuxWriteResult_QTree_Int_onehotd[35]};
  assign writeQTree_IntlizzieLet9_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                demuxWriteResult_QTree_Int_onehotd[36]};
  assign dummy_write_QTree_Int_sink_d = {demuxWriteResult_QTree_Int_d[16:1],
                                         demuxWriteResult_QTree_Int_onehotd[37]};
  assign demuxWriteResult_QTree_Int_r = (| (demuxWriteResult_QTree_Int_onehotd & {dummy_write_QTree_Int_sink_r,
                                                                                  writeQTree_IntlizzieLet9_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet8_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet71_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet66_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet55_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet54_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet53_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet51_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet50_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet48_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet47_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet46_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet45_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet42_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet41_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet40_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet39_1_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet38_1_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet37_2_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet36_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet34_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet33_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet32_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet31_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet28_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet27_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet26_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet25_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet23_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet22_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet21_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet20_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet16_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet15_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet13_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet11_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet10_1_argbuf_r}));
  assign writeMerge_choice_QTree_Int_r = demuxWriteResult_QTree_Int_r;
  
  /* dcon (Ty MemIn_QTree_Int,
      Dcon WriteIn_QTree_Int) : [(forkHP1_QTree_In3,Word16#),
                                 (writeMerge_data_QTree_Int,QTree_Int)] > (dconWriteIn_QTree_Int,MemIn_QTree_Int) */
  assign dconWriteIn_QTree_Int_d = WriteIn_QTree_Int_dc((& {forkHP1_QTree_In3_d[0],
                                                            writeMerge_data_QTree_Int_d[0]}), forkHP1_QTree_In3_d, writeMerge_data_QTree_Int_d);
  assign {forkHP1_QTree_In3_r,
          writeMerge_data_QTree_Int_r} = {2 {(dconWriteIn_QTree_Int_r && dconWriteIn_QTree_Int_d[0])}};
  
  /* dcon (Ty Pointer_QTree_Int,
      Dcon Pointer_QTree_Int) : [(forkHP1_QTree_In4,Word16#)] > (dconPtr_QTree_Int,Pointer_QTree_Int) */
  assign dconPtr_QTree_Int_d = Pointer_QTree_Int_dc((& {forkHP1_QTree_In4_d[0]}), forkHP1_QTree_In4_d);
  assign {forkHP1_QTree_In4_r} = {1 {(dconPtr_QTree_Int_r && dconPtr_QTree_Int_d[0])}};
  
  /* demux (Ty MemOut_QTree_Int,
       Ty Pointer_QTree_Int) : (memWriteOut_QTree_Int,MemOut_QTree_Int) (dconPtr_QTree_Int,Pointer_QTree_Int) > [(_258,Pointer_QTree_Int),
                                                                                                                 (demuxWriteResult_QTree_Int,Pointer_QTree_Int)] */
  logic [1:0] dconPtr_QTree_Int_onehotd;
  always_comb
    if ((memWriteOut_QTree_Int_d[0] && dconPtr_QTree_Int_d[0]))
      unique case (memWriteOut_QTree_Int_d[1:1])
        1'd0: dconPtr_QTree_Int_onehotd = 2'd1;
        1'd1: dconPtr_QTree_Int_onehotd = 2'd2;
        default: dconPtr_QTree_Int_onehotd = 2'd0;
      endcase
    else dconPtr_QTree_Int_onehotd = 2'd0;
  assign _258_d = {dconPtr_QTree_Int_d[16:1],
                   dconPtr_QTree_Int_onehotd[0]};
  assign demuxWriteResult_QTree_Int_d = {dconPtr_QTree_Int_d[16:1],
                                         dconPtr_QTree_Int_onehotd[1]};
  assign dconPtr_QTree_Int_r = (| (dconPtr_QTree_Int_onehotd & {demuxWriteResult_QTree_Int_r,
                                                                _258_r}));
  assign memWriteOut_QTree_Int_r = dconPtr_QTree_Int_r;
  
  /* const (Ty Word16#,
       Lit 0) : (go__7,Go) > (initHP_CTf''''''''''''_f''''''''''''_Int,Word16#) */
  assign \initHP_CTf''''''''''''_f''''''''''''_Int_d  = {16'd0,
                                                         go__7_d[0]};
  assign go__7_r = \initHP_CTf''''''''''''_f''''''''''''_Int_r ;
  
  /* const (Ty Word16#,
       Lit 1) : (incrHP_CTf''''''''''''_f''''''''''''_Int1,Go) > (incrHP_CTf''''''''''''_f''''''''''''_Int,Word16#) */
  assign \incrHP_CTf''''''''''''_f''''''''''''_Int_d  = {16'd1,
                                                         \incrHP_CTf''''''''''''_f''''''''''''_Int1_d [0]};
  assign \incrHP_CTf''''''''''''_f''''''''''''_Int1_r  = \incrHP_CTf''''''''''''_f''''''''''''_Int_r ;
  
  /* merge (Ty Go) : [(go__8,Go),
                 (incrHP_CTf''''''''''''_f''''''''''''_Int2,Go)] > (incrHP_mergeCTf''''''''''''_f''''''''''''_Int,Go) */
  logic [1:0] \incrHP_mergeCTf''''''''''''_f''''''''''''_Int_selected ;
  logic [1:0] \incrHP_mergeCTf''''''''''''_f''''''''''''_Int_select ;
  always_comb
    begin
      \incrHP_mergeCTf''''''''''''_f''''''''''''_Int_selected  = 2'd0;
      if ((| \incrHP_mergeCTf''''''''''''_f''''''''''''_Int_select ))
        \incrHP_mergeCTf''''''''''''_f''''''''''''_Int_selected  = \incrHP_mergeCTf''''''''''''_f''''''''''''_Int_select ;
      else
        if (go__8_d[0])
          \incrHP_mergeCTf''''''''''''_f''''''''''''_Int_selected [0] = 1'd1;
        else if (\incrHP_CTf''''''''''''_f''''''''''''_Int2_d [0])
          \incrHP_mergeCTf''''''''''''_f''''''''''''_Int_selected [1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \incrHP_mergeCTf''''''''''''_f''''''''''''_Int_select  <= 2'd0;
    else
      \incrHP_mergeCTf''''''''''''_f''''''''''''_Int_select  <= (\incrHP_mergeCTf''''''''''''_f''''''''''''_Int_r  ? 2'd0 :
                                                                 \incrHP_mergeCTf''''''''''''_f''''''''''''_Int_selected );
  always_comb
    if (\incrHP_mergeCTf''''''''''''_f''''''''''''_Int_selected [0])
      \incrHP_mergeCTf''''''''''''_f''''''''''''_Int_d  = go__8_d;
    else if (\incrHP_mergeCTf''''''''''''_f''''''''''''_Int_selected [1])
      \incrHP_mergeCTf''''''''''''_f''''''''''''_Int_d  = \incrHP_CTf''''''''''''_f''''''''''''_Int2_d ;
    else \incrHP_mergeCTf''''''''''''_f''''''''''''_Int_d  = 1'd0;
  assign {\incrHP_CTf''''''''''''_f''''''''''''_Int2_r ,
          go__8_r} = (\incrHP_mergeCTf''''''''''''_f''''''''''''_Int_r  ? \incrHP_mergeCTf''''''''''''_f''''''''''''_Int_selected  :
                      2'd0);
  
  /* fork (Ty Go) : (incrHP_mergeCTf''''''''''''_f''''''''''''_Int_buf,Go) > [(incrHP_CTf''''''''''''_f''''''''''''_Int1,Go),
                                                                         (incrHP_CTf''''''''''''_f''''''''''''_Int2,Go)] */
  logic [1:0] \incrHP_mergeCTf''''''''''''_f''''''''''''_Int_buf_emitted ;
  logic [1:0] \incrHP_mergeCTf''''''''''''_f''''''''''''_Int_buf_done ;
  assign \incrHP_CTf''''''''''''_f''''''''''''_Int1_d  = (\incrHP_mergeCTf''''''''''''_f''''''''''''_Int_buf_d [0] && (! \incrHP_mergeCTf''''''''''''_f''''''''''''_Int_buf_emitted [0]));
  assign \incrHP_CTf''''''''''''_f''''''''''''_Int2_d  = (\incrHP_mergeCTf''''''''''''_f''''''''''''_Int_buf_d [0] && (! \incrHP_mergeCTf''''''''''''_f''''''''''''_Int_buf_emitted [1]));
  assign \incrHP_mergeCTf''''''''''''_f''''''''''''_Int_buf_done  = (\incrHP_mergeCTf''''''''''''_f''''''''''''_Int_buf_emitted  | ({\incrHP_CTf''''''''''''_f''''''''''''_Int2_d [0],
                                                                                                                                     \incrHP_CTf''''''''''''_f''''''''''''_Int1_d [0]} & {\incrHP_CTf''''''''''''_f''''''''''''_Int2_r ,
                                                                                                                                                                                          \incrHP_CTf''''''''''''_f''''''''''''_Int1_r }));
  assign \incrHP_mergeCTf''''''''''''_f''''''''''''_Int_buf_r  = (& \incrHP_mergeCTf''''''''''''_f''''''''''''_Int_buf_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \incrHP_mergeCTf''''''''''''_f''''''''''''_Int_buf_emitted  <= 2'd0;
    else
      \incrHP_mergeCTf''''''''''''_f''''''''''''_Int_buf_emitted  <= (\incrHP_mergeCTf''''''''''''_f''''''''''''_Int_buf_r  ? 2'd0 :
                                                                      \incrHP_mergeCTf''''''''''''_f''''''''''''_Int_buf_done );
  
  /* op_add (Ty Word16#) : (incrHP_CTf''''''''''''_f''''''''''''_Int,Word16#) (forkHP1_CTf''''''''''''_f''''''''''''_Int,Word16#) > (addHP_CTf''''''''''''_f''''''''''''_Int,Word16#) */
  assign \addHP_CTf''''''''''''_f''''''''''''_Int_d  = {(\incrHP_CTf''''''''''''_f''''''''''''_Int_d [16:1] + \forkHP1_CTf''''''''''''_f''''''''''''_Int_d [16:1]),
                                                        (\incrHP_CTf''''''''''''_f''''''''''''_Int_d [0] && \forkHP1_CTf''''''''''''_f''''''''''''_Int_d [0])};
  assign {\incrHP_CTf''''''''''''_f''''''''''''_Int_r ,
          \forkHP1_CTf''''''''''''_f''''''''''''_Int_r } = {2 {(\addHP_CTf''''''''''''_f''''''''''''_Int_r  && \addHP_CTf''''''''''''_f''''''''''''_Int_d [0])}};
  
  /* merge (Ty Word16#) : [(initHP_CTf''''''''''''_f''''''''''''_Int,Word16#),
                      (addHP_CTf''''''''''''_f''''''''''''_Int,Word16#)] > (mergeHP_CTf''''''''''''_f''''''''''''_Int,Word16#) */
  logic [1:0] \mergeHP_CTf''''''''''''_f''''''''''''_Int_selected ;
  logic [1:0] \mergeHP_CTf''''''''''''_f''''''''''''_Int_select ;
  always_comb
    begin
      \mergeHP_CTf''''''''''''_f''''''''''''_Int_selected  = 2'd0;
      if ((| \mergeHP_CTf''''''''''''_f''''''''''''_Int_select ))
        \mergeHP_CTf''''''''''''_f''''''''''''_Int_selected  = \mergeHP_CTf''''''''''''_f''''''''''''_Int_select ;
      else
        if (\initHP_CTf''''''''''''_f''''''''''''_Int_d [0])
          \mergeHP_CTf''''''''''''_f''''''''''''_Int_selected [0] = 1'd1;
        else if (\addHP_CTf''''''''''''_f''''''''''''_Int_d [0])
          \mergeHP_CTf''''''''''''_f''''''''''''_Int_selected [1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \mergeHP_CTf''''''''''''_f''''''''''''_Int_select  <= 2'd0;
    else
      \mergeHP_CTf''''''''''''_f''''''''''''_Int_select  <= (\mergeHP_CTf''''''''''''_f''''''''''''_Int_r  ? 2'd0 :
                                                             \mergeHP_CTf''''''''''''_f''''''''''''_Int_selected );
  always_comb
    if (\mergeHP_CTf''''''''''''_f''''''''''''_Int_selected [0])
      \mergeHP_CTf''''''''''''_f''''''''''''_Int_d  = \initHP_CTf''''''''''''_f''''''''''''_Int_d ;
    else if (\mergeHP_CTf''''''''''''_f''''''''''''_Int_selected [1])
      \mergeHP_CTf''''''''''''_f''''''''''''_Int_d  = \addHP_CTf''''''''''''_f''''''''''''_Int_d ;
    else \mergeHP_CTf''''''''''''_f''''''''''''_Int_d  = {16'd0, 1'd0};
  assign {\addHP_CTf''''''''''''_f''''''''''''_Int_r ,
          \initHP_CTf''''''''''''_f''''''''''''_Int_r } = (\mergeHP_CTf''''''''''''_f''''''''''''_Int_r  ? \mergeHP_CTf''''''''''''_f''''''''''''_Int_selected  :
                                                           2'd0);
  
  /* buf (Ty Go) : (incrHP_mergeCTf''''''''''''_f''''''''''''_Int,Go) > (incrHP_mergeCTf''''''''''''_f''''''''''''_Int_buf,Go) */
  Go_t \incrHP_mergeCTf''''''''''''_f''''''''''''_Int_bufchan_d ;
  logic \incrHP_mergeCTf''''''''''''_f''''''''''''_Int_bufchan_r ;
  assign \incrHP_mergeCTf''''''''''''_f''''''''''''_Int_r  = ((! \incrHP_mergeCTf''''''''''''_f''''''''''''_Int_bufchan_d [0]) || \incrHP_mergeCTf''''''''''''_f''''''''''''_Int_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \incrHP_mergeCTf''''''''''''_f''''''''''''_Int_bufchan_d  <= 1'd0;
    else
      if (\incrHP_mergeCTf''''''''''''_f''''''''''''_Int_r )
        \incrHP_mergeCTf''''''''''''_f''''''''''''_Int_bufchan_d  <= \incrHP_mergeCTf''''''''''''_f''''''''''''_Int_d ;
  Go_t \incrHP_mergeCTf''''''''''''_f''''''''''''_Int_bufchan_buf ;
  assign \incrHP_mergeCTf''''''''''''_f''''''''''''_Int_bufchan_r  = (! \incrHP_mergeCTf''''''''''''_f''''''''''''_Int_bufchan_buf [0]);
  assign \incrHP_mergeCTf''''''''''''_f''''''''''''_Int_buf_d  = (\incrHP_mergeCTf''''''''''''_f''''''''''''_Int_bufchan_buf [0] ? \incrHP_mergeCTf''''''''''''_f''''''''''''_Int_bufchan_buf  :
                                                                  \incrHP_mergeCTf''''''''''''_f''''''''''''_Int_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \incrHP_mergeCTf''''''''''''_f''''''''''''_Int_bufchan_buf  <= 1'd0;
    else
      if ((\incrHP_mergeCTf''''''''''''_f''''''''''''_Int_buf_r  && \incrHP_mergeCTf''''''''''''_f''''''''''''_Int_bufchan_buf [0]))
        \incrHP_mergeCTf''''''''''''_f''''''''''''_Int_bufchan_buf  <= 1'd0;
      else if (((! \incrHP_mergeCTf''''''''''''_f''''''''''''_Int_buf_r ) && (! \incrHP_mergeCTf''''''''''''_f''''''''''''_Int_bufchan_buf [0])))
        \incrHP_mergeCTf''''''''''''_f''''''''''''_Int_bufchan_buf  <= \incrHP_mergeCTf''''''''''''_f''''''''''''_Int_bufchan_d ;
  
  /* buf (Ty Word16#) : (mergeHP_CTf''''''''''''_f''''''''''''_Int,Word16#) > (mergeHP_CTf''''''''''''_f''''''''''''_Int_buf,Word16#) */
  \Word16#_t  \mergeHP_CTf''''''''''''_f''''''''''''_Int_bufchan_d ;
  logic \mergeHP_CTf''''''''''''_f''''''''''''_Int_bufchan_r ;
  assign \mergeHP_CTf''''''''''''_f''''''''''''_Int_r  = ((! \mergeHP_CTf''''''''''''_f''''''''''''_Int_bufchan_d [0]) || \mergeHP_CTf''''''''''''_f''''''''''''_Int_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \mergeHP_CTf''''''''''''_f''''''''''''_Int_bufchan_d  <= {16'd0,
                                                                1'd0};
    else
      if (\mergeHP_CTf''''''''''''_f''''''''''''_Int_r )
        \mergeHP_CTf''''''''''''_f''''''''''''_Int_bufchan_d  <= \mergeHP_CTf''''''''''''_f''''''''''''_Int_d ;
  \Word16#_t  \mergeHP_CTf''''''''''''_f''''''''''''_Int_bufchan_buf ;
  assign \mergeHP_CTf''''''''''''_f''''''''''''_Int_bufchan_r  = (! \mergeHP_CTf''''''''''''_f''''''''''''_Int_bufchan_buf [0]);
  assign \mergeHP_CTf''''''''''''_f''''''''''''_Int_buf_d  = (\mergeHP_CTf''''''''''''_f''''''''''''_Int_bufchan_buf [0] ? \mergeHP_CTf''''''''''''_f''''''''''''_Int_bufchan_buf  :
                                                              \mergeHP_CTf''''''''''''_f''''''''''''_Int_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \mergeHP_CTf''''''''''''_f''''''''''''_Int_bufchan_buf  <= {16'd0,
                                                                  1'd0};
    else
      if ((\mergeHP_CTf''''''''''''_f''''''''''''_Int_buf_r  && \mergeHP_CTf''''''''''''_f''''''''''''_Int_bufchan_buf [0]))
        \mergeHP_CTf''''''''''''_f''''''''''''_Int_bufchan_buf  <= {16'd0,
                                                                    1'd0};
      else if (((! \mergeHP_CTf''''''''''''_f''''''''''''_Int_buf_r ) && (! \mergeHP_CTf''''''''''''_f''''''''''''_Int_bufchan_buf [0])))
        \mergeHP_CTf''''''''''''_f''''''''''''_Int_bufchan_buf  <= \mergeHP_CTf''''''''''''_f''''''''''''_Int_bufchan_d ;
  
  /* fork (Ty Word16#) : (mergeHP_CTf''''''''''''_f''''''''''''_Int_buf,Word16#) > [(forkHP1_CTf''''''''''''_f''''''''''''_Int,Word16#),
                                                                               (forkHP1_CTf''''''''''''_f''''''''''''_In2,Word16#),
                                                                               (forkHP1_CTf''''''''''''_f''''''''''''_In3,Word16#)] */
  logic [2:0] \mergeHP_CTf''''''''''''_f''''''''''''_Int_buf_emitted ;
  logic [2:0] \mergeHP_CTf''''''''''''_f''''''''''''_Int_buf_done ;
  assign \forkHP1_CTf''''''''''''_f''''''''''''_Int_d  = {\mergeHP_CTf''''''''''''_f''''''''''''_Int_buf_d [16:1],
                                                          (\mergeHP_CTf''''''''''''_f''''''''''''_Int_buf_d [0] && (! \mergeHP_CTf''''''''''''_f''''''''''''_Int_buf_emitted [0]))};
  assign \forkHP1_CTf''''''''''''_f''''''''''''_In2_d  = {\mergeHP_CTf''''''''''''_f''''''''''''_Int_buf_d [16:1],
                                                          (\mergeHP_CTf''''''''''''_f''''''''''''_Int_buf_d [0] && (! \mergeHP_CTf''''''''''''_f''''''''''''_Int_buf_emitted [1]))};
  assign \forkHP1_CTf''''''''''''_f''''''''''''_In3_d  = {\mergeHP_CTf''''''''''''_f''''''''''''_Int_buf_d [16:1],
                                                          (\mergeHP_CTf''''''''''''_f''''''''''''_Int_buf_d [0] && (! \mergeHP_CTf''''''''''''_f''''''''''''_Int_buf_emitted [2]))};
  assign \mergeHP_CTf''''''''''''_f''''''''''''_Int_buf_done  = (\mergeHP_CTf''''''''''''_f''''''''''''_Int_buf_emitted  | ({\forkHP1_CTf''''''''''''_f''''''''''''_In3_d [0],
                                                                                                                             \forkHP1_CTf''''''''''''_f''''''''''''_In2_d [0],
                                                                                                                             \forkHP1_CTf''''''''''''_f''''''''''''_Int_d [0]} & {\forkHP1_CTf''''''''''''_f''''''''''''_In3_r ,
                                                                                                                                                                                  \forkHP1_CTf''''''''''''_f''''''''''''_In2_r ,
                                                                                                                                                                                  \forkHP1_CTf''''''''''''_f''''''''''''_Int_r }));
  assign \mergeHP_CTf''''''''''''_f''''''''''''_Int_buf_r  = (& \mergeHP_CTf''''''''''''_f''''''''''''_Int_buf_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \mergeHP_CTf''''''''''''_f''''''''''''_Int_buf_emitted  <= 3'd0;
    else
      \mergeHP_CTf''''''''''''_f''''''''''''_Int_buf_emitted  <= (\mergeHP_CTf''''''''''''_f''''''''''''_Int_buf_r  ? 3'd0 :
                                                                  \mergeHP_CTf''''''''''''_f''''''''''''_Int_buf_done );
  
  /* mergectrl (Ty C2,
           Ty MemIn_CTf''''''''''''_f''''''''''''_Int) : [(dconReadIn_CTf''''''''''''_f''''''''''''_Int,MemIn_CTf''''''''''''_f''''''''''''_Int),
                                                          (dconWriteIn_CTf''''''''''''_f''''''''''''_Int,MemIn_CTf''''''''''''_f''''''''''''_Int)] > (memMergeChoice_CTf''''''''''''_f''''''''''''_Int,C2) (memMergeIn_CTf''''''''''''_f''''''''''''_Int,MemIn_CTf''''''''''''_f''''''''''''_Int) */
  logic [1:0] \dconReadIn_CTf''''''''''''_f''''''''''''_Int_select_d ;
  assign \dconReadIn_CTf''''''''''''_f''''''''''''_Int_select_d  = ((| \dconReadIn_CTf''''''''''''_f''''''''''''_Int_select_q ) ? \dconReadIn_CTf''''''''''''_f''''''''''''_Int_select_q  :
                                                                    (\dconReadIn_CTf''''''''''''_f''''''''''''_Int_d [0] ? 2'd1 :
                                                                     (\dconWriteIn_CTf''''''''''''_f''''''''''''_Int_d [0] ? 2'd2 :
                                                                      2'd0)));
  logic [1:0] \dconReadIn_CTf''''''''''''_f''''''''''''_Int_select_q ;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \dconReadIn_CTf''''''''''''_f''''''''''''_Int_select_q  <= 2'd0;
    else
      \dconReadIn_CTf''''''''''''_f''''''''''''_Int_select_q  <= (\dconReadIn_CTf''''''''''''_f''''''''''''_Int_done  ? 2'd0 :
                                                                  \dconReadIn_CTf''''''''''''_f''''''''''''_Int_select_d );
  logic [1:0] \dconReadIn_CTf''''''''''''_f''''''''''''_Int_emit_q ;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \dconReadIn_CTf''''''''''''_f''''''''''''_Int_emit_q  <= 2'd0;
    else
      \dconReadIn_CTf''''''''''''_f''''''''''''_Int_emit_q  <= (\dconReadIn_CTf''''''''''''_f''''''''''''_Int_done  ? 2'd0 :
                                                                \dconReadIn_CTf''''''''''''_f''''''''''''_Int_emit_d );
  logic [1:0] \dconReadIn_CTf''''''''''''_f''''''''''''_Int_emit_d ;
  assign \dconReadIn_CTf''''''''''''_f''''''''''''_Int_emit_d  = (\dconReadIn_CTf''''''''''''_f''''''''''''_Int_emit_q  | ({\memMergeChoice_CTf''''''''''''_f''''''''''''_Int_d [0],
                                                                                                                            \memMergeIn_CTf''''''''''''_f''''''''''''_Int_d [0]} & {\memMergeChoice_CTf''''''''''''_f''''''''''''_Int_r ,
                                                                                                                                                                                    \memMergeIn_CTf''''''''''''_f''''''''''''_Int_r }));
  logic \dconReadIn_CTf''''''''''''_f''''''''''''_Int_done ;
  assign \dconReadIn_CTf''''''''''''_f''''''''''''_Int_done  = (& \dconReadIn_CTf''''''''''''_f''''''''''''_Int_emit_d );
  assign {\dconWriteIn_CTf''''''''''''_f''''''''''''_Int_r ,
          \dconReadIn_CTf''''''''''''_f''''''''''''_Int_r } = (\dconReadIn_CTf''''''''''''_f''''''''''''_Int_done  ? \dconReadIn_CTf''''''''''''_f''''''''''''_Int_select_d  :
                                                               2'd0);
  assign \memMergeIn_CTf''''''''''''_f''''''''''''_Int_d  = ((\dconReadIn_CTf''''''''''''_f''''''''''''_Int_select_d [0] && (! \dconReadIn_CTf''''''''''''_f''''''''''''_Int_emit_q [0])) ? \dconReadIn_CTf''''''''''''_f''''''''''''_Int_d  :
                                                             ((\dconReadIn_CTf''''''''''''_f''''''''''''_Int_select_d [1] && (! \dconReadIn_CTf''''''''''''_f''''''''''''_Int_emit_q [0])) ? \dconWriteIn_CTf''''''''''''_f''''''''''''_Int_d  :
                                                              {132'd0, 1'd0}));
  assign \memMergeChoice_CTf''''''''''''_f''''''''''''_Int_d  = ((\dconReadIn_CTf''''''''''''_f''''''''''''_Int_select_d [0] && (! \dconReadIn_CTf''''''''''''_f''''''''''''_Int_emit_q [1])) ? C1_2_dc(1'd1) :
                                                                 ((\dconReadIn_CTf''''''''''''_f''''''''''''_Int_select_d [1] && (! \dconReadIn_CTf''''''''''''_f''''''''''''_Int_emit_q [1])) ? C2_2_dc(1'd1) :
                                                                  {1'd0, 1'd0}));
  
  /* bram (Ty MemIn_CTf''''''''''''_f''''''''''''_Int,
      Ty MemOut_CTf''''''''''''_f''''''''''''_Int) : (memMergeIn_CTf''''''''''''_f''''''''''''_Int_dbuf,MemIn_CTf''''''''''''_f''''''''''''_Int) > (memOut_CTf''''''''''''_f''''''''''''_Int,MemOut_CTf''''''''''''_f''''''''''''_Int) */
  logic [114:0] \memMergeIn_CTf''''''''''''_f''''''''''''_Int_dbuf_mem [65535:0];
  logic [15:0] \memMergeIn_CTf''''''''''''_f''''''''''''_Int_dbuf_address ;
  logic [114:0] \memMergeIn_CTf''''''''''''_f''''''''''''_Int_dbuf_din ;
  logic [114:0] \memOut_CTf''''''''''''_f''''''''''''_Int_q ;
  logic \memOut_CTf''''''''''''_f''''''''''''_Int_valid ;
  logic \memMergeIn_CTf''''''''''''_f''''''''''''_Int_dbuf_we ;
  logic \memOut_CTf''''''''''''_f''''''''''''_Int_we ;
  assign \memMergeIn_CTf''''''''''''_f''''''''''''_Int_dbuf_din  = \memMergeIn_CTf''''''''''''_f''''''''''''_Int_dbuf_d [132:18];
  assign \memMergeIn_CTf''''''''''''_f''''''''''''_Int_dbuf_address  = \memMergeIn_CTf''''''''''''_f''''''''''''_Int_dbuf_d [17:2];
  assign \memMergeIn_CTf''''''''''''_f''''''''''''_Int_dbuf_we  = (\memMergeIn_CTf''''''''''''_f''''''''''''_Int_dbuf_d [1:1] && \memMergeIn_CTf''''''''''''_f''''''''''''_Int_dbuf_d [0]);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        \memOut_CTf''''''''''''_f''''''''''''_Int_we  <= 1'd0;
        \memOut_CTf''''''''''''_f''''''''''''_Int_valid  <= 1'd0;
      end
    else
      begin
        \memOut_CTf''''''''''''_f''''''''''''_Int_we  <= \memMergeIn_CTf''''''''''''_f''''''''''''_Int_dbuf_we ;
        \memOut_CTf''''''''''''_f''''''''''''_Int_valid  <= \memMergeIn_CTf''''''''''''_f''''''''''''_Int_dbuf_d [0];
        if (\memMergeIn_CTf''''''''''''_f''''''''''''_Int_dbuf_we )
          begin
            \memMergeIn_CTf''''''''''''_f''''''''''''_Int_dbuf_mem [\memMergeIn_CTf''''''''''''_f''''''''''''_Int_dbuf_address ] <= \memMergeIn_CTf''''''''''''_f''''''''''''_Int_dbuf_din ;
            \memOut_CTf''''''''''''_f''''''''''''_Int_q  <= \memMergeIn_CTf''''''''''''_f''''''''''''_Int_dbuf_din ;
          end
        else
          \memOut_CTf''''''''''''_f''''''''''''_Int_q  <= \memMergeIn_CTf''''''''''''_f''''''''''''_Int_dbuf_mem [\memMergeIn_CTf''''''''''''_f''''''''''''_Int_dbuf_address ];
      end
  assign \memOut_CTf''''''''''''_f''''''''''''_Int_d  = {\memOut_CTf''''''''''''_f''''''''''''_Int_q ,
                                                         \memOut_CTf''''''''''''_f''''''''''''_Int_we ,
                                                         \memOut_CTf''''''''''''_f''''''''''''_Int_valid };
  assign \memMergeIn_CTf''''''''''''_f''''''''''''_Int_dbuf_r  = ((! \memOut_CTf''''''''''''_f''''''''''''_Int_valid ) || \memOut_CTf''''''''''''_f''''''''''''_Int_r );
  logic [31:0] \profiling_MemIn_CTf''''''''''''_f''''''''''''_Int_read ;
  logic [31:0] \profiling_MemIn_CTf''''''''''''_f''''''''''''_Int_write ;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        \profiling_MemIn_CTf''''''''''''_f''''''''''''_Int_write  <= 0;
        \profiling_MemIn_CTf''''''''''''_f''''''''''''_Int_read  <= 0;
      end
    else
      if ((\memMergeIn_CTf''''''''''''_f''''''''''''_Int_dbuf_we  == 1'd1))
        \profiling_MemIn_CTf''''''''''''_f''''''''''''_Int_write  <= (\profiling_MemIn_CTf''''''''''''_f''''''''''''_Int_write  + 1);
      else
        if ((\memOut_CTf''''''''''''_f''''''''''''_Int_valid  == 1'd1))
          \profiling_MemIn_CTf''''''''''''_f''''''''''''_Int_read  <= (\profiling_MemIn_CTf''''''''''''_f''''''''''''_Int_read  + 1);
  
  /* demux (Ty C2,
       Ty MemOut_CTf''''''''''''_f''''''''''''_Int) : (memMergeChoice_CTf''''''''''''_f''''''''''''_Int,C2) (memOut_CTf''''''''''''_f''''''''''''_Int_dbuf,MemOut_CTf''''''''''''_f''''''''''''_Int) > [(memReadOut_CTf''''''''''''_f''''''''''''_Int,MemOut_CTf''''''''''''_f''''''''''''_Int),
                                                                                                                                                                                                        (memWriteOut_CTf''''''''''''_f''''''''''''_Int,MemOut_CTf''''''''''''_f''''''''''''_Int)] */
  logic [1:0] \memOut_CTf''''''''''''_f''''''''''''_Int_dbuf_onehotd ;
  always_comb
    if ((\memMergeChoice_CTf''''''''''''_f''''''''''''_Int_d [0] && \memOut_CTf''''''''''''_f''''''''''''_Int_dbuf_d [0]))
      unique case (\memMergeChoice_CTf''''''''''''_f''''''''''''_Int_d [1:1])
        1'd0:
          \memOut_CTf''''''''''''_f''''''''''''_Int_dbuf_onehotd  = 2'd1;
        1'd1:
          \memOut_CTf''''''''''''_f''''''''''''_Int_dbuf_onehotd  = 2'd2;
        default:
          \memOut_CTf''''''''''''_f''''''''''''_Int_dbuf_onehotd  = 2'd0;
      endcase
    else
      \memOut_CTf''''''''''''_f''''''''''''_Int_dbuf_onehotd  = 2'd0;
  assign \memReadOut_CTf''''''''''''_f''''''''''''_Int_d  = {\memOut_CTf''''''''''''_f''''''''''''_Int_dbuf_d [116:1],
                                                             \memOut_CTf''''''''''''_f''''''''''''_Int_dbuf_onehotd [0]};
  assign \memWriteOut_CTf''''''''''''_f''''''''''''_Int_d  = {\memOut_CTf''''''''''''_f''''''''''''_Int_dbuf_d [116:1],
                                                              \memOut_CTf''''''''''''_f''''''''''''_Int_dbuf_onehotd [1]};
  assign \memOut_CTf''''''''''''_f''''''''''''_Int_dbuf_r  = (| (\memOut_CTf''''''''''''_f''''''''''''_Int_dbuf_onehotd  & {\memWriteOut_CTf''''''''''''_f''''''''''''_Int_r ,
                                                                                                                            \memReadOut_CTf''''''''''''_f''''''''''''_Int_r }));
  assign \memMergeChoice_CTf''''''''''''_f''''''''''''_Int_r  = \memOut_CTf''''''''''''_f''''''''''''_Int_dbuf_r ;
  
  /* dbuf (Ty MemIn_CTf''''''''''''_f''''''''''''_Int) : (memMergeIn_CTf''''''''''''_f''''''''''''_Int_rbuf,MemIn_CTf''''''''''''_f''''''''''''_Int) > (memMergeIn_CTf''''''''''''_f''''''''''''_Int_dbuf,MemIn_CTf''''''''''''_f''''''''''''_Int) */
  assign \memMergeIn_CTf''''''''''''_f''''''''''''_Int_rbuf_r  = ((! \memMergeIn_CTf''''''''''''_f''''''''''''_Int_dbuf_d [0]) || \memMergeIn_CTf''''''''''''_f''''''''''''_Int_dbuf_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \memMergeIn_CTf''''''''''''_f''''''''''''_Int_dbuf_d  <= {132'd0,
                                                                1'd0};
    else
      if (\memMergeIn_CTf''''''''''''_f''''''''''''_Int_rbuf_r )
        \memMergeIn_CTf''''''''''''_f''''''''''''_Int_dbuf_d  <= \memMergeIn_CTf''''''''''''_f''''''''''''_Int_rbuf_d ;
  
  /* rbuf (Ty MemIn_CTf''''''''''''_f''''''''''''_Int) : (memMergeIn_CTf''''''''''''_f''''''''''''_Int,MemIn_CTf''''''''''''_f''''''''''''_Int) > (memMergeIn_CTf''''''''''''_f''''''''''''_Int_rbuf,MemIn_CTf''''''''''''_f''''''''''''_Int) */
  \MemIn_CTf''''''''''''_f''''''''''''_Int_t  \memMergeIn_CTf''''''''''''_f''''''''''''_Int_buf ;
  assign \memMergeIn_CTf''''''''''''_f''''''''''''_Int_r  = (! \memMergeIn_CTf''''''''''''_f''''''''''''_Int_buf [0]);
  assign \memMergeIn_CTf''''''''''''_f''''''''''''_Int_rbuf_d  = (\memMergeIn_CTf''''''''''''_f''''''''''''_Int_buf [0] ? \memMergeIn_CTf''''''''''''_f''''''''''''_Int_buf  :
                                                                  \memMergeIn_CTf''''''''''''_f''''''''''''_Int_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \memMergeIn_CTf''''''''''''_f''''''''''''_Int_buf  <= {132'd0,
                                                             1'd0};
    else
      if ((\memMergeIn_CTf''''''''''''_f''''''''''''_Int_rbuf_r  && \memMergeIn_CTf''''''''''''_f''''''''''''_Int_buf [0]))
        \memMergeIn_CTf''''''''''''_f''''''''''''_Int_buf  <= {132'd0,
                                                               1'd0};
      else if (((! \memMergeIn_CTf''''''''''''_f''''''''''''_Int_rbuf_r ) && (! \memMergeIn_CTf''''''''''''_f''''''''''''_Int_buf [0])))
        \memMergeIn_CTf''''''''''''_f''''''''''''_Int_buf  <= \memMergeIn_CTf''''''''''''_f''''''''''''_Int_d ;
  
  /* dbuf (Ty MemOut_CTf''''''''''''_f''''''''''''_Int) : (memOut_CTf''''''''''''_f''''''''''''_Int_rbuf,MemOut_CTf''''''''''''_f''''''''''''_Int) > (memOut_CTf''''''''''''_f''''''''''''_Int_dbuf,MemOut_CTf''''''''''''_f''''''''''''_Int) */
  assign \memOut_CTf''''''''''''_f''''''''''''_Int_rbuf_r  = ((! \memOut_CTf''''''''''''_f''''''''''''_Int_dbuf_d [0]) || \memOut_CTf''''''''''''_f''''''''''''_Int_dbuf_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \memOut_CTf''''''''''''_f''''''''''''_Int_dbuf_d  <= {116'd0,
                                                            1'd0};
    else
      if (\memOut_CTf''''''''''''_f''''''''''''_Int_rbuf_r )
        \memOut_CTf''''''''''''_f''''''''''''_Int_dbuf_d  <= \memOut_CTf''''''''''''_f''''''''''''_Int_rbuf_d ;
  
  /* rbuf (Ty MemOut_CTf''''''''''''_f''''''''''''_Int) : (memOut_CTf''''''''''''_f''''''''''''_Int,MemOut_CTf''''''''''''_f''''''''''''_Int) > (memOut_CTf''''''''''''_f''''''''''''_Int_rbuf,MemOut_CTf''''''''''''_f''''''''''''_Int) */
  \MemOut_CTf''''''''''''_f''''''''''''_Int_t  \memOut_CTf''''''''''''_f''''''''''''_Int_buf ;
  assign \memOut_CTf''''''''''''_f''''''''''''_Int_r  = (! \memOut_CTf''''''''''''_f''''''''''''_Int_buf [0]);
  assign \memOut_CTf''''''''''''_f''''''''''''_Int_rbuf_d  = (\memOut_CTf''''''''''''_f''''''''''''_Int_buf [0] ? \memOut_CTf''''''''''''_f''''''''''''_Int_buf  :
                                                              \memOut_CTf''''''''''''_f''''''''''''_Int_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \memOut_CTf''''''''''''_f''''''''''''_Int_buf  <= {116'd0, 1'd0};
    else
      if ((\memOut_CTf''''''''''''_f''''''''''''_Int_rbuf_r  && \memOut_CTf''''''''''''_f''''''''''''_Int_buf [0]))
        \memOut_CTf''''''''''''_f''''''''''''_Int_buf  <= {116'd0, 1'd0};
      else if (((! \memOut_CTf''''''''''''_f''''''''''''_Int_rbuf_r ) && (! \memOut_CTf''''''''''''_f''''''''''''_Int_buf [0])))
        \memOut_CTf''''''''''''_f''''''''''''_Int_buf  <= \memOut_CTf''''''''''''_f''''''''''''_Int_d ;
  
  /* destruct (Ty Pointer_CTf''''''''''''_f''''''''''''_Int,
          Dcon Pointer_CTf''''''''''''_f''''''''''''_Int) : (scfarg_0_1_1_argbuf,Pointer_CTf''''''''''''_f''''''''''''_Int) > [(destructReadIn_CTf''''''''''''_f''''''''''''_Int,Word16#)] */
  assign \destructReadIn_CTf''''''''''''_f''''''''''''_Int_d  = {scfarg_0_1_1_argbuf_d[16:1],
                                                                 scfarg_0_1_1_argbuf_d[0]};
  assign scfarg_0_1_1_argbuf_r = \destructReadIn_CTf''''''''''''_f''''''''''''_Int_r ;
  
  /* dcon (Ty MemIn_CTf''''''''''''_f''''''''''''_Int,
      Dcon ReadIn_CTf''''''''''''_f''''''''''''_Int) : [(destructReadIn_CTf''''''''''''_f''''''''''''_Int,Word16#)] > (dconReadIn_CTf''''''''''''_f''''''''''''_Int,MemIn_CTf''''''''''''_f''''''''''''_Int) */
  assign \dconReadIn_CTf''''''''''''_f''''''''''''_Int_d  = \ReadIn_CTf''''''''''''_f''''''''''''_Int_dc ((& {\destructReadIn_CTf''''''''''''_f''''''''''''_Int_d [0]}), \destructReadIn_CTf''''''''''''_f''''''''''''_Int_d );
  assign {\destructReadIn_CTf''''''''''''_f''''''''''''_Int_r } = {1 {(\dconReadIn_CTf''''''''''''_f''''''''''''_Int_r  && \dconReadIn_CTf''''''''''''_f''''''''''''_Int_d [0])}};
  
  /* destruct (Ty MemOut_CTf''''''''''''_f''''''''''''_Int,
          Dcon ReadOut_CTf''''''''''''_f''''''''''''_Int) : (memReadOut_CTf''''''''''''_f''''''''''''_Int,MemOut_CTf''''''''''''_f''''''''''''_Int) > [(readPointer_CTf''''''''''''_f''''''''''''_Intscfarg_0_1_1_argbuf,CTf''''''''''''_f''''''''''''_Int)] */
  assign \readPointer_CTf''''''''''''_f''''''''''''_Intscfarg_0_1_1_argbuf_d  = {\memReadOut_CTf''''''''''''_f''''''''''''_Int_d [116:2],
                                                                                 \memReadOut_CTf''''''''''''_f''''''''''''_Int_d [0]};
  assign \memReadOut_CTf''''''''''''_f''''''''''''_Int_r  = \readPointer_CTf''''''''''''_f''''''''''''_Intscfarg_0_1_1_argbuf_r ;
  
  /* mergectrl (Ty C5,
           Ty CTf''''''''''''_f''''''''''''_Int) : [(lizzieLet14_1_argbuf,CTf''''''''''''_f''''''''''''_Int),
                                                    (lizzieLet56_1_argbuf,CTf''''''''''''_f''''''''''''_Int),
                                                    (lizzieLet63_1_argbuf,CTf''''''''''''_f''''''''''''_Int),
                                                    (lizzieLet64_1_argbuf,CTf''''''''''''_f''''''''''''_Int),
                                                    (lizzieLet65_1_argbuf,CTf''''''''''''_f''''''''''''_Int)] > (writeMerge_choice_CTf''''''''''''_f''''''''''''_Int,C5) (writeMerge_data_CTf''''''''''''_f''''''''''''_Int,CTf''''''''''''_f''''''''''''_Int) */
  logic [4:0] lizzieLet14_1_argbuf_select_d;
  assign lizzieLet14_1_argbuf_select_d = ((| lizzieLet14_1_argbuf_select_q) ? lizzieLet14_1_argbuf_select_q :
                                          (lizzieLet14_1_argbuf_d[0] ? 5'd1 :
                                           (lizzieLet56_1_argbuf_d[0] ? 5'd2 :
                                            (lizzieLet63_1_argbuf_d[0] ? 5'd4 :
                                             (lizzieLet64_1_argbuf_d[0] ? 5'd8 :
                                              (lizzieLet65_1_argbuf_d[0] ? 5'd16 :
                                               5'd0))))));
  logic [4:0] lizzieLet14_1_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet14_1_argbuf_select_q <= 5'd0;
    else
      lizzieLet14_1_argbuf_select_q <= (lizzieLet14_1_argbuf_done ? 5'd0 :
                                        lizzieLet14_1_argbuf_select_d);
  logic [1:0] lizzieLet14_1_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet14_1_argbuf_emit_q <= 2'd0;
    else
      lizzieLet14_1_argbuf_emit_q <= (lizzieLet14_1_argbuf_done ? 2'd0 :
                                      lizzieLet14_1_argbuf_emit_d);
  logic [1:0] lizzieLet14_1_argbuf_emit_d;
  assign lizzieLet14_1_argbuf_emit_d = (lizzieLet14_1_argbuf_emit_q | ({\writeMerge_choice_CTf''''''''''''_f''''''''''''_Int_d [0],
                                                                        \writeMerge_data_CTf''''''''''''_f''''''''''''_Int_d [0]} & {\writeMerge_choice_CTf''''''''''''_f''''''''''''_Int_r ,
                                                                                                                                     \writeMerge_data_CTf''''''''''''_f''''''''''''_Int_r }));
  logic lizzieLet14_1_argbuf_done;
  assign lizzieLet14_1_argbuf_done = (& lizzieLet14_1_argbuf_emit_d);
  assign {lizzieLet65_1_argbuf_r,
          lizzieLet64_1_argbuf_r,
          lizzieLet63_1_argbuf_r,
          lizzieLet56_1_argbuf_r,
          lizzieLet14_1_argbuf_r} = (lizzieLet14_1_argbuf_done ? lizzieLet14_1_argbuf_select_d :
                                     5'd0);
  assign \writeMerge_data_CTf''''''''''''_f''''''''''''_Int_d  = ((lizzieLet14_1_argbuf_select_d[0] && (! lizzieLet14_1_argbuf_emit_q[0])) ? lizzieLet14_1_argbuf_d :
                                                                  ((lizzieLet14_1_argbuf_select_d[1] && (! lizzieLet14_1_argbuf_emit_q[0])) ? lizzieLet56_1_argbuf_d :
                                                                   ((lizzieLet14_1_argbuf_select_d[2] && (! lizzieLet14_1_argbuf_emit_q[0])) ? lizzieLet63_1_argbuf_d :
                                                                    ((lizzieLet14_1_argbuf_select_d[3] && (! lizzieLet14_1_argbuf_emit_q[0])) ? lizzieLet64_1_argbuf_d :
                                                                     ((lizzieLet14_1_argbuf_select_d[4] && (! lizzieLet14_1_argbuf_emit_q[0])) ? lizzieLet65_1_argbuf_d :
                                                                      {115'd0, 1'd0})))));
  assign \writeMerge_choice_CTf''''''''''''_f''''''''''''_Int_d  = ((lizzieLet14_1_argbuf_select_d[0] && (! lizzieLet14_1_argbuf_emit_q[1])) ? C1_5_dc(1'd1) :
                                                                    ((lizzieLet14_1_argbuf_select_d[1] && (! lizzieLet14_1_argbuf_emit_q[1])) ? C2_5_dc(1'd1) :
                                                                     ((lizzieLet14_1_argbuf_select_d[2] && (! lizzieLet14_1_argbuf_emit_q[1])) ? C3_5_dc(1'd1) :
                                                                      ((lizzieLet14_1_argbuf_select_d[3] && (! lizzieLet14_1_argbuf_emit_q[1])) ? C4_5_dc(1'd1) :
                                                                       ((lizzieLet14_1_argbuf_select_d[4] && (! lizzieLet14_1_argbuf_emit_q[1])) ? C5_5_dc(1'd1) :
                                                                        {3'd0, 1'd0})))));
  
  /* demux (Ty C5,
       Ty Pointer_CTf''''''''''''_f''''''''''''_Int) : (writeMerge_choice_CTf''''''''''''_f''''''''''''_Int,C5) (demuxWriteResult_CTf''''''''''''_f''''''''''''_Int,Pointer_CTf''''''''''''_f''''''''''''_Int) > [(writeCTf''''''''''''_f''''''''''''_IntlizzieLet14_1_argbuf,Pointer_CTf''''''''''''_f''''''''''''_Int),
                                                                                                                                                                                                                  (writeCTf''''''''''''_f''''''''''''_IntlizzieLet56_1_argbuf,Pointer_CTf''''''''''''_f''''''''''''_Int),
                                                                                                                                                                                                                  (writeCTf''''''''''''_f''''''''''''_IntlizzieLet63_1_argbuf,Pointer_CTf''''''''''''_f''''''''''''_Int),
                                                                                                                                                                                                                  (writeCTf''''''''''''_f''''''''''''_IntlizzieLet64_1_argbuf,Pointer_CTf''''''''''''_f''''''''''''_Int),
                                                                                                                                                                                                                  (writeCTf''''''''''''_f''''''''''''_IntlizzieLet65_1_argbuf,Pointer_CTf''''''''''''_f''''''''''''_Int)] */
  logic [4:0] \demuxWriteResult_CTf''''''''''''_f''''''''''''_Int_onehotd ;
  always_comb
    if ((\writeMerge_choice_CTf''''''''''''_f''''''''''''_Int_d [0] && \demuxWriteResult_CTf''''''''''''_f''''''''''''_Int_d [0]))
      unique case (\writeMerge_choice_CTf''''''''''''_f''''''''''''_Int_d [3:1])
        3'd0:
          \demuxWriteResult_CTf''''''''''''_f''''''''''''_Int_onehotd  = 5'd1;
        3'd1:
          \demuxWriteResult_CTf''''''''''''_f''''''''''''_Int_onehotd  = 5'd2;
        3'd2:
          \demuxWriteResult_CTf''''''''''''_f''''''''''''_Int_onehotd  = 5'd4;
        3'd3:
          \demuxWriteResult_CTf''''''''''''_f''''''''''''_Int_onehotd  = 5'd8;
        3'd4:
          \demuxWriteResult_CTf''''''''''''_f''''''''''''_Int_onehotd  = 5'd16;
        default:
          \demuxWriteResult_CTf''''''''''''_f''''''''''''_Int_onehotd  = 5'd0;
      endcase
    else
      \demuxWriteResult_CTf''''''''''''_f''''''''''''_Int_onehotd  = 5'd0;
  assign \writeCTf''''''''''''_f''''''''''''_IntlizzieLet14_1_argbuf_d  = {\demuxWriteResult_CTf''''''''''''_f''''''''''''_Int_d [16:1],
                                                                           \demuxWriteResult_CTf''''''''''''_f''''''''''''_Int_onehotd [0]};
  assign \writeCTf''''''''''''_f''''''''''''_IntlizzieLet56_1_argbuf_d  = {\demuxWriteResult_CTf''''''''''''_f''''''''''''_Int_d [16:1],
                                                                           \demuxWriteResult_CTf''''''''''''_f''''''''''''_Int_onehotd [1]};
  assign \writeCTf''''''''''''_f''''''''''''_IntlizzieLet63_1_argbuf_d  = {\demuxWriteResult_CTf''''''''''''_f''''''''''''_Int_d [16:1],
                                                                           \demuxWriteResult_CTf''''''''''''_f''''''''''''_Int_onehotd [2]};
  assign \writeCTf''''''''''''_f''''''''''''_IntlizzieLet64_1_argbuf_d  = {\demuxWriteResult_CTf''''''''''''_f''''''''''''_Int_d [16:1],
                                                                           \demuxWriteResult_CTf''''''''''''_f''''''''''''_Int_onehotd [3]};
  assign \writeCTf''''''''''''_f''''''''''''_IntlizzieLet65_1_argbuf_d  = {\demuxWriteResult_CTf''''''''''''_f''''''''''''_Int_d [16:1],
                                                                           \demuxWriteResult_CTf''''''''''''_f''''''''''''_Int_onehotd [4]};
  assign \demuxWriteResult_CTf''''''''''''_f''''''''''''_Int_r  = (| (\demuxWriteResult_CTf''''''''''''_f''''''''''''_Int_onehotd  & {\writeCTf''''''''''''_f''''''''''''_IntlizzieLet65_1_argbuf_r ,
                                                                                                                                      \writeCTf''''''''''''_f''''''''''''_IntlizzieLet64_1_argbuf_r ,
                                                                                                                                      \writeCTf''''''''''''_f''''''''''''_IntlizzieLet63_1_argbuf_r ,
                                                                                                                                      \writeCTf''''''''''''_f''''''''''''_IntlizzieLet56_1_argbuf_r ,
                                                                                                                                      \writeCTf''''''''''''_f''''''''''''_IntlizzieLet14_1_argbuf_r }));
  assign \writeMerge_choice_CTf''''''''''''_f''''''''''''_Int_r  = \demuxWriteResult_CTf''''''''''''_f''''''''''''_Int_r ;
  
  /* dcon (Ty MemIn_CTf''''''''''''_f''''''''''''_Int,
      Dcon WriteIn_CTf''''''''''''_f''''''''''''_Int) : [(forkHP1_CTf''''''''''''_f''''''''''''_In2,Word16#),
                                                         (writeMerge_data_CTf''''''''''''_f''''''''''''_Int,CTf''''''''''''_f''''''''''''_Int)] > (dconWriteIn_CTf''''''''''''_f''''''''''''_Int,MemIn_CTf''''''''''''_f''''''''''''_Int) */
  assign \dconWriteIn_CTf''''''''''''_f''''''''''''_Int_d  = \WriteIn_CTf''''''''''''_f''''''''''''_Int_dc ((& {\forkHP1_CTf''''''''''''_f''''''''''''_In2_d [0],
                                                                                                                \writeMerge_data_CTf''''''''''''_f''''''''''''_Int_d [0]}), \forkHP1_CTf''''''''''''_f''''''''''''_In2_d , \writeMerge_data_CTf''''''''''''_f''''''''''''_Int_d );
  assign {\forkHP1_CTf''''''''''''_f''''''''''''_In2_r ,
          \writeMerge_data_CTf''''''''''''_f''''''''''''_Int_r } = {2 {(\dconWriteIn_CTf''''''''''''_f''''''''''''_Int_r  && \dconWriteIn_CTf''''''''''''_f''''''''''''_Int_d [0])}};
  
  /* dcon (Ty Pointer_CTf''''''''''''_f''''''''''''_Int,
      Dcon Pointer_CTf''''''''''''_f''''''''''''_Int) : [(forkHP1_CTf''''''''''''_f''''''''''''_In3,Word16#)] > (dconPtr_CTf''''''''''''_f''''''''''''_Int,Pointer_CTf''''''''''''_f''''''''''''_Int) */
  assign \dconPtr_CTf''''''''''''_f''''''''''''_Int_d  = \Pointer_CTf''''''''''''_f''''''''''''_Int_dc ((& {\forkHP1_CTf''''''''''''_f''''''''''''_In3_d [0]}), \forkHP1_CTf''''''''''''_f''''''''''''_In3_d );
  assign {\forkHP1_CTf''''''''''''_f''''''''''''_In3_r } = {1 {(\dconPtr_CTf''''''''''''_f''''''''''''_Int_r  && \dconPtr_CTf''''''''''''_f''''''''''''_Int_d [0])}};
  
  /* demux (Ty MemOut_CTf''''''''''''_f''''''''''''_Int,
       Ty Pointer_CTf''''''''''''_f''''''''''''_Int) : (memWriteOut_CTf''''''''''''_f''''''''''''_Int,MemOut_CTf''''''''''''_f''''''''''''_Int) (dconPtr_CTf''''''''''''_f''''''''''''_Int,Pointer_CTf''''''''''''_f''''''''''''_Int) > [(_257,Pointer_CTf''''''''''''_f''''''''''''_Int),
                                                                                                                                                                                                                                         (demuxWriteResult_CTf''''''''''''_f''''''''''''_Int,Pointer_CTf''''''''''''_f''''''''''''_Int)] */
  logic [1:0] \dconPtr_CTf''''''''''''_f''''''''''''_Int_onehotd ;
  always_comb
    if ((\memWriteOut_CTf''''''''''''_f''''''''''''_Int_d [0] && \dconPtr_CTf''''''''''''_f''''''''''''_Int_d [0]))
      unique case (\memWriteOut_CTf''''''''''''_f''''''''''''_Int_d [1:1])
        1'd0: \dconPtr_CTf''''''''''''_f''''''''''''_Int_onehotd  = 2'd1;
        1'd1: \dconPtr_CTf''''''''''''_f''''''''''''_Int_onehotd  = 2'd2;
        default:
          \dconPtr_CTf''''''''''''_f''''''''''''_Int_onehotd  = 2'd0;
      endcase
    else \dconPtr_CTf''''''''''''_f''''''''''''_Int_onehotd  = 2'd0;
  assign _257_d = {\dconPtr_CTf''''''''''''_f''''''''''''_Int_d [16:1],
                   \dconPtr_CTf''''''''''''_f''''''''''''_Int_onehotd [0]};
  assign \demuxWriteResult_CTf''''''''''''_f''''''''''''_Int_d  = {\dconPtr_CTf''''''''''''_f''''''''''''_Int_d [16:1],
                                                                   \dconPtr_CTf''''''''''''_f''''''''''''_Int_onehotd [1]};
  assign \dconPtr_CTf''''''''''''_f''''''''''''_Int_r  = (| (\dconPtr_CTf''''''''''''_f''''''''''''_Int_onehotd  & {\demuxWriteResult_CTf''''''''''''_f''''''''''''_Int_r ,
                                                                                                                    _257_r}));
  assign \memWriteOut_CTf''''''''''''_f''''''''''''_Int_r  = \dconPtr_CTf''''''''''''_f''''''''''''_Int_r ;
  
  /* const (Ty Word16#,Lit 0) : (go__9,Go) > (initHP_CTf_f_Int,Word16#) */
  assign initHP_CTf_f_Int_d = {16'd0, go__9_d[0]};
  assign go__9_r = initHP_CTf_f_Int_r;
  
  /* const (Ty Word16#,
       Lit 1) : (incrHP_CTf_f_Int1,Go) > (incrHP_CTf_f_Int,Word16#) */
  assign incrHP_CTf_f_Int_d = {16'd1, incrHP_CTf_f_Int1_d[0]};
  assign incrHP_CTf_f_Int1_r = incrHP_CTf_f_Int_r;
  
  /* merge (Ty Go) : [(go__10,Go),
                 (incrHP_CTf_f_Int2,Go)] > (incrHP_mergeCTf_f_Int,Go) */
  logic [1:0] incrHP_mergeCTf_f_Int_selected;
  logic [1:0] incrHP_mergeCTf_f_Int_select;
  always_comb
    begin
      incrHP_mergeCTf_f_Int_selected = 2'd0;
      if ((| incrHP_mergeCTf_f_Int_select))
        incrHP_mergeCTf_f_Int_selected = incrHP_mergeCTf_f_Int_select;
      else
        if (go__10_d[0]) incrHP_mergeCTf_f_Int_selected[0] = 1'd1;
        else if (incrHP_CTf_f_Int2_d[0])
          incrHP_mergeCTf_f_Int_selected[1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeCTf_f_Int_select <= 2'd0;
    else
      incrHP_mergeCTf_f_Int_select <= (incrHP_mergeCTf_f_Int_r ? 2'd0 :
                                       incrHP_mergeCTf_f_Int_selected);
  always_comb
    if (incrHP_mergeCTf_f_Int_selected[0])
      incrHP_mergeCTf_f_Int_d = go__10_d;
    else if (incrHP_mergeCTf_f_Int_selected[1])
      incrHP_mergeCTf_f_Int_d = incrHP_CTf_f_Int2_d;
    else incrHP_mergeCTf_f_Int_d = 1'd0;
  assign {incrHP_CTf_f_Int2_r,
          go__10_r} = (incrHP_mergeCTf_f_Int_r ? incrHP_mergeCTf_f_Int_selected :
                       2'd0);
  
  /* fork (Ty Go) : (incrHP_mergeCTf_f_Int_buf,Go) > [(incrHP_CTf_f_Int1,Go),
                                                 (incrHP_CTf_f_Int2,Go)] */
  logic [1:0] incrHP_mergeCTf_f_Int_buf_emitted;
  logic [1:0] incrHP_mergeCTf_f_Int_buf_done;
  assign incrHP_CTf_f_Int1_d = (incrHP_mergeCTf_f_Int_buf_d[0] && (! incrHP_mergeCTf_f_Int_buf_emitted[0]));
  assign incrHP_CTf_f_Int2_d = (incrHP_mergeCTf_f_Int_buf_d[0] && (! incrHP_mergeCTf_f_Int_buf_emitted[1]));
  assign incrHP_mergeCTf_f_Int_buf_done = (incrHP_mergeCTf_f_Int_buf_emitted | ({incrHP_CTf_f_Int2_d[0],
                                                                                 incrHP_CTf_f_Int1_d[0]} & {incrHP_CTf_f_Int2_r,
                                                                                                            incrHP_CTf_f_Int1_r}));
  assign incrHP_mergeCTf_f_Int_buf_r = (& incrHP_mergeCTf_f_Int_buf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeCTf_f_Int_buf_emitted <= 2'd0;
    else
      incrHP_mergeCTf_f_Int_buf_emitted <= (incrHP_mergeCTf_f_Int_buf_r ? 2'd0 :
                                            incrHP_mergeCTf_f_Int_buf_done);
  
  /* op_add (Ty Word16#) : (incrHP_CTf_f_Int,Word16#) (forkHP1_CTf_f_Int,Word16#) > (addHP_CTf_f_Int,Word16#) */
  assign addHP_CTf_f_Int_d = {(incrHP_CTf_f_Int_d[16:1] + forkHP1_CTf_f_Int_d[16:1]),
                              (incrHP_CTf_f_Int_d[0] && forkHP1_CTf_f_Int_d[0])};
  assign {incrHP_CTf_f_Int_r,
          forkHP1_CTf_f_Int_r} = {2 {(addHP_CTf_f_Int_r && addHP_CTf_f_Int_d[0])}};
  
  /* merge (Ty Word16#) : [(initHP_CTf_f_Int,Word16#),
                      (addHP_CTf_f_Int,Word16#)] > (mergeHP_CTf_f_Int,Word16#) */
  logic [1:0] mergeHP_CTf_f_Int_selected;
  logic [1:0] mergeHP_CTf_f_Int_select;
  always_comb
    begin
      mergeHP_CTf_f_Int_selected = 2'd0;
      if ((| mergeHP_CTf_f_Int_select))
        mergeHP_CTf_f_Int_selected = mergeHP_CTf_f_Int_select;
      else
        if (initHP_CTf_f_Int_d[0]) mergeHP_CTf_f_Int_selected[0] = 1'd1;
        else if (addHP_CTf_f_Int_d[0])
          mergeHP_CTf_f_Int_selected[1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_CTf_f_Int_select <= 2'd0;
    else
      mergeHP_CTf_f_Int_select <= (mergeHP_CTf_f_Int_r ? 2'd0 :
                                   mergeHP_CTf_f_Int_selected);
  always_comb
    if (mergeHP_CTf_f_Int_selected[0])
      mergeHP_CTf_f_Int_d = initHP_CTf_f_Int_d;
    else if (mergeHP_CTf_f_Int_selected[1])
      mergeHP_CTf_f_Int_d = addHP_CTf_f_Int_d;
    else mergeHP_CTf_f_Int_d = {16'd0, 1'd0};
  assign {addHP_CTf_f_Int_r,
          initHP_CTf_f_Int_r} = (mergeHP_CTf_f_Int_r ? mergeHP_CTf_f_Int_selected :
                                 2'd0);
  
  /* buf (Ty Go) : (incrHP_mergeCTf_f_Int,Go) > (incrHP_mergeCTf_f_Int_buf,Go) */
  Go_t incrHP_mergeCTf_f_Int_bufchan_d;
  logic incrHP_mergeCTf_f_Int_bufchan_r;
  assign incrHP_mergeCTf_f_Int_r = ((! incrHP_mergeCTf_f_Int_bufchan_d[0]) || incrHP_mergeCTf_f_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeCTf_f_Int_bufchan_d <= 1'd0;
    else
      if (incrHP_mergeCTf_f_Int_r)
        incrHP_mergeCTf_f_Int_bufchan_d <= incrHP_mergeCTf_f_Int_d;
  Go_t incrHP_mergeCTf_f_Int_bufchan_buf;
  assign incrHP_mergeCTf_f_Int_bufchan_r = (! incrHP_mergeCTf_f_Int_bufchan_buf[0]);
  assign incrHP_mergeCTf_f_Int_buf_d = (incrHP_mergeCTf_f_Int_bufchan_buf[0] ? incrHP_mergeCTf_f_Int_bufchan_buf :
                                        incrHP_mergeCTf_f_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeCTf_f_Int_bufchan_buf <= 1'd0;
    else
      if ((incrHP_mergeCTf_f_Int_buf_r && incrHP_mergeCTf_f_Int_bufchan_buf[0]))
        incrHP_mergeCTf_f_Int_bufchan_buf <= 1'd0;
      else if (((! incrHP_mergeCTf_f_Int_buf_r) && (! incrHP_mergeCTf_f_Int_bufchan_buf[0])))
        incrHP_mergeCTf_f_Int_bufchan_buf <= incrHP_mergeCTf_f_Int_bufchan_d;
  
  /* buf (Ty Word16#) : (mergeHP_CTf_f_Int,Word16#) > (mergeHP_CTf_f_Int_buf,Word16#) */
  \Word16#_t  mergeHP_CTf_f_Int_bufchan_d;
  logic mergeHP_CTf_f_Int_bufchan_r;
  assign mergeHP_CTf_f_Int_r = ((! mergeHP_CTf_f_Int_bufchan_d[0]) || mergeHP_CTf_f_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_CTf_f_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (mergeHP_CTf_f_Int_r)
        mergeHP_CTf_f_Int_bufchan_d <= mergeHP_CTf_f_Int_d;
  \Word16#_t  mergeHP_CTf_f_Int_bufchan_buf;
  assign mergeHP_CTf_f_Int_bufchan_r = (! mergeHP_CTf_f_Int_bufchan_buf[0]);
  assign mergeHP_CTf_f_Int_buf_d = (mergeHP_CTf_f_Int_bufchan_buf[0] ? mergeHP_CTf_f_Int_bufchan_buf :
                                    mergeHP_CTf_f_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      mergeHP_CTf_f_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((mergeHP_CTf_f_Int_buf_r && mergeHP_CTf_f_Int_bufchan_buf[0]))
        mergeHP_CTf_f_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! mergeHP_CTf_f_Int_buf_r) && (! mergeHP_CTf_f_Int_bufchan_buf[0])))
        mergeHP_CTf_f_Int_bufchan_buf <= mergeHP_CTf_f_Int_bufchan_d;
  
  /* fork (Ty Word16#) : (mergeHP_CTf_f_Int_buf,Word16#) > [(forkHP1_CTf_f_Int,Word16#),
                                                       (forkHP1_CTf_f_In2,Word16#),
                                                       (forkHP1_CTf_f_In3,Word16#)] */
  logic [2:0] mergeHP_CTf_f_Int_buf_emitted;
  logic [2:0] mergeHP_CTf_f_Int_buf_done;
  assign forkHP1_CTf_f_Int_d = {mergeHP_CTf_f_Int_buf_d[16:1],
                                (mergeHP_CTf_f_Int_buf_d[0] && (! mergeHP_CTf_f_Int_buf_emitted[0]))};
  assign forkHP1_CTf_f_In2_d = {mergeHP_CTf_f_Int_buf_d[16:1],
                                (mergeHP_CTf_f_Int_buf_d[0] && (! mergeHP_CTf_f_Int_buf_emitted[1]))};
  assign forkHP1_CTf_f_In3_d = {mergeHP_CTf_f_Int_buf_d[16:1],
                                (mergeHP_CTf_f_Int_buf_d[0] && (! mergeHP_CTf_f_Int_buf_emitted[2]))};
  assign mergeHP_CTf_f_Int_buf_done = (mergeHP_CTf_f_Int_buf_emitted | ({forkHP1_CTf_f_In3_d[0],
                                                                         forkHP1_CTf_f_In2_d[0],
                                                                         forkHP1_CTf_f_Int_d[0]} & {forkHP1_CTf_f_In3_r,
                                                                                                    forkHP1_CTf_f_In2_r,
                                                                                                    forkHP1_CTf_f_Int_r}));
  assign mergeHP_CTf_f_Int_buf_r = (& mergeHP_CTf_f_Int_buf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_CTf_f_Int_buf_emitted <= 3'd0;
    else
      mergeHP_CTf_f_Int_buf_emitted <= (mergeHP_CTf_f_Int_buf_r ? 3'd0 :
                                        mergeHP_CTf_f_Int_buf_done);
  
  /* mergectrl (Ty C2,
           Ty MemIn_CTf_f_Int) : [(dconReadIn_CTf_f_Int,MemIn_CTf_f_Int),
                                  (dconWriteIn_CTf_f_Int,MemIn_CTf_f_Int)] > (memMergeChoice_CTf_f_Int,C2) (memMergeIn_CTf_f_Int,MemIn_CTf_f_Int) */
  logic [1:0] dconReadIn_CTf_f_Int_select_d;
  assign dconReadIn_CTf_f_Int_select_d = ((| dconReadIn_CTf_f_Int_select_q) ? dconReadIn_CTf_f_Int_select_q :
                                          (dconReadIn_CTf_f_Int_d[0] ? 2'd1 :
                                           (dconWriteIn_CTf_f_Int_d[0] ? 2'd2 :
                                            2'd0)));
  logic [1:0] dconReadIn_CTf_f_Int_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) dconReadIn_CTf_f_Int_select_q <= 2'd0;
    else
      dconReadIn_CTf_f_Int_select_q <= (dconReadIn_CTf_f_Int_done ? 2'd0 :
                                        dconReadIn_CTf_f_Int_select_d);
  logic [1:0] dconReadIn_CTf_f_Int_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) dconReadIn_CTf_f_Int_emit_q <= 2'd0;
    else
      dconReadIn_CTf_f_Int_emit_q <= (dconReadIn_CTf_f_Int_done ? 2'd0 :
                                      dconReadIn_CTf_f_Int_emit_d);
  logic [1:0] dconReadIn_CTf_f_Int_emit_d;
  assign dconReadIn_CTf_f_Int_emit_d = (dconReadIn_CTf_f_Int_emit_q | ({memMergeChoice_CTf_f_Int_d[0],
                                                                        memMergeIn_CTf_f_Int_d[0]} & {memMergeChoice_CTf_f_Int_r,
                                                                                                      memMergeIn_CTf_f_Int_r}));
  logic dconReadIn_CTf_f_Int_done;
  assign dconReadIn_CTf_f_Int_done = (& dconReadIn_CTf_f_Int_emit_d);
  assign {dconWriteIn_CTf_f_Int_r,
          dconReadIn_CTf_f_Int_r} = (dconReadIn_CTf_f_Int_done ? dconReadIn_CTf_f_Int_select_d :
                                     2'd0);
  assign memMergeIn_CTf_f_Int_d = ((dconReadIn_CTf_f_Int_select_d[0] && (! dconReadIn_CTf_f_Int_emit_q[0])) ? dconReadIn_CTf_f_Int_d :
                                   ((dconReadIn_CTf_f_Int_select_d[1] && (! dconReadIn_CTf_f_Int_emit_q[0])) ? dconWriteIn_CTf_f_Int_d :
                                    {180'd0, 1'd0}));
  assign memMergeChoice_CTf_f_Int_d = ((dconReadIn_CTf_f_Int_select_d[0] && (! dconReadIn_CTf_f_Int_emit_q[1])) ? C1_2_dc(1'd1) :
                                       ((dconReadIn_CTf_f_Int_select_d[1] && (! dconReadIn_CTf_f_Int_emit_q[1])) ? C2_2_dc(1'd1) :
                                        {1'd0, 1'd0}));
  
  /* bram (Ty MemIn_CTf_f_Int,
      Ty MemOut_CTf_f_Int) : (memMergeIn_CTf_f_Int_dbuf,MemIn_CTf_f_Int) > (memOut_CTf_f_Int,MemOut_CTf_f_Int) */
  logic [162:0] memMergeIn_CTf_f_Int_dbuf_mem[65535:0];
  logic [15:0] memMergeIn_CTf_f_Int_dbuf_address;
  logic [162:0] memMergeIn_CTf_f_Int_dbuf_din;
  logic [162:0] memOut_CTf_f_Int_q;
  logic memOut_CTf_f_Int_valid;
  logic memMergeIn_CTf_f_Int_dbuf_we;
  logic memOut_CTf_f_Int_we;
  assign memMergeIn_CTf_f_Int_dbuf_din = memMergeIn_CTf_f_Int_dbuf_d[180:18];
  assign memMergeIn_CTf_f_Int_dbuf_address = memMergeIn_CTf_f_Int_dbuf_d[17:2];
  assign memMergeIn_CTf_f_Int_dbuf_we = (memMergeIn_CTf_f_Int_dbuf_d[1:1] && memMergeIn_CTf_f_Int_dbuf_d[0]);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        memOut_CTf_f_Int_we <= 1'd0;
        memOut_CTf_f_Int_valid <= 1'd0;
      end
    else
      begin
        memOut_CTf_f_Int_we <= memMergeIn_CTf_f_Int_dbuf_we;
        memOut_CTf_f_Int_valid <= memMergeIn_CTf_f_Int_dbuf_d[0];
        if (memMergeIn_CTf_f_Int_dbuf_we)
          begin
            memMergeIn_CTf_f_Int_dbuf_mem[memMergeIn_CTf_f_Int_dbuf_address] <= memMergeIn_CTf_f_Int_dbuf_din;
            memOut_CTf_f_Int_q <= memMergeIn_CTf_f_Int_dbuf_din;
          end
        else
          memOut_CTf_f_Int_q <= memMergeIn_CTf_f_Int_dbuf_mem[memMergeIn_CTf_f_Int_dbuf_address];
      end
  assign memOut_CTf_f_Int_d = {memOut_CTf_f_Int_q,
                               memOut_CTf_f_Int_we,
                               memOut_CTf_f_Int_valid};
  assign memMergeIn_CTf_f_Int_dbuf_r = ((! memOut_CTf_f_Int_valid) || memOut_CTf_f_Int_r);
  logic [31:0] profiling_MemIn_CTf_f_Int_read;
  logic [31:0] profiling_MemIn_CTf_f_Int_write;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        profiling_MemIn_CTf_f_Int_write <= 0;
        profiling_MemIn_CTf_f_Int_read <= 0;
      end
    else
      if ((memMergeIn_CTf_f_Int_dbuf_we == 1'd1))
        profiling_MemIn_CTf_f_Int_write <= (profiling_MemIn_CTf_f_Int_write + 1);
      else
        if ((memOut_CTf_f_Int_valid == 1'd1))
          profiling_MemIn_CTf_f_Int_read <= (profiling_MemIn_CTf_f_Int_read + 1);
  
  /* demux (Ty C2,
       Ty MemOut_CTf_f_Int) : (memMergeChoice_CTf_f_Int,C2) (memOut_CTf_f_Int_dbuf,MemOut_CTf_f_Int) > [(memReadOut_CTf_f_Int,MemOut_CTf_f_Int),
                                                                                                        (memWriteOut_CTf_f_Int,MemOut_CTf_f_Int)] */
  logic [1:0] memOut_CTf_f_Int_dbuf_onehotd;
  always_comb
    if ((memMergeChoice_CTf_f_Int_d[0] && memOut_CTf_f_Int_dbuf_d[0]))
      unique case (memMergeChoice_CTf_f_Int_d[1:1])
        1'd0: memOut_CTf_f_Int_dbuf_onehotd = 2'd1;
        1'd1: memOut_CTf_f_Int_dbuf_onehotd = 2'd2;
        default: memOut_CTf_f_Int_dbuf_onehotd = 2'd0;
      endcase
    else memOut_CTf_f_Int_dbuf_onehotd = 2'd0;
  assign memReadOut_CTf_f_Int_d = {memOut_CTf_f_Int_dbuf_d[164:1],
                                   memOut_CTf_f_Int_dbuf_onehotd[0]};
  assign memWriteOut_CTf_f_Int_d = {memOut_CTf_f_Int_dbuf_d[164:1],
                                    memOut_CTf_f_Int_dbuf_onehotd[1]};
  assign memOut_CTf_f_Int_dbuf_r = (| (memOut_CTf_f_Int_dbuf_onehotd & {memWriteOut_CTf_f_Int_r,
                                                                        memReadOut_CTf_f_Int_r}));
  assign memMergeChoice_CTf_f_Int_r = memOut_CTf_f_Int_dbuf_r;
  
  /* dbuf (Ty MemIn_CTf_f_Int) : (memMergeIn_CTf_f_Int_rbuf,MemIn_CTf_f_Int) > (memMergeIn_CTf_f_Int_dbuf,MemIn_CTf_f_Int) */
  assign memMergeIn_CTf_f_Int_rbuf_r = ((! memMergeIn_CTf_f_Int_dbuf_d[0]) || memMergeIn_CTf_f_Int_dbuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memMergeIn_CTf_f_Int_dbuf_d <= {180'd0, 1'd0};
    else
      if (memMergeIn_CTf_f_Int_rbuf_r)
        memMergeIn_CTf_f_Int_dbuf_d <= memMergeIn_CTf_f_Int_rbuf_d;
  
  /* rbuf (Ty MemIn_CTf_f_Int) : (memMergeIn_CTf_f_Int,MemIn_CTf_f_Int) > (memMergeIn_CTf_f_Int_rbuf,MemIn_CTf_f_Int) */
  MemIn_CTf_f_Int_t memMergeIn_CTf_f_Int_buf;
  assign memMergeIn_CTf_f_Int_r = (! memMergeIn_CTf_f_Int_buf[0]);
  assign memMergeIn_CTf_f_Int_rbuf_d = (memMergeIn_CTf_f_Int_buf[0] ? memMergeIn_CTf_f_Int_buf :
                                        memMergeIn_CTf_f_Int_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memMergeIn_CTf_f_Int_buf <= {180'd0, 1'd0};
    else
      if ((memMergeIn_CTf_f_Int_rbuf_r && memMergeIn_CTf_f_Int_buf[0]))
        memMergeIn_CTf_f_Int_buf <= {180'd0, 1'd0};
      else if (((! memMergeIn_CTf_f_Int_rbuf_r) && (! memMergeIn_CTf_f_Int_buf[0])))
        memMergeIn_CTf_f_Int_buf <= memMergeIn_CTf_f_Int_d;
  
  /* dbuf (Ty MemOut_CTf_f_Int) : (memOut_CTf_f_Int_rbuf,MemOut_CTf_f_Int) > (memOut_CTf_f_Int_dbuf,MemOut_CTf_f_Int) */
  assign memOut_CTf_f_Int_rbuf_r = ((! memOut_CTf_f_Int_dbuf_d[0]) || memOut_CTf_f_Int_dbuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memOut_CTf_f_Int_dbuf_d <= {164'd0, 1'd0};
    else
      if (memOut_CTf_f_Int_rbuf_r)
        memOut_CTf_f_Int_dbuf_d <= memOut_CTf_f_Int_rbuf_d;
  
  /* rbuf (Ty MemOut_CTf_f_Int) : (memOut_CTf_f_Int,MemOut_CTf_f_Int) > (memOut_CTf_f_Int_rbuf,MemOut_CTf_f_Int) */
  MemOut_CTf_f_Int_t memOut_CTf_f_Int_buf;
  assign memOut_CTf_f_Int_r = (! memOut_CTf_f_Int_buf[0]);
  assign memOut_CTf_f_Int_rbuf_d = (memOut_CTf_f_Int_buf[0] ? memOut_CTf_f_Int_buf :
                                    memOut_CTf_f_Int_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memOut_CTf_f_Int_buf <= {164'd0, 1'd0};
    else
      if ((memOut_CTf_f_Int_rbuf_r && memOut_CTf_f_Int_buf[0]))
        memOut_CTf_f_Int_buf <= {164'd0, 1'd0};
      else if (((! memOut_CTf_f_Int_rbuf_r) && (! memOut_CTf_f_Int_buf[0])))
        memOut_CTf_f_Int_buf <= memOut_CTf_f_Int_d;
  
  /* destruct (Ty Pointer_CTf_f_Int,
          Dcon Pointer_CTf_f_Int) : (scfarg_0_2_1_argbuf,Pointer_CTf_f_Int) > [(destructReadIn_CTf_f_Int,Word16#)] */
  assign destructReadIn_CTf_f_Int_d = {scfarg_0_2_1_argbuf_d[16:1],
                                       scfarg_0_2_1_argbuf_d[0]};
  assign scfarg_0_2_1_argbuf_r = destructReadIn_CTf_f_Int_r;
  
  /* dcon (Ty MemIn_CTf_f_Int,
      Dcon ReadIn_CTf_f_Int) : [(destructReadIn_CTf_f_Int,Word16#)] > (dconReadIn_CTf_f_Int,MemIn_CTf_f_Int) */
  assign dconReadIn_CTf_f_Int_d = ReadIn_CTf_f_Int_dc((& {destructReadIn_CTf_f_Int_d[0]}), destructReadIn_CTf_f_Int_d);
  assign {destructReadIn_CTf_f_Int_r} = {1 {(dconReadIn_CTf_f_Int_r && dconReadIn_CTf_f_Int_d[0])}};
  
  /* destruct (Ty MemOut_CTf_f_Int,
          Dcon ReadOut_CTf_f_Int) : (memReadOut_CTf_f_Int,MemOut_CTf_f_Int) > [(readPointer_CTf_f_Intscfarg_0_2_1_argbuf,CTf_f_Int)] */
  assign readPointer_CTf_f_Intscfarg_0_2_1_argbuf_d = {memReadOut_CTf_f_Int_d[164:2],
                                                       memReadOut_CTf_f_Int_d[0]};
  assign memReadOut_CTf_f_Int_r = readPointer_CTf_f_Intscfarg_0_2_1_argbuf_r;
  
  /* mergectrl (Ty C5,Ty CTf_f_Int) : [(lizzieLet52_1_argbuf,CTf_f_Int),
                                  (lizzieLet57_1_argbuf,CTf_f_Int),
                                  (lizzieLet68_1_argbuf,CTf_f_Int),
                                  (lizzieLet69_1_argbuf,CTf_f_Int),
                                  (lizzieLet70_1_argbuf,CTf_f_Int)] > (writeMerge_choice_CTf_f_Int,C5) (writeMerge_data_CTf_f_Int,CTf_f_Int) */
  logic [4:0] lizzieLet52_1_argbuf_select_d;
  assign lizzieLet52_1_argbuf_select_d = ((| lizzieLet52_1_argbuf_select_q) ? lizzieLet52_1_argbuf_select_q :
                                          (lizzieLet52_1_argbuf_d[0] ? 5'd1 :
                                           (lizzieLet57_1_argbuf_d[0] ? 5'd2 :
                                            (lizzieLet68_1_argbuf_d[0] ? 5'd4 :
                                             (lizzieLet69_1_argbuf_d[0] ? 5'd8 :
                                              (lizzieLet70_1_argbuf_d[0] ? 5'd16 :
                                               5'd0))))));
  logic [4:0] lizzieLet52_1_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet52_1_argbuf_select_q <= 5'd0;
    else
      lizzieLet52_1_argbuf_select_q <= (lizzieLet52_1_argbuf_done ? 5'd0 :
                                        lizzieLet52_1_argbuf_select_d);
  logic [1:0] lizzieLet52_1_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet52_1_argbuf_emit_q <= 2'd0;
    else
      lizzieLet52_1_argbuf_emit_q <= (lizzieLet52_1_argbuf_done ? 2'd0 :
                                      lizzieLet52_1_argbuf_emit_d);
  logic [1:0] lizzieLet52_1_argbuf_emit_d;
  assign lizzieLet52_1_argbuf_emit_d = (lizzieLet52_1_argbuf_emit_q | ({writeMerge_choice_CTf_f_Int_d[0],
                                                                        writeMerge_data_CTf_f_Int_d[0]} & {writeMerge_choice_CTf_f_Int_r,
                                                                                                           writeMerge_data_CTf_f_Int_r}));
  logic lizzieLet52_1_argbuf_done;
  assign lizzieLet52_1_argbuf_done = (& lizzieLet52_1_argbuf_emit_d);
  assign {lizzieLet70_1_argbuf_r,
          lizzieLet69_1_argbuf_r,
          lizzieLet68_1_argbuf_r,
          lizzieLet57_1_argbuf_r,
          lizzieLet52_1_argbuf_r} = (lizzieLet52_1_argbuf_done ? lizzieLet52_1_argbuf_select_d :
                                     5'd0);
  assign writeMerge_data_CTf_f_Int_d = ((lizzieLet52_1_argbuf_select_d[0] && (! lizzieLet52_1_argbuf_emit_q[0])) ? lizzieLet52_1_argbuf_d :
                                        ((lizzieLet52_1_argbuf_select_d[1] && (! lizzieLet52_1_argbuf_emit_q[0])) ? lizzieLet57_1_argbuf_d :
                                         ((lizzieLet52_1_argbuf_select_d[2] && (! lizzieLet52_1_argbuf_emit_q[0])) ? lizzieLet68_1_argbuf_d :
                                          ((lizzieLet52_1_argbuf_select_d[3] && (! lizzieLet52_1_argbuf_emit_q[0])) ? lizzieLet69_1_argbuf_d :
                                           ((lizzieLet52_1_argbuf_select_d[4] && (! lizzieLet52_1_argbuf_emit_q[0])) ? lizzieLet70_1_argbuf_d :
                                            {163'd0, 1'd0})))));
  assign writeMerge_choice_CTf_f_Int_d = ((lizzieLet52_1_argbuf_select_d[0] && (! lizzieLet52_1_argbuf_emit_q[1])) ? C1_5_dc(1'd1) :
                                          ((lizzieLet52_1_argbuf_select_d[1] && (! lizzieLet52_1_argbuf_emit_q[1])) ? C2_5_dc(1'd1) :
                                           ((lizzieLet52_1_argbuf_select_d[2] && (! lizzieLet52_1_argbuf_emit_q[1])) ? C3_5_dc(1'd1) :
                                            ((lizzieLet52_1_argbuf_select_d[3] && (! lizzieLet52_1_argbuf_emit_q[1])) ? C4_5_dc(1'd1) :
                                             ((lizzieLet52_1_argbuf_select_d[4] && (! lizzieLet52_1_argbuf_emit_q[1])) ? C5_5_dc(1'd1) :
                                              {3'd0, 1'd0})))));
  
  /* demux (Ty C5,
       Ty Pointer_CTf_f_Int) : (writeMerge_choice_CTf_f_Int,C5) (demuxWriteResult_CTf_f_Int,Pointer_CTf_f_Int) > [(writeCTf_f_IntlizzieLet52_1_argbuf,Pointer_CTf_f_Int),
                                                                                                                  (writeCTf_f_IntlizzieLet57_1_argbuf,Pointer_CTf_f_Int),
                                                                                                                  (writeCTf_f_IntlizzieLet68_1_argbuf,Pointer_CTf_f_Int),
                                                                                                                  (writeCTf_f_IntlizzieLet69_1_argbuf,Pointer_CTf_f_Int),
                                                                                                                  (writeCTf_f_IntlizzieLet70_1_argbuf,Pointer_CTf_f_Int)] */
  logic [4:0] demuxWriteResult_CTf_f_Int_onehotd;
  always_comb
    if ((writeMerge_choice_CTf_f_Int_d[0] && demuxWriteResult_CTf_f_Int_d[0]))
      unique case (writeMerge_choice_CTf_f_Int_d[3:1])
        3'd0: demuxWriteResult_CTf_f_Int_onehotd = 5'd1;
        3'd1: demuxWriteResult_CTf_f_Int_onehotd = 5'd2;
        3'd2: demuxWriteResult_CTf_f_Int_onehotd = 5'd4;
        3'd3: demuxWriteResult_CTf_f_Int_onehotd = 5'd8;
        3'd4: demuxWriteResult_CTf_f_Int_onehotd = 5'd16;
        default: demuxWriteResult_CTf_f_Int_onehotd = 5'd0;
      endcase
    else demuxWriteResult_CTf_f_Int_onehotd = 5'd0;
  assign writeCTf_f_IntlizzieLet52_1_argbuf_d = {demuxWriteResult_CTf_f_Int_d[16:1],
                                                 demuxWriteResult_CTf_f_Int_onehotd[0]};
  assign writeCTf_f_IntlizzieLet57_1_argbuf_d = {demuxWriteResult_CTf_f_Int_d[16:1],
                                                 demuxWriteResult_CTf_f_Int_onehotd[1]};
  assign writeCTf_f_IntlizzieLet68_1_argbuf_d = {demuxWriteResult_CTf_f_Int_d[16:1],
                                                 demuxWriteResult_CTf_f_Int_onehotd[2]};
  assign writeCTf_f_IntlizzieLet69_1_argbuf_d = {demuxWriteResult_CTf_f_Int_d[16:1],
                                                 demuxWriteResult_CTf_f_Int_onehotd[3]};
  assign writeCTf_f_IntlizzieLet70_1_argbuf_d = {demuxWriteResult_CTf_f_Int_d[16:1],
                                                 demuxWriteResult_CTf_f_Int_onehotd[4]};
  assign demuxWriteResult_CTf_f_Int_r = (| (demuxWriteResult_CTf_f_Int_onehotd & {writeCTf_f_IntlizzieLet70_1_argbuf_r,
                                                                                  writeCTf_f_IntlizzieLet69_1_argbuf_r,
                                                                                  writeCTf_f_IntlizzieLet68_1_argbuf_r,
                                                                                  writeCTf_f_IntlizzieLet57_1_argbuf_r,
                                                                                  writeCTf_f_IntlizzieLet52_1_argbuf_r}));
  assign writeMerge_choice_CTf_f_Int_r = demuxWriteResult_CTf_f_Int_r;
  
  /* dcon (Ty MemIn_CTf_f_Int,
      Dcon WriteIn_CTf_f_Int) : [(forkHP1_CTf_f_In2,Word16#),
                                 (writeMerge_data_CTf_f_Int,CTf_f_Int)] > (dconWriteIn_CTf_f_Int,MemIn_CTf_f_Int) */
  assign dconWriteIn_CTf_f_Int_d = WriteIn_CTf_f_Int_dc((& {forkHP1_CTf_f_In2_d[0],
                                                            writeMerge_data_CTf_f_Int_d[0]}), forkHP1_CTf_f_In2_d, writeMerge_data_CTf_f_Int_d);
  assign {forkHP1_CTf_f_In2_r,
          writeMerge_data_CTf_f_Int_r} = {2 {(dconWriteIn_CTf_f_Int_r && dconWriteIn_CTf_f_Int_d[0])}};
  
  /* dcon (Ty Pointer_CTf_f_Int,
      Dcon Pointer_CTf_f_Int) : [(forkHP1_CTf_f_In3,Word16#)] > (dconPtr_CTf_f_Int,Pointer_CTf_f_Int) */
  assign dconPtr_CTf_f_Int_d = Pointer_CTf_f_Int_dc((& {forkHP1_CTf_f_In3_d[0]}), forkHP1_CTf_f_In3_d);
  assign {forkHP1_CTf_f_In3_r} = {1 {(dconPtr_CTf_f_Int_r && dconPtr_CTf_f_Int_d[0])}};
  
  /* demux (Ty MemOut_CTf_f_Int,
       Ty Pointer_CTf_f_Int) : (memWriteOut_CTf_f_Int,MemOut_CTf_f_Int) (dconPtr_CTf_f_Int,Pointer_CTf_f_Int) > [(_256,Pointer_CTf_f_Int),
                                                                                                                 (demuxWriteResult_CTf_f_Int,Pointer_CTf_f_Int)] */
  logic [1:0] dconPtr_CTf_f_Int_onehotd;
  always_comb
    if ((memWriteOut_CTf_f_Int_d[0] && dconPtr_CTf_f_Int_d[0]))
      unique case (memWriteOut_CTf_f_Int_d[1:1])
        1'd0: dconPtr_CTf_f_Int_onehotd = 2'd1;
        1'd1: dconPtr_CTf_f_Int_onehotd = 2'd2;
        default: dconPtr_CTf_f_Int_onehotd = 2'd0;
      endcase
    else dconPtr_CTf_f_Int_onehotd = 2'd0;
  assign _256_d = {dconPtr_CTf_f_Int_d[16:1],
                   dconPtr_CTf_f_Int_onehotd[0]};
  assign demuxWriteResult_CTf_f_Int_d = {dconPtr_CTf_f_Int_d[16:1],
                                         dconPtr_CTf_f_Int_onehotd[1]};
  assign dconPtr_CTf_f_Int_r = (| (dconPtr_CTf_f_Int_onehotd & {demuxWriteResult_CTf_f_Int_r,
                                                                _256_r}));
  assign memWriteOut_CTf_f_Int_r = dconPtr_CTf_f_Int_r;
  
  /* source (Ty Go) : > (sourceGo,Go) */
  
  /* source (Ty Pointer_QTree_Int) : > (m1aen_0,Pointer_QTree_Int) */
  
  /* source (Ty Pointer_QTree_Int) : > (m2aeo_1,Pointer_QTree_Int) */
  
  /* source (Ty Pointer_QTree_Int) : > (m3aep_2,Pointer_QTree_Int) */
  
  /* destruct (Ty TupGo___Pointer_QTree_Int,
          Dcon TupGo___Pointer_QTree_Int) : ($wnnzTupGo___Pointer_QTree_Int_1,TupGo___Pointer_QTree_Int) > [($wnnzTupGo___Pointer_QTree_Intgo_6,Go),
                                                                                                            ($wnnzTupGo___Pointer_QTree_Intwsmk,Pointer_QTree_Int)] */
  logic [1:0] \$wnnzTupGo___Pointer_QTree_Int_1_emitted ;
  logic [1:0] \$wnnzTupGo___Pointer_QTree_Int_1_done ;
  assign \$wnnzTupGo___Pointer_QTree_Intgo_6_d  = (\$wnnzTupGo___Pointer_QTree_Int_1_d [0] && (! \$wnnzTupGo___Pointer_QTree_Int_1_emitted [0]));
  assign \$wnnzTupGo___Pointer_QTree_Intwsmk_d  = {\$wnnzTupGo___Pointer_QTree_Int_1_d [16:1],
                                                   (\$wnnzTupGo___Pointer_QTree_Int_1_d [0] && (! \$wnnzTupGo___Pointer_QTree_Int_1_emitted [1]))};
  assign \$wnnzTupGo___Pointer_QTree_Int_1_done  = (\$wnnzTupGo___Pointer_QTree_Int_1_emitted  | ({\$wnnzTupGo___Pointer_QTree_Intwsmk_d [0],
                                                                                                   \$wnnzTupGo___Pointer_QTree_Intgo_6_d [0]} & {\$wnnzTupGo___Pointer_QTree_Intwsmk_r ,
                                                                                                                                                 \$wnnzTupGo___Pointer_QTree_Intgo_6_r }));
  assign \$wnnzTupGo___Pointer_QTree_Int_1_r  = (& \$wnnzTupGo___Pointer_QTree_Int_1_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \$wnnzTupGo___Pointer_QTree_Int_1_emitted  <= 2'd0;
    else
      \$wnnzTupGo___Pointer_QTree_Int_1_emitted  <= (\$wnnzTupGo___Pointer_QTree_Int_1_r  ? 2'd0 :
                                                     \$wnnzTupGo___Pointer_QTree_Int_1_done );
  
  /* fork (Ty Go) : ($wnnzTupGo___Pointer_QTree_Intgo_6,Go) > [(go_6_1,Go),
                                                          (go_6_2,Go)] */
  logic [1:0] \$wnnzTupGo___Pointer_QTree_Intgo_6_emitted ;
  logic [1:0] \$wnnzTupGo___Pointer_QTree_Intgo_6_done ;
  assign go_6_1_d = (\$wnnzTupGo___Pointer_QTree_Intgo_6_d [0] && (! \$wnnzTupGo___Pointer_QTree_Intgo_6_emitted [0]));
  assign go_6_2_d = (\$wnnzTupGo___Pointer_QTree_Intgo_6_d [0] && (! \$wnnzTupGo___Pointer_QTree_Intgo_6_emitted [1]));
  assign \$wnnzTupGo___Pointer_QTree_Intgo_6_done  = (\$wnnzTupGo___Pointer_QTree_Intgo_6_emitted  | ({go_6_2_d[0],
                                                                                                       go_6_1_d[0]} & {go_6_2_r,
                                                                                                                       go_6_1_r}));
  assign \$wnnzTupGo___Pointer_QTree_Intgo_6_r  = (& \$wnnzTupGo___Pointer_QTree_Intgo_6_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \$wnnzTupGo___Pointer_QTree_Intgo_6_emitted  <= 2'd0;
    else
      \$wnnzTupGo___Pointer_QTree_Intgo_6_emitted  <= (\$wnnzTupGo___Pointer_QTree_Intgo_6_r  ? 2'd0 :
                                                       \$wnnzTupGo___Pointer_QTree_Intgo_6_done );
  
  /* buf (Ty Pointer_QTree_Int) : ($wnnzTupGo___Pointer_QTree_Intwsmk,Pointer_QTree_Int) > (wsmk_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t \$wnnzTupGo___Pointer_QTree_Intwsmk_bufchan_d ;
  logic \$wnnzTupGo___Pointer_QTree_Intwsmk_bufchan_r ;
  assign \$wnnzTupGo___Pointer_QTree_Intwsmk_r  = ((! \$wnnzTupGo___Pointer_QTree_Intwsmk_bufchan_d [0]) || \$wnnzTupGo___Pointer_QTree_Intwsmk_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \$wnnzTupGo___Pointer_QTree_Intwsmk_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\$wnnzTupGo___Pointer_QTree_Intwsmk_r )
        \$wnnzTupGo___Pointer_QTree_Intwsmk_bufchan_d  <= \$wnnzTupGo___Pointer_QTree_Intwsmk_d ;
  Pointer_QTree_Int_t \$wnnzTupGo___Pointer_QTree_Intwsmk_bufchan_buf ;
  assign \$wnnzTupGo___Pointer_QTree_Intwsmk_bufchan_r  = (! \$wnnzTupGo___Pointer_QTree_Intwsmk_bufchan_buf [0]);
  assign wsmk_1_argbuf_d = (\$wnnzTupGo___Pointer_QTree_Intwsmk_bufchan_buf [0] ? \$wnnzTupGo___Pointer_QTree_Intwsmk_bufchan_buf  :
                            \$wnnzTupGo___Pointer_QTree_Intwsmk_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \$wnnzTupGo___Pointer_QTree_Intwsmk_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((wsmk_1_argbuf_r && \$wnnzTupGo___Pointer_QTree_Intwsmk_bufchan_buf [0]))
        \$wnnzTupGo___Pointer_QTree_Intwsmk_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! wsmk_1_argbuf_r) && (! \$wnnzTupGo___Pointer_QTree_Intwsmk_bufchan_buf [0])))
        \$wnnzTupGo___Pointer_QTree_Intwsmk_bufchan_buf  <= \$wnnzTupGo___Pointer_QTree_Intwsmk_bufchan_d ;
  
  /* dcon (Ty Int,Dcon I#) : [($wnnz_resbuf,Int#)] > (es_6_1I#,Int) */
  assign \es_6_1I#_d  = \I#_dc ((& {\$wnnz_resbuf_d [0]}), \$wnnz_resbuf_d );
  assign {\$wnnz_resbuf_r } = {1 {(\es_6_1I#_r  && \es_6_1I#_d [0])}};
  
  /* mergectrl (Ty C5,
           Ty TupGo___MyDTInt_Bool___Int) : [(applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1,TupGo___MyDTInt_Bool___Int),
                                             (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int2,TupGo___MyDTInt_Bool___Int),
                                             (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int3,TupGo___MyDTInt_Bool___Int),
                                             (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int4,TupGo___MyDTInt_Bool___Int),
                                             (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int5,TupGo___MyDTInt_Bool___Int)] > (applyfnInt_Bool_5_choice,C5) (applyfnInt_Bool_5_data,TupGo___MyDTInt_Bool___Int) */
  logic [4:0] applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_select_d;
  assign applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_select_d = ((| applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_select_q) ? applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_select_q :
                                                                   (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_d[0] ? 5'd1 :
                                                                    (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int2_d[0] ? 5'd2 :
                                                                     (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int3_d[0] ? 5'd4 :
                                                                      (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int4_d[0] ? 5'd8 :
                                                                       (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int5_d[0] ? 5'd16 :
                                                                        5'd0))))));
  logic [4:0] applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_select_q <= 5'd0;
    else
      applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_select_q <= (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_done ? 5'd0 :
                                                                 applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_select_d);
  logic [1:0] applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_emit_q <= 2'd0;
    else
      applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_emit_q <= (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_done ? 2'd0 :
                                                               applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_emit_d);
  logic [1:0] applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_emit_d;
  assign applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_emit_d = (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_emit_q | ({applyfnInt_Bool_5_choice_d[0],
                                                                                                                          applyfnInt_Bool_5_data_d[0]} & {applyfnInt_Bool_5_choice_r,
                                                                                                                                                          applyfnInt_Bool_5_data_r}));
  logic applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_done;
  assign applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_done = (& applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_emit_d);
  assign {applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int5_r,
          applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int4_r,
          applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int3_r,
          applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int2_r,
          applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_r} = (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_done ? applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_select_d :
                                                              5'd0);
  assign applyfnInt_Bool_5_data_d = ((applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_select_d[0] && (! applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_emit_q[0])) ? applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_d :
                                     ((applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_select_d[1] && (! applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_emit_q[0])) ? applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int2_d :
                                      ((applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_select_d[2] && (! applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_emit_q[0])) ? applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int3_d :
                                       ((applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_select_d[3] && (! applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_emit_q[0])) ? applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int4_d :
                                        ((applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_select_d[4] && (! applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_emit_q[0])) ? applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int5_d :
                                         {32'd0, 1'd0})))));
  assign applyfnInt_Bool_5_choice_d = ((applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_select_d[0] && (! applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_emit_q[1])) ? C1_5_dc(1'd1) :
                                       ((applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_select_d[1] && (! applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_emit_q[1])) ? C2_5_dc(1'd1) :
                                        ((applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_select_d[2] && (! applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_emit_q[1])) ? C3_5_dc(1'd1) :
                                         ((applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_select_d[3] && (! applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_emit_q[1])) ? C4_5_dc(1'd1) :
                                          ((applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_select_d[4] && (! applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_emit_q[1])) ? C5_5_dc(1'd1) :
                                           {3'd0, 1'd0})))));
  
  /* fork (Ty MyDTInt_Bool) : (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0,MyDTInt_Bool) > [(arg0_1,MyDTInt_Bool),
                                                                                           (arg0_2,MyDTInt_Bool),
                                                                                           (arg0_3,MyDTInt_Bool)] */
  logic [2:0] applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_emitted;
  logic [2:0] applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_done;
  assign arg0_1_d = (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_d[0] && (! applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_emitted[0]));
  assign arg0_2_d = (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_d[0] && (! applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_emitted[1]));
  assign arg0_3_d = (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_d[0] && (! applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_emitted[2]));
  assign applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_done = (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_emitted | ({arg0_3_d[0],
                                                                                                                             arg0_2_d[0],
                                                                                                                             arg0_1_d[0]} & {arg0_3_r,
                                                                                                                                             arg0_2_r,
                                                                                                                                             arg0_1_r}));
  assign applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_r = (& applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_emitted <= 3'd0;
    else
      applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_emitted <= (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_r ? 3'd0 :
                                                                  applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_done);
  
  /* buf (Ty MyBool) : (applyfnInt_Bool_5_1,MyBool) > (applyfnInt_Bool_5_resbuf,MyBool) */
  MyBool_t applyfnInt_Bool_5_1_bufchan_d;
  logic applyfnInt_Bool_5_1_bufchan_r;
  assign applyfnInt_Bool_5_1_r = ((! applyfnInt_Bool_5_1_bufchan_d[0]) || applyfnInt_Bool_5_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) applyfnInt_Bool_5_1_bufchan_d <= {1'd0, 1'd0};
    else
      if (applyfnInt_Bool_5_1_r)
        applyfnInt_Bool_5_1_bufchan_d <= applyfnInt_Bool_5_1_d;
  MyBool_t applyfnInt_Bool_5_1_bufchan_buf;
  assign applyfnInt_Bool_5_1_bufchan_r = (! applyfnInt_Bool_5_1_bufchan_buf[0]);
  assign applyfnInt_Bool_5_resbuf_d = (applyfnInt_Bool_5_1_bufchan_buf[0] ? applyfnInt_Bool_5_1_bufchan_buf :
                                       applyfnInt_Bool_5_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Bool_5_1_bufchan_buf <= {1'd0, 1'd0};
    else
      if ((applyfnInt_Bool_5_resbuf_r && applyfnInt_Bool_5_1_bufchan_buf[0]))
        applyfnInt_Bool_5_1_bufchan_buf <= {1'd0, 1'd0};
      else if (((! applyfnInt_Bool_5_resbuf_r) && (! applyfnInt_Bool_5_1_bufchan_buf[0])))
        applyfnInt_Bool_5_1_bufchan_buf <= applyfnInt_Bool_5_1_bufchan_d;
  
  /* buf (Ty MyBool) : (applyfnInt_Bool_5_2,MyBool) > (applyfnInt_Bool_5_2_argbuf,MyBool) */
  MyBool_t applyfnInt_Bool_5_2_bufchan_d;
  logic applyfnInt_Bool_5_2_bufchan_r;
  assign applyfnInt_Bool_5_2_r = ((! applyfnInt_Bool_5_2_bufchan_d[0]) || applyfnInt_Bool_5_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) applyfnInt_Bool_5_2_bufchan_d <= {1'd0, 1'd0};
    else
      if (applyfnInt_Bool_5_2_r)
        applyfnInt_Bool_5_2_bufchan_d <= applyfnInt_Bool_5_2_d;
  MyBool_t applyfnInt_Bool_5_2_bufchan_buf;
  assign applyfnInt_Bool_5_2_bufchan_r = (! applyfnInt_Bool_5_2_bufchan_buf[0]);
  assign applyfnInt_Bool_5_2_argbuf_d = (applyfnInt_Bool_5_2_bufchan_buf[0] ? applyfnInt_Bool_5_2_bufchan_buf :
                                         applyfnInt_Bool_5_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Bool_5_2_bufchan_buf <= {1'd0, 1'd0};
    else
      if ((applyfnInt_Bool_5_2_argbuf_r && applyfnInt_Bool_5_2_bufchan_buf[0]))
        applyfnInt_Bool_5_2_bufchan_buf <= {1'd0, 1'd0};
      else if (((! applyfnInt_Bool_5_2_argbuf_r) && (! applyfnInt_Bool_5_2_bufchan_buf[0])))
        applyfnInt_Bool_5_2_bufchan_buf <= applyfnInt_Bool_5_2_bufchan_d;
  
  /* fork (Ty MyBool) : (applyfnInt_Bool_5_2_argbuf,MyBool) > [(es_2_1,MyBool),
                                                          (es_2_2,MyBool),
                                                          (es_2_3,MyBool),
                                                          (es_2_4,MyBool),
                                                          (es_2_5,MyBool)] */
  logic [4:0] applyfnInt_Bool_5_2_argbuf_emitted;
  logic [4:0] applyfnInt_Bool_5_2_argbuf_done;
  assign es_2_1_d = {applyfnInt_Bool_5_2_argbuf_d[1:1],
                     (applyfnInt_Bool_5_2_argbuf_d[0] && (! applyfnInt_Bool_5_2_argbuf_emitted[0]))};
  assign es_2_2_d = {applyfnInt_Bool_5_2_argbuf_d[1:1],
                     (applyfnInt_Bool_5_2_argbuf_d[0] && (! applyfnInt_Bool_5_2_argbuf_emitted[1]))};
  assign es_2_3_d = {applyfnInt_Bool_5_2_argbuf_d[1:1],
                     (applyfnInt_Bool_5_2_argbuf_d[0] && (! applyfnInt_Bool_5_2_argbuf_emitted[2]))};
  assign es_2_4_d = {applyfnInt_Bool_5_2_argbuf_d[1:1],
                     (applyfnInt_Bool_5_2_argbuf_d[0] && (! applyfnInt_Bool_5_2_argbuf_emitted[3]))};
  assign es_2_5_d = {applyfnInt_Bool_5_2_argbuf_d[1:1],
                     (applyfnInt_Bool_5_2_argbuf_d[0] && (! applyfnInt_Bool_5_2_argbuf_emitted[4]))};
  assign applyfnInt_Bool_5_2_argbuf_done = (applyfnInt_Bool_5_2_argbuf_emitted | ({es_2_5_d[0],
                                                                                   es_2_4_d[0],
                                                                                   es_2_3_d[0],
                                                                                   es_2_2_d[0],
                                                                                   es_2_1_d[0]} & {es_2_5_r,
                                                                                                   es_2_4_r,
                                                                                                   es_2_3_r,
                                                                                                   es_2_2_r,
                                                                                                   es_2_1_r}));
  assign applyfnInt_Bool_5_2_argbuf_r = (& applyfnInt_Bool_5_2_argbuf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) applyfnInt_Bool_5_2_argbuf_emitted <= 5'd0;
    else
      applyfnInt_Bool_5_2_argbuf_emitted <= (applyfnInt_Bool_5_2_argbuf_r ? 5'd0 :
                                             applyfnInt_Bool_5_2_argbuf_done);
  
  /* buf (Ty MyBool) : (applyfnInt_Bool_5_3,MyBool) > (applyfnInt_Bool_5_3_argbuf,MyBool) */
  MyBool_t applyfnInt_Bool_5_3_bufchan_d;
  logic applyfnInt_Bool_5_3_bufchan_r;
  assign applyfnInt_Bool_5_3_r = ((! applyfnInt_Bool_5_3_bufchan_d[0]) || applyfnInt_Bool_5_3_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) applyfnInt_Bool_5_3_bufchan_d <= {1'd0, 1'd0};
    else
      if (applyfnInt_Bool_5_3_r)
        applyfnInt_Bool_5_3_bufchan_d <= applyfnInt_Bool_5_3_d;
  MyBool_t applyfnInt_Bool_5_3_bufchan_buf;
  assign applyfnInt_Bool_5_3_bufchan_r = (! applyfnInt_Bool_5_3_bufchan_buf[0]);
  assign applyfnInt_Bool_5_3_argbuf_d = (applyfnInt_Bool_5_3_bufchan_buf[0] ? applyfnInt_Bool_5_3_bufchan_buf :
                                         applyfnInt_Bool_5_3_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Bool_5_3_bufchan_buf <= {1'd0, 1'd0};
    else
      if ((applyfnInt_Bool_5_3_argbuf_r && applyfnInt_Bool_5_3_bufchan_buf[0]))
        applyfnInt_Bool_5_3_bufchan_buf <= {1'd0, 1'd0};
      else if (((! applyfnInt_Bool_5_3_argbuf_r) && (! applyfnInt_Bool_5_3_bufchan_buf[0])))
        applyfnInt_Bool_5_3_bufchan_buf <= applyfnInt_Bool_5_3_bufchan_d;
  
  /* fork (Ty MyBool) : (applyfnInt_Bool_5_3_argbuf,MyBool) > [(es_10_1,MyBool),
                                                          (es_10_2,MyBool),
                                                          (es_10_3,MyBool),
                                                          (es_10_4,MyBool),
                                                          (es_10_5,MyBool)] */
  logic [4:0] applyfnInt_Bool_5_3_argbuf_emitted;
  logic [4:0] applyfnInt_Bool_5_3_argbuf_done;
  assign es_10_1_d = {applyfnInt_Bool_5_3_argbuf_d[1:1],
                      (applyfnInt_Bool_5_3_argbuf_d[0] && (! applyfnInt_Bool_5_3_argbuf_emitted[0]))};
  assign es_10_2_d = {applyfnInt_Bool_5_3_argbuf_d[1:1],
                      (applyfnInt_Bool_5_3_argbuf_d[0] && (! applyfnInt_Bool_5_3_argbuf_emitted[1]))};
  assign es_10_3_d = {applyfnInt_Bool_5_3_argbuf_d[1:1],
                      (applyfnInt_Bool_5_3_argbuf_d[0] && (! applyfnInt_Bool_5_3_argbuf_emitted[2]))};
  assign es_10_4_d = {applyfnInt_Bool_5_3_argbuf_d[1:1],
                      (applyfnInt_Bool_5_3_argbuf_d[0] && (! applyfnInt_Bool_5_3_argbuf_emitted[3]))};
  assign es_10_5_d = {applyfnInt_Bool_5_3_argbuf_d[1:1],
                      (applyfnInt_Bool_5_3_argbuf_d[0] && (! applyfnInt_Bool_5_3_argbuf_emitted[4]))};
  assign applyfnInt_Bool_5_3_argbuf_done = (applyfnInt_Bool_5_3_argbuf_emitted | ({es_10_5_d[0],
                                                                                   es_10_4_d[0],
                                                                                   es_10_3_d[0],
                                                                                   es_10_2_d[0],
                                                                                   es_10_1_d[0]} & {es_10_5_r,
                                                                                                    es_10_4_r,
                                                                                                    es_10_3_r,
                                                                                                    es_10_2_r,
                                                                                                    es_10_1_r}));
  assign applyfnInt_Bool_5_3_argbuf_r = (& applyfnInt_Bool_5_3_argbuf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) applyfnInt_Bool_5_3_argbuf_emitted <= 5'd0;
    else
      applyfnInt_Bool_5_3_argbuf_emitted <= (applyfnInt_Bool_5_3_argbuf_r ? 5'd0 :
                                             applyfnInt_Bool_5_3_argbuf_done);
  
  /* buf (Ty MyBool) : (applyfnInt_Bool_5_4,MyBool) > (applyfnInt_Bool_5_4_argbuf,MyBool) */
  MyBool_t applyfnInt_Bool_5_4_bufchan_d;
  logic applyfnInt_Bool_5_4_bufchan_r;
  assign applyfnInt_Bool_5_4_r = ((! applyfnInt_Bool_5_4_bufchan_d[0]) || applyfnInt_Bool_5_4_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) applyfnInt_Bool_5_4_bufchan_d <= {1'd0, 1'd0};
    else
      if (applyfnInt_Bool_5_4_r)
        applyfnInt_Bool_5_4_bufchan_d <= applyfnInt_Bool_5_4_d;
  MyBool_t applyfnInt_Bool_5_4_bufchan_buf;
  assign applyfnInt_Bool_5_4_bufchan_r = (! applyfnInt_Bool_5_4_bufchan_buf[0]);
  assign applyfnInt_Bool_5_4_argbuf_d = (applyfnInt_Bool_5_4_bufchan_buf[0] ? applyfnInt_Bool_5_4_bufchan_buf :
                                         applyfnInt_Bool_5_4_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Bool_5_4_bufchan_buf <= {1'd0, 1'd0};
    else
      if ((applyfnInt_Bool_5_4_argbuf_r && applyfnInt_Bool_5_4_bufchan_buf[0]))
        applyfnInt_Bool_5_4_bufchan_buf <= {1'd0, 1'd0};
      else if (((! applyfnInt_Bool_5_4_argbuf_r) && (! applyfnInt_Bool_5_4_bufchan_buf[0])))
        applyfnInt_Bool_5_4_bufchan_buf <= applyfnInt_Bool_5_4_bufchan_d;
  
  /* fork (Ty MyBool) : (applyfnInt_Bool_5_4_argbuf,MyBool) > [(es_14_1,MyBool),
                                                          (es_14_2,MyBool),
                                                          (es_14_3,MyBool),
                                                          (es_14_4,MyBool),
                                                          (es_14_5,MyBool),
                                                          (es_14_6,MyBool),
                                                          (es_14_7,MyBool),
                                                          (es_14_8,MyBool)] */
  logic [7:0] applyfnInt_Bool_5_4_argbuf_emitted;
  logic [7:0] applyfnInt_Bool_5_4_argbuf_done;
  assign es_14_1_d = {applyfnInt_Bool_5_4_argbuf_d[1:1],
                      (applyfnInt_Bool_5_4_argbuf_d[0] && (! applyfnInt_Bool_5_4_argbuf_emitted[0]))};
  assign es_14_2_d = {applyfnInt_Bool_5_4_argbuf_d[1:1],
                      (applyfnInt_Bool_5_4_argbuf_d[0] && (! applyfnInt_Bool_5_4_argbuf_emitted[1]))};
  assign es_14_3_d = {applyfnInt_Bool_5_4_argbuf_d[1:1],
                      (applyfnInt_Bool_5_4_argbuf_d[0] && (! applyfnInt_Bool_5_4_argbuf_emitted[2]))};
  assign es_14_4_d = {applyfnInt_Bool_5_4_argbuf_d[1:1],
                      (applyfnInt_Bool_5_4_argbuf_d[0] && (! applyfnInt_Bool_5_4_argbuf_emitted[3]))};
  assign es_14_5_d = {applyfnInt_Bool_5_4_argbuf_d[1:1],
                      (applyfnInt_Bool_5_4_argbuf_d[0] && (! applyfnInt_Bool_5_4_argbuf_emitted[4]))};
  assign es_14_6_d = {applyfnInt_Bool_5_4_argbuf_d[1:1],
                      (applyfnInt_Bool_5_4_argbuf_d[0] && (! applyfnInt_Bool_5_4_argbuf_emitted[5]))};
  assign es_14_7_d = {applyfnInt_Bool_5_4_argbuf_d[1:1],
                      (applyfnInt_Bool_5_4_argbuf_d[0] && (! applyfnInt_Bool_5_4_argbuf_emitted[6]))};
  assign es_14_8_d = {applyfnInt_Bool_5_4_argbuf_d[1:1],
                      (applyfnInt_Bool_5_4_argbuf_d[0] && (! applyfnInt_Bool_5_4_argbuf_emitted[7]))};
  assign applyfnInt_Bool_5_4_argbuf_done = (applyfnInt_Bool_5_4_argbuf_emitted | ({es_14_8_d[0],
                                                                                   es_14_7_d[0],
                                                                                   es_14_6_d[0],
                                                                                   es_14_5_d[0],
                                                                                   es_14_4_d[0],
                                                                                   es_14_3_d[0],
                                                                                   es_14_2_d[0],
                                                                                   es_14_1_d[0]} & {es_14_8_r,
                                                                                                    es_14_7_r,
                                                                                                    es_14_6_r,
                                                                                                    es_14_5_r,
                                                                                                    es_14_4_r,
                                                                                                    es_14_3_r,
                                                                                                    es_14_2_r,
                                                                                                    es_14_1_r}));
  assign applyfnInt_Bool_5_4_argbuf_r = (& applyfnInt_Bool_5_4_argbuf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) applyfnInt_Bool_5_4_argbuf_emitted <= 8'd0;
    else
      applyfnInt_Bool_5_4_argbuf_emitted <= (applyfnInt_Bool_5_4_argbuf_r ? 8'd0 :
                                             applyfnInt_Bool_5_4_argbuf_done);
  
  /* buf (Ty MyBool) : (applyfnInt_Bool_5_5,MyBool) > (applyfnInt_Bool_5_5_argbuf,MyBool) */
  MyBool_t applyfnInt_Bool_5_5_bufchan_d;
  logic applyfnInt_Bool_5_5_bufchan_r;
  assign applyfnInt_Bool_5_5_r = ((! applyfnInt_Bool_5_5_bufchan_d[0]) || applyfnInt_Bool_5_5_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) applyfnInt_Bool_5_5_bufchan_d <= {1'd0, 1'd0};
    else
      if (applyfnInt_Bool_5_5_r)
        applyfnInt_Bool_5_5_bufchan_d <= applyfnInt_Bool_5_5_d;
  MyBool_t applyfnInt_Bool_5_5_bufchan_buf;
  assign applyfnInt_Bool_5_5_bufchan_r = (! applyfnInt_Bool_5_5_bufchan_buf[0]);
  assign applyfnInt_Bool_5_5_argbuf_d = (applyfnInt_Bool_5_5_bufchan_buf[0] ? applyfnInt_Bool_5_5_bufchan_buf :
                                         applyfnInt_Bool_5_5_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Bool_5_5_bufchan_buf <= {1'd0, 1'd0};
    else
      if ((applyfnInt_Bool_5_5_argbuf_r && applyfnInt_Bool_5_5_bufchan_buf[0]))
        applyfnInt_Bool_5_5_bufchan_buf <= {1'd0, 1'd0};
      else if (((! applyfnInt_Bool_5_5_argbuf_r) && (! applyfnInt_Bool_5_5_bufchan_buf[0])))
        applyfnInt_Bool_5_5_bufchan_buf <= applyfnInt_Bool_5_5_bufchan_d;
  
  /* fork (Ty MyBool) : (applyfnInt_Bool_5_5_argbuf,MyBool) > [(es_21_1,MyBool),
                                                          (es_21_2,MyBool),
                                                          (es_21_3,MyBool),
                                                          (es_21_4,MyBool),
                                                          (es_21_5,MyBool),
                                                          (es_21_6,MyBool)] */
  logic [5:0] applyfnInt_Bool_5_5_argbuf_emitted;
  logic [5:0] applyfnInt_Bool_5_5_argbuf_done;
  assign es_21_1_d = {applyfnInt_Bool_5_5_argbuf_d[1:1],
                      (applyfnInt_Bool_5_5_argbuf_d[0] && (! applyfnInt_Bool_5_5_argbuf_emitted[0]))};
  assign es_21_2_d = {applyfnInt_Bool_5_5_argbuf_d[1:1],
                      (applyfnInt_Bool_5_5_argbuf_d[0] && (! applyfnInt_Bool_5_5_argbuf_emitted[1]))};
  assign es_21_3_d = {applyfnInt_Bool_5_5_argbuf_d[1:1],
                      (applyfnInt_Bool_5_5_argbuf_d[0] && (! applyfnInt_Bool_5_5_argbuf_emitted[2]))};
  assign es_21_4_d = {applyfnInt_Bool_5_5_argbuf_d[1:1],
                      (applyfnInt_Bool_5_5_argbuf_d[0] && (! applyfnInt_Bool_5_5_argbuf_emitted[3]))};
  assign es_21_5_d = {applyfnInt_Bool_5_5_argbuf_d[1:1],
                      (applyfnInt_Bool_5_5_argbuf_d[0] && (! applyfnInt_Bool_5_5_argbuf_emitted[4]))};
  assign es_21_6_d = {applyfnInt_Bool_5_5_argbuf_d[1:1],
                      (applyfnInt_Bool_5_5_argbuf_d[0] && (! applyfnInt_Bool_5_5_argbuf_emitted[5]))};
  assign applyfnInt_Bool_5_5_argbuf_done = (applyfnInt_Bool_5_5_argbuf_emitted | ({es_21_6_d[0],
                                                                                   es_21_5_d[0],
                                                                                   es_21_4_d[0],
                                                                                   es_21_3_d[0],
                                                                                   es_21_2_d[0],
                                                                                   es_21_1_d[0]} & {es_21_6_r,
                                                                                                    es_21_5_r,
                                                                                                    es_21_4_r,
                                                                                                    es_21_3_r,
                                                                                                    es_21_2_r,
                                                                                                    es_21_1_r}));
  assign applyfnInt_Bool_5_5_argbuf_r = (& applyfnInt_Bool_5_5_argbuf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) applyfnInt_Bool_5_5_argbuf_emitted <= 6'd0;
    else
      applyfnInt_Bool_5_5_argbuf_emitted <= (applyfnInt_Bool_5_5_argbuf_r ? 6'd0 :
                                             applyfnInt_Bool_5_5_argbuf_done);
  
  /* demux (Ty C5,
       Ty MyBool) : (applyfnInt_Bool_5_choice,C5) (lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux,MyBool) > [(applyfnInt_Bool_5_1,MyBool),
                                                                                                                                 (applyfnInt_Bool_5_2,MyBool),
                                                                                                                                 (applyfnInt_Bool_5_3,MyBool),
                                                                                                                                 (applyfnInt_Bool_5_4,MyBool),
                                                                                                                                 (applyfnInt_Bool_5_5,MyBool)] */
  logic [4:0] lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_onehotd;
  always_comb
    if ((applyfnInt_Bool_5_choice_d[0] && lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_d[0]))
      unique case (applyfnInt_Bool_5_choice_d[3:1])
        3'd0:
          lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_onehotd = 5'd1;
        3'd1:
          lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_onehotd = 5'd2;
        3'd2:
          lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_onehotd = 5'd4;
        3'd3:
          lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_onehotd = 5'd8;
        3'd4:
          lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_onehotd = 5'd16;
        default:
          lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_onehotd = 5'd0;
      endcase
    else
      lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_onehotd = 5'd0;
  assign applyfnInt_Bool_5_1_d = {lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_d[1:1],
                                  lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_onehotd[0]};
  assign applyfnInt_Bool_5_2_d = {lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_d[1:1],
                                  lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_onehotd[1]};
  assign applyfnInt_Bool_5_3_d = {lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_d[1:1],
                                  lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_onehotd[2]};
  assign applyfnInt_Bool_5_4_d = {lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_d[1:1],
                                  lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_onehotd[3]};
  assign applyfnInt_Bool_5_5_d = {lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_d[1:1],
                                  lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_onehotd[4]};
  assign lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_r = (| (lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_onehotd & {applyfnInt_Bool_5_5_r,
                                                                                                                                                                  applyfnInt_Bool_5_4_r,
                                                                                                                                                                  applyfnInt_Bool_5_3_r,
                                                                                                                                                                  applyfnInt_Bool_5_2_r,
                                                                                                                                                                  applyfnInt_Bool_5_1_r}));
  assign applyfnInt_Bool_5_choice_r = lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_r;
  
  /* destruct (Ty TupGo___MyDTInt_Bool___Int,
          Dcon TupGo___MyDTInt_Bool___Int) : (applyfnInt_Bool_5_data,TupGo___MyDTInt_Bool___Int) > [(applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intgo_7,Go),
                                                                                                    (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0,MyDTInt_Bool),
                                                                                                    (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg1,Int)] */
  logic [2:0] applyfnInt_Bool_5_data_emitted;
  logic [2:0] applyfnInt_Bool_5_data_done;
  assign applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intgo_7_d = (applyfnInt_Bool_5_data_d[0] && (! applyfnInt_Bool_5_data_emitted[0]));
  assign applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_d = (applyfnInt_Bool_5_data_d[0] && (! applyfnInt_Bool_5_data_emitted[1]));
  assign applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg1_d = {applyfnInt_Bool_5_data_d[32:1],
                                                              (applyfnInt_Bool_5_data_d[0] && (! applyfnInt_Bool_5_data_emitted[2]))};
  assign applyfnInt_Bool_5_data_done = (applyfnInt_Bool_5_data_emitted | ({applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg1_d[0],
                                                                           applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_d[0],
                                                                           applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intgo_7_d[0]} & {applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg1_r,
                                                                                                                                    applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_r,
                                                                                                                                    applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intgo_7_r}));
  assign applyfnInt_Bool_5_data_r = (& applyfnInt_Bool_5_data_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) applyfnInt_Bool_5_data_emitted <= 3'd0;
    else
      applyfnInt_Bool_5_data_emitted <= (applyfnInt_Bool_5_data_r ? 3'd0 :
                                         applyfnInt_Bool_5_data_done);
  
  /* fork (Ty MyBool) : (applyfnInt_Bool_5_resbuf,MyBool) > [(es_2_1_1,MyBool),
                                                        (es_2_1_2,MyBool),
                                                        (es_2_1_3,MyBool),
                                                        (es_2_1_4,MyBool),
                                                        (es_2_1_5,MyBool)] */
  logic [4:0] applyfnInt_Bool_5_resbuf_emitted;
  logic [4:0] applyfnInt_Bool_5_resbuf_done;
  assign es_2_1_1_d = {applyfnInt_Bool_5_resbuf_d[1:1],
                       (applyfnInt_Bool_5_resbuf_d[0] && (! applyfnInt_Bool_5_resbuf_emitted[0]))};
  assign es_2_1_2_d = {applyfnInt_Bool_5_resbuf_d[1:1],
                       (applyfnInt_Bool_5_resbuf_d[0] && (! applyfnInt_Bool_5_resbuf_emitted[1]))};
  assign es_2_1_3_d = {applyfnInt_Bool_5_resbuf_d[1:1],
                       (applyfnInt_Bool_5_resbuf_d[0] && (! applyfnInt_Bool_5_resbuf_emitted[2]))};
  assign es_2_1_4_d = {applyfnInt_Bool_5_resbuf_d[1:1],
                       (applyfnInt_Bool_5_resbuf_d[0] && (! applyfnInt_Bool_5_resbuf_emitted[3]))};
  assign es_2_1_5_d = {applyfnInt_Bool_5_resbuf_d[1:1],
                       (applyfnInt_Bool_5_resbuf_d[0] && (! applyfnInt_Bool_5_resbuf_emitted[4]))};
  assign applyfnInt_Bool_5_resbuf_done = (applyfnInt_Bool_5_resbuf_emitted | ({es_2_1_5_d[0],
                                                                               es_2_1_4_d[0],
                                                                               es_2_1_3_d[0],
                                                                               es_2_1_2_d[0],
                                                                               es_2_1_1_d[0]} & {es_2_1_5_r,
                                                                                                 es_2_1_4_r,
                                                                                                 es_2_1_3_r,
                                                                                                 es_2_1_2_r,
                                                                                                 es_2_1_1_r}));
  assign applyfnInt_Bool_5_resbuf_r = (& applyfnInt_Bool_5_resbuf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) applyfnInt_Bool_5_resbuf_emitted <= 5'd0;
    else
      applyfnInt_Bool_5_resbuf_emitted <= (applyfnInt_Bool_5_resbuf_r ? 5'd0 :
                                           applyfnInt_Bool_5_resbuf_done);
  
  /* mergectrl (Ty C12,
           Ty TupMyDTInt_Int_Int___Int___Int) : [(applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1,TupMyDTInt_Int_Int___Int___Int),
                                                 (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int2,TupMyDTInt_Int_Int___Int___Int),
                                                 (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int3,TupMyDTInt_Int_Int___Int___Int),
                                                 (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int4,TupMyDTInt_Int_Int___Int___Int),
                                                 (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int5,TupMyDTInt_Int_Int___Int___Int),
                                                 (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int6,TupMyDTInt_Int_Int___Int___Int),
                                                 (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int7,TupMyDTInt_Int_Int___Int___Int),
                                                 (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int8,TupMyDTInt_Int_Int___Int___Int),
                                                 (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int9,TupMyDTInt_Int_Int___Int___Int),
                                                 (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int10,TupMyDTInt_Int_Int___Int___Int),
                                                 (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int11,TupMyDTInt_Int_Int___Int___Int),
                                                 (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int12,TupMyDTInt_Int_Int___Int___Int)] > (applyfnInt_Int_Int_5_choice,C12) (applyfnInt_Int_Int_5_data,TupMyDTInt_Int_Int___Int___Int) */
  logic [11:0] applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_select_d;
  assign applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_select_d = ((| applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_select_q) ? applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_select_q :
                                                                          (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_d[0] ? 12'd1 :
                                                                           (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int2_d[0] ? 12'd2 :
                                                                            (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int3_d[0] ? 12'd4 :
                                                                             (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int4_d[0] ? 12'd8 :
                                                                              (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int5_d[0] ? 12'd16 :
                                                                               (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int6_d[0] ? 12'd32 :
                                                                                (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int7_d[0] ? 12'd64 :
                                                                                 (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int8_d[0] ? 12'd128 :
                                                                                  (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int9_d[0] ? 12'd256 :
                                                                                   (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int10_d[0] ? 12'd512 :
                                                                                    (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int11_d[0] ? 12'd1024 :
                                                                                     (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int12_d[0] ? 12'd2048 :
                                                                                      12'd0)))))))))))));
  logic [11:0] applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_select_q <= 12'd0;
    else
      applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_select_q <= (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_done ? 12'd0 :
                                                                        applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_select_d);
  logic [1:0] applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_emit_q <= 2'd0;
    else
      applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_emit_q <= (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_done ? 2'd0 :
                                                                      applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_emit_d);
  logic [1:0] applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_emit_d;
  assign applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_emit_d = (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_emit_q | ({applyfnInt_Int_Int_5_choice_d[0],
                                                                                                                                        applyfnInt_Int_Int_5_data_d[0]} & {applyfnInt_Int_Int_5_choice_r,
                                                                                                                                                                           applyfnInt_Int_Int_5_data_r}));
  logic applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_done;
  assign applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_done = (& applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_emit_d);
  assign {applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int12_r,
          applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int11_r,
          applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int10_r,
          applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int9_r,
          applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int8_r,
          applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int7_r,
          applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int6_r,
          applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int5_r,
          applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int4_r,
          applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int3_r,
          applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int2_r,
          applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_r} = (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_done ? applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_select_d :
                                                                     12'd0);
  assign applyfnInt_Int_Int_5_data_d = ((applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_select_d[0] && (! applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_emit_q[0])) ? applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_d :
                                        ((applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_select_d[1] && (! applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_emit_q[0])) ? applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int2_d :
                                         ((applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_select_d[2] && (! applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_emit_q[0])) ? applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int3_d :
                                          ((applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_select_d[3] && (! applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_emit_q[0])) ? applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int4_d :
                                           ((applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_select_d[4] && (! applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_emit_q[0])) ? applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int5_d :
                                            ((applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_select_d[5] && (! applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_emit_q[0])) ? applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int6_d :
                                             ((applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_select_d[6] && (! applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_emit_q[0])) ? applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int7_d :
                                              ((applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_select_d[7] && (! applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_emit_q[0])) ? applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int8_d :
                                               ((applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_select_d[8] && (! applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_emit_q[0])) ? applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int9_d :
                                                ((applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_select_d[9] && (! applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_emit_q[0])) ? applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int10_d :
                                                 ((applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_select_d[10] && (! applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_emit_q[0])) ? applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int11_d :
                                                  ((applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_select_d[11] && (! applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_emit_q[0])) ? applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int12_d :
                                                   {64'd0, 1'd0}))))))))))));
  assign applyfnInt_Int_Int_5_choice_d = ((applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_select_d[0] && (! applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_emit_q[1])) ? C1_12_dc(1'd1) :
                                          ((applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_select_d[1] && (! applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_emit_q[1])) ? C2_12_dc(1'd1) :
                                           ((applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_select_d[2] && (! applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_emit_q[1])) ? C3_12_dc(1'd1) :
                                            ((applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_select_d[3] && (! applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_emit_q[1])) ? C4_12_dc(1'd1) :
                                             ((applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_select_d[4] && (! applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_emit_q[1])) ? C5_12_dc(1'd1) :
                                              ((applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_select_d[5] && (! applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_emit_q[1])) ? C6_12_dc(1'd1) :
                                               ((applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_select_d[6] && (! applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_emit_q[1])) ? C7_12_dc(1'd1) :
                                                ((applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_select_d[7] && (! applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_emit_q[1])) ? C8_12_dc(1'd1) :
                                                 ((applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_select_d[8] && (! applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_emit_q[1])) ? C9_12_dc(1'd1) :
                                                  ((applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_select_d[9] && (! applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_emit_q[1])) ? C10_12_dc(1'd1) :
                                                   ((applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_select_d[10] && (! applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_emit_q[1])) ? C11_12_dc(1'd1) :
                                                    ((applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_select_d[11] && (! applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_emit_q[1])) ? C12_12_dc(1'd1) :
                                                     {4'd0, 1'd0}))))))))))));
  
  /* fork (Ty MyDTInt_Int_Int) : (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_2,MyDTInt_Int_Int) > [(arg0_2_1,MyDTInt_Int_Int),
                                                                                                          (arg0_2_2,MyDTInt_Int_Int),
                                                                                                          (arg0_2_3,MyDTInt_Int_Int)] */
  logic [2:0] applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_2_emitted;
  logic [2:0] applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_2_done;
  assign arg0_2_1_d = (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_2_d[0] && (! applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_2_emitted[0]));
  assign arg0_2_2_d = (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_2_d[0] && (! applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_2_emitted[1]));
  assign arg0_2_3_d = (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_2_d[0] && (! applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_2_emitted[2]));
  assign applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_2_done = (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_2_emitted | ({arg0_2_3_d[0],
                                                                                                                                               arg0_2_2_d[0],
                                                                                                                                               arg0_2_1_d[0]} & {arg0_2_3_r,
                                                                                                                                                                 arg0_2_2_r,
                                                                                                                                                                 arg0_2_1_r}));
  assign applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_2_r = (& applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_2_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_2_emitted <= 3'd0;
    else
      applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_2_emitted <= (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_2_r ? 3'd0 :
                                                                           applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_2_done);
  
  /* buf (Ty Int) : (applyfnInt_Int_Int_5_1,Int) > (applyfnInt_Int_Int_5_resbuf,Int) */
  Int_t applyfnInt_Int_Int_5_1_bufchan_d;
  logic applyfnInt_Int_Int_5_1_bufchan_r;
  assign applyfnInt_Int_Int_5_1_r = ((! applyfnInt_Int_Int_5_1_bufchan_d[0]) || applyfnInt_Int_Int_5_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_Int_5_1_bufchan_d <= {32'd0, 1'd0};
    else
      if (applyfnInt_Int_Int_5_1_r)
        applyfnInt_Int_Int_5_1_bufchan_d <= applyfnInt_Int_Int_5_1_d;
  Int_t applyfnInt_Int_Int_5_1_bufchan_buf;
  assign applyfnInt_Int_Int_5_1_bufchan_r = (! applyfnInt_Int_Int_5_1_bufchan_buf[0]);
  assign applyfnInt_Int_Int_5_resbuf_d = (applyfnInt_Int_Int_5_1_bufchan_buf[0] ? applyfnInt_Int_Int_5_1_bufchan_buf :
                                          applyfnInt_Int_Int_5_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_Int_5_1_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((applyfnInt_Int_Int_5_resbuf_r && applyfnInt_Int_Int_5_1_bufchan_buf[0]))
        applyfnInt_Int_Int_5_1_bufchan_buf <= {32'd0, 1'd0};
      else if (((! applyfnInt_Int_Int_5_resbuf_r) && (! applyfnInt_Int_Int_5_1_bufchan_buf[0])))
        applyfnInt_Int_Int_5_1_bufchan_buf <= applyfnInt_Int_Int_5_1_bufchan_d;
  
  /* buf (Ty Int) : (applyfnInt_Int_Int_5_10,Int) > (applyfnInt_Int_Int_5_10_argbuf,Int) */
  Int_t applyfnInt_Int_Int_5_10_bufchan_d;
  logic applyfnInt_Int_Int_5_10_bufchan_r;
  assign applyfnInt_Int_Int_5_10_r = ((! applyfnInt_Int_Int_5_10_bufchan_d[0]) || applyfnInt_Int_Int_5_10_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_Int_5_10_bufchan_d <= {32'd0, 1'd0};
    else
      if (applyfnInt_Int_Int_5_10_r)
        applyfnInt_Int_Int_5_10_bufchan_d <= applyfnInt_Int_Int_5_10_d;
  Int_t applyfnInt_Int_Int_5_10_bufchan_buf;
  assign applyfnInt_Int_Int_5_10_bufchan_r = (! applyfnInt_Int_Int_5_10_bufchan_buf[0]);
  assign applyfnInt_Int_Int_5_10_argbuf_d = (applyfnInt_Int_Int_5_10_bufchan_buf[0] ? applyfnInt_Int_Int_5_10_bufchan_buf :
                                             applyfnInt_Int_Int_5_10_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_Int_5_10_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((applyfnInt_Int_Int_5_10_argbuf_r && applyfnInt_Int_Int_5_10_bufchan_buf[0]))
        applyfnInt_Int_Int_5_10_bufchan_buf <= {32'd0, 1'd0};
      else if (((! applyfnInt_Int_Int_5_10_argbuf_r) && (! applyfnInt_Int_Int_5_10_bufchan_buf[0])))
        applyfnInt_Int_Int_5_10_bufchan_buf <= applyfnInt_Int_Int_5_10_bufchan_d;
  
  /* buf (Ty Int) : (applyfnInt_Int_Int_5_10_argbuf,Int) > (es_17_1_argbuf,Int) */
  Int_t applyfnInt_Int_Int_5_10_argbuf_bufchan_d;
  logic applyfnInt_Int_Int_5_10_argbuf_bufchan_r;
  assign applyfnInt_Int_Int_5_10_argbuf_r = ((! applyfnInt_Int_Int_5_10_argbuf_bufchan_d[0]) || applyfnInt_Int_Int_5_10_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_Int_5_10_argbuf_bufchan_d <= {32'd0, 1'd0};
    else
      if (applyfnInt_Int_Int_5_10_argbuf_r)
        applyfnInt_Int_Int_5_10_argbuf_bufchan_d <= applyfnInt_Int_Int_5_10_argbuf_d;
  Int_t applyfnInt_Int_Int_5_10_argbuf_bufchan_buf;
  assign applyfnInt_Int_Int_5_10_argbuf_bufchan_r = (! applyfnInt_Int_Int_5_10_argbuf_bufchan_buf[0]);
  assign es_17_1_argbuf_d = (applyfnInt_Int_Int_5_10_argbuf_bufchan_buf[0] ? applyfnInt_Int_Int_5_10_argbuf_bufchan_buf :
                             applyfnInt_Int_Int_5_10_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_Int_5_10_argbuf_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((es_17_1_argbuf_r && applyfnInt_Int_Int_5_10_argbuf_bufchan_buf[0]))
        applyfnInt_Int_Int_5_10_argbuf_bufchan_buf <= {32'd0, 1'd0};
      else if (((! es_17_1_argbuf_r) && (! applyfnInt_Int_Int_5_10_argbuf_bufchan_buf[0])))
        applyfnInt_Int_Int_5_10_argbuf_bufchan_buf <= applyfnInt_Int_Int_5_10_argbuf_bufchan_d;
  
  /* buf (Ty Int) : (applyfnInt_Int_Int_5_11,Int) > (applyfnInt_Int_Int_5_11_argbuf,Int) */
  Int_t applyfnInt_Int_Int_5_11_bufchan_d;
  logic applyfnInt_Int_Int_5_11_bufchan_r;
  assign applyfnInt_Int_Int_5_11_r = ((! applyfnInt_Int_Int_5_11_bufchan_d[0]) || applyfnInt_Int_Int_5_11_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_Int_5_11_bufchan_d <= {32'd0, 1'd0};
    else
      if (applyfnInt_Int_Int_5_11_r)
        applyfnInt_Int_Int_5_11_bufchan_d <= applyfnInt_Int_Int_5_11_d;
  Int_t applyfnInt_Int_Int_5_11_bufchan_buf;
  assign applyfnInt_Int_Int_5_11_bufchan_r = (! applyfnInt_Int_Int_5_11_bufchan_buf[0]);
  assign applyfnInt_Int_Int_5_11_argbuf_d = (applyfnInt_Int_Int_5_11_bufchan_buf[0] ? applyfnInt_Int_Int_5_11_bufchan_buf :
                                             applyfnInt_Int_Int_5_11_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_Int_5_11_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((applyfnInt_Int_Int_5_11_argbuf_r && applyfnInt_Int_Int_5_11_bufchan_buf[0]))
        applyfnInt_Int_Int_5_11_bufchan_buf <= {32'd0, 1'd0};
      else if (((! applyfnInt_Int_Int_5_11_argbuf_r) && (! applyfnInt_Int_Int_5_11_bufchan_buf[0])))
        applyfnInt_Int_Int_5_11_bufchan_buf <= applyfnInt_Int_Int_5_11_bufchan_d;
  
  /* buf (Ty Int) : (applyfnInt_Int_Int_5_11_argbuf,Int) > (es_24_1_argbuf,Int) */
  Int_t applyfnInt_Int_Int_5_11_argbuf_bufchan_d;
  logic applyfnInt_Int_Int_5_11_argbuf_bufchan_r;
  assign applyfnInt_Int_Int_5_11_argbuf_r = ((! applyfnInt_Int_Int_5_11_argbuf_bufchan_d[0]) || applyfnInt_Int_Int_5_11_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_Int_5_11_argbuf_bufchan_d <= {32'd0, 1'd0};
    else
      if (applyfnInt_Int_Int_5_11_argbuf_r)
        applyfnInt_Int_Int_5_11_argbuf_bufchan_d <= applyfnInt_Int_Int_5_11_argbuf_d;
  Int_t applyfnInt_Int_Int_5_11_argbuf_bufchan_buf;
  assign applyfnInt_Int_Int_5_11_argbuf_bufchan_r = (! applyfnInt_Int_Int_5_11_argbuf_bufchan_buf[0]);
  assign es_24_1_argbuf_d = (applyfnInt_Int_Int_5_11_argbuf_bufchan_buf[0] ? applyfnInt_Int_Int_5_11_argbuf_bufchan_buf :
                             applyfnInt_Int_Int_5_11_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_Int_5_11_argbuf_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((es_24_1_argbuf_r && applyfnInt_Int_Int_5_11_argbuf_bufchan_buf[0]))
        applyfnInt_Int_Int_5_11_argbuf_bufchan_buf <= {32'd0, 1'd0};
      else if (((! es_24_1_argbuf_r) && (! applyfnInt_Int_Int_5_11_argbuf_bufchan_buf[0])))
        applyfnInt_Int_Int_5_11_argbuf_bufchan_buf <= applyfnInt_Int_Int_5_11_argbuf_bufchan_d;
  
  /* buf (Ty Int) : (applyfnInt_Int_Int_5_12,Int) > (applyfnInt_Int_Int_5_12_argbuf,Int) */
  Int_t applyfnInt_Int_Int_5_12_bufchan_d;
  logic applyfnInt_Int_Int_5_12_bufchan_r;
  assign applyfnInt_Int_Int_5_12_r = ((! applyfnInt_Int_Int_5_12_bufchan_d[0]) || applyfnInt_Int_Int_5_12_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_Int_5_12_bufchan_d <= {32'd0, 1'd0};
    else
      if (applyfnInt_Int_Int_5_12_r)
        applyfnInt_Int_Int_5_12_bufchan_d <= applyfnInt_Int_Int_5_12_d;
  Int_t applyfnInt_Int_Int_5_12_bufchan_buf;
  assign applyfnInt_Int_Int_5_12_bufchan_r = (! applyfnInt_Int_Int_5_12_bufchan_buf[0]);
  assign applyfnInt_Int_Int_5_12_argbuf_d = (applyfnInt_Int_Int_5_12_bufchan_buf[0] ? applyfnInt_Int_Int_5_12_bufchan_buf :
                                             applyfnInt_Int_Int_5_12_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_Int_5_12_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((applyfnInt_Int_Int_5_12_argbuf_r && applyfnInt_Int_Int_5_12_bufchan_buf[0]))
        applyfnInt_Int_Int_5_12_bufchan_buf <= {32'd0, 1'd0};
      else if (((! applyfnInt_Int_Int_5_12_argbuf_r) && (! applyfnInt_Int_Int_5_12_bufchan_buf[0])))
        applyfnInt_Int_Int_5_12_bufchan_buf <= applyfnInt_Int_Int_5_12_bufchan_d;
  
  /* dcon (Ty QTree_Int,
      Dcon QVal_Int) : [(applyfnInt_Int_Int_5_12_argbuf,Int)] > (es_22_1QVal_Int,QTree_Int) */
  assign es_22_1QVal_Int_d = QVal_Int_dc((& {applyfnInt_Int_Int_5_12_argbuf_d[0]}), applyfnInt_Int_Int_5_12_argbuf_d);
  assign {applyfnInt_Int_Int_5_12_argbuf_r} = {1 {(es_22_1QVal_Int_r && es_22_1QVal_Int_d[0])}};
  
  /* buf (Ty Int) : (applyfnInt_Int_Int_5_2,Int) > (applyfnInt_Int_Int_5_2_argbuf,Int) */
  Int_t applyfnInt_Int_Int_5_2_bufchan_d;
  logic applyfnInt_Int_Int_5_2_bufchan_r;
  assign applyfnInt_Int_Int_5_2_r = ((! applyfnInt_Int_Int_5_2_bufchan_d[0]) || applyfnInt_Int_Int_5_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_Int_5_2_bufchan_d <= {32'd0, 1'd0};
    else
      if (applyfnInt_Int_Int_5_2_r)
        applyfnInt_Int_Int_5_2_bufchan_d <= applyfnInt_Int_Int_5_2_d;
  Int_t applyfnInt_Int_Int_5_2_bufchan_buf;
  assign applyfnInt_Int_Int_5_2_bufchan_r = (! applyfnInt_Int_Int_5_2_bufchan_buf[0]);
  assign applyfnInt_Int_Int_5_2_argbuf_d = (applyfnInt_Int_Int_5_2_bufchan_buf[0] ? applyfnInt_Int_Int_5_2_bufchan_buf :
                                            applyfnInt_Int_Int_5_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_Int_5_2_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((applyfnInt_Int_Int_5_2_argbuf_r && applyfnInt_Int_Int_5_2_bufchan_buf[0]))
        applyfnInt_Int_Int_5_2_bufchan_buf <= {32'd0, 1'd0};
      else if (((! applyfnInt_Int_Int_5_2_argbuf_r) && (! applyfnInt_Int_Int_5_2_bufchan_buf[0])))
        applyfnInt_Int_Int_5_2_bufchan_buf <= applyfnInt_Int_Int_5_2_bufchan_d;
  
  /* dcon (Ty QTree_Int,
      Dcon QVal_Int) : [(applyfnInt_Int_Int_5_2_argbuf,Int)] > (es_3_1_1QVal_Int,QTree_Int) */
  assign es_3_1_1QVal_Int_d = QVal_Int_dc((& {applyfnInt_Int_Int_5_2_argbuf_d[0]}), applyfnInt_Int_Int_5_2_argbuf_d);
  assign {applyfnInt_Int_Int_5_2_argbuf_r} = {1 {(es_3_1_1QVal_Int_r && es_3_1_1QVal_Int_d[0])}};
  
  /* buf (Ty Int) : (applyfnInt_Int_Int_5_3,Int) > (applyfnInt_Int_Int_5_3_argbuf,Int) */
  Int_t applyfnInt_Int_Int_5_3_bufchan_d;
  logic applyfnInt_Int_Int_5_3_bufchan_r;
  assign applyfnInt_Int_Int_5_3_r = ((! applyfnInt_Int_Int_5_3_bufchan_d[0]) || applyfnInt_Int_Int_5_3_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_Int_5_3_bufchan_d <= {32'd0, 1'd0};
    else
      if (applyfnInt_Int_Int_5_3_r)
        applyfnInt_Int_Int_5_3_bufchan_d <= applyfnInt_Int_Int_5_3_d;
  Int_t applyfnInt_Int_Int_5_3_bufchan_buf;
  assign applyfnInt_Int_Int_5_3_bufchan_r = (! applyfnInt_Int_Int_5_3_bufchan_buf[0]);
  assign applyfnInt_Int_Int_5_3_argbuf_d = (applyfnInt_Int_Int_5_3_bufchan_buf[0] ? applyfnInt_Int_Int_5_3_bufchan_buf :
                                            applyfnInt_Int_Int_5_3_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_Int_5_3_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((applyfnInt_Int_Int_5_3_argbuf_r && applyfnInt_Int_Int_5_3_bufchan_buf[0]))
        applyfnInt_Int_Int_5_3_bufchan_buf <= {32'd0, 1'd0};
      else if (((! applyfnInt_Int_Int_5_3_argbuf_r) && (! applyfnInt_Int_Int_5_3_bufchan_buf[0])))
        applyfnInt_Int_Int_5_3_bufchan_buf <= applyfnInt_Int_Int_5_3_bufchan_d;
  
  /* buf (Ty Int) : (applyfnInt_Int_Int_5_3_argbuf,Int) > (es_1_1_argbuf,Int) */
  Int_t applyfnInt_Int_Int_5_3_argbuf_bufchan_d;
  logic applyfnInt_Int_Int_5_3_argbuf_bufchan_r;
  assign applyfnInt_Int_Int_5_3_argbuf_r = ((! applyfnInt_Int_Int_5_3_argbuf_bufchan_d[0]) || applyfnInt_Int_Int_5_3_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_Int_5_3_argbuf_bufchan_d <= {32'd0, 1'd0};
    else
      if (applyfnInt_Int_Int_5_3_argbuf_r)
        applyfnInt_Int_Int_5_3_argbuf_bufchan_d <= applyfnInt_Int_Int_5_3_argbuf_d;
  Int_t applyfnInt_Int_Int_5_3_argbuf_bufchan_buf;
  assign applyfnInt_Int_Int_5_3_argbuf_bufchan_r = (! applyfnInt_Int_Int_5_3_argbuf_bufchan_buf[0]);
  assign es_1_1_argbuf_d = (applyfnInt_Int_Int_5_3_argbuf_bufchan_buf[0] ? applyfnInt_Int_Int_5_3_argbuf_bufchan_buf :
                            applyfnInt_Int_Int_5_3_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_Int_5_3_argbuf_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((es_1_1_argbuf_r && applyfnInt_Int_Int_5_3_argbuf_bufchan_buf[0]))
        applyfnInt_Int_Int_5_3_argbuf_bufchan_buf <= {32'd0, 1'd0};
      else if (((! es_1_1_argbuf_r) && (! applyfnInt_Int_Int_5_3_argbuf_bufchan_buf[0])))
        applyfnInt_Int_Int_5_3_argbuf_bufchan_buf <= applyfnInt_Int_Int_5_3_argbuf_bufchan_d;
  
  /* buf (Ty Int) : (applyfnInt_Int_Int_5_4,Int) > (applyfnInt_Int_Int_5_4_argbuf,Int) */
  Int_t applyfnInt_Int_Int_5_4_bufchan_d;
  logic applyfnInt_Int_Int_5_4_bufchan_r;
  assign applyfnInt_Int_Int_5_4_r = ((! applyfnInt_Int_Int_5_4_bufchan_d[0]) || applyfnInt_Int_Int_5_4_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_Int_5_4_bufchan_d <= {32'd0, 1'd0};
    else
      if (applyfnInt_Int_Int_5_4_r)
        applyfnInt_Int_Int_5_4_bufchan_d <= applyfnInt_Int_Int_5_4_d;
  Int_t applyfnInt_Int_Int_5_4_bufchan_buf;
  assign applyfnInt_Int_Int_5_4_bufchan_r = (! applyfnInt_Int_Int_5_4_bufchan_buf[0]);
  assign applyfnInt_Int_Int_5_4_argbuf_d = (applyfnInt_Int_Int_5_4_bufchan_buf[0] ? applyfnInt_Int_Int_5_4_bufchan_buf :
                                            applyfnInt_Int_Int_5_4_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_Int_5_4_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((applyfnInt_Int_Int_5_4_argbuf_r && applyfnInt_Int_Int_5_4_bufchan_buf[0]))
        applyfnInt_Int_Int_5_4_bufchan_buf <= {32'd0, 1'd0};
      else if (((! applyfnInt_Int_Int_5_4_argbuf_r) && (! applyfnInt_Int_Int_5_4_bufchan_buf[0])))
        applyfnInt_Int_Int_5_4_bufchan_buf <= applyfnInt_Int_Int_5_4_bufchan_d;
  
  /* dcon (Ty QTree_Int,
      Dcon QVal_Int) : [(applyfnInt_Int_Int_5_4_argbuf,Int)] > (es_3_1QVal_Int,QTree_Int) */
  assign es_3_1QVal_Int_d = QVal_Int_dc((& {applyfnInt_Int_Int_5_4_argbuf_d[0]}), applyfnInt_Int_Int_5_4_argbuf_d);
  assign {applyfnInt_Int_Int_5_4_argbuf_r} = {1 {(es_3_1QVal_Int_r && es_3_1QVal_Int_d[0])}};
  
  /* buf (Ty Int) : (applyfnInt_Int_Int_5_5,Int) > (applyfnInt_Int_Int_5_5_argbuf,Int) */
  Int_t applyfnInt_Int_Int_5_5_bufchan_d;
  logic applyfnInt_Int_Int_5_5_bufchan_r;
  assign applyfnInt_Int_Int_5_5_r = ((! applyfnInt_Int_Int_5_5_bufchan_d[0]) || applyfnInt_Int_Int_5_5_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_Int_5_5_bufchan_d <= {32'd0, 1'd0};
    else
      if (applyfnInt_Int_Int_5_5_r)
        applyfnInt_Int_Int_5_5_bufchan_d <= applyfnInt_Int_Int_5_5_d;
  Int_t applyfnInt_Int_Int_5_5_bufchan_buf;
  assign applyfnInt_Int_Int_5_5_bufchan_r = (! applyfnInt_Int_Int_5_5_bufchan_buf[0]);
  assign applyfnInt_Int_Int_5_5_argbuf_d = (applyfnInt_Int_Int_5_5_bufchan_buf[0] ? applyfnInt_Int_Int_5_5_bufchan_buf :
                                            applyfnInt_Int_Int_5_5_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_Int_5_5_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((applyfnInt_Int_Int_5_5_argbuf_r && applyfnInt_Int_Int_5_5_bufchan_buf[0]))
        applyfnInt_Int_Int_5_5_bufchan_buf <= {32'd0, 1'd0};
      else if (((! applyfnInt_Int_Int_5_5_argbuf_r) && (! applyfnInt_Int_Int_5_5_bufchan_buf[0])))
        applyfnInt_Int_Int_5_5_bufchan_buf <= applyfnInt_Int_Int_5_5_bufchan_d;
  
  /* buf (Ty Int) : (applyfnInt_Int_Int_5_5_argbuf,Int) > (es_9_1_argbuf,Int) */
  Int_t applyfnInt_Int_Int_5_5_argbuf_bufchan_d;
  logic applyfnInt_Int_Int_5_5_argbuf_bufchan_r;
  assign applyfnInt_Int_Int_5_5_argbuf_r = ((! applyfnInt_Int_Int_5_5_argbuf_bufchan_d[0]) || applyfnInt_Int_Int_5_5_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_Int_5_5_argbuf_bufchan_d <= {32'd0, 1'd0};
    else
      if (applyfnInt_Int_Int_5_5_argbuf_r)
        applyfnInt_Int_Int_5_5_argbuf_bufchan_d <= applyfnInt_Int_Int_5_5_argbuf_d;
  Int_t applyfnInt_Int_Int_5_5_argbuf_bufchan_buf;
  assign applyfnInt_Int_Int_5_5_argbuf_bufchan_r = (! applyfnInt_Int_Int_5_5_argbuf_bufchan_buf[0]);
  assign es_9_1_argbuf_d = (applyfnInt_Int_Int_5_5_argbuf_bufchan_buf[0] ? applyfnInt_Int_Int_5_5_argbuf_bufchan_buf :
                            applyfnInt_Int_Int_5_5_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_Int_5_5_argbuf_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((es_9_1_argbuf_r && applyfnInt_Int_Int_5_5_argbuf_bufchan_buf[0]))
        applyfnInt_Int_Int_5_5_argbuf_bufchan_buf <= {32'd0, 1'd0};
      else if (((! es_9_1_argbuf_r) && (! applyfnInt_Int_Int_5_5_argbuf_bufchan_buf[0])))
        applyfnInt_Int_Int_5_5_argbuf_bufchan_buf <= applyfnInt_Int_Int_5_5_argbuf_bufchan_d;
  
  /* buf (Ty Int) : (applyfnInt_Int_Int_5_6,Int) > (applyfnInt_Int_Int_5_6_argbuf,Int) */
  Int_t applyfnInt_Int_Int_5_6_bufchan_d;
  logic applyfnInt_Int_Int_5_6_bufchan_r;
  assign applyfnInt_Int_Int_5_6_r = ((! applyfnInt_Int_Int_5_6_bufchan_d[0]) || applyfnInt_Int_Int_5_6_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_Int_5_6_bufchan_d <= {32'd0, 1'd0};
    else
      if (applyfnInt_Int_Int_5_6_r)
        applyfnInt_Int_Int_5_6_bufchan_d <= applyfnInt_Int_Int_5_6_d;
  Int_t applyfnInt_Int_Int_5_6_bufchan_buf;
  assign applyfnInt_Int_Int_5_6_bufchan_r = (! applyfnInt_Int_Int_5_6_bufchan_buf[0]);
  assign applyfnInt_Int_Int_5_6_argbuf_d = (applyfnInt_Int_Int_5_6_bufchan_buf[0] ? applyfnInt_Int_Int_5_6_bufchan_buf :
                                            applyfnInt_Int_Int_5_6_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_Int_5_6_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((applyfnInt_Int_Int_5_6_argbuf_r && applyfnInt_Int_Int_5_6_bufchan_buf[0]))
        applyfnInt_Int_Int_5_6_bufchan_buf <= {32'd0, 1'd0};
      else if (((! applyfnInt_Int_Int_5_6_argbuf_r) && (! applyfnInt_Int_Int_5_6_bufchan_buf[0])))
        applyfnInt_Int_Int_5_6_bufchan_buf <= applyfnInt_Int_Int_5_6_bufchan_d;
  
  /* dcon (Ty QTree_Int,
      Dcon QVal_Int) : [(applyfnInt_Int_Int_5_6_argbuf,Int)] > (es_11_1QVal_Int,QTree_Int) */
  assign es_11_1QVal_Int_d = QVal_Int_dc((& {applyfnInt_Int_Int_5_6_argbuf_d[0]}), applyfnInt_Int_Int_5_6_argbuf_d);
  assign {applyfnInt_Int_Int_5_6_argbuf_r} = {1 {(es_11_1QVal_Int_r && es_11_1QVal_Int_d[0])}};
  
  /* buf (Ty Int) : (applyfnInt_Int_Int_5_7,Int) > (applyfnInt_Int_Int_5_7_argbuf,Int) */
  Int_t applyfnInt_Int_Int_5_7_bufchan_d;
  logic applyfnInt_Int_Int_5_7_bufchan_r;
  assign applyfnInt_Int_Int_5_7_r = ((! applyfnInt_Int_Int_5_7_bufchan_d[0]) || applyfnInt_Int_Int_5_7_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_Int_5_7_bufchan_d <= {32'd0, 1'd0};
    else
      if (applyfnInt_Int_Int_5_7_r)
        applyfnInt_Int_Int_5_7_bufchan_d <= applyfnInt_Int_Int_5_7_d;
  Int_t applyfnInt_Int_Int_5_7_bufchan_buf;
  assign applyfnInt_Int_Int_5_7_bufchan_r = (! applyfnInt_Int_Int_5_7_bufchan_buf[0]);
  assign applyfnInt_Int_Int_5_7_argbuf_d = (applyfnInt_Int_Int_5_7_bufchan_buf[0] ? applyfnInt_Int_Int_5_7_bufchan_buf :
                                            applyfnInt_Int_Int_5_7_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_Int_5_7_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((applyfnInt_Int_Int_5_7_argbuf_r && applyfnInt_Int_Int_5_7_bufchan_buf[0]))
        applyfnInt_Int_Int_5_7_bufchan_buf <= {32'd0, 1'd0};
      else if (((! applyfnInt_Int_Int_5_7_argbuf_r) && (! applyfnInt_Int_Int_5_7_bufchan_buf[0])))
        applyfnInt_Int_Int_5_7_bufchan_buf <= applyfnInt_Int_Int_5_7_bufchan_d;
  
  /* buf (Ty Int) : (applyfnInt_Int_Int_5_7_argbuf,Int) > (es_13_1_argbuf,Int) */
  Int_t applyfnInt_Int_Int_5_7_argbuf_bufchan_d;
  logic applyfnInt_Int_Int_5_7_argbuf_bufchan_r;
  assign applyfnInt_Int_Int_5_7_argbuf_r = ((! applyfnInt_Int_Int_5_7_argbuf_bufchan_d[0]) || applyfnInt_Int_Int_5_7_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_Int_5_7_argbuf_bufchan_d <= {32'd0, 1'd0};
    else
      if (applyfnInt_Int_Int_5_7_argbuf_r)
        applyfnInt_Int_Int_5_7_argbuf_bufchan_d <= applyfnInt_Int_Int_5_7_argbuf_d;
  Int_t applyfnInt_Int_Int_5_7_argbuf_bufchan_buf;
  assign applyfnInt_Int_Int_5_7_argbuf_bufchan_r = (! applyfnInt_Int_Int_5_7_argbuf_bufchan_buf[0]);
  assign es_13_1_argbuf_d = (applyfnInt_Int_Int_5_7_argbuf_bufchan_buf[0] ? applyfnInt_Int_Int_5_7_argbuf_bufchan_buf :
                             applyfnInt_Int_Int_5_7_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_Int_5_7_argbuf_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((es_13_1_argbuf_r && applyfnInt_Int_Int_5_7_argbuf_bufchan_buf[0]))
        applyfnInt_Int_Int_5_7_argbuf_bufchan_buf <= {32'd0, 1'd0};
      else if (((! es_13_1_argbuf_r) && (! applyfnInt_Int_Int_5_7_argbuf_bufchan_buf[0])))
        applyfnInt_Int_Int_5_7_argbuf_bufchan_buf <= applyfnInt_Int_Int_5_7_argbuf_bufchan_d;
  
  /* buf (Ty Int) : (applyfnInt_Int_Int_5_8,Int) > (applyfnInt_Int_Int_5_8_argbuf,Int) */
  Int_t applyfnInt_Int_Int_5_8_bufchan_d;
  logic applyfnInt_Int_Int_5_8_bufchan_r;
  assign applyfnInt_Int_Int_5_8_r = ((! applyfnInt_Int_Int_5_8_bufchan_d[0]) || applyfnInt_Int_Int_5_8_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_Int_5_8_bufchan_d <= {32'd0, 1'd0};
    else
      if (applyfnInt_Int_Int_5_8_r)
        applyfnInt_Int_Int_5_8_bufchan_d <= applyfnInt_Int_Int_5_8_d;
  Int_t applyfnInt_Int_Int_5_8_bufchan_buf;
  assign applyfnInt_Int_Int_5_8_bufchan_r = (! applyfnInt_Int_Int_5_8_bufchan_buf[0]);
  assign applyfnInt_Int_Int_5_8_argbuf_d = (applyfnInt_Int_Int_5_8_bufchan_buf[0] ? applyfnInt_Int_Int_5_8_bufchan_buf :
                                            applyfnInt_Int_Int_5_8_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_Int_5_8_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((applyfnInt_Int_Int_5_8_argbuf_r && applyfnInt_Int_Int_5_8_bufchan_buf[0]))
        applyfnInt_Int_Int_5_8_bufchan_buf <= {32'd0, 1'd0};
      else if (((! applyfnInt_Int_Int_5_8_argbuf_r) && (! applyfnInt_Int_Int_5_8_bufchan_buf[0])))
        applyfnInt_Int_Int_5_8_bufchan_buf <= applyfnInt_Int_Int_5_8_bufchan_d;
  
  /* dcon (Ty QTree_Int,
      Dcon QVal_Int) : [(applyfnInt_Int_Int_5_8_argbuf,Int)] > (es_15_1QVal_Int,QTree_Int) */
  assign es_15_1QVal_Int_d = QVal_Int_dc((& {applyfnInt_Int_Int_5_8_argbuf_d[0]}), applyfnInt_Int_Int_5_8_argbuf_d);
  assign {applyfnInt_Int_Int_5_8_argbuf_r} = {1 {(es_15_1QVal_Int_r && es_15_1QVal_Int_d[0])}};
  
  /* buf (Ty Int) : (applyfnInt_Int_Int_5_9,Int) > (applyfnInt_Int_Int_5_9_argbuf,Int) */
  Int_t applyfnInt_Int_Int_5_9_bufchan_d;
  logic applyfnInt_Int_Int_5_9_bufchan_r;
  assign applyfnInt_Int_Int_5_9_r = ((! applyfnInt_Int_Int_5_9_bufchan_d[0]) || applyfnInt_Int_Int_5_9_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_Int_5_9_bufchan_d <= {32'd0, 1'd0};
    else
      if (applyfnInt_Int_Int_5_9_r)
        applyfnInt_Int_Int_5_9_bufchan_d <= applyfnInt_Int_Int_5_9_d;
  Int_t applyfnInt_Int_Int_5_9_bufchan_buf;
  assign applyfnInt_Int_Int_5_9_bufchan_r = (! applyfnInt_Int_Int_5_9_bufchan_buf[0]);
  assign applyfnInt_Int_Int_5_9_argbuf_d = (applyfnInt_Int_Int_5_9_bufchan_buf[0] ? applyfnInt_Int_Int_5_9_bufchan_buf :
                                            applyfnInt_Int_Int_5_9_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_Int_5_9_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((applyfnInt_Int_Int_5_9_argbuf_r && applyfnInt_Int_Int_5_9_bufchan_buf[0]))
        applyfnInt_Int_Int_5_9_bufchan_buf <= {32'd0, 1'd0};
      else if (((! applyfnInt_Int_Int_5_9_argbuf_r) && (! applyfnInt_Int_Int_5_9_bufchan_buf[0])))
        applyfnInt_Int_Int_5_9_bufchan_buf <= applyfnInt_Int_Int_5_9_bufchan_d;
  
  /* buf (Ty Int) : (applyfnInt_Int_Int_5_9_argbuf,Int) > (es_19_1_argbuf,Int) */
  Int_t applyfnInt_Int_Int_5_9_argbuf_bufchan_d;
  logic applyfnInt_Int_Int_5_9_argbuf_bufchan_r;
  assign applyfnInt_Int_Int_5_9_argbuf_r = ((! applyfnInt_Int_Int_5_9_argbuf_bufchan_d[0]) || applyfnInt_Int_Int_5_9_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_Int_5_9_argbuf_bufchan_d <= {32'd0, 1'd0};
    else
      if (applyfnInt_Int_Int_5_9_argbuf_r)
        applyfnInt_Int_Int_5_9_argbuf_bufchan_d <= applyfnInt_Int_Int_5_9_argbuf_d;
  Int_t applyfnInt_Int_Int_5_9_argbuf_bufchan_buf;
  assign applyfnInt_Int_Int_5_9_argbuf_bufchan_r = (! applyfnInt_Int_Int_5_9_argbuf_bufchan_buf[0]);
  assign es_19_1_argbuf_d = (applyfnInt_Int_Int_5_9_argbuf_bufchan_buf[0] ? applyfnInt_Int_Int_5_9_argbuf_bufchan_buf :
                             applyfnInt_Int_Int_5_9_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_Int_5_9_argbuf_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((es_19_1_argbuf_r && applyfnInt_Int_Int_5_9_argbuf_bufchan_buf[0]))
        applyfnInt_Int_Int_5_9_argbuf_bufchan_buf <= {32'd0, 1'd0};
      else if (((! es_19_1_argbuf_r) && (! applyfnInt_Int_Int_5_9_argbuf_bufchan_buf[0])))
        applyfnInt_Int_Int_5_9_argbuf_bufchan_buf <= applyfnInt_Int_Int_5_9_argbuf_bufchan_d;
  
  /* demux (Ty C12,
       Ty Int) : (applyfnInt_Int_Int_5_choice,C12) (es_0_1_1I#_mux_mux_mux,Int) > [(applyfnInt_Int_Int_5_1,Int),
                                                                                   (applyfnInt_Int_Int_5_2,Int),
                                                                                   (applyfnInt_Int_Int_5_3,Int),
                                                                                   (applyfnInt_Int_Int_5_4,Int),
                                                                                   (applyfnInt_Int_Int_5_5,Int),
                                                                                   (applyfnInt_Int_Int_5_6,Int),
                                                                                   (applyfnInt_Int_Int_5_7,Int),
                                                                                   (applyfnInt_Int_Int_5_8,Int),
                                                                                   (applyfnInt_Int_Int_5_9,Int),
                                                                                   (applyfnInt_Int_Int_5_10,Int),
                                                                                   (applyfnInt_Int_Int_5_11,Int),
                                                                                   (applyfnInt_Int_Int_5_12,Int)] */
  logic [11:0] \es_0_1_1I#_mux_mux_mux_onehotd ;
  always_comb
    if ((applyfnInt_Int_Int_5_choice_d[0] && \es_0_1_1I#_mux_mux_mux_d [0]))
      unique case (applyfnInt_Int_Int_5_choice_d[4:1])
        4'd0: \es_0_1_1I#_mux_mux_mux_onehotd  = 12'd1;
        4'd1: \es_0_1_1I#_mux_mux_mux_onehotd  = 12'd2;
        4'd2: \es_0_1_1I#_mux_mux_mux_onehotd  = 12'd4;
        4'd3: \es_0_1_1I#_mux_mux_mux_onehotd  = 12'd8;
        4'd4: \es_0_1_1I#_mux_mux_mux_onehotd  = 12'd16;
        4'd5: \es_0_1_1I#_mux_mux_mux_onehotd  = 12'd32;
        4'd6: \es_0_1_1I#_mux_mux_mux_onehotd  = 12'd64;
        4'd7: \es_0_1_1I#_mux_mux_mux_onehotd  = 12'd128;
        4'd8: \es_0_1_1I#_mux_mux_mux_onehotd  = 12'd256;
        4'd9: \es_0_1_1I#_mux_mux_mux_onehotd  = 12'd512;
        4'd10: \es_0_1_1I#_mux_mux_mux_onehotd  = 12'd1024;
        4'd11: \es_0_1_1I#_mux_mux_mux_onehotd  = 12'd2048;
        default: \es_0_1_1I#_mux_mux_mux_onehotd  = 12'd0;
      endcase
    else \es_0_1_1I#_mux_mux_mux_onehotd  = 12'd0;
  assign applyfnInt_Int_Int_5_1_d = {\es_0_1_1I#_mux_mux_mux_d [32:1],
                                     \es_0_1_1I#_mux_mux_mux_onehotd [0]};
  assign applyfnInt_Int_Int_5_2_d = {\es_0_1_1I#_mux_mux_mux_d [32:1],
                                     \es_0_1_1I#_mux_mux_mux_onehotd [1]};
  assign applyfnInt_Int_Int_5_3_d = {\es_0_1_1I#_mux_mux_mux_d [32:1],
                                     \es_0_1_1I#_mux_mux_mux_onehotd [2]};
  assign applyfnInt_Int_Int_5_4_d = {\es_0_1_1I#_mux_mux_mux_d [32:1],
                                     \es_0_1_1I#_mux_mux_mux_onehotd [3]};
  assign applyfnInt_Int_Int_5_5_d = {\es_0_1_1I#_mux_mux_mux_d [32:1],
                                     \es_0_1_1I#_mux_mux_mux_onehotd [4]};
  assign applyfnInt_Int_Int_5_6_d = {\es_0_1_1I#_mux_mux_mux_d [32:1],
                                     \es_0_1_1I#_mux_mux_mux_onehotd [5]};
  assign applyfnInt_Int_Int_5_7_d = {\es_0_1_1I#_mux_mux_mux_d [32:1],
                                     \es_0_1_1I#_mux_mux_mux_onehotd [6]};
  assign applyfnInt_Int_Int_5_8_d = {\es_0_1_1I#_mux_mux_mux_d [32:1],
                                     \es_0_1_1I#_mux_mux_mux_onehotd [7]};
  assign applyfnInt_Int_Int_5_9_d = {\es_0_1_1I#_mux_mux_mux_d [32:1],
                                     \es_0_1_1I#_mux_mux_mux_onehotd [8]};
  assign applyfnInt_Int_Int_5_10_d = {\es_0_1_1I#_mux_mux_mux_d [32:1],
                                      \es_0_1_1I#_mux_mux_mux_onehotd [9]};
  assign applyfnInt_Int_Int_5_11_d = {\es_0_1_1I#_mux_mux_mux_d [32:1],
                                      \es_0_1_1I#_mux_mux_mux_onehotd [10]};
  assign applyfnInt_Int_Int_5_12_d = {\es_0_1_1I#_mux_mux_mux_d [32:1],
                                      \es_0_1_1I#_mux_mux_mux_onehotd [11]};
  assign \es_0_1_1I#_mux_mux_mux_r  = (| (\es_0_1_1I#_mux_mux_mux_onehotd  & {applyfnInt_Int_Int_5_12_r,
                                                                              applyfnInt_Int_Int_5_11_r,
                                                                              applyfnInt_Int_Int_5_10_r,
                                                                              applyfnInt_Int_Int_5_9_r,
                                                                              applyfnInt_Int_Int_5_8_r,
                                                                              applyfnInt_Int_Int_5_7_r,
                                                                              applyfnInt_Int_Int_5_6_r,
                                                                              applyfnInt_Int_Int_5_5_r,
                                                                              applyfnInt_Int_Int_5_4_r,
                                                                              applyfnInt_Int_Int_5_3_r,
                                                                              applyfnInt_Int_Int_5_2_r,
                                                                              applyfnInt_Int_Int_5_1_r}));
  assign applyfnInt_Int_Int_5_choice_r = \es_0_1_1I#_mux_mux_mux_r ;
  
  /* destruct (Ty TupMyDTInt_Int_Int___Int___Int,
          Dcon TupMyDTInt_Int_Int___Int___Int) : (applyfnInt_Int_Int_5_data,TupMyDTInt_Int_Int___Int___Int) > [(applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_2,MyDTInt_Int_Int),
                                                                                                               (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg2,Int),
                                                                                                               (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg1_1,Int)] */
  logic [2:0] applyfnInt_Int_Int_5_data_emitted;
  logic [2:0] applyfnInt_Int_Int_5_data_done;
  assign applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_2_d = (applyfnInt_Int_Int_5_data_d[0] && (! applyfnInt_Int_Int_5_data_emitted[0]));
  assign applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg2_d = {applyfnInt_Int_Int_5_data_d[32:1],
                                                                     (applyfnInt_Int_Int_5_data_d[0] && (! applyfnInt_Int_Int_5_data_emitted[1]))};
  assign applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg1_1_d = {applyfnInt_Int_Int_5_data_d[64:33],
                                                                       (applyfnInt_Int_Int_5_data_d[0] && (! applyfnInt_Int_Int_5_data_emitted[2]))};
  assign applyfnInt_Int_Int_5_data_done = (applyfnInt_Int_Int_5_data_emitted | ({applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg1_1_d[0],
                                                                                 applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg2_d[0],
                                                                                 applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_2_d[0]} & {applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg1_1_r,
                                                                                                                                                   applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg2_r,
                                                                                                                                                   applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_2_r}));
  assign applyfnInt_Int_Int_5_data_r = (& applyfnInt_Int_Int_5_data_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) applyfnInt_Int_Int_5_data_emitted <= 3'd0;
    else
      applyfnInt_Int_Int_5_data_emitted <= (applyfnInt_Int_Int_5_data_r ? 3'd0 :
                                            applyfnInt_Int_Int_5_data_done);
  
  /* buf (Ty Int) : (applyfnInt_Int_Int_5_resbuf,Int) > (es_1_1_1_argbuf,Int) */
  Int_t applyfnInt_Int_Int_5_resbuf_bufchan_d;
  logic applyfnInt_Int_Int_5_resbuf_bufchan_r;
  assign applyfnInt_Int_Int_5_resbuf_r = ((! applyfnInt_Int_Int_5_resbuf_bufchan_d[0]) || applyfnInt_Int_Int_5_resbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_Int_5_resbuf_bufchan_d <= {32'd0, 1'd0};
    else
      if (applyfnInt_Int_Int_5_resbuf_r)
        applyfnInt_Int_Int_5_resbuf_bufchan_d <= applyfnInt_Int_Int_5_resbuf_d;
  Int_t applyfnInt_Int_Int_5_resbuf_bufchan_buf;
  assign applyfnInt_Int_Int_5_resbuf_bufchan_r = (! applyfnInt_Int_Int_5_resbuf_bufchan_buf[0]);
  assign es_1_1_1_argbuf_d = (applyfnInt_Int_Int_5_resbuf_bufchan_buf[0] ? applyfnInt_Int_Int_5_resbuf_bufchan_buf :
                              applyfnInt_Int_Int_5_resbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_Int_5_resbuf_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((es_1_1_1_argbuf_r && applyfnInt_Int_Int_5_resbuf_bufchan_buf[0]))
        applyfnInt_Int_Int_5_resbuf_bufchan_buf <= {32'd0, 1'd0};
      else if (((! es_1_1_1_argbuf_r) && (! applyfnInt_Int_Int_5_resbuf_bufchan_buf[0])))
        applyfnInt_Int_Int_5_resbuf_bufchan_buf <= applyfnInt_Int_Int_5_resbuf_bufchan_d;
  
  /* demux (Ty MyDTInt_Bool,
       Ty Int) : (arg0_1,MyDTInt_Bool) (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg1,Int) > [(arg0_1Dcon_isZ,Int)] */
  assign arg0_1Dcon_isZ_d = {applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg1_d[32:1],
                             (arg0_1_d[0] && applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg1_d[0])};
  assign applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg1_r = (arg0_1Dcon_isZ_r && (arg0_1_d[0] && applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg1_d[0]));
  assign arg0_1_r = (arg0_1Dcon_isZ_r && (arg0_1_d[0] && applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg1_d[0]));
  
  /* fork (Ty Int) : (arg0_1Dcon_isZ,Int) > [(arg0_1Dcon_isZ_1,Int),
                                        (arg0_1Dcon_isZ_2,Int),
                                        (arg0_1Dcon_isZ_3,Int),
                                        (arg0_1Dcon_isZ_4,Int)] */
  logic [3:0] arg0_1Dcon_isZ_emitted;
  logic [3:0] arg0_1Dcon_isZ_done;
  assign arg0_1Dcon_isZ_1_d = {arg0_1Dcon_isZ_d[32:1],
                               (arg0_1Dcon_isZ_d[0] && (! arg0_1Dcon_isZ_emitted[0]))};
  assign arg0_1Dcon_isZ_2_d = {arg0_1Dcon_isZ_d[32:1],
                               (arg0_1Dcon_isZ_d[0] && (! arg0_1Dcon_isZ_emitted[1]))};
  assign arg0_1Dcon_isZ_3_d = {arg0_1Dcon_isZ_d[32:1],
                               (arg0_1Dcon_isZ_d[0] && (! arg0_1Dcon_isZ_emitted[2]))};
  assign arg0_1Dcon_isZ_4_d = {arg0_1Dcon_isZ_d[32:1],
                               (arg0_1Dcon_isZ_d[0] && (! arg0_1Dcon_isZ_emitted[3]))};
  assign arg0_1Dcon_isZ_done = (arg0_1Dcon_isZ_emitted | ({arg0_1Dcon_isZ_4_d[0],
                                                           arg0_1Dcon_isZ_3_d[0],
                                                           arg0_1Dcon_isZ_2_d[0],
                                                           arg0_1Dcon_isZ_1_d[0]} & {arg0_1Dcon_isZ_4_r,
                                                                                     arg0_1Dcon_isZ_3_r,
                                                                                     arg0_1Dcon_isZ_2_r,
                                                                                     arg0_1Dcon_isZ_1_r}));
  assign arg0_1Dcon_isZ_r = (& arg0_1Dcon_isZ_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) arg0_1Dcon_isZ_emitted <= 4'd0;
    else
      arg0_1Dcon_isZ_emitted <= (arg0_1Dcon_isZ_r ? 4'd0 :
                                 arg0_1Dcon_isZ_done);
  
  /* destruct (Ty Int,
          Dcon I#) : (arg0_1Dcon_isZ_1I#,Int) > [(x1ajq_destruct,Int#)] */
  assign x1ajq_destruct_d = {\arg0_1Dcon_isZ_1I#_d [32:1],
                             \arg0_1Dcon_isZ_1I#_d [0]};
  assign \arg0_1Dcon_isZ_1I#_r  = x1ajq_destruct_r;
  
  /* demux (Ty Int,
       Ty Int) : (arg0_1Dcon_isZ_2,Int) (arg0_1Dcon_isZ_1,Int) > [(arg0_1Dcon_isZ_1I#,Int)] */
  assign \arg0_1Dcon_isZ_1I#_d  = {arg0_1Dcon_isZ_1_d[32:1],
                                   (arg0_1Dcon_isZ_2_d[0] && arg0_1Dcon_isZ_1_d[0])};
  assign arg0_1Dcon_isZ_1_r = (\arg0_1Dcon_isZ_1I#_r  && (arg0_1Dcon_isZ_2_d[0] && arg0_1Dcon_isZ_1_d[0]));
  assign arg0_1Dcon_isZ_2_r = (\arg0_1Dcon_isZ_1I#_r  && (arg0_1Dcon_isZ_2_d[0] && arg0_1Dcon_isZ_1_d[0]));
  
  /* demux (Ty Int,
       Ty Go) : (arg0_1Dcon_isZ_3,Int) (arg0_2Dcon_isZ,Go) > [(arg0_1Dcon_isZ_3I#,Go)] */
  assign \arg0_1Dcon_isZ_3I#_d  = (arg0_1Dcon_isZ_3_d[0] && arg0_2Dcon_isZ_d[0]);
  assign arg0_2Dcon_isZ_r = (\arg0_1Dcon_isZ_3I#_r  && (arg0_1Dcon_isZ_3_d[0] && arg0_2Dcon_isZ_d[0]));
  assign arg0_1Dcon_isZ_3_r = (\arg0_1Dcon_isZ_3I#_r  && (arg0_1Dcon_isZ_3_d[0] && arg0_2Dcon_isZ_d[0]));
  
  /* fork (Ty Go) : (arg0_1Dcon_isZ_3I#,Go) > [(arg0_1Dcon_isZ_3I#_1,Go),
                                          (arg0_1Dcon_isZ_3I#_2,Go),
                                          (arg0_1Dcon_isZ_3I#_3,Go)] */
  logic [2:0] \arg0_1Dcon_isZ_3I#_emitted ;
  logic [2:0] \arg0_1Dcon_isZ_3I#_done ;
  assign \arg0_1Dcon_isZ_3I#_1_d  = (\arg0_1Dcon_isZ_3I#_d [0] && (! \arg0_1Dcon_isZ_3I#_emitted [0]));
  assign \arg0_1Dcon_isZ_3I#_2_d  = (\arg0_1Dcon_isZ_3I#_d [0] && (! \arg0_1Dcon_isZ_3I#_emitted [1]));
  assign \arg0_1Dcon_isZ_3I#_3_d  = (\arg0_1Dcon_isZ_3I#_d [0] && (! \arg0_1Dcon_isZ_3I#_emitted [2]));
  assign \arg0_1Dcon_isZ_3I#_done  = (\arg0_1Dcon_isZ_3I#_emitted  | ({\arg0_1Dcon_isZ_3I#_3_d [0],
                                                                       \arg0_1Dcon_isZ_3I#_2_d [0],
                                                                       \arg0_1Dcon_isZ_3I#_1_d [0]} & {\arg0_1Dcon_isZ_3I#_3_r ,
                                                                                                       \arg0_1Dcon_isZ_3I#_2_r ,
                                                                                                       \arg0_1Dcon_isZ_3I#_1_r }));
  assign \arg0_1Dcon_isZ_3I#_r  = (& \arg0_1Dcon_isZ_3I#_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \arg0_1Dcon_isZ_3I#_emitted  <= 3'd0;
    else
      \arg0_1Dcon_isZ_3I#_emitted  <= (\arg0_1Dcon_isZ_3I#_r  ? 3'd0 :
                                       \arg0_1Dcon_isZ_3I#_done );
  
  /* buf (Ty Go) : (arg0_1Dcon_isZ_3I#_1,Go) > (arg0_1Dcon_isZ_3I#_1_argbuf,Go) */
  Go_t \arg0_1Dcon_isZ_3I#_1_bufchan_d ;
  logic \arg0_1Dcon_isZ_3I#_1_bufchan_r ;
  assign \arg0_1Dcon_isZ_3I#_1_r  = ((! \arg0_1Dcon_isZ_3I#_1_bufchan_d [0]) || \arg0_1Dcon_isZ_3I#_1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \arg0_1Dcon_isZ_3I#_1_bufchan_d  <= 1'd0;
    else
      if (\arg0_1Dcon_isZ_3I#_1_r )
        \arg0_1Dcon_isZ_3I#_1_bufchan_d  <= \arg0_1Dcon_isZ_3I#_1_d ;
  Go_t \arg0_1Dcon_isZ_3I#_1_bufchan_buf ;
  assign \arg0_1Dcon_isZ_3I#_1_bufchan_r  = (! \arg0_1Dcon_isZ_3I#_1_bufchan_buf [0]);
  assign \arg0_1Dcon_isZ_3I#_1_argbuf_d  = (\arg0_1Dcon_isZ_3I#_1_bufchan_buf [0] ? \arg0_1Dcon_isZ_3I#_1_bufchan_buf  :
                                            \arg0_1Dcon_isZ_3I#_1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \arg0_1Dcon_isZ_3I#_1_bufchan_buf  <= 1'd0;
    else
      if ((\arg0_1Dcon_isZ_3I#_1_argbuf_r  && \arg0_1Dcon_isZ_3I#_1_bufchan_buf [0]))
        \arg0_1Dcon_isZ_3I#_1_bufchan_buf  <= 1'd0;
      else if (((! \arg0_1Dcon_isZ_3I#_1_argbuf_r ) && (! \arg0_1Dcon_isZ_3I#_1_bufchan_buf [0])))
        \arg0_1Dcon_isZ_3I#_1_bufchan_buf  <= \arg0_1Dcon_isZ_3I#_1_bufchan_d ;
  
  /* const (Ty Int#,
       Lit 0) : (arg0_1Dcon_isZ_3I#_1_argbuf,Go) > (arg0_1Dcon_isZ_3I#_1_argbuf_0,Int#) */
  assign \arg0_1Dcon_isZ_3I#_1_argbuf_0_d  = {32'd0,
                                              \arg0_1Dcon_isZ_3I#_1_argbuf_d [0]};
  assign \arg0_1Dcon_isZ_3I#_1_argbuf_r  = \arg0_1Dcon_isZ_3I#_1_argbuf_0_r ;
  
  /* op_eq (Ty Int#) : (arg0_1Dcon_isZ_3I#_1_argbuf_0,Int#) (x1ajq_destruct,Int#) > (lizzieLet1_1wild1Xv_1_Eq,Bool) */
  assign lizzieLet1_1wild1Xv_1_Eq_d = {(\arg0_1Dcon_isZ_3I#_1_argbuf_0_d [32:1] == x1ajq_destruct_d[32:1]),
                                       (\arg0_1Dcon_isZ_3I#_1_argbuf_0_d [0] && x1ajq_destruct_d[0])};
  assign {\arg0_1Dcon_isZ_3I#_1_argbuf_0_r ,
          x1ajq_destruct_r} = {2 {(lizzieLet1_1wild1Xv_1_Eq_r && lizzieLet1_1wild1Xv_1_Eq_d[0])}};
  
  /* buf (Ty Go) : (arg0_1Dcon_isZ_3I#_2,Go) > (arg0_1Dcon_isZ_3I#_2_argbuf,Go) */
  Go_t \arg0_1Dcon_isZ_3I#_2_bufchan_d ;
  logic \arg0_1Dcon_isZ_3I#_2_bufchan_r ;
  assign \arg0_1Dcon_isZ_3I#_2_r  = ((! \arg0_1Dcon_isZ_3I#_2_bufchan_d [0]) || \arg0_1Dcon_isZ_3I#_2_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \arg0_1Dcon_isZ_3I#_2_bufchan_d  <= 1'd0;
    else
      if (\arg0_1Dcon_isZ_3I#_2_r )
        \arg0_1Dcon_isZ_3I#_2_bufchan_d  <= \arg0_1Dcon_isZ_3I#_2_d ;
  Go_t \arg0_1Dcon_isZ_3I#_2_bufchan_buf ;
  assign \arg0_1Dcon_isZ_3I#_2_bufchan_r  = (! \arg0_1Dcon_isZ_3I#_2_bufchan_buf [0]);
  assign \arg0_1Dcon_isZ_3I#_2_argbuf_d  = (\arg0_1Dcon_isZ_3I#_2_bufchan_buf [0] ? \arg0_1Dcon_isZ_3I#_2_bufchan_buf  :
                                            \arg0_1Dcon_isZ_3I#_2_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \arg0_1Dcon_isZ_3I#_2_bufchan_buf  <= 1'd0;
    else
      if ((\arg0_1Dcon_isZ_3I#_2_argbuf_r  && \arg0_1Dcon_isZ_3I#_2_bufchan_buf [0]))
        \arg0_1Dcon_isZ_3I#_2_bufchan_buf  <= 1'd0;
      else if (((! \arg0_1Dcon_isZ_3I#_2_argbuf_r ) && (! \arg0_1Dcon_isZ_3I#_2_bufchan_buf [0])))
        \arg0_1Dcon_isZ_3I#_2_bufchan_buf  <= \arg0_1Dcon_isZ_3I#_2_bufchan_d ;
  
  /* dcon (Ty TupGo___Bool,
      Dcon TupGo___Bool) : [(arg0_1Dcon_isZ_3I#_2_argbuf,Go),
                            (lizzieLet2_1_argbuf,Bool)] > (boolConvert_1TupGo___Bool_1,TupGo___Bool) */
  assign boolConvert_1TupGo___Bool_1_d = TupGo___Bool_dc((& {\arg0_1Dcon_isZ_3I#_2_argbuf_d [0],
                                                             lizzieLet2_1_argbuf_d[0]}), \arg0_1Dcon_isZ_3I#_2_argbuf_d , lizzieLet2_1_argbuf_d);
  assign {\arg0_1Dcon_isZ_3I#_2_argbuf_r ,
          lizzieLet2_1_argbuf_r} = {2 {(boolConvert_1TupGo___Bool_1_r && boolConvert_1TupGo___Bool_1_d[0])}};
  
  /* mux (Ty Int,
     Ty MyBool) : (arg0_1Dcon_isZ_4,Int) [(lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux,MyBool)] > (lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux,MyBool) */
  assign lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_d = {lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_d[1:1],
                                                                             (arg0_1Dcon_isZ_4_d[0] && lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_d[0])};
  assign lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_r = (lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_r && (arg0_1Dcon_isZ_4_d[0] && lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_d[0]));
  assign arg0_1Dcon_isZ_4_r = (lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_r && (arg0_1Dcon_isZ_4_d[0] && lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_d[0]));
  
  /* demux (Ty MyDTInt_Bool,
       Ty Go) : (arg0_2,MyDTInt_Bool) (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intgo_7,Go) > [(arg0_2Dcon_isZ,Go)] */
  assign arg0_2Dcon_isZ_d = (arg0_2_d[0] && applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intgo_7_d[0]);
  assign applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intgo_7_r = (arg0_2Dcon_isZ_r && (arg0_2_d[0] && applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intgo_7_d[0]));
  assign arg0_2_r = (arg0_2Dcon_isZ_r && (arg0_2_d[0] && applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intgo_7_d[0]));
  
  /* demux (Ty MyDTInt_Int_Int,
       Ty Int) : (arg0_2_1,MyDTInt_Int_Int) (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg1_1,Int) > [(arg0_2_1Dcon_$fNumInt_$c+,Int)] */
  assign \arg0_2_1Dcon_$fNumInt_$c+_d  = {applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg1_1_d[32:1],
                                          (arg0_2_1_d[0] && applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg1_1_d[0])};
  assign applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg1_1_r = (\arg0_2_1Dcon_$fNumInt_$c+_r  && (arg0_2_1_d[0] && applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg1_1_d[0]));
  assign arg0_2_1_r = (\arg0_2_1Dcon_$fNumInt_$c+_r  && (arg0_2_1_d[0] && applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg1_1_d[0]));
  
  /* demux (Ty MyDTInt_Int_Int,
       Ty Int) : (arg0_2_2,MyDTInt_Int_Int) (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg2,Int) > [(arg0_2_2Dcon_$fNumInt_$c+,Int)] */
  assign \arg0_2_2Dcon_$fNumInt_$c+_d  = {applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg2_d[32:1],
                                          (arg0_2_2_d[0] && applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg2_d[0])};
  assign applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg2_r = (\arg0_2_2Dcon_$fNumInt_$c+_r  && (arg0_2_2_d[0] && applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg2_d[0]));
  assign arg0_2_2_r = (\arg0_2_2Dcon_$fNumInt_$c+_r  && (arg0_2_2_d[0] && applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg2_d[0]));
  
  /* fork (Ty Int) : (arg0_2_2Dcon_$fNumInt_$c+,Int) > [(arg0_2_2Dcon_$fNumInt_$c+_1,Int),
                                                   (arg0_2_2Dcon_$fNumInt_$c+_2,Int),
                                                   (arg0_2_2Dcon_$fNumInt_$c+_3,Int),
                                                   (arg0_2_2Dcon_$fNumInt_$c+_4,Int)] */
  logic [3:0] \arg0_2_2Dcon_$fNumInt_$c+_emitted ;
  logic [3:0] \arg0_2_2Dcon_$fNumInt_$c+_done ;
  assign \arg0_2_2Dcon_$fNumInt_$c+_1_d  = {\arg0_2_2Dcon_$fNumInt_$c+_d [32:1],
                                            (\arg0_2_2Dcon_$fNumInt_$c+_d [0] && (! \arg0_2_2Dcon_$fNumInt_$c+_emitted [0]))};
  assign \arg0_2_2Dcon_$fNumInt_$c+_2_d  = {\arg0_2_2Dcon_$fNumInt_$c+_d [32:1],
                                            (\arg0_2_2Dcon_$fNumInt_$c+_d [0] && (! \arg0_2_2Dcon_$fNumInt_$c+_emitted [1]))};
  assign \arg0_2_2Dcon_$fNumInt_$c+_3_d  = {\arg0_2_2Dcon_$fNumInt_$c+_d [32:1],
                                            (\arg0_2_2Dcon_$fNumInt_$c+_d [0] && (! \arg0_2_2Dcon_$fNumInt_$c+_emitted [2]))};
  assign \arg0_2_2Dcon_$fNumInt_$c+_4_d  = {\arg0_2_2Dcon_$fNumInt_$c+_d [32:1],
                                            (\arg0_2_2Dcon_$fNumInt_$c+_d [0] && (! \arg0_2_2Dcon_$fNumInt_$c+_emitted [3]))};
  assign \arg0_2_2Dcon_$fNumInt_$c+_done  = (\arg0_2_2Dcon_$fNumInt_$c+_emitted  | ({\arg0_2_2Dcon_$fNumInt_$c+_4_d [0],
                                                                                     \arg0_2_2Dcon_$fNumInt_$c+_3_d [0],
                                                                                     \arg0_2_2Dcon_$fNumInt_$c+_2_d [0],
                                                                                     \arg0_2_2Dcon_$fNumInt_$c+_1_d [0]} & {\arg0_2_2Dcon_$fNumInt_$c+_4_r ,
                                                                                                                            \arg0_2_2Dcon_$fNumInt_$c+_3_r ,
                                                                                                                            \arg0_2_2Dcon_$fNumInt_$c+_2_r ,
                                                                                                                            \arg0_2_2Dcon_$fNumInt_$c+_1_r }));
  assign \arg0_2_2Dcon_$fNumInt_$c+_r  = (& \arg0_2_2Dcon_$fNumInt_$c+_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \arg0_2_2Dcon_$fNumInt_$c+_emitted  <= 4'd0;
    else
      \arg0_2_2Dcon_$fNumInt_$c+_emitted  <= (\arg0_2_2Dcon_$fNumInt_$c+_r  ? 4'd0 :
                                              \arg0_2_2Dcon_$fNumInt_$c+_done );
  
  /* destruct (Ty Int,
          Dcon I#) : (arg0_2_2Dcon_$fNumInt_$c+_1I#,Int) > [(xa1lV_destruct,Int#)] */
  assign xa1lV_destruct_d = {\arg0_2_2Dcon_$fNumInt_$c+_1I#_d [32:1],
                             \arg0_2_2Dcon_$fNumInt_$c+_1I#_d [0]};
  assign \arg0_2_2Dcon_$fNumInt_$c+_1I#_r  = xa1lV_destruct_r;
  
  /* demux (Ty Int,
       Ty Int) : (arg0_2_2Dcon_$fNumInt_$c+_2,Int) (arg0_2_2Dcon_$fNumInt_$c+_1,Int) > [(arg0_2_2Dcon_$fNumInt_$c+_1I#,Int)] */
  assign \arg0_2_2Dcon_$fNumInt_$c+_1I#_d  = {\arg0_2_2Dcon_$fNumInt_$c+_1_d [32:1],
                                              (\arg0_2_2Dcon_$fNumInt_$c+_2_d [0] && \arg0_2_2Dcon_$fNumInt_$c+_1_d [0])};
  assign \arg0_2_2Dcon_$fNumInt_$c+_1_r  = (\arg0_2_2Dcon_$fNumInt_$c+_1I#_r  && (\arg0_2_2Dcon_$fNumInt_$c+_2_d [0] && \arg0_2_2Dcon_$fNumInt_$c+_1_d [0]));
  assign \arg0_2_2Dcon_$fNumInt_$c+_2_r  = (\arg0_2_2Dcon_$fNumInt_$c+_1I#_r  && (\arg0_2_2Dcon_$fNumInt_$c+_2_d [0] && \arg0_2_2Dcon_$fNumInt_$c+_1_d [0]));
  
  /* demux (Ty Int,
       Ty Int) : (arg0_2_2Dcon_$fNumInt_$c+_3,Int) (arg0_2_1Dcon_$fNumInt_$c+,Int) > [(arg0_2_2Dcon_$fNumInt_$c+_3I#,Int)] */
  assign \arg0_2_2Dcon_$fNumInt_$c+_3I#_d  = {\arg0_2_1Dcon_$fNumInt_$c+_d [32:1],
                                              (\arg0_2_2Dcon_$fNumInt_$c+_3_d [0] && \arg0_2_1Dcon_$fNumInt_$c+_d [0])};
  assign \arg0_2_1Dcon_$fNumInt_$c+_r  = (\arg0_2_2Dcon_$fNumInt_$c+_3I#_r  && (\arg0_2_2Dcon_$fNumInt_$c+_3_d [0] && \arg0_2_1Dcon_$fNumInt_$c+_d [0]));
  assign \arg0_2_2Dcon_$fNumInt_$c+_3_r  = (\arg0_2_2Dcon_$fNumInt_$c+_3I#_r  && (\arg0_2_2Dcon_$fNumInt_$c+_3_d [0] && \arg0_2_1Dcon_$fNumInt_$c+_d [0]));
  
  /* fork (Ty Int) : (arg0_2_2Dcon_$fNumInt_$c+_3I#,Int) > [(arg0_2_2Dcon_$fNumInt_$c+_3I#_1,Int),
                                                       (arg0_2_2Dcon_$fNumInt_$c+_3I#_2,Int),
                                                       (arg0_2_2Dcon_$fNumInt_$c+_3I#_3,Int),
                                                       (arg0_2_2Dcon_$fNumInt_$c+_3I#_4,Int)] */
  logic [3:0] \arg0_2_2Dcon_$fNumInt_$c+_3I#_emitted ;
  logic [3:0] \arg0_2_2Dcon_$fNumInt_$c+_3I#_done ;
  assign \arg0_2_2Dcon_$fNumInt_$c+_3I#_1_d  = {\arg0_2_2Dcon_$fNumInt_$c+_3I#_d [32:1],
                                                (\arg0_2_2Dcon_$fNumInt_$c+_3I#_d [0] && (! \arg0_2_2Dcon_$fNumInt_$c+_3I#_emitted [0]))};
  assign \arg0_2_2Dcon_$fNumInt_$c+_3I#_2_d  = {\arg0_2_2Dcon_$fNumInt_$c+_3I#_d [32:1],
                                                (\arg0_2_2Dcon_$fNumInt_$c+_3I#_d [0] && (! \arg0_2_2Dcon_$fNumInt_$c+_3I#_emitted [1]))};
  assign \arg0_2_2Dcon_$fNumInt_$c+_3I#_3_d  = {\arg0_2_2Dcon_$fNumInt_$c+_3I#_d [32:1],
                                                (\arg0_2_2Dcon_$fNumInt_$c+_3I#_d [0] && (! \arg0_2_2Dcon_$fNumInt_$c+_3I#_emitted [2]))};
  assign \arg0_2_2Dcon_$fNumInt_$c+_3I#_4_d  = {\arg0_2_2Dcon_$fNumInt_$c+_3I#_d [32:1],
                                                (\arg0_2_2Dcon_$fNumInt_$c+_3I#_d [0] && (! \arg0_2_2Dcon_$fNumInt_$c+_3I#_emitted [3]))};
  assign \arg0_2_2Dcon_$fNumInt_$c+_3I#_done  = (\arg0_2_2Dcon_$fNumInt_$c+_3I#_emitted  | ({\arg0_2_2Dcon_$fNumInt_$c+_3I#_4_d [0],
                                                                                             \arg0_2_2Dcon_$fNumInt_$c+_3I#_3_d [0],
                                                                                             \arg0_2_2Dcon_$fNumInt_$c+_3I#_2_d [0],
                                                                                             \arg0_2_2Dcon_$fNumInt_$c+_3I#_1_d [0]} & {\arg0_2_2Dcon_$fNumInt_$c+_3I#_4_r ,
                                                                                                                                        \arg0_2_2Dcon_$fNumInt_$c+_3I#_3_r ,
                                                                                                                                        \arg0_2_2Dcon_$fNumInt_$c+_3I#_2_r ,
                                                                                                                                        \arg0_2_2Dcon_$fNumInt_$c+_3I#_1_r }));
  assign \arg0_2_2Dcon_$fNumInt_$c+_3I#_r  = (& \arg0_2_2Dcon_$fNumInt_$c+_3I#_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \arg0_2_2Dcon_$fNumInt_$c+_3I#_emitted  <= 4'd0;
    else
      \arg0_2_2Dcon_$fNumInt_$c+_3I#_emitted  <= (\arg0_2_2Dcon_$fNumInt_$c+_3I#_r  ? 4'd0 :
                                                  \arg0_2_2Dcon_$fNumInt_$c+_3I#_done );
  
  /* destruct (Ty Int,
          Dcon I#) : (arg0_2_2Dcon_$fNumInt_$c+_3I#_1I#,Int) > [(ya1lW_destruct,Int#)] */
  assign ya1lW_destruct_d = {\arg0_2_2Dcon_$fNumInt_$c+_3I#_1I#_d [32:1],
                             \arg0_2_2Dcon_$fNumInt_$c+_3I#_1I#_d [0]};
  assign \arg0_2_2Dcon_$fNumInt_$c+_3I#_1I#_r  = ya1lW_destruct_r;
  
  /* demux (Ty Int,
       Ty Int) : (arg0_2_2Dcon_$fNumInt_$c+_3I#_2,Int) (arg0_2_2Dcon_$fNumInt_$c+_3I#_1,Int) > [(arg0_2_2Dcon_$fNumInt_$c+_3I#_1I#,Int)] */
  assign \arg0_2_2Dcon_$fNumInt_$c+_3I#_1I#_d  = {\arg0_2_2Dcon_$fNumInt_$c+_3I#_1_d [32:1],
                                                  (\arg0_2_2Dcon_$fNumInt_$c+_3I#_2_d [0] && \arg0_2_2Dcon_$fNumInt_$c+_3I#_1_d [0])};
  assign \arg0_2_2Dcon_$fNumInt_$c+_3I#_1_r  = (\arg0_2_2Dcon_$fNumInt_$c+_3I#_1I#_r  && (\arg0_2_2Dcon_$fNumInt_$c+_3I#_2_d [0] && \arg0_2_2Dcon_$fNumInt_$c+_3I#_1_d [0]));
  assign \arg0_2_2Dcon_$fNumInt_$c+_3I#_2_r  = (\arg0_2_2Dcon_$fNumInt_$c+_3I#_1I#_r  && (\arg0_2_2Dcon_$fNumInt_$c+_3I#_2_d [0] && \arg0_2_2Dcon_$fNumInt_$c+_3I#_1_d [0]));
  
  /* demux (Ty Int,
       Ty Int#) : (arg0_2_2Dcon_$fNumInt_$c+_3I#_3,Int) (xa1lV_destruct,Int#) > [(arg0_2_2Dcon_$fNumInt_$c+_3I#_3I#,Int#)] */
  assign \arg0_2_2Dcon_$fNumInt_$c+_3I#_3I#_d  = {xa1lV_destruct_d[32:1],
                                                  (\arg0_2_2Dcon_$fNumInt_$c+_3I#_3_d [0] && xa1lV_destruct_d[0])};
  assign xa1lV_destruct_r = (\arg0_2_2Dcon_$fNumInt_$c+_3I#_3I#_r  && (\arg0_2_2Dcon_$fNumInt_$c+_3I#_3_d [0] && xa1lV_destruct_d[0]));
  assign \arg0_2_2Dcon_$fNumInt_$c+_3I#_3_r  = (\arg0_2_2Dcon_$fNumInt_$c+_3I#_3I#_r  && (\arg0_2_2Dcon_$fNumInt_$c+_3I#_3_d [0] && xa1lV_destruct_d[0]));
  
  /* op_add (Ty Int#) : (arg0_2_2Dcon_$fNumInt_$c+_3I#_3I#,Int#) (ya1lW_destruct,Int#) > (arg0_2_2Dcon_$fNumInt_$c+_3I#_3I#_1ya1lW_1_Add32,Int#) */
  assign \arg0_2_2Dcon_$fNumInt_$c+_3I#_3I#_1ya1lW_1_Add32_d  = {(\arg0_2_2Dcon_$fNumInt_$c+_3I#_3I#_d [32:1] + ya1lW_destruct_d[32:1]),
                                                                 (\arg0_2_2Dcon_$fNumInt_$c+_3I#_3I#_d [0] && ya1lW_destruct_d[0])};
  assign {\arg0_2_2Dcon_$fNumInt_$c+_3I#_3I#_r ,
          ya1lW_destruct_r} = {2 {(\arg0_2_2Dcon_$fNumInt_$c+_3I#_3I#_1ya1lW_1_Add32_r  && \arg0_2_2Dcon_$fNumInt_$c+_3I#_3I#_1ya1lW_1_Add32_d [0])}};
  
  /* dcon (Ty Int,
      Dcon I#) : [(arg0_2_2Dcon_$fNumInt_$c+_3I#_3I#_1ya1lW_1_Add32,Int#)] > (es_0_1_1I#,Int) */
  assign \es_0_1_1I#_d  = \I#_dc ((& {\arg0_2_2Dcon_$fNumInt_$c+_3I#_3I#_1ya1lW_1_Add32_d [0]}), \arg0_2_2Dcon_$fNumInt_$c+_3I#_3I#_1ya1lW_1_Add32_d );
  assign {\arg0_2_2Dcon_$fNumInt_$c+_3I#_3I#_1ya1lW_1_Add32_r } = {1 {(\es_0_1_1I#_r  && \es_0_1_1I#_d [0])}};
  
  /* mux (Ty Int,
     Ty Int) : (arg0_2_2Dcon_$fNumInt_$c+_3I#_4,Int) [(es_0_1_1I#,Int)] > (es_0_1_1I#_mux,Int) */
  assign \es_0_1_1I#_mux_d  = {\es_0_1_1I#_d [32:1],
                               (\arg0_2_2Dcon_$fNumInt_$c+_3I#_4_d [0] && \es_0_1_1I#_d [0])};
  assign \es_0_1_1I#_r  = (\es_0_1_1I#_mux_r  && (\arg0_2_2Dcon_$fNumInt_$c+_3I#_4_d [0] && \es_0_1_1I#_d [0]));
  assign \arg0_2_2Dcon_$fNumInt_$c+_3I#_4_r  = (\es_0_1_1I#_mux_r  && (\arg0_2_2Dcon_$fNumInt_$c+_3I#_4_d [0] && \es_0_1_1I#_d [0]));
  
  /* mux (Ty Int,
     Ty Int) : (arg0_2_2Dcon_$fNumInt_$c+_4,Int) [(es_0_1_1I#_mux,Int)] > (es_0_1_1I#_mux_mux,Int) */
  assign \es_0_1_1I#_mux_mux_d  = {\es_0_1_1I#_mux_d [32:1],
                                   (\arg0_2_2Dcon_$fNumInt_$c+_4_d [0] && \es_0_1_1I#_mux_d [0])};
  assign \es_0_1_1I#_mux_r  = (\es_0_1_1I#_mux_mux_r  && (\arg0_2_2Dcon_$fNumInt_$c+_4_d [0] && \es_0_1_1I#_mux_d [0]));
  assign \arg0_2_2Dcon_$fNumInt_$c+_4_r  = (\es_0_1_1I#_mux_mux_r  && (\arg0_2_2Dcon_$fNumInt_$c+_4_d [0] && \es_0_1_1I#_mux_d [0]));
  
  /* mux (Ty MyDTInt_Int_Int,
     Ty Int) : (arg0_2_3,MyDTInt_Int_Int) [(es_0_1_1I#_mux_mux,Int)] > (es_0_1_1I#_mux_mux_mux,Int) */
  assign \es_0_1_1I#_mux_mux_mux_d  = {\es_0_1_1I#_mux_mux_d [32:1],
                                       (arg0_2_3_d[0] && \es_0_1_1I#_mux_mux_d [0])};
  assign \es_0_1_1I#_mux_mux_r  = (\es_0_1_1I#_mux_mux_mux_r  && (arg0_2_3_d[0] && \es_0_1_1I#_mux_mux_d [0]));
  assign arg0_2_3_r = (\es_0_1_1I#_mux_mux_mux_r  && (arg0_2_3_d[0] && \es_0_1_1I#_mux_mux_d [0]));
  
  /* mux (Ty MyDTInt_Bool,
     Ty MyBool) : (arg0_3,MyDTInt_Bool) [(lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux,MyBool)] > (lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux,MyBool) */
  assign lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_d = {lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_d[1:1],
                                                                                 (arg0_3_d[0] && lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_d[0])};
  assign lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_r = (lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_r && (arg0_3_d[0] && lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_d[0]));
  assign arg0_3_r = (lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_r && (arg0_3_d[0] && lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_d[0]));
  
  /* destruct (Ty TupGo___Bool,
          Dcon TupGo___Bool) : (boolConvert_1TupGo___Bool_1,TupGo___Bool) > [(boolConvert_1TupGo___Boolgo_1,Go),
                                                                             (boolConvert_1TupGo___Boolbool,Bool)] */
  logic [1:0] boolConvert_1TupGo___Bool_1_emitted;
  logic [1:0] boolConvert_1TupGo___Bool_1_done;
  assign boolConvert_1TupGo___Boolgo_1_d = (boolConvert_1TupGo___Bool_1_d[0] && (! boolConvert_1TupGo___Bool_1_emitted[0]));
  assign boolConvert_1TupGo___Boolbool_d = {boolConvert_1TupGo___Bool_1_d[1:1],
                                            (boolConvert_1TupGo___Bool_1_d[0] && (! boolConvert_1TupGo___Bool_1_emitted[1]))};
  assign boolConvert_1TupGo___Bool_1_done = (boolConvert_1TupGo___Bool_1_emitted | ({boolConvert_1TupGo___Boolbool_d[0],
                                                                                     boolConvert_1TupGo___Boolgo_1_d[0]} & {boolConvert_1TupGo___Boolbool_r,
                                                                                                                            boolConvert_1TupGo___Boolgo_1_r}));
  assign boolConvert_1TupGo___Bool_1_r = (& boolConvert_1TupGo___Bool_1_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) boolConvert_1TupGo___Bool_1_emitted <= 2'd0;
    else
      boolConvert_1TupGo___Bool_1_emitted <= (boolConvert_1TupGo___Bool_1_r ? 2'd0 :
                                              boolConvert_1TupGo___Bool_1_done);
  
  /* fork (Ty Bool) : (boolConvert_1TupGo___Boolbool,Bool) > [(bool_1,Bool),
                                                         (bool_2,Bool)] */
  logic [1:0] boolConvert_1TupGo___Boolbool_emitted;
  logic [1:0] boolConvert_1TupGo___Boolbool_done;
  assign bool_1_d = {boolConvert_1TupGo___Boolbool_d[1:1],
                     (boolConvert_1TupGo___Boolbool_d[0] && (! boolConvert_1TupGo___Boolbool_emitted[0]))};
  assign bool_2_d = {boolConvert_1TupGo___Boolbool_d[1:1],
                     (boolConvert_1TupGo___Boolbool_d[0] && (! boolConvert_1TupGo___Boolbool_emitted[1]))};
  assign boolConvert_1TupGo___Boolbool_done = (boolConvert_1TupGo___Boolbool_emitted | ({bool_2_d[0],
                                                                                         bool_1_d[0]} & {bool_2_r,
                                                                                                         bool_1_r}));
  assign boolConvert_1TupGo___Boolbool_r = (& boolConvert_1TupGo___Boolbool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) boolConvert_1TupGo___Boolbool_emitted <= 2'd0;
    else
      boolConvert_1TupGo___Boolbool_emitted <= (boolConvert_1TupGo___Boolbool_r ? 2'd0 :
                                                boolConvert_1TupGo___Boolbool_done);
  
  /* fork (Ty MyBool) : (boolConvert_1_resbuf,MyBool) > [(lizzieLet3_1,MyBool),
                                                    (lizzieLet3_2,MyBool)] */
  logic [1:0] boolConvert_1_resbuf_emitted;
  logic [1:0] boolConvert_1_resbuf_done;
  assign lizzieLet3_1_d = {boolConvert_1_resbuf_d[1:1],
                           (boolConvert_1_resbuf_d[0] && (! boolConvert_1_resbuf_emitted[0]))};
  assign lizzieLet3_2_d = {boolConvert_1_resbuf_d[1:1],
                           (boolConvert_1_resbuf_d[0] && (! boolConvert_1_resbuf_emitted[1]))};
  assign boolConvert_1_resbuf_done = (boolConvert_1_resbuf_emitted | ({lizzieLet3_2_d[0],
                                                                       lizzieLet3_1_d[0]} & {lizzieLet3_2_r,
                                                                                             lizzieLet3_1_r}));
  assign boolConvert_1_resbuf_r = (& boolConvert_1_resbuf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) boolConvert_1_resbuf_emitted <= 2'd0;
    else
      boolConvert_1_resbuf_emitted <= (boolConvert_1_resbuf_r ? 2'd0 :
                                       boolConvert_1_resbuf_done);
  
  /* demux (Ty Bool,
       Ty Go) : (bool_1,Bool) (boolConvert_1TupGo___Boolgo_1,Go) > [(bool_1False,Go),
                                                                    (bool_1True,Go)] */
  logic [1:0] boolConvert_1TupGo___Boolgo_1_onehotd;
  always_comb
    if ((bool_1_d[0] && boolConvert_1TupGo___Boolgo_1_d[0]))
      unique case (bool_1_d[1:1])
        1'd0: boolConvert_1TupGo___Boolgo_1_onehotd = 2'd1;
        1'd1: boolConvert_1TupGo___Boolgo_1_onehotd = 2'd2;
        default: boolConvert_1TupGo___Boolgo_1_onehotd = 2'd0;
      endcase
    else boolConvert_1TupGo___Boolgo_1_onehotd = 2'd0;
  assign bool_1False_d = boolConvert_1TupGo___Boolgo_1_onehotd[0];
  assign bool_1True_d = boolConvert_1TupGo___Boolgo_1_onehotd[1];
  assign boolConvert_1TupGo___Boolgo_1_r = (| (boolConvert_1TupGo___Boolgo_1_onehotd & {bool_1True_r,
                                                                                        bool_1False_r}));
  assign bool_1_r = boolConvert_1TupGo___Boolgo_1_r;
  
  /* dcon (Ty MyBool,
      Dcon MyFalse) : [(bool_1False,Go)] > (bool_1False_1MyFalse,MyBool) */
  assign bool_1False_1MyFalse_d = MyFalse_dc((& {bool_1False_d[0]}), bool_1False_d);
  assign {bool_1False_r} = {1 {(bool_1False_1MyFalse_r && bool_1False_1MyFalse_d[0])}};
  
  /* buf (Ty MyBool) : (bool_1False_1MyFalsebool_1True_1MyTrue_mux,MyBool) > (boolConvert_1_resbuf,MyBool) */
  MyBool_t bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_d;
  logic bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_r;
  assign bool_1False_1MyFalsebool_1True_1MyTrue_mux_r = ((! bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_d[0]) || bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_d <= {1'd0,
                                                               1'd0};
    else
      if (bool_1False_1MyFalsebool_1True_1MyTrue_mux_r)
        bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_d <= bool_1False_1MyFalsebool_1True_1MyTrue_mux_d;
  MyBool_t bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_buf;
  assign bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_r = (! bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_buf[0]);
  assign boolConvert_1_resbuf_d = (bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_buf[0] ? bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_buf :
                                   bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_buf <= {1'd0,
                                                                 1'd0};
    else
      if ((boolConvert_1_resbuf_r && bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_buf[0]))
        bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_buf <= {1'd0,
                                                                   1'd0};
      else if (((! boolConvert_1_resbuf_r) && (! bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_buf[0])))
        bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_buf <= bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_d;
  
  /* dcon (Ty MyBool,
      Dcon MyTrue) : [(bool_1True,Go)] > (bool_1True_1MyTrue,MyBool) */
  assign bool_1True_1MyTrue_d = MyTrue_dc((& {bool_1True_d[0]}), bool_1True_d);
  assign {bool_1True_r} = {1 {(bool_1True_1MyTrue_r && bool_1True_1MyTrue_d[0])}};
  
  /* mux (Ty Bool,
     Ty MyBool) : (bool_2,Bool) [(bool_1False_1MyFalse,MyBool),
                                 (bool_1True_1MyTrue,MyBool)] > (bool_1False_1MyFalsebool_1True_1MyTrue_mux,MyBool) */
  logic [1:0] bool_1False_1MyFalsebool_1True_1MyTrue_mux_mux;
  logic [1:0] bool_1False_1MyFalsebool_1True_1MyTrue_mux_onehot;
  always_comb
    unique case (bool_2_d[1:1])
      1'd0:
        {bool_1False_1MyFalsebool_1True_1MyTrue_mux_onehot,
         bool_1False_1MyFalsebool_1True_1MyTrue_mux_mux} = {2'd1,
                                                            bool_1False_1MyFalse_d};
      1'd1:
        {bool_1False_1MyFalsebool_1True_1MyTrue_mux_onehot,
         bool_1False_1MyFalsebool_1True_1MyTrue_mux_mux} = {2'd2,
                                                            bool_1True_1MyTrue_d};
      default:
        {bool_1False_1MyFalsebool_1True_1MyTrue_mux_onehot,
         bool_1False_1MyFalsebool_1True_1MyTrue_mux_mux} = {2'd0,
                                                            {1'd0, 1'd0}};
    endcase
  assign bool_1False_1MyFalsebool_1True_1MyTrue_mux_d = {bool_1False_1MyFalsebool_1True_1MyTrue_mux_mux[1:1],
                                                         (bool_1False_1MyFalsebool_1True_1MyTrue_mux_mux[0] && bool_2_d[0])};
  assign bool_2_r = (bool_1False_1MyFalsebool_1True_1MyTrue_mux_d[0] && bool_1False_1MyFalsebool_1True_1MyTrue_mux_r);
  assign {bool_1True_1MyTrue_r,
          bool_1False_1MyFalse_r} = (bool_2_r ? bool_1False_1MyFalsebool_1True_1MyTrue_mux_onehot :
                                     2'd0);
  
  /* destruct (Ty TupGo___Pointer_QTree_Int___Pointer_CT$wnnz,
          Dcon TupGo___Pointer_QTree_Int___Pointer_CT$wnnz) : (call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_1,TupGo___Pointer_QTree_Int___Pointer_CT$wnnz) > [(call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnzgo_8,Go),
                                                                                                                                                                       (call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnzwsmk_1,Pointer_QTree_Int),
                                                                                                                                                                       (call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnzsc_0,Pointer_CT$wnnz)] */
  logic [2:0] call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_1_emitted;
  logic [2:0] call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_1_done;
  assign call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnzgo_8_d = (call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_1_d[0] && (! call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_1_emitted[0]));
  assign call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnzwsmk_1_d = {call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_1_d[16:1],
                                                                          (call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_1_d[0] && (! call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_1_emitted[1]))};
  assign call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnzsc_0_d = {call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_1_d[32:17],
                                                                        (call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_1_d[0] && (! call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_1_emitted[2]))};
  assign call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_1_done = (call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_1_emitted | ({call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnzsc_0_d[0],
                                                                                                                                             call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnzwsmk_1_d[0],
                                                                                                                                             call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnzgo_8_d[0]} & {call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnzsc_0_r,
                                                                                                                                                                                                                call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnzwsmk_1_r,
                                                                                                                                                                                                                call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnzgo_8_r}));
  assign call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_1_r = (& call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_1_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_1_emitted <= 3'd0;
    else
      call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_1_emitted <= (call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_1_r ? 3'd0 :
                                                                          call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_1_done);
  
  /* rbuf (Ty Go) : (call_$wnnz_goConst,Go) > (call_$wnnz_initBufi,Go) */
  Go_t call_$wnnz_goConst_buf;
  assign call_$wnnz_goConst_r = (! call_$wnnz_goConst_buf[0]);
  assign call_$wnnz_initBufi_d = (call_$wnnz_goConst_buf[0] ? call_$wnnz_goConst_buf :
                                  call_$wnnz_goConst_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_$wnnz_goConst_buf <= 1'd0;
    else
      if ((call_$wnnz_initBufi_r && call_$wnnz_goConst_buf[0]))
        call_$wnnz_goConst_buf <= 1'd0;
      else if (((! call_$wnnz_initBufi_r) && (! call_$wnnz_goConst_buf[0])))
        call_$wnnz_goConst_buf <= call_$wnnz_goConst_d;
  
  /* mergectrl (Ty C5,Ty Go) : [(call_$wnnz_goMux1,Go),
                           (lizzieLet58_3Lcall_$wnnz3_1_argbuf,Go),
                           (lizzieLet58_3Lcall_$wnnz2_1_argbuf,Go),
                           (lizzieLet58_3Lcall_$wnnz1_1_argbuf,Go),
                           (lizzieLet4_3QNode_Int_1_argbuf,Go)] > (go_8_goMux_choice,C5) (go_8_goMux_data,Go) */
  logic [4:0] call_$wnnz_goMux1_select_d;
  assign call_$wnnz_goMux1_select_d = ((| call_$wnnz_goMux1_select_q) ? call_$wnnz_goMux1_select_q :
                                       (call_$wnnz_goMux1_d[0] ? 5'd1 :
                                        (lizzieLet58_3Lcall_$wnnz3_1_argbuf_d[0] ? 5'd2 :
                                         (lizzieLet58_3Lcall_$wnnz2_1_argbuf_d[0] ? 5'd4 :
                                          (lizzieLet58_3Lcall_$wnnz1_1_argbuf_d[0] ? 5'd8 :
                                           (lizzieLet4_3QNode_Int_1_argbuf_d[0] ? 5'd16 :
                                            5'd0))))));
  logic [4:0] call_$wnnz_goMux1_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_$wnnz_goMux1_select_q <= 5'd0;
    else
      call_$wnnz_goMux1_select_q <= (call_$wnnz_goMux1_done ? 5'd0 :
                                     call_$wnnz_goMux1_select_d);
  logic [1:0] call_$wnnz_goMux1_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_$wnnz_goMux1_emit_q <= 2'd0;
    else
      call_$wnnz_goMux1_emit_q <= (call_$wnnz_goMux1_done ? 2'd0 :
                                   call_$wnnz_goMux1_emit_d);
  logic [1:0] call_$wnnz_goMux1_emit_d;
  assign call_$wnnz_goMux1_emit_d = (call_$wnnz_goMux1_emit_q | ({go_8_goMux_choice_d[0],
                                                                  go_8_goMux_data_d[0]} & {go_8_goMux_choice_r,
                                                                                           go_8_goMux_data_r}));
  logic call_$wnnz_goMux1_done;
  assign call_$wnnz_goMux1_done = (& call_$wnnz_goMux1_emit_d);
  assign {lizzieLet4_3QNode_Int_1_argbuf_r,
          lizzieLet58_3Lcall_$wnnz1_1_argbuf_r,
          lizzieLet58_3Lcall_$wnnz2_1_argbuf_r,
          lizzieLet58_3Lcall_$wnnz3_1_argbuf_r,
          call_$wnnz_goMux1_r} = (call_$wnnz_goMux1_done ? call_$wnnz_goMux1_select_d :
                                  5'd0);
  assign go_8_goMux_data_d = ((call_$wnnz_goMux1_select_d[0] && (! call_$wnnz_goMux1_emit_q[0])) ? call_$wnnz_goMux1_d :
                              ((call_$wnnz_goMux1_select_d[1] && (! call_$wnnz_goMux1_emit_q[0])) ? lizzieLet58_3Lcall_$wnnz3_1_argbuf_d :
                               ((call_$wnnz_goMux1_select_d[2] && (! call_$wnnz_goMux1_emit_q[0])) ? lizzieLet58_3Lcall_$wnnz2_1_argbuf_d :
                                ((call_$wnnz_goMux1_select_d[3] && (! call_$wnnz_goMux1_emit_q[0])) ? lizzieLet58_3Lcall_$wnnz1_1_argbuf_d :
                                 ((call_$wnnz_goMux1_select_d[4] && (! call_$wnnz_goMux1_emit_q[0])) ? lizzieLet4_3QNode_Int_1_argbuf_d :
                                  1'd0)))));
  assign go_8_goMux_choice_d = ((call_$wnnz_goMux1_select_d[0] && (! call_$wnnz_goMux1_emit_q[1])) ? C1_5_dc(1'd1) :
                                ((call_$wnnz_goMux1_select_d[1] && (! call_$wnnz_goMux1_emit_q[1])) ? C2_5_dc(1'd1) :
                                 ((call_$wnnz_goMux1_select_d[2] && (! call_$wnnz_goMux1_emit_q[1])) ? C3_5_dc(1'd1) :
                                  ((call_$wnnz_goMux1_select_d[3] && (! call_$wnnz_goMux1_emit_q[1])) ? C4_5_dc(1'd1) :
                                   ((call_$wnnz_goMux1_select_d[4] && (! call_$wnnz_goMux1_emit_q[1])) ? C5_5_dc(1'd1) :
                                    {3'd0, 1'd0})))));
  
  /* fork (Ty Go) : (call_$wnnz_initBuf,Go) > [(call_$wnnz_unlockFork1,Go),
                                          (call_$wnnz_unlockFork2,Go),
                                          (call_$wnnz_unlockFork3,Go)] */
  logic [2:0] call_$wnnz_initBuf_emitted;
  logic [2:0] call_$wnnz_initBuf_done;
  assign call_$wnnz_unlockFork1_d = (call_$wnnz_initBuf_d[0] && (! call_$wnnz_initBuf_emitted[0]));
  assign call_$wnnz_unlockFork2_d = (call_$wnnz_initBuf_d[0] && (! call_$wnnz_initBuf_emitted[1]));
  assign call_$wnnz_unlockFork3_d = (call_$wnnz_initBuf_d[0] && (! call_$wnnz_initBuf_emitted[2]));
  assign call_$wnnz_initBuf_done = (call_$wnnz_initBuf_emitted | ({call_$wnnz_unlockFork3_d[0],
                                                                   call_$wnnz_unlockFork2_d[0],
                                                                   call_$wnnz_unlockFork1_d[0]} & {call_$wnnz_unlockFork3_r,
                                                                                                   call_$wnnz_unlockFork2_r,
                                                                                                   call_$wnnz_unlockFork1_r}));
  assign call_$wnnz_initBuf_r = (& call_$wnnz_initBuf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_$wnnz_initBuf_emitted <= 3'd0;
    else
      call_$wnnz_initBuf_emitted <= (call_$wnnz_initBuf_r ? 3'd0 :
                                     call_$wnnz_initBuf_done);
  
  /* initbuf (Ty Go,
         Dcon Go) : (call_$wnnz_initBufi,Go) > (call_$wnnz_initBuf,Go) */
  assign call_$wnnz_initBufi_r = ((! call_$wnnz_initBuf_d[0]) || call_$wnnz_initBuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_$wnnz_initBuf_d <= Go_dc(1'd1);
    else
      if (call_$wnnz_initBufi_r)
        call_$wnnz_initBuf_d <= call_$wnnz_initBufi_d;
  
  /* mux (Ty Go,
     Ty Go) : (call_$wnnz_unlockFork1,Go) [(call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnzgo_8,Go)] > (call_$wnnz_goMux1,Go) */
  assign call_$wnnz_goMux1_d = (call_$wnnz_unlockFork1_d[0] && call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnzgo_8_d[0]);
  assign call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnzgo_8_r = (call_$wnnz_goMux1_r && (call_$wnnz_unlockFork1_d[0] && call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnzgo_8_d[0]));
  assign call_$wnnz_unlockFork1_r = (call_$wnnz_goMux1_r && (call_$wnnz_unlockFork1_d[0] && call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnzgo_8_d[0]));
  
  /* mux (Ty Go,
     Ty Pointer_QTree_Int) : (call_$wnnz_unlockFork2,Go) [(call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnzwsmk_1,Pointer_QTree_Int)] > (call_$wnnz_goMux2,Pointer_QTree_Int) */
  assign call_$wnnz_goMux2_d = {call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnzwsmk_1_d[16:1],
                                (call_$wnnz_unlockFork2_d[0] && call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnzwsmk_1_d[0])};
  assign call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnzwsmk_1_r = (call_$wnnz_goMux2_r && (call_$wnnz_unlockFork2_d[0] && call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnzwsmk_1_d[0]));
  assign call_$wnnz_unlockFork2_r = (call_$wnnz_goMux2_r && (call_$wnnz_unlockFork2_d[0] && call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnzwsmk_1_d[0]));
  
  /* mux (Ty Go,
     Ty Pointer_CT$wnnz) : (call_$wnnz_unlockFork3,Go) [(call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnzsc_0,Pointer_CT$wnnz)] > (call_$wnnz_goMux3,Pointer_CT$wnnz) */
  assign call_$wnnz_goMux3_d = {call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnzsc_0_d[16:1],
                                (call_$wnnz_unlockFork3_d[0] && call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnzsc_0_d[0])};
  assign call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnzsc_0_r = (call_$wnnz_goMux3_r && (call_$wnnz_unlockFork3_d[0] && call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnzsc_0_d[0]));
  assign call_$wnnz_unlockFork3_r = (call_$wnnz_goMux3_r && (call_$wnnz_unlockFork3_d[0] && call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnzsc_0_d[0]));
  
  /* destruct (Ty TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf''''''''''''_f''''''''''''_Int,
          Dcon TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf''''''''''''_f''''''''''''_Int) : (call_f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf''''''''''''_f''''''''''''_Int_1,TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf''''''''''''_f''''''''''''_Int) > [(call_f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf''''''''''''_f''''''''''''_Intgo_9,Go),
                                                                                                                                                                                                                                                                                                                                                                                                                                              (call_f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf''''''''''''_f''''''''''''_Intq4afj,Pointer_QTree_Int),
                                                                                                                                                                                                                                                                                                                                                                                                                                              (call_f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf''''''''''''_f''''''''''''_Intt4afk,Pointer_QTree_Int),
                                                                                                                                                                                                                                                                                                                                                                                                                                              (call_f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf''''''''''''_f''''''''''''_Intis_zafl,MyDTInt_Bool),
                                                                                                                                                                                                                                                                                                                                                                                                                                              (call_f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf''''''''''''_f''''''''''''_Intop_addafm,MyDTInt_Int_Int),
                                                                                                                                                                                                                                                                                                                                                                                                                                              (call_f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf''''''''''''_f''''''''''''_Intsc_0_1,Pointer_CTf''''''''''''_f''''''''''''_Int)] */
  logic [5:0] \call_f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf''''''''''''_f''''''''''''_Int_1_emitted ;
  logic [5:0] \call_f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf''''''''''''_f''''''''''''_Int_1_done ;
  assign \call_f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf''''''''''''_f''''''''''''_Intgo_9_d  = (\call_f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf''''''''''''_f''''''''''''_Int_1_d [0] && (! \call_f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf''''''''''''_f''''''''''''_Int_1_emitted [0]));
  assign \call_f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf''''''''''''_f''''''''''''_Intq4afj_d  = {\call_f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf''''''''''''_f''''''''''''_Int_1_d [16:1],
                                                                                                                                                                                    (\call_f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf''''''''''''_f''''''''''''_Int_1_d [0] && (! \call_f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf''''''''''''_f''''''''''''_Int_1_emitted [1]))};
  assign \call_f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf''''''''''''_f''''''''''''_Intt4afk_d  = {\call_f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf''''''''''''_f''''''''''''_Int_1_d [32:17],
                                                                                                                                                                                    (\call_f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf''''''''''''_f''''''''''''_Int_1_d [0] && (! \call_f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf''''''''''''_f''''''''''''_Int_1_emitted [2]))};
  assign \call_f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf''''''''''''_f''''''''''''_Intis_zafl_d  = (\call_f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf''''''''''''_f''''''''''''_Int_1_d [0] && (! \call_f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf''''''''''''_f''''''''''''_Int_1_emitted [3]));
  assign \call_f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf''''''''''''_f''''''''''''_Intop_addafm_d  = (\call_f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf''''''''''''_f''''''''''''_Int_1_d [0] && (! \call_f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf''''''''''''_f''''''''''''_Int_1_emitted [4]));
  assign \call_f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf''''''''''''_f''''''''''''_Intsc_0_1_d  = {\call_f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf''''''''''''_f''''''''''''_Int_1_d [48:33],
                                                                                                                                                                                     (\call_f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf''''''''''''_f''''''''''''_Int_1_d [0] && (! \call_f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf''''''''''''_f''''''''''''_Int_1_emitted [5]))};
  assign \call_f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf''''''''''''_f''''''''''''_Int_1_done  = (\call_f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf''''''''''''_f''''''''''''_Int_1_emitted  | ({\call_f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf''''''''''''_f''''''''''''_Intsc_0_1_d [0],
                                                                                                                                                                                                                                                                                                                                                                   \call_f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf''''''''''''_f''''''''''''_Intop_addafm_d [0],
                                                                                                                                                                                                                                                                                                                                                                   \call_f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf''''''''''''_f''''''''''''_Intis_zafl_d [0],
                                                                                                                                                                                                                                                                                                                                                                   \call_f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf''''''''''''_f''''''''''''_Intt4afk_d [0],
                                                                                                                                                                                                                                                                                                                                                                   \call_f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf''''''''''''_f''''''''''''_Intq4afj_d [0],
                                                                                                                                                                                                                                                                                                                                                                   \call_f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf''''''''''''_f''''''''''''_Intgo_9_d [0]} & {\call_f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf''''''''''''_f''''''''''''_Intsc_0_1_r ,
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 \call_f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf''''''''''''_f''''''''''''_Intop_addafm_r ,
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 \call_f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf''''''''''''_f''''''''''''_Intis_zafl_r ,
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 \call_f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf''''''''''''_f''''''''''''_Intt4afk_r ,
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 \call_f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf''''''''''''_f''''''''''''_Intq4afj_r ,
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 \call_f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf''''''''''''_f''''''''''''_Intgo_9_r }));
  assign \call_f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf''''''''''''_f''''''''''''_Int_1_r  = (& \call_f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf''''''''''''_f''''''''''''_Int_1_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \call_f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf''''''''''''_f''''''''''''_Int_1_emitted  <= 6'd0;
    else
      \call_f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf''''''''''''_f''''''''''''_Int_1_emitted  <= (\call_f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf''''''''''''_f''''''''''''_Int_1_r  ? 6'd0 :
                                                                                                                                                                                     \call_f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf''''''''''''_f''''''''''''_Int_1_done );
  
  /* rbuf (Ty Go) : (call_f''''''''''''_f''''''''''''_Int_goConst,Go) > (call_f''''''''''''_f''''''''''''_Int_initBufi,Go) */
  Go_t \call_f''''''''''''_f''''''''''''_Int_goConst_buf ;
  assign \call_f''''''''''''_f''''''''''''_Int_goConst_r  = (! \call_f''''''''''''_f''''''''''''_Int_goConst_buf [0]);
  assign \call_f''''''''''''_f''''''''''''_Int_initBufi_d  = (\call_f''''''''''''_f''''''''''''_Int_goConst_buf [0] ? \call_f''''''''''''_f''''''''''''_Int_goConst_buf  :
                                                              \call_f''''''''''''_f''''''''''''_Int_goConst_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \call_f''''''''''''_f''''''''''''_Int_goConst_buf  <= 1'd0;
    else
      if ((\call_f''''''''''''_f''''''''''''_Int_initBufi_r  && \call_f''''''''''''_f''''''''''''_Int_goConst_buf [0]))
        \call_f''''''''''''_f''''''''''''_Int_goConst_buf  <= 1'd0;
      else if (((! \call_f''''''''''''_f''''''''''''_Int_initBufi_r ) && (! \call_f''''''''''''_f''''''''''''_Int_goConst_buf [0])))
        \call_f''''''''''''_f''''''''''''_Int_goConst_buf  <= \call_f''''''''''''_f''''''''''''_Int_goConst_d ;
  
  /* mergectrl (Ty C5,
           Ty Go) : [(call_f''''''''''''_f''''''''''''_Int_goMux1,Go),
                     (lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int3_1_argbuf,Go),
                     (lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int2_1_argbuf,Go),
                     (lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int1_1_argbuf,Go),
                     (lizzieLet6_5QNode_Int_3QNode_Int_1_argbuf,Go)] > (go_9_goMux_choice,C5) (go_9_goMux_data,Go) */
  logic [4:0] \call_f''''''''''''_f''''''''''''_Int_goMux1_select_d ;
  assign \call_f''''''''''''_f''''''''''''_Int_goMux1_select_d  = ((| \call_f''''''''''''_f''''''''''''_Int_goMux1_select_q ) ? \call_f''''''''''''_f''''''''''''_Int_goMux1_select_q  :
                                                                   (\call_f''''''''''''_f''''''''''''_Int_goMux1_d [0] ? 5'd1 :
                                                                    (\lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int3_1_argbuf_d [0] ? 5'd2 :
                                                                     (\lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int2_1_argbuf_d [0] ? 5'd4 :
                                                                      (\lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int1_1_argbuf_d [0] ? 5'd8 :
                                                                       (lizzieLet6_5QNode_Int_3QNode_Int_1_argbuf_d[0] ? 5'd16 :
                                                                        5'd0))))));
  logic [4:0] \call_f''''''''''''_f''''''''''''_Int_goMux1_select_q ;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \call_f''''''''''''_f''''''''''''_Int_goMux1_select_q  <= 5'd0;
    else
      \call_f''''''''''''_f''''''''''''_Int_goMux1_select_q  <= (\call_f''''''''''''_f''''''''''''_Int_goMux1_done  ? 5'd0 :
                                                                 \call_f''''''''''''_f''''''''''''_Int_goMux1_select_d );
  logic [1:0] \call_f''''''''''''_f''''''''''''_Int_goMux1_emit_q ;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \call_f''''''''''''_f''''''''''''_Int_goMux1_emit_q  <= 2'd0;
    else
      \call_f''''''''''''_f''''''''''''_Int_goMux1_emit_q  <= (\call_f''''''''''''_f''''''''''''_Int_goMux1_done  ? 2'd0 :
                                                               \call_f''''''''''''_f''''''''''''_Int_goMux1_emit_d );
  logic [1:0] \call_f''''''''''''_f''''''''''''_Int_goMux1_emit_d ;
  assign \call_f''''''''''''_f''''''''''''_Int_goMux1_emit_d  = (\call_f''''''''''''_f''''''''''''_Int_goMux1_emit_q  | ({go_9_goMux_choice_d[0],
                                                                                                                          go_9_goMux_data_d[0]} & {go_9_goMux_choice_r,
                                                                                                                                                   go_9_goMux_data_r}));
  logic \call_f''''''''''''_f''''''''''''_Int_goMux1_done ;
  assign \call_f''''''''''''_f''''''''''''_Int_goMux1_done  = (& \call_f''''''''''''_f''''''''''''_Int_goMux1_emit_d );
  assign {lizzieLet6_5QNode_Int_3QNode_Int_1_argbuf_r,
          \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int1_1_argbuf_r ,
          \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int2_1_argbuf_r ,
          \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int3_1_argbuf_r ,
          \call_f''''''''''''_f''''''''''''_Int_goMux1_r } = (\call_f''''''''''''_f''''''''''''_Int_goMux1_done  ? \call_f''''''''''''_f''''''''''''_Int_goMux1_select_d  :
                                                              5'd0);
  assign go_9_goMux_data_d = ((\call_f''''''''''''_f''''''''''''_Int_goMux1_select_d [0] && (! \call_f''''''''''''_f''''''''''''_Int_goMux1_emit_q [0])) ? \call_f''''''''''''_f''''''''''''_Int_goMux1_d  :
                              ((\call_f''''''''''''_f''''''''''''_Int_goMux1_select_d [1] && (! \call_f''''''''''''_f''''''''''''_Int_goMux1_emit_q [0])) ? \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int3_1_argbuf_d  :
                               ((\call_f''''''''''''_f''''''''''''_Int_goMux1_select_d [2] && (! \call_f''''''''''''_f''''''''''''_Int_goMux1_emit_q [0])) ? \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int2_1_argbuf_d  :
                                ((\call_f''''''''''''_f''''''''''''_Int_goMux1_select_d [3] && (! \call_f''''''''''''_f''''''''''''_Int_goMux1_emit_q [0])) ? \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int1_1_argbuf_d  :
                                 ((\call_f''''''''''''_f''''''''''''_Int_goMux1_select_d [4] && (! \call_f''''''''''''_f''''''''''''_Int_goMux1_emit_q [0])) ? lizzieLet6_5QNode_Int_3QNode_Int_1_argbuf_d :
                                  1'd0)))));
  assign go_9_goMux_choice_d = ((\call_f''''''''''''_f''''''''''''_Int_goMux1_select_d [0] && (! \call_f''''''''''''_f''''''''''''_Int_goMux1_emit_q [1])) ? C1_5_dc(1'd1) :
                                ((\call_f''''''''''''_f''''''''''''_Int_goMux1_select_d [1] && (! \call_f''''''''''''_f''''''''''''_Int_goMux1_emit_q [1])) ? C2_5_dc(1'd1) :
                                 ((\call_f''''''''''''_f''''''''''''_Int_goMux1_select_d [2] && (! \call_f''''''''''''_f''''''''''''_Int_goMux1_emit_q [1])) ? C3_5_dc(1'd1) :
                                  ((\call_f''''''''''''_f''''''''''''_Int_goMux1_select_d [3] && (! \call_f''''''''''''_f''''''''''''_Int_goMux1_emit_q [1])) ? C4_5_dc(1'd1) :
                                   ((\call_f''''''''''''_f''''''''''''_Int_goMux1_select_d [4] && (! \call_f''''''''''''_f''''''''''''_Int_goMux1_emit_q [1])) ? C5_5_dc(1'd1) :
                                    {3'd0, 1'd0})))));
  
  /* fork (Ty Go) : (call_f''''''''''''_f''''''''''''_Int_initBuf,Go) > [(call_f''''''''''''_f''''''''''''_Int_unlockFork1,Go),
                                                                    (call_f''''''''''''_f''''''''''''_Int_unlockFork2,Go),
                                                                    (call_f''''''''''''_f''''''''''''_Int_unlockFork3,Go),
                                                                    (call_f''''''''''''_f''''''''''''_Int_unlockFork4,Go),
                                                                    (call_f''''''''''''_f''''''''''''_Int_unlockFork5,Go),
                                                                    (call_f''''''''''''_f''''''''''''_Int_unlockFork6,Go)] */
  logic [5:0] \call_f''''''''''''_f''''''''''''_Int_initBuf_emitted ;
  logic [5:0] \call_f''''''''''''_f''''''''''''_Int_initBuf_done ;
  assign \call_f''''''''''''_f''''''''''''_Int_unlockFork1_d  = (\call_f''''''''''''_f''''''''''''_Int_initBuf_d [0] && (! \call_f''''''''''''_f''''''''''''_Int_initBuf_emitted [0]));
  assign \call_f''''''''''''_f''''''''''''_Int_unlockFork2_d  = (\call_f''''''''''''_f''''''''''''_Int_initBuf_d [0] && (! \call_f''''''''''''_f''''''''''''_Int_initBuf_emitted [1]));
  assign \call_f''''''''''''_f''''''''''''_Int_unlockFork3_d  = (\call_f''''''''''''_f''''''''''''_Int_initBuf_d [0] && (! \call_f''''''''''''_f''''''''''''_Int_initBuf_emitted [2]));
  assign \call_f''''''''''''_f''''''''''''_Int_unlockFork4_d  = (\call_f''''''''''''_f''''''''''''_Int_initBuf_d [0] && (! \call_f''''''''''''_f''''''''''''_Int_initBuf_emitted [3]));
  assign \call_f''''''''''''_f''''''''''''_Int_unlockFork5_d  = (\call_f''''''''''''_f''''''''''''_Int_initBuf_d [0] && (! \call_f''''''''''''_f''''''''''''_Int_initBuf_emitted [4]));
  assign \call_f''''''''''''_f''''''''''''_Int_unlockFork6_d  = (\call_f''''''''''''_f''''''''''''_Int_initBuf_d [0] && (! \call_f''''''''''''_f''''''''''''_Int_initBuf_emitted [5]));
  assign \call_f''''''''''''_f''''''''''''_Int_initBuf_done  = (\call_f''''''''''''_f''''''''''''_Int_initBuf_emitted  | ({\call_f''''''''''''_f''''''''''''_Int_unlockFork6_d [0],
                                                                                                                           \call_f''''''''''''_f''''''''''''_Int_unlockFork5_d [0],
                                                                                                                           \call_f''''''''''''_f''''''''''''_Int_unlockFork4_d [0],
                                                                                                                           \call_f''''''''''''_f''''''''''''_Int_unlockFork3_d [0],
                                                                                                                           \call_f''''''''''''_f''''''''''''_Int_unlockFork2_d [0],
                                                                                                                           \call_f''''''''''''_f''''''''''''_Int_unlockFork1_d [0]} & {\call_f''''''''''''_f''''''''''''_Int_unlockFork6_r ,
                                                                                                                                                                                       \call_f''''''''''''_f''''''''''''_Int_unlockFork5_r ,
                                                                                                                                                                                       \call_f''''''''''''_f''''''''''''_Int_unlockFork4_r ,
                                                                                                                                                                                       \call_f''''''''''''_f''''''''''''_Int_unlockFork3_r ,
                                                                                                                                                                                       \call_f''''''''''''_f''''''''''''_Int_unlockFork2_r ,
                                                                                                                                                                                       \call_f''''''''''''_f''''''''''''_Int_unlockFork1_r }));
  assign \call_f''''''''''''_f''''''''''''_Int_initBuf_r  = (& \call_f''''''''''''_f''''''''''''_Int_initBuf_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \call_f''''''''''''_f''''''''''''_Int_initBuf_emitted  <= 6'd0;
    else
      \call_f''''''''''''_f''''''''''''_Int_initBuf_emitted  <= (\call_f''''''''''''_f''''''''''''_Int_initBuf_r  ? 6'd0 :
                                                                 \call_f''''''''''''_f''''''''''''_Int_initBuf_done );
  
  /* initbuf (Ty Go,
         Dcon Go) : (call_f''''''''''''_f''''''''''''_Int_initBufi,Go) > (call_f''''''''''''_f''''''''''''_Int_initBuf,Go) */
  assign \call_f''''''''''''_f''''''''''''_Int_initBufi_r  = ((! \call_f''''''''''''_f''''''''''''_Int_initBuf_d [0]) || \call_f''''''''''''_f''''''''''''_Int_initBuf_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \call_f''''''''''''_f''''''''''''_Int_initBuf_d  <= Go_dc(1'd1);
    else
      if (\call_f''''''''''''_f''''''''''''_Int_initBufi_r )
        \call_f''''''''''''_f''''''''''''_Int_initBuf_d  <= \call_f''''''''''''_f''''''''''''_Int_initBufi_d ;
  
  /* mux (Ty Go,
     Ty Go) : (call_f''''''''''''_f''''''''''''_Int_unlockFork1,Go) [(call_f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf''''''''''''_f''''''''''''_Intgo_9,Go)] > (call_f''''''''''''_f''''''''''''_Int_goMux1,Go) */
  assign \call_f''''''''''''_f''''''''''''_Int_goMux1_d  = (\call_f''''''''''''_f''''''''''''_Int_unlockFork1_d [0] && \call_f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf''''''''''''_f''''''''''''_Intgo_9_d [0]);
  assign \call_f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf''''''''''''_f''''''''''''_Intgo_9_r  = (\call_f''''''''''''_f''''''''''''_Int_goMux1_r  && (\call_f''''''''''''_f''''''''''''_Int_unlockFork1_d [0] && \call_f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf''''''''''''_f''''''''''''_Intgo_9_d [0]));
  assign \call_f''''''''''''_f''''''''''''_Int_unlockFork1_r  = (\call_f''''''''''''_f''''''''''''_Int_goMux1_r  && (\call_f''''''''''''_f''''''''''''_Int_unlockFork1_d [0] && \call_f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf''''''''''''_f''''''''''''_Intgo_9_d [0]));
  
  /* mux (Ty Go,
     Ty Pointer_QTree_Int) : (call_f''''''''''''_f''''''''''''_Int_unlockFork2,Go) [(call_f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf''''''''''''_f''''''''''''_Intq4afj,Pointer_QTree_Int)] > (call_f''''''''''''_f''''''''''''_Int_goMux2,Pointer_QTree_Int) */
  assign \call_f''''''''''''_f''''''''''''_Int_goMux2_d  = {\call_f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf''''''''''''_f''''''''''''_Intq4afj_d [16:1],
                                                            (\call_f''''''''''''_f''''''''''''_Int_unlockFork2_d [0] && \call_f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf''''''''''''_f''''''''''''_Intq4afj_d [0])};
  assign \call_f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf''''''''''''_f''''''''''''_Intq4afj_r  = (\call_f''''''''''''_f''''''''''''_Int_goMux2_r  && (\call_f''''''''''''_f''''''''''''_Int_unlockFork2_d [0] && \call_f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf''''''''''''_f''''''''''''_Intq4afj_d [0]));
  assign \call_f''''''''''''_f''''''''''''_Int_unlockFork2_r  = (\call_f''''''''''''_f''''''''''''_Int_goMux2_r  && (\call_f''''''''''''_f''''''''''''_Int_unlockFork2_d [0] && \call_f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf''''''''''''_f''''''''''''_Intq4afj_d [0]));
  
  /* mux (Ty Go,
     Ty Pointer_QTree_Int) : (call_f''''''''''''_f''''''''''''_Int_unlockFork3,Go) [(call_f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf''''''''''''_f''''''''''''_Intt4afk,Pointer_QTree_Int)] > (call_f''''''''''''_f''''''''''''_Int_goMux3,Pointer_QTree_Int) */
  assign \call_f''''''''''''_f''''''''''''_Int_goMux3_d  = {\call_f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf''''''''''''_f''''''''''''_Intt4afk_d [16:1],
                                                            (\call_f''''''''''''_f''''''''''''_Int_unlockFork3_d [0] && \call_f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf''''''''''''_f''''''''''''_Intt4afk_d [0])};
  assign \call_f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf''''''''''''_f''''''''''''_Intt4afk_r  = (\call_f''''''''''''_f''''''''''''_Int_goMux3_r  && (\call_f''''''''''''_f''''''''''''_Int_unlockFork3_d [0] && \call_f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf''''''''''''_f''''''''''''_Intt4afk_d [0]));
  assign \call_f''''''''''''_f''''''''''''_Int_unlockFork3_r  = (\call_f''''''''''''_f''''''''''''_Int_goMux3_r  && (\call_f''''''''''''_f''''''''''''_Int_unlockFork3_d [0] && \call_f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf''''''''''''_f''''''''''''_Intt4afk_d [0]));
  
  /* mux (Ty Go,
     Ty MyDTInt_Bool) : (call_f''''''''''''_f''''''''''''_Int_unlockFork4,Go) [(call_f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf''''''''''''_f''''''''''''_Intis_zafl,MyDTInt_Bool)] > (call_f''''''''''''_f''''''''''''_Int_goMux4,MyDTInt_Bool) */
  assign \call_f''''''''''''_f''''''''''''_Int_goMux4_d  = (\call_f''''''''''''_f''''''''''''_Int_unlockFork4_d [0] && \call_f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf''''''''''''_f''''''''''''_Intis_zafl_d [0]);
  assign \call_f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf''''''''''''_f''''''''''''_Intis_zafl_r  = (\call_f''''''''''''_f''''''''''''_Int_goMux4_r  && (\call_f''''''''''''_f''''''''''''_Int_unlockFork4_d [0] && \call_f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf''''''''''''_f''''''''''''_Intis_zafl_d [0]));
  assign \call_f''''''''''''_f''''''''''''_Int_unlockFork4_r  = (\call_f''''''''''''_f''''''''''''_Int_goMux4_r  && (\call_f''''''''''''_f''''''''''''_Int_unlockFork4_d [0] && \call_f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf''''''''''''_f''''''''''''_Intis_zafl_d [0]));
  
  /* mux (Ty Go,
     Ty MyDTInt_Int_Int) : (call_f''''''''''''_f''''''''''''_Int_unlockFork5,Go) [(call_f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf''''''''''''_f''''''''''''_Intop_addafm,MyDTInt_Int_Int)] > (call_f''''''''''''_f''''''''''''_Int_goMux5,MyDTInt_Int_Int) */
  assign \call_f''''''''''''_f''''''''''''_Int_goMux5_d  = (\call_f''''''''''''_f''''''''''''_Int_unlockFork5_d [0] && \call_f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf''''''''''''_f''''''''''''_Intop_addafm_d [0]);
  assign \call_f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf''''''''''''_f''''''''''''_Intop_addafm_r  = (\call_f''''''''''''_f''''''''''''_Int_goMux5_r  && (\call_f''''''''''''_f''''''''''''_Int_unlockFork5_d [0] && \call_f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf''''''''''''_f''''''''''''_Intop_addafm_d [0]));
  assign \call_f''''''''''''_f''''''''''''_Int_unlockFork5_r  = (\call_f''''''''''''_f''''''''''''_Int_goMux5_r  && (\call_f''''''''''''_f''''''''''''_Int_unlockFork5_d [0] && \call_f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf''''''''''''_f''''''''''''_Intop_addafm_d [0]));
  
  /* mux (Ty Go,
     Ty Pointer_CTf''''''''''''_f''''''''''''_Int) : (call_f''''''''''''_f''''''''''''_Int_unlockFork6,Go) [(call_f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf''''''''''''_f''''''''''''_Intsc_0_1,Pointer_CTf''''''''''''_f''''''''''''_Int)] > (call_f''''''''''''_f''''''''''''_Int_goMux6,Pointer_CTf''''''''''''_f''''''''''''_Int) */
  assign \call_f''''''''''''_f''''''''''''_Int_goMux6_d  = {\call_f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf''''''''''''_f''''''''''''_Intsc_0_1_d [16:1],
                                                            (\call_f''''''''''''_f''''''''''''_Int_unlockFork6_d [0] && \call_f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf''''''''''''_f''''''''''''_Intsc_0_1_d [0])};
  assign \call_f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf''''''''''''_f''''''''''''_Intsc_0_1_r  = (\call_f''''''''''''_f''''''''''''_Int_goMux6_r  && (\call_f''''''''''''_f''''''''''''_Int_unlockFork6_d [0] && \call_f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf''''''''''''_f''''''''''''_Intsc_0_1_d [0]));
  assign \call_f''''''''''''_f''''''''''''_Int_unlockFork6_r  = (\call_f''''''''''''_f''''''''''''_Int_goMux6_r  && (\call_f''''''''''''_f''''''''''''_Int_unlockFork6_d [0] && \call_f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf''''''''''''_f''''''''''''_Intsc_0_1_d [0]));
  
  /* destruct (Ty TupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int,
          Dcon TupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int) : (call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_1,TupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int) > [(call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intgo_10,Go),
                                                                                                                                                                                                                                                                                                                                                                                                          (call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intm1aeq,Pointer_QTree_Int),
                                                                                                                                                                                                                                                                                                                                                                                                          (call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intm2aer,Pointer_QTree_Int),
                                                                                                                                                                                                                                                                                                                                                                                                          (call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intm3aes,Pointer_QTree_Int),
                                                                                                                                                                                                                                                                                                                                                                                                          (call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intis_zaet,MyDTInt_Bool),
                                                                                                                                                                                                                                                                                                                                                                                                          (call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intop_addaeu,MyDTInt_Int_Int),
                                                                                                                                                                                                                                                                                                                                                                                                          (call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intsc_0_2,Pointer_CTf_f_Int)] */
  logic [6:0] call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_1_emitted;
  logic [6:0] call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_1_done;
  assign call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intgo_10_d = (call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_1_d[0] && (! call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_1_emitted[0]));
  assign call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intm1aeq_d = {call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_1_d[16:1],
                                                                                                                                                      (call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_1_d[0] && (! call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_1_emitted[1]))};
  assign call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intm2aer_d = {call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_1_d[32:17],
                                                                                                                                                      (call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_1_d[0] && (! call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_1_emitted[2]))};
  assign call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intm3aes_d = {call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_1_d[48:33],
                                                                                                                                                      (call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_1_d[0] && (! call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_1_emitted[3]))};
  assign call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intis_zaet_d = (call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_1_d[0] && (! call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_1_emitted[4]));
  assign call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intop_addaeu_d = (call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_1_d[0] && (! call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_1_emitted[5]));
  assign call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intsc_0_2_d = {call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_1_d[64:49],
                                                                                                                                                       (call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_1_d[0] && (! call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_1_emitted[6]))};
  assign call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_1_done = (call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_1_emitted | ({call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intsc_0_2_d[0],
                                                                                                                                                                                                                                                                                                       call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intop_addaeu_d[0],
                                                                                                                                                                                                                                                                                                       call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intis_zaet_d[0],
                                                                                                                                                                                                                                                                                                       call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intm3aes_d[0],
                                                                                                                                                                                                                                                                                                       call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intm2aer_d[0],
                                                                                                                                                                                                                                                                                                       call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intm1aeq_d[0],
                                                                                                                                                                                                                                                                                                       call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intgo_10_d[0]} & {call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intsc_0_2_r,
                                                                                                                                                                                                                                                                                                                                                                                                                                                        call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intop_addaeu_r,
                                                                                                                                                                                                                                                                                                                                                                                                                                                        call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intis_zaet_r,
                                                                                                                                                                                                                                                                                                                                                                                                                                                        call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intm3aes_r,
                                                                                                                                                                                                                                                                                                                                                                                                                                                        call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intm2aer_r,
                                                                                                                                                                                                                                                                                                                                                                                                                                                        call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intm1aeq_r,
                                                                                                                                                                                                                                                                                                                                                                                                                                                        call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intgo_10_r}));
  assign call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_1_r = (& call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_1_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_1_emitted <= 7'd0;
    else
      call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_1_emitted <= (call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_1_r ? 7'd0 :
                                                                                                                                                       call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_1_done);
  
  /* rbuf (Ty Go) : (call_f_f_Int_goConst,Go) > (call_f_f_Int_initBufi,Go) */
  Go_t call_f_f_Int_goConst_buf;
  assign call_f_f_Int_goConst_r = (! call_f_f_Int_goConst_buf[0]);
  assign call_f_f_Int_initBufi_d = (call_f_f_Int_goConst_buf[0] ? call_f_f_Int_goConst_buf :
                                    call_f_f_Int_goConst_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_f_f_Int_goConst_buf <= 1'd0;
    else
      if ((call_f_f_Int_initBufi_r && call_f_f_Int_goConst_buf[0]))
        call_f_f_Int_goConst_buf <= 1'd0;
      else if (((! call_f_f_Int_initBufi_r) && (! call_f_f_Int_goConst_buf[0])))
        call_f_f_Int_goConst_buf <= call_f_f_Int_goConst_d;
  
  /* mergectrl (Ty C5,Ty Go) : [(call_f_f_Int_goMux1,Go),
                           (lizzieLet67_3Lcall_f_f_Int3_1_argbuf,Go),
                           (lizzieLet67_3Lcall_f_f_Int2_1_argbuf,Go),
                           (lizzieLet67_3Lcall_f_f_Int1_1_argbuf,Go),
                           (lizzieLet17_5QNode_Int_7QNode_Int_8QNode_Int_1_argbuf,Go)] > (go_10_goMux_choice,C5) (go_10_goMux_data,Go) */
  logic [4:0] call_f_f_Int_goMux1_select_d;
  assign call_f_f_Int_goMux1_select_d = ((| call_f_f_Int_goMux1_select_q) ? call_f_f_Int_goMux1_select_q :
                                         (call_f_f_Int_goMux1_d[0] ? 5'd1 :
                                          (lizzieLet67_3Lcall_f_f_Int3_1_argbuf_d[0] ? 5'd2 :
                                           (lizzieLet67_3Lcall_f_f_Int2_1_argbuf_d[0] ? 5'd4 :
                                            (lizzieLet67_3Lcall_f_f_Int1_1_argbuf_d[0] ? 5'd8 :
                                             (lizzieLet17_5QNode_Int_7QNode_Int_8QNode_Int_1_argbuf_d[0] ? 5'd16 :
                                              5'd0))))));
  logic [4:0] call_f_f_Int_goMux1_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_f_f_Int_goMux1_select_q <= 5'd0;
    else
      call_f_f_Int_goMux1_select_q <= (call_f_f_Int_goMux1_done ? 5'd0 :
                                       call_f_f_Int_goMux1_select_d);
  logic [1:0] call_f_f_Int_goMux1_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_f_f_Int_goMux1_emit_q <= 2'd0;
    else
      call_f_f_Int_goMux1_emit_q <= (call_f_f_Int_goMux1_done ? 2'd0 :
                                     call_f_f_Int_goMux1_emit_d);
  logic [1:0] call_f_f_Int_goMux1_emit_d;
  assign call_f_f_Int_goMux1_emit_d = (call_f_f_Int_goMux1_emit_q | ({go_10_goMux_choice_d[0],
                                                                      go_10_goMux_data_d[0]} & {go_10_goMux_choice_r,
                                                                                                go_10_goMux_data_r}));
  logic call_f_f_Int_goMux1_done;
  assign call_f_f_Int_goMux1_done = (& call_f_f_Int_goMux1_emit_d);
  assign {lizzieLet17_5QNode_Int_7QNode_Int_8QNode_Int_1_argbuf_r,
          lizzieLet67_3Lcall_f_f_Int1_1_argbuf_r,
          lizzieLet67_3Lcall_f_f_Int2_1_argbuf_r,
          lizzieLet67_3Lcall_f_f_Int3_1_argbuf_r,
          call_f_f_Int_goMux1_r} = (call_f_f_Int_goMux1_done ? call_f_f_Int_goMux1_select_d :
                                    5'd0);
  assign go_10_goMux_data_d = ((call_f_f_Int_goMux1_select_d[0] && (! call_f_f_Int_goMux1_emit_q[0])) ? call_f_f_Int_goMux1_d :
                               ((call_f_f_Int_goMux1_select_d[1] && (! call_f_f_Int_goMux1_emit_q[0])) ? lizzieLet67_3Lcall_f_f_Int3_1_argbuf_d :
                                ((call_f_f_Int_goMux1_select_d[2] && (! call_f_f_Int_goMux1_emit_q[0])) ? lizzieLet67_3Lcall_f_f_Int2_1_argbuf_d :
                                 ((call_f_f_Int_goMux1_select_d[3] && (! call_f_f_Int_goMux1_emit_q[0])) ? lizzieLet67_3Lcall_f_f_Int1_1_argbuf_d :
                                  ((call_f_f_Int_goMux1_select_d[4] && (! call_f_f_Int_goMux1_emit_q[0])) ? lizzieLet17_5QNode_Int_7QNode_Int_8QNode_Int_1_argbuf_d :
                                   1'd0)))));
  assign go_10_goMux_choice_d = ((call_f_f_Int_goMux1_select_d[0] && (! call_f_f_Int_goMux1_emit_q[1])) ? C1_5_dc(1'd1) :
                                 ((call_f_f_Int_goMux1_select_d[1] && (! call_f_f_Int_goMux1_emit_q[1])) ? C2_5_dc(1'd1) :
                                  ((call_f_f_Int_goMux1_select_d[2] && (! call_f_f_Int_goMux1_emit_q[1])) ? C3_5_dc(1'd1) :
                                   ((call_f_f_Int_goMux1_select_d[3] && (! call_f_f_Int_goMux1_emit_q[1])) ? C4_5_dc(1'd1) :
                                    ((call_f_f_Int_goMux1_select_d[4] && (! call_f_f_Int_goMux1_emit_q[1])) ? C5_5_dc(1'd1) :
                                     {3'd0, 1'd0})))));
  
  /* fork (Ty Go) : (call_f_f_Int_initBuf,Go) > [(call_f_f_Int_unlockFork1,Go),
                                            (call_f_f_Int_unlockFork2,Go),
                                            (call_f_f_Int_unlockFork3,Go),
                                            (call_f_f_Int_unlockFork4,Go),
                                            (call_f_f_Int_unlockFork5,Go),
                                            (call_f_f_Int_unlockFork6,Go),
                                            (call_f_f_Int_unlockFork7,Go)] */
  logic [6:0] call_f_f_Int_initBuf_emitted;
  logic [6:0] call_f_f_Int_initBuf_done;
  assign call_f_f_Int_unlockFork1_d = (call_f_f_Int_initBuf_d[0] && (! call_f_f_Int_initBuf_emitted[0]));
  assign call_f_f_Int_unlockFork2_d = (call_f_f_Int_initBuf_d[0] && (! call_f_f_Int_initBuf_emitted[1]));
  assign call_f_f_Int_unlockFork3_d = (call_f_f_Int_initBuf_d[0] && (! call_f_f_Int_initBuf_emitted[2]));
  assign call_f_f_Int_unlockFork4_d = (call_f_f_Int_initBuf_d[0] && (! call_f_f_Int_initBuf_emitted[3]));
  assign call_f_f_Int_unlockFork5_d = (call_f_f_Int_initBuf_d[0] && (! call_f_f_Int_initBuf_emitted[4]));
  assign call_f_f_Int_unlockFork6_d = (call_f_f_Int_initBuf_d[0] && (! call_f_f_Int_initBuf_emitted[5]));
  assign call_f_f_Int_unlockFork7_d = (call_f_f_Int_initBuf_d[0] && (! call_f_f_Int_initBuf_emitted[6]));
  assign call_f_f_Int_initBuf_done = (call_f_f_Int_initBuf_emitted | ({call_f_f_Int_unlockFork7_d[0],
                                                                       call_f_f_Int_unlockFork6_d[0],
                                                                       call_f_f_Int_unlockFork5_d[0],
                                                                       call_f_f_Int_unlockFork4_d[0],
                                                                       call_f_f_Int_unlockFork3_d[0],
                                                                       call_f_f_Int_unlockFork2_d[0],
                                                                       call_f_f_Int_unlockFork1_d[0]} & {call_f_f_Int_unlockFork7_r,
                                                                                                         call_f_f_Int_unlockFork6_r,
                                                                                                         call_f_f_Int_unlockFork5_r,
                                                                                                         call_f_f_Int_unlockFork4_r,
                                                                                                         call_f_f_Int_unlockFork3_r,
                                                                                                         call_f_f_Int_unlockFork2_r,
                                                                                                         call_f_f_Int_unlockFork1_r}));
  assign call_f_f_Int_initBuf_r = (& call_f_f_Int_initBuf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_f_f_Int_initBuf_emitted <= 7'd0;
    else
      call_f_f_Int_initBuf_emitted <= (call_f_f_Int_initBuf_r ? 7'd0 :
                                       call_f_f_Int_initBuf_done);
  
  /* initbuf (Ty Go,
         Dcon Go) : (call_f_f_Int_initBufi,Go) > (call_f_f_Int_initBuf,Go) */
  assign call_f_f_Int_initBufi_r = ((! call_f_f_Int_initBuf_d[0]) || call_f_f_Int_initBuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_f_f_Int_initBuf_d <= Go_dc(1'd1);
    else
      if (call_f_f_Int_initBufi_r)
        call_f_f_Int_initBuf_d <= call_f_f_Int_initBufi_d;
  
  /* mux (Ty Go,
     Ty Go) : (call_f_f_Int_unlockFork1,Go) [(call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intgo_10,Go)] > (call_f_f_Int_goMux1,Go) */
  assign call_f_f_Int_goMux1_d = (call_f_f_Int_unlockFork1_d[0] && call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intgo_10_d[0]);
  assign call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intgo_10_r = (call_f_f_Int_goMux1_r && (call_f_f_Int_unlockFork1_d[0] && call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intgo_10_d[0]));
  assign call_f_f_Int_unlockFork1_r = (call_f_f_Int_goMux1_r && (call_f_f_Int_unlockFork1_d[0] && call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intgo_10_d[0]));
  
  /* mux (Ty Go,
     Ty Pointer_QTree_Int) : (call_f_f_Int_unlockFork2,Go) [(call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intm1aeq,Pointer_QTree_Int)] > (call_f_f_Int_goMux2,Pointer_QTree_Int) */
  assign call_f_f_Int_goMux2_d = {call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intm1aeq_d[16:1],
                                  (call_f_f_Int_unlockFork2_d[0] && call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intm1aeq_d[0])};
  assign call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intm1aeq_r = (call_f_f_Int_goMux2_r && (call_f_f_Int_unlockFork2_d[0] && call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intm1aeq_d[0]));
  assign call_f_f_Int_unlockFork2_r = (call_f_f_Int_goMux2_r && (call_f_f_Int_unlockFork2_d[0] && call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intm1aeq_d[0]));
  
  /* mux (Ty Go,
     Ty Pointer_QTree_Int) : (call_f_f_Int_unlockFork3,Go) [(call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intm2aer,Pointer_QTree_Int)] > (call_f_f_Int_goMux3,Pointer_QTree_Int) */
  assign call_f_f_Int_goMux3_d = {call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intm2aer_d[16:1],
                                  (call_f_f_Int_unlockFork3_d[0] && call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intm2aer_d[0])};
  assign call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intm2aer_r = (call_f_f_Int_goMux3_r && (call_f_f_Int_unlockFork3_d[0] && call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intm2aer_d[0]));
  assign call_f_f_Int_unlockFork3_r = (call_f_f_Int_goMux3_r && (call_f_f_Int_unlockFork3_d[0] && call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intm2aer_d[0]));
  
  /* mux (Ty Go,
     Ty Pointer_QTree_Int) : (call_f_f_Int_unlockFork4,Go) [(call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intm3aes,Pointer_QTree_Int)] > (call_f_f_Int_goMux4,Pointer_QTree_Int) */
  assign call_f_f_Int_goMux4_d = {call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intm3aes_d[16:1],
                                  (call_f_f_Int_unlockFork4_d[0] && call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intm3aes_d[0])};
  assign call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intm3aes_r = (call_f_f_Int_goMux4_r && (call_f_f_Int_unlockFork4_d[0] && call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intm3aes_d[0]));
  assign call_f_f_Int_unlockFork4_r = (call_f_f_Int_goMux4_r && (call_f_f_Int_unlockFork4_d[0] && call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intm3aes_d[0]));
  
  /* mux (Ty Go,
     Ty MyDTInt_Bool) : (call_f_f_Int_unlockFork5,Go) [(call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intis_zaet,MyDTInt_Bool)] > (call_f_f_Int_goMux5,MyDTInt_Bool) */
  assign call_f_f_Int_goMux5_d = (call_f_f_Int_unlockFork5_d[0] && call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intis_zaet_d[0]);
  assign call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intis_zaet_r = (call_f_f_Int_goMux5_r && (call_f_f_Int_unlockFork5_d[0] && call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intis_zaet_d[0]));
  assign call_f_f_Int_unlockFork5_r = (call_f_f_Int_goMux5_r && (call_f_f_Int_unlockFork5_d[0] && call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intis_zaet_d[0]));
  
  /* mux (Ty Go,
     Ty MyDTInt_Int_Int) : (call_f_f_Int_unlockFork6,Go) [(call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intop_addaeu,MyDTInt_Int_Int)] > (call_f_f_Int_goMux6,MyDTInt_Int_Int) */
  assign call_f_f_Int_goMux6_d = (call_f_f_Int_unlockFork6_d[0] && call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intop_addaeu_d[0]);
  assign call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intop_addaeu_r = (call_f_f_Int_goMux6_r && (call_f_f_Int_unlockFork6_d[0] && call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intop_addaeu_d[0]));
  assign call_f_f_Int_unlockFork6_r = (call_f_f_Int_goMux6_r && (call_f_f_Int_unlockFork6_d[0] && call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intop_addaeu_d[0]));
  
  /* mux (Ty Go,
     Ty Pointer_CTf_f_Int) : (call_f_f_Int_unlockFork7,Go) [(call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intsc_0_2,Pointer_CTf_f_Int)] > (call_f_f_Int_goMux7,Pointer_CTf_f_Int) */
  assign call_f_f_Int_goMux7_d = {call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intsc_0_2_d[16:1],
                                  (call_f_f_Int_unlockFork7_d[0] && call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intsc_0_2_d[0])};
  assign call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intsc_0_2_r = (call_f_f_Int_goMux7_r && (call_f_f_Int_unlockFork7_d[0] && call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intsc_0_2_d[0]));
  assign call_f_f_Int_unlockFork7_r = (call_f_f_Int_goMux7_r && (call_f_f_Int_unlockFork7_d[0] && call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intsc_0_2_d[0]));
  
  /* demux (Ty MyBool,
       Ty Int) : (es_10_1,MyBool) (lizzieLet17_5QVal_Int_7QNone_Int_3QVal_Int_2,Int) > [(es_10_1MyFalse,Int),
                                                                                        (_255,Int)] */
  logic [1:0] lizzieLet17_5QVal_Int_7QNone_Int_3QVal_Int_2_onehotd;
  always_comb
    if ((es_10_1_d[0] && lizzieLet17_5QVal_Int_7QNone_Int_3QVal_Int_2_d[0]))
      unique case (es_10_1_d[1:1])
        1'd0: lizzieLet17_5QVal_Int_7QNone_Int_3QVal_Int_2_onehotd = 2'd1;
        1'd1: lizzieLet17_5QVal_Int_7QNone_Int_3QVal_Int_2_onehotd = 2'd2;
        default:
          lizzieLet17_5QVal_Int_7QNone_Int_3QVal_Int_2_onehotd = 2'd0;
      endcase
    else lizzieLet17_5QVal_Int_7QNone_Int_3QVal_Int_2_onehotd = 2'd0;
  assign es_10_1MyFalse_d = {lizzieLet17_5QVal_Int_7QNone_Int_3QVal_Int_2_d[32:1],
                             lizzieLet17_5QVal_Int_7QNone_Int_3QVal_Int_2_onehotd[0]};
  assign _255_d = {lizzieLet17_5QVal_Int_7QNone_Int_3QVal_Int_2_d[32:1],
                   lizzieLet17_5QVal_Int_7QNone_Int_3QVal_Int_2_onehotd[1]};
  assign lizzieLet17_5QVal_Int_7QNone_Int_3QVal_Int_2_r = (| (lizzieLet17_5QVal_Int_7QNone_Int_3QVal_Int_2_onehotd & {_255_r,
                                                                                                                      es_10_1MyFalse_r}));
  assign es_10_1_r = lizzieLet17_5QVal_Int_7QNone_Int_3QVal_Int_2_r;
  
  /* buf (Ty Int) : (es_10_1MyFalse,Int) > (es_10_1MyFalse_1_argbuf,Int) */
  Int_t es_10_1MyFalse_bufchan_d;
  logic es_10_1MyFalse_bufchan_r;
  assign es_10_1MyFalse_r = ((! es_10_1MyFalse_bufchan_d[0]) || es_10_1MyFalse_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_10_1MyFalse_bufchan_d <= {32'd0, 1'd0};
    else
      if (es_10_1MyFalse_r) es_10_1MyFalse_bufchan_d <= es_10_1MyFalse_d;
  Int_t es_10_1MyFalse_bufchan_buf;
  assign es_10_1MyFalse_bufchan_r = (! es_10_1MyFalse_bufchan_buf[0]);
  assign es_10_1MyFalse_1_argbuf_d = (es_10_1MyFalse_bufchan_buf[0] ? es_10_1MyFalse_bufchan_buf :
                                      es_10_1MyFalse_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_10_1MyFalse_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((es_10_1MyFalse_1_argbuf_r && es_10_1MyFalse_bufchan_buf[0]))
        es_10_1MyFalse_bufchan_buf <= {32'd0, 1'd0};
      else if (((! es_10_1MyFalse_1_argbuf_r) && (! es_10_1MyFalse_bufchan_buf[0])))
        es_10_1MyFalse_bufchan_buf <= es_10_1MyFalse_bufchan_d;
  
  /* demux (Ty MyBool,
       Ty MyDTInt_Int_Int) : (es_10_2,MyBool) (lizzieLet17_5QVal_Int_7QNone_Int_4QVal_Int_2,MyDTInt_Int_Int) > [(es_10_2MyFalse,MyDTInt_Int_Int),
                                                                                                                (_254,MyDTInt_Int_Int)] */
  logic [1:0] lizzieLet17_5QVal_Int_7QNone_Int_4QVal_Int_2_onehotd;
  always_comb
    if ((es_10_2_d[0] && lizzieLet17_5QVal_Int_7QNone_Int_4QVal_Int_2_d[0]))
      unique case (es_10_2_d[1:1])
        1'd0: lizzieLet17_5QVal_Int_7QNone_Int_4QVal_Int_2_onehotd = 2'd1;
        1'd1: lizzieLet17_5QVal_Int_7QNone_Int_4QVal_Int_2_onehotd = 2'd2;
        default:
          lizzieLet17_5QVal_Int_7QNone_Int_4QVal_Int_2_onehotd = 2'd0;
      endcase
    else lizzieLet17_5QVal_Int_7QNone_Int_4QVal_Int_2_onehotd = 2'd0;
  assign es_10_2MyFalse_d = lizzieLet17_5QVal_Int_7QNone_Int_4QVal_Int_2_onehotd[0];
  assign _254_d = lizzieLet17_5QVal_Int_7QNone_Int_4QVal_Int_2_onehotd[1];
  assign lizzieLet17_5QVal_Int_7QNone_Int_4QVal_Int_2_r = (| (lizzieLet17_5QVal_Int_7QNone_Int_4QVal_Int_2_onehotd & {_254_r,
                                                                                                                      es_10_2MyFalse_r}));
  assign es_10_2_r = lizzieLet17_5QVal_Int_7QNone_Int_4QVal_Int_2_r;
  
  /* buf (Ty MyDTInt_Int_Int) : (es_10_2MyFalse,MyDTInt_Int_Int) > (es_10_2MyFalse_1_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t es_10_2MyFalse_bufchan_d;
  logic es_10_2MyFalse_bufchan_r;
  assign es_10_2MyFalse_r = ((! es_10_2MyFalse_bufchan_d[0]) || es_10_2MyFalse_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_10_2MyFalse_bufchan_d <= 1'd0;
    else
      if (es_10_2MyFalse_r) es_10_2MyFalse_bufchan_d <= es_10_2MyFalse_d;
  MyDTInt_Int_Int_t es_10_2MyFalse_bufchan_buf;
  assign es_10_2MyFalse_bufchan_r = (! es_10_2MyFalse_bufchan_buf[0]);
  assign es_10_2MyFalse_1_argbuf_d = (es_10_2MyFalse_bufchan_buf[0] ? es_10_2MyFalse_bufchan_buf :
                                      es_10_2MyFalse_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_10_2MyFalse_bufchan_buf <= 1'd0;
    else
      if ((es_10_2MyFalse_1_argbuf_r && es_10_2MyFalse_bufchan_buf[0]))
        es_10_2MyFalse_bufchan_buf <= 1'd0;
      else if (((! es_10_2MyFalse_1_argbuf_r) && (! es_10_2MyFalse_bufchan_buf[0])))
        es_10_2MyFalse_bufchan_buf <= es_10_2MyFalse_bufchan_d;
  
  /* dcon (Ty TupMyDTInt_Int_Int___Int___Int,
      Dcon TupMyDTInt_Int_Int___Int___Int) : [(es_10_2MyFalse_1_argbuf,MyDTInt_Int_Int),
                                              (es_10_1MyFalse_1_argbuf,Int),
                                              (es_10_5MyFalse_1_argbuf,Int)] > (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int6,TupMyDTInt_Int_Int___Int___Int) */
  assign applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int6_d = TupMyDTInt_Int_Int___Int___Int_dc((& {es_10_2MyFalse_1_argbuf_d[0],
                                                                                                       es_10_1MyFalse_1_argbuf_d[0],
                                                                                                       es_10_5MyFalse_1_argbuf_d[0]}), es_10_2MyFalse_1_argbuf_d, es_10_1MyFalse_1_argbuf_d, es_10_5MyFalse_1_argbuf_d);
  assign {es_10_2MyFalse_1_argbuf_r,
          es_10_1MyFalse_1_argbuf_r,
          es_10_5MyFalse_1_argbuf_r} = {3 {(applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int6_r && applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int6_d[0])}};
  
  /* demux (Ty MyBool,
       Ty Pointer_CTf_f_Int) : (es_10_3,MyBool) (lizzieLet17_5QVal_Int_7QNone_Int_5QVal_Int,Pointer_CTf_f_Int) > [(es_10_3MyFalse,Pointer_CTf_f_Int),
                                                                                                                  (es_10_3MyTrue,Pointer_CTf_f_Int)] */
  logic [1:0] lizzieLet17_5QVal_Int_7QNone_Int_5QVal_Int_onehotd;
  always_comb
    if ((es_10_3_d[0] && lizzieLet17_5QVal_Int_7QNone_Int_5QVal_Int_d[0]))
      unique case (es_10_3_d[1:1])
        1'd0: lizzieLet17_5QVal_Int_7QNone_Int_5QVal_Int_onehotd = 2'd1;
        1'd1: lizzieLet17_5QVal_Int_7QNone_Int_5QVal_Int_onehotd = 2'd2;
        default: lizzieLet17_5QVal_Int_7QNone_Int_5QVal_Int_onehotd = 2'd0;
      endcase
    else lizzieLet17_5QVal_Int_7QNone_Int_5QVal_Int_onehotd = 2'd0;
  assign es_10_3MyFalse_d = {lizzieLet17_5QVal_Int_7QNone_Int_5QVal_Int_d[16:1],
                             lizzieLet17_5QVal_Int_7QNone_Int_5QVal_Int_onehotd[0]};
  assign es_10_3MyTrue_d = {lizzieLet17_5QVal_Int_7QNone_Int_5QVal_Int_d[16:1],
                            lizzieLet17_5QVal_Int_7QNone_Int_5QVal_Int_onehotd[1]};
  assign lizzieLet17_5QVal_Int_7QNone_Int_5QVal_Int_r = (| (lizzieLet17_5QVal_Int_7QNone_Int_5QVal_Int_onehotd & {es_10_3MyTrue_r,
                                                                                                                  es_10_3MyFalse_r}));
  assign es_10_3_r = lizzieLet17_5QVal_Int_7QNone_Int_5QVal_Int_r;
  
  /* buf (Ty Pointer_CTf_f_Int) : (es_10_3MyFalse,Pointer_CTf_f_Int) > (es_10_3MyFalse_1_argbuf,Pointer_CTf_f_Int) */
  Pointer_CTf_f_Int_t es_10_3MyFalse_bufchan_d;
  logic es_10_3MyFalse_bufchan_r;
  assign es_10_3MyFalse_r = ((! es_10_3MyFalse_bufchan_d[0]) || es_10_3MyFalse_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_10_3MyFalse_bufchan_d <= {16'd0, 1'd0};
    else
      if (es_10_3MyFalse_r) es_10_3MyFalse_bufchan_d <= es_10_3MyFalse_d;
  Pointer_CTf_f_Int_t es_10_3MyFalse_bufchan_buf;
  assign es_10_3MyFalse_bufchan_r = (! es_10_3MyFalse_bufchan_buf[0]);
  assign es_10_3MyFalse_1_argbuf_d = (es_10_3MyFalse_bufchan_buf[0] ? es_10_3MyFalse_bufchan_buf :
                                      es_10_3MyFalse_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_10_3MyFalse_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((es_10_3MyFalse_1_argbuf_r && es_10_3MyFalse_bufchan_buf[0]))
        es_10_3MyFalse_bufchan_buf <= {16'd0, 1'd0};
      else if (((! es_10_3MyFalse_1_argbuf_r) && (! es_10_3MyFalse_bufchan_buf[0])))
        es_10_3MyFalse_bufchan_buf <= es_10_3MyFalse_bufchan_d;
  
  /* buf (Ty Pointer_CTf_f_Int) : (es_10_3MyTrue,Pointer_CTf_f_Int) > (es_10_3MyTrue_1_argbuf,Pointer_CTf_f_Int) */
  Pointer_CTf_f_Int_t es_10_3MyTrue_bufchan_d;
  logic es_10_3MyTrue_bufchan_r;
  assign es_10_3MyTrue_r = ((! es_10_3MyTrue_bufchan_d[0]) || es_10_3MyTrue_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_10_3MyTrue_bufchan_d <= {16'd0, 1'd0};
    else
      if (es_10_3MyTrue_r) es_10_3MyTrue_bufchan_d <= es_10_3MyTrue_d;
  Pointer_CTf_f_Int_t es_10_3MyTrue_bufchan_buf;
  assign es_10_3MyTrue_bufchan_r = (! es_10_3MyTrue_bufchan_buf[0]);
  assign es_10_3MyTrue_1_argbuf_d = (es_10_3MyTrue_bufchan_buf[0] ? es_10_3MyTrue_bufchan_buf :
                                     es_10_3MyTrue_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_10_3MyTrue_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((es_10_3MyTrue_1_argbuf_r && es_10_3MyTrue_bufchan_buf[0]))
        es_10_3MyTrue_bufchan_buf <= {16'd0, 1'd0};
      else if (((! es_10_3MyTrue_1_argbuf_r) && (! es_10_3MyTrue_bufchan_buf[0])))
        es_10_3MyTrue_bufchan_buf <= es_10_3MyTrue_bufchan_d;
  
  /* demux (Ty MyBool,
       Ty Go) : (es_10_4,MyBool) (lizzieLet17_5QVal_Int_7QNone_Int_6QVal_Int_2,Go) > [(es_10_4MyFalse,Go),
                                                                                      (es_10_4MyTrue,Go)] */
  logic [1:0] lizzieLet17_5QVal_Int_7QNone_Int_6QVal_Int_2_onehotd;
  always_comb
    if ((es_10_4_d[0] && lizzieLet17_5QVal_Int_7QNone_Int_6QVal_Int_2_d[0]))
      unique case (es_10_4_d[1:1])
        1'd0: lizzieLet17_5QVal_Int_7QNone_Int_6QVal_Int_2_onehotd = 2'd1;
        1'd1: lizzieLet17_5QVal_Int_7QNone_Int_6QVal_Int_2_onehotd = 2'd2;
        default:
          lizzieLet17_5QVal_Int_7QNone_Int_6QVal_Int_2_onehotd = 2'd0;
      endcase
    else lizzieLet17_5QVal_Int_7QNone_Int_6QVal_Int_2_onehotd = 2'd0;
  assign es_10_4MyFalse_d = lizzieLet17_5QVal_Int_7QNone_Int_6QVal_Int_2_onehotd[0];
  assign es_10_4MyTrue_d = lizzieLet17_5QVal_Int_7QNone_Int_6QVal_Int_2_onehotd[1];
  assign lizzieLet17_5QVal_Int_7QNone_Int_6QVal_Int_2_r = (| (lizzieLet17_5QVal_Int_7QNone_Int_6QVal_Int_2_onehotd & {es_10_4MyTrue_r,
                                                                                                                      es_10_4MyFalse_r}));
  assign es_10_4_r = lizzieLet17_5QVal_Int_7QNone_Int_6QVal_Int_2_r;
  
  /* buf (Ty Go) : (es_10_4MyFalse,Go) > (es_10_4MyFalse_1_argbuf,Go) */
  Go_t es_10_4MyFalse_bufchan_d;
  logic es_10_4MyFalse_bufchan_r;
  assign es_10_4MyFalse_r = ((! es_10_4MyFalse_bufchan_d[0]) || es_10_4MyFalse_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_10_4MyFalse_bufchan_d <= 1'd0;
    else
      if (es_10_4MyFalse_r) es_10_4MyFalse_bufchan_d <= es_10_4MyFalse_d;
  Go_t es_10_4MyFalse_bufchan_buf;
  assign es_10_4MyFalse_bufchan_r = (! es_10_4MyFalse_bufchan_buf[0]);
  assign es_10_4MyFalse_1_argbuf_d = (es_10_4MyFalse_bufchan_buf[0] ? es_10_4MyFalse_bufchan_buf :
                                      es_10_4MyFalse_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_10_4MyFalse_bufchan_buf <= 1'd0;
    else
      if ((es_10_4MyFalse_1_argbuf_r && es_10_4MyFalse_bufchan_buf[0]))
        es_10_4MyFalse_bufchan_buf <= 1'd0;
      else if (((! es_10_4MyFalse_1_argbuf_r) && (! es_10_4MyFalse_bufchan_buf[0])))
        es_10_4MyFalse_bufchan_buf <= es_10_4MyFalse_bufchan_d;
  
  /* fork (Ty Go) : (es_10_4MyTrue,Go) > [(es_10_4MyTrue_1,Go),
                                     (es_10_4MyTrue_2,Go)] */
  logic [1:0] es_10_4MyTrue_emitted;
  logic [1:0] es_10_4MyTrue_done;
  assign es_10_4MyTrue_1_d = (es_10_4MyTrue_d[0] && (! es_10_4MyTrue_emitted[0]));
  assign es_10_4MyTrue_2_d = (es_10_4MyTrue_d[0] && (! es_10_4MyTrue_emitted[1]));
  assign es_10_4MyTrue_done = (es_10_4MyTrue_emitted | ({es_10_4MyTrue_2_d[0],
                                                         es_10_4MyTrue_1_d[0]} & {es_10_4MyTrue_2_r,
                                                                                  es_10_4MyTrue_1_r}));
  assign es_10_4MyTrue_r = (& es_10_4MyTrue_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_10_4MyTrue_emitted <= 2'd0;
    else
      es_10_4MyTrue_emitted <= (es_10_4MyTrue_r ? 2'd0 :
                                es_10_4MyTrue_done);
  
  /* dcon (Ty QTree_Int,
      Dcon QNone_Int) : [(es_10_4MyTrue_1,Go)] > (es_10_4MyTrue_1QNone_Int,QTree_Int) */
  assign es_10_4MyTrue_1QNone_Int_d = QNone_Int_dc((& {es_10_4MyTrue_1_d[0]}), es_10_4MyTrue_1_d);
  assign {es_10_4MyTrue_1_r} = {1 {(es_10_4MyTrue_1QNone_Int_r && es_10_4MyTrue_1QNone_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (es_10_4MyTrue_1QNone_Int,QTree_Int) > (lizzieLet32_1_argbuf,QTree_Int) */
  QTree_Int_t es_10_4MyTrue_1QNone_Int_bufchan_d;
  logic es_10_4MyTrue_1QNone_Int_bufchan_r;
  assign es_10_4MyTrue_1QNone_Int_r = ((! es_10_4MyTrue_1QNone_Int_bufchan_d[0]) || es_10_4MyTrue_1QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_10_4MyTrue_1QNone_Int_bufchan_d <= {66'd0, 1'd0};
    else
      if (es_10_4MyTrue_1QNone_Int_r)
        es_10_4MyTrue_1QNone_Int_bufchan_d <= es_10_4MyTrue_1QNone_Int_d;
  QTree_Int_t es_10_4MyTrue_1QNone_Int_bufchan_buf;
  assign es_10_4MyTrue_1QNone_Int_bufchan_r = (! es_10_4MyTrue_1QNone_Int_bufchan_buf[0]);
  assign lizzieLet32_1_argbuf_d = (es_10_4MyTrue_1QNone_Int_bufchan_buf[0] ? es_10_4MyTrue_1QNone_Int_bufchan_buf :
                                   es_10_4MyTrue_1QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_10_4MyTrue_1QNone_Int_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((lizzieLet32_1_argbuf_r && es_10_4MyTrue_1QNone_Int_bufchan_buf[0]))
        es_10_4MyTrue_1QNone_Int_bufchan_buf <= {66'd0, 1'd0};
      else if (((! lizzieLet32_1_argbuf_r) && (! es_10_4MyTrue_1QNone_Int_bufchan_buf[0])))
        es_10_4MyTrue_1QNone_Int_bufchan_buf <= es_10_4MyTrue_1QNone_Int_bufchan_d;
  
  /* buf (Ty Go) : (es_10_4MyTrue_2,Go) > (es_10_4MyTrue_2_argbuf,Go) */
  Go_t es_10_4MyTrue_2_bufchan_d;
  logic es_10_4MyTrue_2_bufchan_r;
  assign es_10_4MyTrue_2_r = ((! es_10_4MyTrue_2_bufchan_d[0]) || es_10_4MyTrue_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_10_4MyTrue_2_bufchan_d <= 1'd0;
    else
      if (es_10_4MyTrue_2_r)
        es_10_4MyTrue_2_bufchan_d <= es_10_4MyTrue_2_d;
  Go_t es_10_4MyTrue_2_bufchan_buf;
  assign es_10_4MyTrue_2_bufchan_r = (! es_10_4MyTrue_2_bufchan_buf[0]);
  assign es_10_4MyTrue_2_argbuf_d = (es_10_4MyTrue_2_bufchan_buf[0] ? es_10_4MyTrue_2_bufchan_buf :
                                     es_10_4MyTrue_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_10_4MyTrue_2_bufchan_buf <= 1'd0;
    else
      if ((es_10_4MyTrue_2_argbuf_r && es_10_4MyTrue_2_bufchan_buf[0]))
        es_10_4MyTrue_2_bufchan_buf <= 1'd0;
      else if (((! es_10_4MyTrue_2_argbuf_r) && (! es_10_4MyTrue_2_bufchan_buf[0])))
        es_10_4MyTrue_2_bufchan_buf <= es_10_4MyTrue_2_bufchan_d;
  
  /* demux (Ty MyBool,
       Ty Int) : (es_10_5,MyBool) (vaeL_2,Int) > [(es_10_5MyFalse,Int),
                                                  (_253,Int)] */
  logic [1:0] vaeL_2_onehotd;
  always_comb
    if ((es_10_5_d[0] && vaeL_2_d[0]))
      unique case (es_10_5_d[1:1])
        1'd0: vaeL_2_onehotd = 2'd1;
        1'd1: vaeL_2_onehotd = 2'd2;
        default: vaeL_2_onehotd = 2'd0;
      endcase
    else vaeL_2_onehotd = 2'd0;
  assign es_10_5MyFalse_d = {vaeL_2_d[32:1], vaeL_2_onehotd[0]};
  assign _253_d = {vaeL_2_d[32:1], vaeL_2_onehotd[1]};
  assign vaeL_2_r = (| (vaeL_2_onehotd & {_253_r,
                                          es_10_5MyFalse_r}));
  assign es_10_5_r = vaeL_2_r;
  
  /* buf (Ty Int) : (es_10_5MyFalse,Int) > (es_10_5MyFalse_1_argbuf,Int) */
  Int_t es_10_5MyFalse_bufchan_d;
  logic es_10_5MyFalse_bufchan_r;
  assign es_10_5MyFalse_r = ((! es_10_5MyFalse_bufchan_d[0]) || es_10_5MyFalse_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_10_5MyFalse_bufchan_d <= {32'd0, 1'd0};
    else
      if (es_10_5MyFalse_r) es_10_5MyFalse_bufchan_d <= es_10_5MyFalse_d;
  Int_t es_10_5MyFalse_bufchan_buf;
  assign es_10_5MyFalse_bufchan_r = (! es_10_5MyFalse_bufchan_buf[0]);
  assign es_10_5MyFalse_1_argbuf_d = (es_10_5MyFalse_bufchan_buf[0] ? es_10_5MyFalse_bufchan_buf :
                                      es_10_5MyFalse_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_10_5MyFalse_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((es_10_5MyFalse_1_argbuf_r && es_10_5MyFalse_bufchan_buf[0]))
        es_10_5MyFalse_bufchan_buf <= {32'd0, 1'd0};
      else if (((! es_10_5MyFalse_1_argbuf_r) && (! es_10_5MyFalse_bufchan_buf[0])))
        es_10_5MyFalse_bufchan_buf <= es_10_5MyFalse_bufchan_d;
  
  /* buf (Ty QTree_Int) : (es_11_1QVal_Int,QTree_Int) > (lizzieLet31_1_argbuf,QTree_Int) */
  QTree_Int_t es_11_1QVal_Int_bufchan_d;
  logic es_11_1QVal_Int_bufchan_r;
  assign es_11_1QVal_Int_r = ((! es_11_1QVal_Int_bufchan_d[0]) || es_11_1QVal_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_11_1QVal_Int_bufchan_d <= {66'd0, 1'd0};
    else
      if (es_11_1QVal_Int_r)
        es_11_1QVal_Int_bufchan_d <= es_11_1QVal_Int_d;
  QTree_Int_t es_11_1QVal_Int_bufchan_buf;
  assign es_11_1QVal_Int_bufchan_r = (! es_11_1QVal_Int_bufchan_buf[0]);
  assign lizzieLet31_1_argbuf_d = (es_11_1QVal_Int_bufchan_buf[0] ? es_11_1QVal_Int_bufchan_buf :
                                   es_11_1QVal_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_11_1QVal_Int_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((lizzieLet31_1_argbuf_r && es_11_1QVal_Int_bufchan_buf[0]))
        es_11_1QVal_Int_bufchan_buf <= {66'd0, 1'd0};
      else if (((! lizzieLet31_1_argbuf_r) && (! es_11_1QVal_Int_bufchan_buf[0])))
        es_11_1QVal_Int_bufchan_buf <= es_11_1QVal_Int_bufchan_d;
  
  /* demux (Ty MyBool,
       Ty Int) : (es_14_1,MyBool) (lizzieLet17_5QVal_Int_10QVal_Int_2,Int) > [(es_14_1MyFalse,Int),
                                                                              (_252,Int)] */
  logic [1:0] lizzieLet17_5QVal_Int_10QVal_Int_2_onehotd;
  always_comb
    if ((es_14_1_d[0] && lizzieLet17_5QVal_Int_10QVal_Int_2_d[0]))
      unique case (es_14_1_d[1:1])
        1'd0: lizzieLet17_5QVal_Int_10QVal_Int_2_onehotd = 2'd1;
        1'd1: lizzieLet17_5QVal_Int_10QVal_Int_2_onehotd = 2'd2;
        default: lizzieLet17_5QVal_Int_10QVal_Int_2_onehotd = 2'd0;
      endcase
    else lizzieLet17_5QVal_Int_10QVal_Int_2_onehotd = 2'd0;
  assign es_14_1MyFalse_d = {lizzieLet17_5QVal_Int_10QVal_Int_2_d[32:1],
                             lizzieLet17_5QVal_Int_10QVal_Int_2_onehotd[0]};
  assign _252_d = {lizzieLet17_5QVal_Int_10QVal_Int_2_d[32:1],
                   lizzieLet17_5QVal_Int_10QVal_Int_2_onehotd[1]};
  assign lizzieLet17_5QVal_Int_10QVal_Int_2_r = (| (lizzieLet17_5QVal_Int_10QVal_Int_2_onehotd & {_252_r,
                                                                                                  es_14_1MyFalse_r}));
  assign es_14_1_r = lizzieLet17_5QVal_Int_10QVal_Int_2_r;
  
  /* demux (Ty MyBool,
       Ty MyDTInt_Int_Int) : (es_14_2,MyBool) (lizzieLet17_5QVal_Int_3QVal_Int_2,MyDTInt_Int_Int) > [(es_14_2MyFalse,MyDTInt_Int_Int),
                                                                                                     (_251,MyDTInt_Int_Int)] */
  logic [1:0] lizzieLet17_5QVal_Int_3QVal_Int_2_onehotd;
  always_comb
    if ((es_14_2_d[0] && lizzieLet17_5QVal_Int_3QVal_Int_2_d[0]))
      unique case (es_14_2_d[1:1])
        1'd0: lizzieLet17_5QVal_Int_3QVal_Int_2_onehotd = 2'd1;
        1'd1: lizzieLet17_5QVal_Int_3QVal_Int_2_onehotd = 2'd2;
        default: lizzieLet17_5QVal_Int_3QVal_Int_2_onehotd = 2'd0;
      endcase
    else lizzieLet17_5QVal_Int_3QVal_Int_2_onehotd = 2'd0;
  assign es_14_2MyFalse_d = lizzieLet17_5QVal_Int_3QVal_Int_2_onehotd[0];
  assign _251_d = lizzieLet17_5QVal_Int_3QVal_Int_2_onehotd[1];
  assign lizzieLet17_5QVal_Int_3QVal_Int_2_r = (| (lizzieLet17_5QVal_Int_3QVal_Int_2_onehotd & {_251_r,
                                                                                                es_14_2MyFalse_r}));
  assign es_14_2_r = lizzieLet17_5QVal_Int_3QVal_Int_2_r;
  
  /* demux (Ty MyBool,
       Ty Pointer_CTf_f_Int) : (es_14_3,MyBool) (lizzieLet17_5QVal_Int_4QVal_Int,Pointer_CTf_f_Int) > [(es_14_3MyFalse,Pointer_CTf_f_Int),
                                                                                                       (es_14_3MyTrue,Pointer_CTf_f_Int)] */
  logic [1:0] lizzieLet17_5QVal_Int_4QVal_Int_onehotd;
  always_comb
    if ((es_14_3_d[0] && lizzieLet17_5QVal_Int_4QVal_Int_d[0]))
      unique case (es_14_3_d[1:1])
        1'd0: lizzieLet17_5QVal_Int_4QVal_Int_onehotd = 2'd1;
        1'd1: lizzieLet17_5QVal_Int_4QVal_Int_onehotd = 2'd2;
        default: lizzieLet17_5QVal_Int_4QVal_Int_onehotd = 2'd0;
      endcase
    else lizzieLet17_5QVal_Int_4QVal_Int_onehotd = 2'd0;
  assign es_14_3MyFalse_d = {lizzieLet17_5QVal_Int_4QVal_Int_d[16:1],
                             lizzieLet17_5QVal_Int_4QVal_Int_onehotd[0]};
  assign es_14_3MyTrue_d = {lizzieLet17_5QVal_Int_4QVal_Int_d[16:1],
                            lizzieLet17_5QVal_Int_4QVal_Int_onehotd[1]};
  assign lizzieLet17_5QVal_Int_4QVal_Int_r = (| (lizzieLet17_5QVal_Int_4QVal_Int_onehotd & {es_14_3MyTrue_r,
                                                                                            es_14_3MyFalse_r}));
  assign es_14_3_r = lizzieLet17_5QVal_Int_4QVal_Int_r;
  
  /* buf (Ty Pointer_CTf_f_Int) : (es_14_3MyTrue,Pointer_CTf_f_Int) > (es_14_3MyTrue_1_argbuf,Pointer_CTf_f_Int) */
  Pointer_CTf_f_Int_t es_14_3MyTrue_bufchan_d;
  logic es_14_3MyTrue_bufchan_r;
  assign es_14_3MyTrue_r = ((! es_14_3MyTrue_bufchan_d[0]) || es_14_3MyTrue_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_14_3MyTrue_bufchan_d <= {16'd0, 1'd0};
    else
      if (es_14_3MyTrue_r) es_14_3MyTrue_bufchan_d <= es_14_3MyTrue_d;
  Pointer_CTf_f_Int_t es_14_3MyTrue_bufchan_buf;
  assign es_14_3MyTrue_bufchan_r = (! es_14_3MyTrue_bufchan_buf[0]);
  assign es_14_3MyTrue_1_argbuf_d = (es_14_3MyTrue_bufchan_buf[0] ? es_14_3MyTrue_bufchan_buf :
                                     es_14_3MyTrue_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_14_3MyTrue_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((es_14_3MyTrue_1_argbuf_r && es_14_3MyTrue_bufchan_buf[0]))
        es_14_3MyTrue_bufchan_buf <= {16'd0, 1'd0};
      else if (((! es_14_3MyTrue_1_argbuf_r) && (! es_14_3MyTrue_bufchan_buf[0])))
        es_14_3MyTrue_bufchan_buf <= es_14_3MyTrue_bufchan_d;
  
  /* demux (Ty MyBool,
       Ty Go) : (es_14_4,MyBool) (lizzieLet17_5QVal_Int_5QVal_Int_2,Go) > [(es_14_4MyFalse,Go),
                                                                           (es_14_4MyTrue,Go)] */
  logic [1:0] lizzieLet17_5QVal_Int_5QVal_Int_2_onehotd;
  always_comb
    if ((es_14_4_d[0] && lizzieLet17_5QVal_Int_5QVal_Int_2_d[0]))
      unique case (es_14_4_d[1:1])
        1'd0: lizzieLet17_5QVal_Int_5QVal_Int_2_onehotd = 2'd1;
        1'd1: lizzieLet17_5QVal_Int_5QVal_Int_2_onehotd = 2'd2;
        default: lizzieLet17_5QVal_Int_5QVal_Int_2_onehotd = 2'd0;
      endcase
    else lizzieLet17_5QVal_Int_5QVal_Int_2_onehotd = 2'd0;
  assign es_14_4MyFalse_d = lizzieLet17_5QVal_Int_5QVal_Int_2_onehotd[0];
  assign es_14_4MyTrue_d = lizzieLet17_5QVal_Int_5QVal_Int_2_onehotd[1];
  assign lizzieLet17_5QVal_Int_5QVal_Int_2_r = (| (lizzieLet17_5QVal_Int_5QVal_Int_2_onehotd & {es_14_4MyTrue_r,
                                                                                                es_14_4MyFalse_r}));
  assign es_14_4_r = lizzieLet17_5QVal_Int_5QVal_Int_2_r;
  
  /* buf (Ty Go) : (es_14_4MyTrue,Go) > (es_14_4MyTrue_1_argbuf,Go) */
  Go_t es_14_4MyTrue_bufchan_d;
  logic es_14_4MyTrue_bufchan_r;
  assign es_14_4MyTrue_r = ((! es_14_4MyTrue_bufchan_d[0]) || es_14_4MyTrue_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_14_4MyTrue_bufchan_d <= 1'd0;
    else
      if (es_14_4MyTrue_r) es_14_4MyTrue_bufchan_d <= es_14_4MyTrue_d;
  Go_t es_14_4MyTrue_bufchan_buf;
  assign es_14_4MyTrue_bufchan_r = (! es_14_4MyTrue_bufchan_buf[0]);
  assign es_14_4MyTrue_1_argbuf_d = (es_14_4MyTrue_bufchan_buf[0] ? es_14_4MyTrue_bufchan_buf :
                                     es_14_4MyTrue_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_14_4MyTrue_bufchan_buf <= 1'd0;
    else
      if ((es_14_4MyTrue_1_argbuf_r && es_14_4MyTrue_bufchan_buf[0]))
        es_14_4MyTrue_bufchan_buf <= 1'd0;
      else if (((! es_14_4MyTrue_1_argbuf_r) && (! es_14_4MyTrue_bufchan_buf[0])))
        es_14_4MyTrue_bufchan_buf <= es_14_4MyTrue_bufchan_d;
  
  /* demux (Ty MyBool,
       Ty MyDTInt_Bool) : (es_14_5,MyBool) (lizzieLet17_5QVal_Int_6QVal_Int_2,MyDTInt_Bool) > [(es_14_5MyFalse,MyDTInt_Bool),
                                                                                               (_250,MyDTInt_Bool)] */
  logic [1:0] lizzieLet17_5QVal_Int_6QVal_Int_2_onehotd;
  always_comb
    if ((es_14_5_d[0] && lizzieLet17_5QVal_Int_6QVal_Int_2_d[0]))
      unique case (es_14_5_d[1:1])
        1'd0: lizzieLet17_5QVal_Int_6QVal_Int_2_onehotd = 2'd1;
        1'd1: lizzieLet17_5QVal_Int_6QVal_Int_2_onehotd = 2'd2;
        default: lizzieLet17_5QVal_Int_6QVal_Int_2_onehotd = 2'd0;
      endcase
    else lizzieLet17_5QVal_Int_6QVal_Int_2_onehotd = 2'd0;
  assign es_14_5MyFalse_d = lizzieLet17_5QVal_Int_6QVal_Int_2_onehotd[0];
  assign _250_d = lizzieLet17_5QVal_Int_6QVal_Int_2_onehotd[1];
  assign lizzieLet17_5QVal_Int_6QVal_Int_2_r = (| (lizzieLet17_5QVal_Int_6QVal_Int_2_onehotd & {_250_r,
                                                                                                es_14_5MyFalse_r}));
  assign es_14_5_r = lizzieLet17_5QVal_Int_6QVal_Int_2_r;
  
  /* demux (Ty MyBool,
       Ty QTree_Int) : (es_14_6,MyBool) (lizzieLet17_5QVal_Int_7QVal_Int,QTree_Int) > [(es_14_6MyFalse,QTree_Int),
                                                                                       (_249,QTree_Int)] */
  logic [1:0] lizzieLet17_5QVal_Int_7QVal_Int_onehotd;
  always_comb
    if ((es_14_6_d[0] && lizzieLet17_5QVal_Int_7QVal_Int_d[0]))
      unique case (es_14_6_d[1:1])
        1'd0: lizzieLet17_5QVal_Int_7QVal_Int_onehotd = 2'd1;
        1'd1: lizzieLet17_5QVal_Int_7QVal_Int_onehotd = 2'd2;
        default: lizzieLet17_5QVal_Int_7QVal_Int_onehotd = 2'd0;
      endcase
    else lizzieLet17_5QVal_Int_7QVal_Int_onehotd = 2'd0;
  assign es_14_6MyFalse_d = {lizzieLet17_5QVal_Int_7QVal_Int_d[66:1],
                             lizzieLet17_5QVal_Int_7QVal_Int_onehotd[0]};
  assign _249_d = {lizzieLet17_5QVal_Int_7QVal_Int_d[66:1],
                   lizzieLet17_5QVal_Int_7QVal_Int_onehotd[1]};
  assign lizzieLet17_5QVal_Int_7QVal_Int_r = (| (lizzieLet17_5QVal_Int_7QVal_Int_onehotd & {_249_r,
                                                                                            es_14_6MyFalse_r}));
  assign es_14_6_r = lizzieLet17_5QVal_Int_7QVal_Int_r;
  
  /* fork (Ty QTree_Int) : (es_14_6MyFalse,QTree_Int) > [(es_14_6MyFalse_1,QTree_Int),
                                                    (es_14_6MyFalse_2,QTree_Int),
                                                    (es_14_6MyFalse_3,QTree_Int),
                                                    (es_14_6MyFalse_4,QTree_Int),
                                                    (es_14_6MyFalse_5,QTree_Int),
                                                    (es_14_6MyFalse_6,QTree_Int),
                                                    (es_14_6MyFalse_7,QTree_Int),
                                                    (es_14_6MyFalse_8,QTree_Int)] */
  logic [7:0] es_14_6MyFalse_emitted;
  logic [7:0] es_14_6MyFalse_done;
  assign es_14_6MyFalse_1_d = {es_14_6MyFalse_d[66:1],
                               (es_14_6MyFalse_d[0] && (! es_14_6MyFalse_emitted[0]))};
  assign es_14_6MyFalse_2_d = {es_14_6MyFalse_d[66:1],
                               (es_14_6MyFalse_d[0] && (! es_14_6MyFalse_emitted[1]))};
  assign es_14_6MyFalse_3_d = {es_14_6MyFalse_d[66:1],
                               (es_14_6MyFalse_d[0] && (! es_14_6MyFalse_emitted[2]))};
  assign es_14_6MyFalse_4_d = {es_14_6MyFalse_d[66:1],
                               (es_14_6MyFalse_d[0] && (! es_14_6MyFalse_emitted[3]))};
  assign es_14_6MyFalse_5_d = {es_14_6MyFalse_d[66:1],
                               (es_14_6MyFalse_d[0] && (! es_14_6MyFalse_emitted[4]))};
  assign es_14_6MyFalse_6_d = {es_14_6MyFalse_d[66:1],
                               (es_14_6MyFalse_d[0] && (! es_14_6MyFalse_emitted[5]))};
  assign es_14_6MyFalse_7_d = {es_14_6MyFalse_d[66:1],
                               (es_14_6MyFalse_d[0] && (! es_14_6MyFalse_emitted[6]))};
  assign es_14_6MyFalse_8_d = {es_14_6MyFalse_d[66:1],
                               (es_14_6MyFalse_d[0] && (! es_14_6MyFalse_emitted[7]))};
  assign es_14_6MyFalse_done = (es_14_6MyFalse_emitted | ({es_14_6MyFalse_8_d[0],
                                                           es_14_6MyFalse_7_d[0],
                                                           es_14_6MyFalse_6_d[0],
                                                           es_14_6MyFalse_5_d[0],
                                                           es_14_6MyFalse_4_d[0],
                                                           es_14_6MyFalse_3_d[0],
                                                           es_14_6MyFalse_2_d[0],
                                                           es_14_6MyFalse_1_d[0]} & {es_14_6MyFalse_8_r,
                                                                                     es_14_6MyFalse_7_r,
                                                                                     es_14_6MyFalse_6_r,
                                                                                     es_14_6MyFalse_5_r,
                                                                                     es_14_6MyFalse_4_r,
                                                                                     es_14_6MyFalse_3_r,
                                                                                     es_14_6MyFalse_2_r,
                                                                                     es_14_6MyFalse_1_r}));
  assign es_14_6MyFalse_r = (& es_14_6MyFalse_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_14_6MyFalse_emitted <= 8'd0;
    else
      es_14_6MyFalse_emitted <= (es_14_6MyFalse_r ? 8'd0 :
                                 es_14_6MyFalse_done);
  
  /* destruct (Ty QTree_Int,
          Dcon QVal_Int) : (es_14_6MyFalse_1QVal_Int,QTree_Int) > [(v'aeR_destruct,Int)] */
  assign \v'aeR_destruct_d  = {es_14_6MyFalse_1QVal_Int_d[34:3],
                               es_14_6MyFalse_1QVal_Int_d[0]};
  assign es_14_6MyFalse_1QVal_Int_r = \v'aeR_destruct_r ;
  
  /* demux (Ty QTree_Int,
       Ty QTree_Int) : (es_14_6MyFalse_2,QTree_Int) (es_14_6MyFalse_1,QTree_Int) > [(_248,QTree_Int),
                                                                                    (es_14_6MyFalse_1QVal_Int,QTree_Int),
                                                                                    (_247,QTree_Int),
                                                                                    (_246,QTree_Int)] */
  logic [3:0] es_14_6MyFalse_1_onehotd;
  always_comb
    if ((es_14_6MyFalse_2_d[0] && es_14_6MyFalse_1_d[0]))
      unique case (es_14_6MyFalse_2_d[2:1])
        2'd0: es_14_6MyFalse_1_onehotd = 4'd1;
        2'd1: es_14_6MyFalse_1_onehotd = 4'd2;
        2'd2: es_14_6MyFalse_1_onehotd = 4'd4;
        2'd3: es_14_6MyFalse_1_onehotd = 4'd8;
        default: es_14_6MyFalse_1_onehotd = 4'd0;
      endcase
    else es_14_6MyFalse_1_onehotd = 4'd0;
  assign _248_d = {es_14_6MyFalse_1_d[66:1],
                   es_14_6MyFalse_1_onehotd[0]};
  assign es_14_6MyFalse_1QVal_Int_d = {es_14_6MyFalse_1_d[66:1],
                                       es_14_6MyFalse_1_onehotd[1]};
  assign _247_d = {es_14_6MyFalse_1_d[66:1],
                   es_14_6MyFalse_1_onehotd[2]};
  assign _246_d = {es_14_6MyFalse_1_d[66:1],
                   es_14_6MyFalse_1_onehotd[3]};
  assign es_14_6MyFalse_1_r = (| (es_14_6MyFalse_1_onehotd & {_246_r,
                                                              _247_r,
                                                              es_14_6MyFalse_1QVal_Int_r,
                                                              _248_r}));
  assign es_14_6MyFalse_2_r = es_14_6MyFalse_1_r;
  
  /* demux (Ty QTree_Int,
       Ty Int) : (es_14_6MyFalse_3,QTree_Int) (es_14_1MyFalse,Int) > [(es_14_6MyFalse_3QNone_Int,Int),
                                                                      (es_14_6MyFalse_3QVal_Int,Int),
                                                                      (_245,Int),
                                                                      (_244,Int)] */
  logic [3:0] es_14_1MyFalse_onehotd;
  always_comb
    if ((es_14_6MyFalse_3_d[0] && es_14_1MyFalse_d[0]))
      unique case (es_14_6MyFalse_3_d[2:1])
        2'd0: es_14_1MyFalse_onehotd = 4'd1;
        2'd1: es_14_1MyFalse_onehotd = 4'd2;
        2'd2: es_14_1MyFalse_onehotd = 4'd4;
        2'd3: es_14_1MyFalse_onehotd = 4'd8;
        default: es_14_1MyFalse_onehotd = 4'd0;
      endcase
    else es_14_1MyFalse_onehotd = 4'd0;
  assign es_14_6MyFalse_3QNone_Int_d = {es_14_1MyFalse_d[32:1],
                                        es_14_1MyFalse_onehotd[0]};
  assign es_14_6MyFalse_3QVal_Int_d = {es_14_1MyFalse_d[32:1],
                                       es_14_1MyFalse_onehotd[1]};
  assign _245_d = {es_14_1MyFalse_d[32:1],
                   es_14_1MyFalse_onehotd[2]};
  assign _244_d = {es_14_1MyFalse_d[32:1],
                   es_14_1MyFalse_onehotd[3]};
  assign es_14_1MyFalse_r = (| (es_14_1MyFalse_onehotd & {_244_r,
                                                          _245_r,
                                                          es_14_6MyFalse_3QVal_Int_r,
                                                          es_14_6MyFalse_3QNone_Int_r}));
  assign es_14_6MyFalse_3_r = es_14_1MyFalse_r;
  
  /* buf (Ty Int) : (es_14_6MyFalse_3QNone_Int,Int) > (es_14_6MyFalse_3QNone_Int_1_argbuf,Int) */
  Int_t es_14_6MyFalse_3QNone_Int_bufchan_d;
  logic es_14_6MyFalse_3QNone_Int_bufchan_r;
  assign es_14_6MyFalse_3QNone_Int_r = ((! es_14_6MyFalse_3QNone_Int_bufchan_d[0]) || es_14_6MyFalse_3QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_14_6MyFalse_3QNone_Int_bufchan_d <= {32'd0, 1'd0};
    else
      if (es_14_6MyFalse_3QNone_Int_r)
        es_14_6MyFalse_3QNone_Int_bufchan_d <= es_14_6MyFalse_3QNone_Int_d;
  Int_t es_14_6MyFalse_3QNone_Int_bufchan_buf;
  assign es_14_6MyFalse_3QNone_Int_bufchan_r = (! es_14_6MyFalse_3QNone_Int_bufchan_buf[0]);
  assign es_14_6MyFalse_3QNone_Int_1_argbuf_d = (es_14_6MyFalse_3QNone_Int_bufchan_buf[0] ? es_14_6MyFalse_3QNone_Int_bufchan_buf :
                                                 es_14_6MyFalse_3QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_14_6MyFalse_3QNone_Int_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((es_14_6MyFalse_3QNone_Int_1_argbuf_r && es_14_6MyFalse_3QNone_Int_bufchan_buf[0]))
        es_14_6MyFalse_3QNone_Int_bufchan_buf <= {32'd0, 1'd0};
      else if (((! es_14_6MyFalse_3QNone_Int_1_argbuf_r) && (! es_14_6MyFalse_3QNone_Int_bufchan_buf[0])))
        es_14_6MyFalse_3QNone_Int_bufchan_buf <= es_14_6MyFalse_3QNone_Int_bufchan_d;
  
  /* fork (Ty Int) : (es_14_6MyFalse_3QVal_Int,Int) > [(es_14_6MyFalse_3QVal_Int_1,Int),
                                                  (es_14_6MyFalse_3QVal_Int_2,Int)] */
  logic [1:0] es_14_6MyFalse_3QVal_Int_emitted;
  logic [1:0] es_14_6MyFalse_3QVal_Int_done;
  assign es_14_6MyFalse_3QVal_Int_1_d = {es_14_6MyFalse_3QVal_Int_d[32:1],
                                         (es_14_6MyFalse_3QVal_Int_d[0] && (! es_14_6MyFalse_3QVal_Int_emitted[0]))};
  assign es_14_6MyFalse_3QVal_Int_2_d = {es_14_6MyFalse_3QVal_Int_d[32:1],
                                         (es_14_6MyFalse_3QVal_Int_d[0] && (! es_14_6MyFalse_3QVal_Int_emitted[1]))};
  assign es_14_6MyFalse_3QVal_Int_done = (es_14_6MyFalse_3QVal_Int_emitted | ({es_14_6MyFalse_3QVal_Int_2_d[0],
                                                                               es_14_6MyFalse_3QVal_Int_1_d[0]} & {es_14_6MyFalse_3QVal_Int_2_r,
                                                                                                                   es_14_6MyFalse_3QVal_Int_1_r}));
  assign es_14_6MyFalse_3QVal_Int_r = (& es_14_6MyFalse_3QVal_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_14_6MyFalse_3QVal_Int_emitted <= 2'd0;
    else
      es_14_6MyFalse_3QVal_Int_emitted <= (es_14_6MyFalse_3QVal_Int_r ? 2'd0 :
                                           es_14_6MyFalse_3QVal_Int_done);
  
  /* buf (Ty Int) : (es_14_6MyFalse_3QVal_Int_1,Int) > (es_14_6MyFalse_3QVal_Int_1_argbuf,Int) */
  Int_t es_14_6MyFalse_3QVal_Int_1_bufchan_d;
  logic es_14_6MyFalse_3QVal_Int_1_bufchan_r;
  assign es_14_6MyFalse_3QVal_Int_1_r = ((! es_14_6MyFalse_3QVal_Int_1_bufchan_d[0]) || es_14_6MyFalse_3QVal_Int_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_14_6MyFalse_3QVal_Int_1_bufchan_d <= {32'd0, 1'd0};
    else
      if (es_14_6MyFalse_3QVal_Int_1_r)
        es_14_6MyFalse_3QVal_Int_1_bufchan_d <= es_14_6MyFalse_3QVal_Int_1_d;
  Int_t es_14_6MyFalse_3QVal_Int_1_bufchan_buf;
  assign es_14_6MyFalse_3QVal_Int_1_bufchan_r = (! es_14_6MyFalse_3QVal_Int_1_bufchan_buf[0]);
  assign es_14_6MyFalse_3QVal_Int_1_argbuf_d = (es_14_6MyFalse_3QVal_Int_1_bufchan_buf[0] ? es_14_6MyFalse_3QVal_Int_1_bufchan_buf :
                                                es_14_6MyFalse_3QVal_Int_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_14_6MyFalse_3QVal_Int_1_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((es_14_6MyFalse_3QVal_Int_1_argbuf_r && es_14_6MyFalse_3QVal_Int_1_bufchan_buf[0]))
        es_14_6MyFalse_3QVal_Int_1_bufchan_buf <= {32'd0, 1'd0};
      else if (((! es_14_6MyFalse_3QVal_Int_1_argbuf_r) && (! es_14_6MyFalse_3QVal_Int_1_bufchan_buf[0])))
        es_14_6MyFalse_3QVal_Int_1_bufchan_buf <= es_14_6MyFalse_3QVal_Int_1_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty MyDTInt_Int_Int) : (es_14_6MyFalse_4,QTree_Int) (es_14_2MyFalse,MyDTInt_Int_Int) > [(es_14_6MyFalse_4QNone_Int,MyDTInt_Int_Int),
                                                                                              (es_14_6MyFalse_4QVal_Int,MyDTInt_Int_Int),
                                                                                              (_243,MyDTInt_Int_Int),
                                                                                              (_242,MyDTInt_Int_Int)] */
  logic [3:0] es_14_2MyFalse_onehotd;
  always_comb
    if ((es_14_6MyFalse_4_d[0] && es_14_2MyFalse_d[0]))
      unique case (es_14_6MyFalse_4_d[2:1])
        2'd0: es_14_2MyFalse_onehotd = 4'd1;
        2'd1: es_14_2MyFalse_onehotd = 4'd2;
        2'd2: es_14_2MyFalse_onehotd = 4'd4;
        2'd3: es_14_2MyFalse_onehotd = 4'd8;
        default: es_14_2MyFalse_onehotd = 4'd0;
      endcase
    else es_14_2MyFalse_onehotd = 4'd0;
  assign es_14_6MyFalse_4QNone_Int_d = es_14_2MyFalse_onehotd[0];
  assign es_14_6MyFalse_4QVal_Int_d = es_14_2MyFalse_onehotd[1];
  assign _243_d = es_14_2MyFalse_onehotd[2];
  assign _242_d = es_14_2MyFalse_onehotd[3];
  assign es_14_2MyFalse_r = (| (es_14_2MyFalse_onehotd & {_242_r,
                                                          _243_r,
                                                          es_14_6MyFalse_4QVal_Int_r,
                                                          es_14_6MyFalse_4QNone_Int_r}));
  assign es_14_6MyFalse_4_r = es_14_2MyFalse_r;
  
  /* buf (Ty MyDTInt_Int_Int) : (es_14_6MyFalse_4QNone_Int,MyDTInt_Int_Int) > (es_14_6MyFalse_4QNone_Int_1_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t es_14_6MyFalse_4QNone_Int_bufchan_d;
  logic es_14_6MyFalse_4QNone_Int_bufchan_r;
  assign es_14_6MyFalse_4QNone_Int_r = ((! es_14_6MyFalse_4QNone_Int_bufchan_d[0]) || es_14_6MyFalse_4QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_14_6MyFalse_4QNone_Int_bufchan_d <= 1'd0;
    else
      if (es_14_6MyFalse_4QNone_Int_r)
        es_14_6MyFalse_4QNone_Int_bufchan_d <= es_14_6MyFalse_4QNone_Int_d;
  MyDTInt_Int_Int_t es_14_6MyFalse_4QNone_Int_bufchan_buf;
  assign es_14_6MyFalse_4QNone_Int_bufchan_r = (! es_14_6MyFalse_4QNone_Int_bufchan_buf[0]);
  assign es_14_6MyFalse_4QNone_Int_1_argbuf_d = (es_14_6MyFalse_4QNone_Int_bufchan_buf[0] ? es_14_6MyFalse_4QNone_Int_bufchan_buf :
                                                 es_14_6MyFalse_4QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_14_6MyFalse_4QNone_Int_bufchan_buf <= 1'd0;
    else
      if ((es_14_6MyFalse_4QNone_Int_1_argbuf_r && es_14_6MyFalse_4QNone_Int_bufchan_buf[0]))
        es_14_6MyFalse_4QNone_Int_bufchan_buf <= 1'd0;
      else if (((! es_14_6MyFalse_4QNone_Int_1_argbuf_r) && (! es_14_6MyFalse_4QNone_Int_bufchan_buf[0])))
        es_14_6MyFalse_4QNone_Int_bufchan_buf <= es_14_6MyFalse_4QNone_Int_bufchan_d;
  
  /* dcon (Ty TupMyDTInt_Int_Int___Int___Int,
      Dcon TupMyDTInt_Int_Int___Int___Int) : [(es_14_6MyFalse_4QNone_Int_1_argbuf,MyDTInt_Int_Int),
                                              (es_14_6MyFalse_3QNone_Int_1_argbuf,Int),
                                              (es_14_6MyFalse_8QNone_Int_1_argbuf,Int)] > (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int8,TupMyDTInt_Int_Int___Int___Int) */
  assign applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int8_d = TupMyDTInt_Int_Int___Int___Int_dc((& {es_14_6MyFalse_4QNone_Int_1_argbuf_d[0],
                                                                                                       es_14_6MyFalse_3QNone_Int_1_argbuf_d[0],
                                                                                                       es_14_6MyFalse_8QNone_Int_1_argbuf_d[0]}), es_14_6MyFalse_4QNone_Int_1_argbuf_d, es_14_6MyFalse_3QNone_Int_1_argbuf_d, es_14_6MyFalse_8QNone_Int_1_argbuf_d);
  assign {es_14_6MyFalse_4QNone_Int_1_argbuf_r,
          es_14_6MyFalse_3QNone_Int_1_argbuf_r,
          es_14_6MyFalse_8QNone_Int_1_argbuf_r} = {3 {(applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int8_r && applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int8_d[0])}};
  
  /* fork (Ty MyDTInt_Int_Int) : (es_14_6MyFalse_4QVal_Int,MyDTInt_Int_Int) > [(es_14_6MyFalse_4QVal_Int_1,MyDTInt_Int_Int),
                                                                          (es_14_6MyFalse_4QVal_Int_2,MyDTInt_Int_Int),
                                                                          (es_14_6MyFalse_4QVal_Int_3,MyDTInt_Int_Int)] */
  logic [2:0] es_14_6MyFalse_4QVal_Int_emitted;
  logic [2:0] es_14_6MyFalse_4QVal_Int_done;
  assign es_14_6MyFalse_4QVal_Int_1_d = (es_14_6MyFalse_4QVal_Int_d[0] && (! es_14_6MyFalse_4QVal_Int_emitted[0]));
  assign es_14_6MyFalse_4QVal_Int_2_d = (es_14_6MyFalse_4QVal_Int_d[0] && (! es_14_6MyFalse_4QVal_Int_emitted[1]));
  assign es_14_6MyFalse_4QVal_Int_3_d = (es_14_6MyFalse_4QVal_Int_d[0] && (! es_14_6MyFalse_4QVal_Int_emitted[2]));
  assign es_14_6MyFalse_4QVal_Int_done = (es_14_6MyFalse_4QVal_Int_emitted | ({es_14_6MyFalse_4QVal_Int_3_d[0],
                                                                               es_14_6MyFalse_4QVal_Int_2_d[0],
                                                                               es_14_6MyFalse_4QVal_Int_1_d[0]} & {es_14_6MyFalse_4QVal_Int_3_r,
                                                                                                                   es_14_6MyFalse_4QVal_Int_2_r,
                                                                                                                   es_14_6MyFalse_4QVal_Int_1_r}));
  assign es_14_6MyFalse_4QVal_Int_r = (& es_14_6MyFalse_4QVal_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_14_6MyFalse_4QVal_Int_emitted <= 3'd0;
    else
      es_14_6MyFalse_4QVal_Int_emitted <= (es_14_6MyFalse_4QVal_Int_r ? 3'd0 :
                                           es_14_6MyFalse_4QVal_Int_done);
  
  /* buf (Ty MyDTInt_Int_Int) : (es_14_6MyFalse_4QVal_Int_1,MyDTInt_Int_Int) > (es_14_6MyFalse_4QVal_Int_1_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t es_14_6MyFalse_4QVal_Int_1_bufchan_d;
  logic es_14_6MyFalse_4QVal_Int_1_bufchan_r;
  assign es_14_6MyFalse_4QVal_Int_1_r = ((! es_14_6MyFalse_4QVal_Int_1_bufchan_d[0]) || es_14_6MyFalse_4QVal_Int_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_14_6MyFalse_4QVal_Int_1_bufchan_d <= 1'd0;
    else
      if (es_14_6MyFalse_4QVal_Int_1_r)
        es_14_6MyFalse_4QVal_Int_1_bufchan_d <= es_14_6MyFalse_4QVal_Int_1_d;
  MyDTInt_Int_Int_t es_14_6MyFalse_4QVal_Int_1_bufchan_buf;
  assign es_14_6MyFalse_4QVal_Int_1_bufchan_r = (! es_14_6MyFalse_4QVal_Int_1_bufchan_buf[0]);
  assign es_14_6MyFalse_4QVal_Int_1_argbuf_d = (es_14_6MyFalse_4QVal_Int_1_bufchan_buf[0] ? es_14_6MyFalse_4QVal_Int_1_bufchan_buf :
                                                es_14_6MyFalse_4QVal_Int_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_14_6MyFalse_4QVal_Int_1_bufchan_buf <= 1'd0;
    else
      if ((es_14_6MyFalse_4QVal_Int_1_argbuf_r && es_14_6MyFalse_4QVal_Int_1_bufchan_buf[0]))
        es_14_6MyFalse_4QVal_Int_1_bufchan_buf <= 1'd0;
      else if (((! es_14_6MyFalse_4QVal_Int_1_argbuf_r) && (! es_14_6MyFalse_4QVal_Int_1_bufchan_buf[0])))
        es_14_6MyFalse_4QVal_Int_1_bufchan_buf <= es_14_6MyFalse_4QVal_Int_1_bufchan_d;
  
  /* dcon (Ty TupMyDTInt_Int_Int___Int___Int,
      Dcon TupMyDTInt_Int_Int___Int___Int) : [(es_14_6MyFalse_4QVal_Int_1_argbuf,MyDTInt_Int_Int),
                                              (es_14_6MyFalse_3QVal_Int_1_argbuf,Int),
                                              (es_14_6MyFalse_8QVal_Int_1_argbuf,Int)] > (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int9,TupMyDTInt_Int_Int___Int___Int) */
  assign applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int9_d = TupMyDTInt_Int_Int___Int___Int_dc((& {es_14_6MyFalse_4QVal_Int_1_argbuf_d[0],
                                                                                                       es_14_6MyFalse_3QVal_Int_1_argbuf_d[0],
                                                                                                       es_14_6MyFalse_8QVal_Int_1_argbuf_d[0]}), es_14_6MyFalse_4QVal_Int_1_argbuf_d, es_14_6MyFalse_3QVal_Int_1_argbuf_d, es_14_6MyFalse_8QVal_Int_1_argbuf_d);
  assign {es_14_6MyFalse_4QVal_Int_1_argbuf_r,
          es_14_6MyFalse_3QVal_Int_1_argbuf_r,
          es_14_6MyFalse_8QVal_Int_1_argbuf_r} = {3 {(applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int9_r && applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int9_d[0])}};
  
  /* buf (Ty MyDTInt_Int_Int) : (es_14_6MyFalse_4QVal_Int_2,MyDTInt_Int_Int) > (es_14_6MyFalse_4QVal_Int_2_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t es_14_6MyFalse_4QVal_Int_2_bufchan_d;
  logic es_14_6MyFalse_4QVal_Int_2_bufchan_r;
  assign es_14_6MyFalse_4QVal_Int_2_r = ((! es_14_6MyFalse_4QVal_Int_2_bufchan_d[0]) || es_14_6MyFalse_4QVal_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_14_6MyFalse_4QVal_Int_2_bufchan_d <= 1'd0;
    else
      if (es_14_6MyFalse_4QVal_Int_2_r)
        es_14_6MyFalse_4QVal_Int_2_bufchan_d <= es_14_6MyFalse_4QVal_Int_2_d;
  MyDTInt_Int_Int_t es_14_6MyFalse_4QVal_Int_2_bufchan_buf;
  assign es_14_6MyFalse_4QVal_Int_2_bufchan_r = (! es_14_6MyFalse_4QVal_Int_2_bufchan_buf[0]);
  assign es_14_6MyFalse_4QVal_Int_2_argbuf_d = (es_14_6MyFalse_4QVal_Int_2_bufchan_buf[0] ? es_14_6MyFalse_4QVal_Int_2_bufchan_buf :
                                                es_14_6MyFalse_4QVal_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_14_6MyFalse_4QVal_Int_2_bufchan_buf <= 1'd0;
    else
      if ((es_14_6MyFalse_4QVal_Int_2_argbuf_r && es_14_6MyFalse_4QVal_Int_2_bufchan_buf[0]))
        es_14_6MyFalse_4QVal_Int_2_bufchan_buf <= 1'd0;
      else if (((! es_14_6MyFalse_4QVal_Int_2_argbuf_r) && (! es_14_6MyFalse_4QVal_Int_2_bufchan_buf[0])))
        es_14_6MyFalse_4QVal_Int_2_bufchan_buf <= es_14_6MyFalse_4QVal_Int_2_bufchan_d;
  
  /* dcon (Ty TupMyDTInt_Int_Int___Int___Int,
      Dcon TupMyDTInt_Int_Int___Int___Int) : [(es_14_6MyFalse_4QVal_Int_2_argbuf,MyDTInt_Int_Int),
                                              (es_19_1_argbuf,Int),
                                              (v'aeR_1_argbuf,Int)] > (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int10,TupMyDTInt_Int_Int___Int___Int) */
  assign applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int10_d = TupMyDTInt_Int_Int___Int___Int_dc((& {es_14_6MyFalse_4QVal_Int_2_argbuf_d[0],
                                                                                                        es_19_1_argbuf_d[0],
                                                                                                        \v'aeR_1_argbuf_d [0]}), es_14_6MyFalse_4QVal_Int_2_argbuf_d, es_19_1_argbuf_d, \v'aeR_1_argbuf_d );
  assign {es_14_6MyFalse_4QVal_Int_2_argbuf_r,
          es_19_1_argbuf_r,
          \v'aeR_1_argbuf_r } = {3 {(applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int10_r && applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int10_d[0])}};
  
  /* demux (Ty QTree_Int,
       Ty Pointer_CTf_f_Int) : (es_14_6MyFalse_5,QTree_Int) (es_14_3MyFalse,Pointer_CTf_f_Int) > [(es_14_6MyFalse_5QNone_Int,Pointer_CTf_f_Int),
                                                                                                  (es_14_6MyFalse_5QVal_Int,Pointer_CTf_f_Int),
                                                                                                  (es_14_6MyFalse_5QNode_Int,Pointer_CTf_f_Int),
                                                                                                  (es_14_6MyFalse_5QError_Int,Pointer_CTf_f_Int)] */
  logic [3:0] es_14_3MyFalse_onehotd;
  always_comb
    if ((es_14_6MyFalse_5_d[0] && es_14_3MyFalse_d[0]))
      unique case (es_14_6MyFalse_5_d[2:1])
        2'd0: es_14_3MyFalse_onehotd = 4'd1;
        2'd1: es_14_3MyFalse_onehotd = 4'd2;
        2'd2: es_14_3MyFalse_onehotd = 4'd4;
        2'd3: es_14_3MyFalse_onehotd = 4'd8;
        default: es_14_3MyFalse_onehotd = 4'd0;
      endcase
    else es_14_3MyFalse_onehotd = 4'd0;
  assign es_14_6MyFalse_5QNone_Int_d = {es_14_3MyFalse_d[16:1],
                                        es_14_3MyFalse_onehotd[0]};
  assign es_14_6MyFalse_5QVal_Int_d = {es_14_3MyFalse_d[16:1],
                                       es_14_3MyFalse_onehotd[1]};
  assign es_14_6MyFalse_5QNode_Int_d = {es_14_3MyFalse_d[16:1],
                                        es_14_3MyFalse_onehotd[2]};
  assign es_14_6MyFalse_5QError_Int_d = {es_14_3MyFalse_d[16:1],
                                         es_14_3MyFalse_onehotd[3]};
  assign es_14_3MyFalse_r = (| (es_14_3MyFalse_onehotd & {es_14_6MyFalse_5QError_Int_r,
                                                          es_14_6MyFalse_5QNode_Int_r,
                                                          es_14_6MyFalse_5QVal_Int_r,
                                                          es_14_6MyFalse_5QNone_Int_r}));
  assign es_14_6MyFalse_5_r = es_14_3MyFalse_r;
  
  /* buf (Ty Pointer_CTf_f_Int) : (es_14_6MyFalse_5QError_Int,Pointer_CTf_f_Int) > (es_14_6MyFalse_5QError_Int_1_argbuf,Pointer_CTf_f_Int) */
  Pointer_CTf_f_Int_t es_14_6MyFalse_5QError_Int_bufchan_d;
  logic es_14_6MyFalse_5QError_Int_bufchan_r;
  assign es_14_6MyFalse_5QError_Int_r = ((! es_14_6MyFalse_5QError_Int_bufchan_d[0]) || es_14_6MyFalse_5QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_14_6MyFalse_5QError_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (es_14_6MyFalse_5QError_Int_r)
        es_14_6MyFalse_5QError_Int_bufchan_d <= es_14_6MyFalse_5QError_Int_d;
  Pointer_CTf_f_Int_t es_14_6MyFalse_5QError_Int_bufchan_buf;
  assign es_14_6MyFalse_5QError_Int_bufchan_r = (! es_14_6MyFalse_5QError_Int_bufchan_buf[0]);
  assign es_14_6MyFalse_5QError_Int_1_argbuf_d = (es_14_6MyFalse_5QError_Int_bufchan_buf[0] ? es_14_6MyFalse_5QError_Int_bufchan_buf :
                                                  es_14_6MyFalse_5QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_14_6MyFalse_5QError_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((es_14_6MyFalse_5QError_Int_1_argbuf_r && es_14_6MyFalse_5QError_Int_bufchan_buf[0]))
        es_14_6MyFalse_5QError_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! es_14_6MyFalse_5QError_Int_1_argbuf_r) && (! es_14_6MyFalse_5QError_Int_bufchan_buf[0])))
        es_14_6MyFalse_5QError_Int_bufchan_buf <= es_14_6MyFalse_5QError_Int_bufchan_d;
  
  /* buf (Ty Pointer_CTf_f_Int) : (es_14_6MyFalse_5QNode_Int,Pointer_CTf_f_Int) > (es_14_6MyFalse_5QNode_Int_1_argbuf,Pointer_CTf_f_Int) */
  Pointer_CTf_f_Int_t es_14_6MyFalse_5QNode_Int_bufchan_d;
  logic es_14_6MyFalse_5QNode_Int_bufchan_r;
  assign es_14_6MyFalse_5QNode_Int_r = ((! es_14_6MyFalse_5QNode_Int_bufchan_d[0]) || es_14_6MyFalse_5QNode_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_14_6MyFalse_5QNode_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (es_14_6MyFalse_5QNode_Int_r)
        es_14_6MyFalse_5QNode_Int_bufchan_d <= es_14_6MyFalse_5QNode_Int_d;
  Pointer_CTf_f_Int_t es_14_6MyFalse_5QNode_Int_bufchan_buf;
  assign es_14_6MyFalse_5QNode_Int_bufchan_r = (! es_14_6MyFalse_5QNode_Int_bufchan_buf[0]);
  assign es_14_6MyFalse_5QNode_Int_1_argbuf_d = (es_14_6MyFalse_5QNode_Int_bufchan_buf[0] ? es_14_6MyFalse_5QNode_Int_bufchan_buf :
                                                 es_14_6MyFalse_5QNode_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_14_6MyFalse_5QNode_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((es_14_6MyFalse_5QNode_Int_1_argbuf_r && es_14_6MyFalse_5QNode_Int_bufchan_buf[0]))
        es_14_6MyFalse_5QNode_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! es_14_6MyFalse_5QNode_Int_1_argbuf_r) && (! es_14_6MyFalse_5QNode_Int_bufchan_buf[0])))
        es_14_6MyFalse_5QNode_Int_bufchan_buf <= es_14_6MyFalse_5QNode_Int_bufchan_d;
  
  /* buf (Ty Pointer_CTf_f_Int) : (es_14_6MyFalse_5QNone_Int,Pointer_CTf_f_Int) > (es_14_6MyFalse_5QNone_Int_1_argbuf,Pointer_CTf_f_Int) */
  Pointer_CTf_f_Int_t es_14_6MyFalse_5QNone_Int_bufchan_d;
  logic es_14_6MyFalse_5QNone_Int_bufchan_r;
  assign es_14_6MyFalse_5QNone_Int_r = ((! es_14_6MyFalse_5QNone_Int_bufchan_d[0]) || es_14_6MyFalse_5QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_14_6MyFalse_5QNone_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (es_14_6MyFalse_5QNone_Int_r)
        es_14_6MyFalse_5QNone_Int_bufchan_d <= es_14_6MyFalse_5QNone_Int_d;
  Pointer_CTf_f_Int_t es_14_6MyFalse_5QNone_Int_bufchan_buf;
  assign es_14_6MyFalse_5QNone_Int_bufchan_r = (! es_14_6MyFalse_5QNone_Int_bufchan_buf[0]);
  assign es_14_6MyFalse_5QNone_Int_1_argbuf_d = (es_14_6MyFalse_5QNone_Int_bufchan_buf[0] ? es_14_6MyFalse_5QNone_Int_bufchan_buf :
                                                 es_14_6MyFalse_5QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_14_6MyFalse_5QNone_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((es_14_6MyFalse_5QNone_Int_1_argbuf_r && es_14_6MyFalse_5QNone_Int_bufchan_buf[0]))
        es_14_6MyFalse_5QNone_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! es_14_6MyFalse_5QNone_Int_1_argbuf_r) && (! es_14_6MyFalse_5QNone_Int_bufchan_buf[0])))
        es_14_6MyFalse_5QNone_Int_bufchan_buf <= es_14_6MyFalse_5QNone_Int_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Go) : (es_14_6MyFalse_6,QTree_Int) (es_14_4MyFalse,Go) > [(es_14_6MyFalse_6QNone_Int,Go),
                                                                    (es_14_6MyFalse_6QVal_Int,Go),
                                                                    (es_14_6MyFalse_6QNode_Int,Go),
                                                                    (es_14_6MyFalse_6QError_Int,Go)] */
  logic [3:0] es_14_4MyFalse_onehotd;
  always_comb
    if ((es_14_6MyFalse_6_d[0] && es_14_4MyFalse_d[0]))
      unique case (es_14_6MyFalse_6_d[2:1])
        2'd0: es_14_4MyFalse_onehotd = 4'd1;
        2'd1: es_14_4MyFalse_onehotd = 4'd2;
        2'd2: es_14_4MyFalse_onehotd = 4'd4;
        2'd3: es_14_4MyFalse_onehotd = 4'd8;
        default: es_14_4MyFalse_onehotd = 4'd0;
      endcase
    else es_14_4MyFalse_onehotd = 4'd0;
  assign es_14_6MyFalse_6QNone_Int_d = es_14_4MyFalse_onehotd[0];
  assign es_14_6MyFalse_6QVal_Int_d = es_14_4MyFalse_onehotd[1];
  assign es_14_6MyFalse_6QNode_Int_d = es_14_4MyFalse_onehotd[2];
  assign es_14_6MyFalse_6QError_Int_d = es_14_4MyFalse_onehotd[3];
  assign es_14_4MyFalse_r = (| (es_14_4MyFalse_onehotd & {es_14_6MyFalse_6QError_Int_r,
                                                          es_14_6MyFalse_6QNode_Int_r,
                                                          es_14_6MyFalse_6QVal_Int_r,
                                                          es_14_6MyFalse_6QNone_Int_r}));
  assign es_14_6MyFalse_6_r = es_14_4MyFalse_r;
  
  /* fork (Ty Go) : (es_14_6MyFalse_6QError_Int,Go) > [(es_14_6MyFalse_6QError_Int_1,Go),
                                                  (es_14_6MyFalse_6QError_Int_2,Go)] */
  logic [1:0] es_14_6MyFalse_6QError_Int_emitted;
  logic [1:0] es_14_6MyFalse_6QError_Int_done;
  assign es_14_6MyFalse_6QError_Int_1_d = (es_14_6MyFalse_6QError_Int_d[0] && (! es_14_6MyFalse_6QError_Int_emitted[0]));
  assign es_14_6MyFalse_6QError_Int_2_d = (es_14_6MyFalse_6QError_Int_d[0] && (! es_14_6MyFalse_6QError_Int_emitted[1]));
  assign es_14_6MyFalse_6QError_Int_done = (es_14_6MyFalse_6QError_Int_emitted | ({es_14_6MyFalse_6QError_Int_2_d[0],
                                                                                   es_14_6MyFalse_6QError_Int_1_d[0]} & {es_14_6MyFalse_6QError_Int_2_r,
                                                                                                                         es_14_6MyFalse_6QError_Int_1_r}));
  assign es_14_6MyFalse_6QError_Int_r = (& es_14_6MyFalse_6QError_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_14_6MyFalse_6QError_Int_emitted <= 2'd0;
    else
      es_14_6MyFalse_6QError_Int_emitted <= (es_14_6MyFalse_6QError_Int_r ? 2'd0 :
                                             es_14_6MyFalse_6QError_Int_done);
  
  /* dcon (Ty QTree_Int,
      Dcon QError_Int) : [(es_14_6MyFalse_6QError_Int_1,Go)] > (es_14_6MyFalse_6QError_Int_1QError_Int,QTree_Int) */
  assign es_14_6MyFalse_6QError_Int_1QError_Int_d = QError_Int_dc((& {es_14_6MyFalse_6QError_Int_1_d[0]}), es_14_6MyFalse_6QError_Int_1_d);
  assign {es_14_6MyFalse_6QError_Int_1_r} = {1 {(es_14_6MyFalse_6QError_Int_1QError_Int_r && es_14_6MyFalse_6QError_Int_1QError_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (es_14_6MyFalse_6QError_Int_1QError_Int,QTree_Int) > (lizzieLet40_1_argbuf,QTree_Int) */
  QTree_Int_t es_14_6MyFalse_6QError_Int_1QError_Int_bufchan_d;
  logic es_14_6MyFalse_6QError_Int_1QError_Int_bufchan_r;
  assign es_14_6MyFalse_6QError_Int_1QError_Int_r = ((! es_14_6MyFalse_6QError_Int_1QError_Int_bufchan_d[0]) || es_14_6MyFalse_6QError_Int_1QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_14_6MyFalse_6QError_Int_1QError_Int_bufchan_d <= {66'd0, 1'd0};
    else
      if (es_14_6MyFalse_6QError_Int_1QError_Int_r)
        es_14_6MyFalse_6QError_Int_1QError_Int_bufchan_d <= es_14_6MyFalse_6QError_Int_1QError_Int_d;
  QTree_Int_t es_14_6MyFalse_6QError_Int_1QError_Int_bufchan_buf;
  assign es_14_6MyFalse_6QError_Int_1QError_Int_bufchan_r = (! es_14_6MyFalse_6QError_Int_1QError_Int_bufchan_buf[0]);
  assign lizzieLet40_1_argbuf_d = (es_14_6MyFalse_6QError_Int_1QError_Int_bufchan_buf[0] ? es_14_6MyFalse_6QError_Int_1QError_Int_bufchan_buf :
                                   es_14_6MyFalse_6QError_Int_1QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_14_6MyFalse_6QError_Int_1QError_Int_bufchan_buf <= {66'd0,
                                                             1'd0};
    else
      if ((lizzieLet40_1_argbuf_r && es_14_6MyFalse_6QError_Int_1QError_Int_bufchan_buf[0]))
        es_14_6MyFalse_6QError_Int_1QError_Int_bufchan_buf <= {66'd0,
                                                               1'd0};
      else if (((! lizzieLet40_1_argbuf_r) && (! es_14_6MyFalse_6QError_Int_1QError_Int_bufchan_buf[0])))
        es_14_6MyFalse_6QError_Int_1QError_Int_bufchan_buf <= es_14_6MyFalse_6QError_Int_1QError_Int_bufchan_d;
  
  /* buf (Ty Go) : (es_14_6MyFalse_6QError_Int_2,Go) > (es_14_6MyFalse_6QError_Int_2_argbuf,Go) */
  Go_t es_14_6MyFalse_6QError_Int_2_bufchan_d;
  logic es_14_6MyFalse_6QError_Int_2_bufchan_r;
  assign es_14_6MyFalse_6QError_Int_2_r = ((! es_14_6MyFalse_6QError_Int_2_bufchan_d[0]) || es_14_6MyFalse_6QError_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_14_6MyFalse_6QError_Int_2_bufchan_d <= 1'd0;
    else
      if (es_14_6MyFalse_6QError_Int_2_r)
        es_14_6MyFalse_6QError_Int_2_bufchan_d <= es_14_6MyFalse_6QError_Int_2_d;
  Go_t es_14_6MyFalse_6QError_Int_2_bufchan_buf;
  assign es_14_6MyFalse_6QError_Int_2_bufchan_r = (! es_14_6MyFalse_6QError_Int_2_bufchan_buf[0]);
  assign es_14_6MyFalse_6QError_Int_2_argbuf_d = (es_14_6MyFalse_6QError_Int_2_bufchan_buf[0] ? es_14_6MyFalse_6QError_Int_2_bufchan_buf :
                                                  es_14_6MyFalse_6QError_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_14_6MyFalse_6QError_Int_2_bufchan_buf <= 1'd0;
    else
      if ((es_14_6MyFalse_6QError_Int_2_argbuf_r && es_14_6MyFalse_6QError_Int_2_bufchan_buf[0]))
        es_14_6MyFalse_6QError_Int_2_bufchan_buf <= 1'd0;
      else if (((! es_14_6MyFalse_6QError_Int_2_argbuf_r) && (! es_14_6MyFalse_6QError_Int_2_bufchan_buf[0])))
        es_14_6MyFalse_6QError_Int_2_bufchan_buf <= es_14_6MyFalse_6QError_Int_2_bufchan_d;
  
  /* fork (Ty Go) : (es_14_6MyFalse_6QNode_Int,Go) > [(es_14_6MyFalse_6QNode_Int_1,Go),
                                                 (es_14_6MyFalse_6QNode_Int_2,Go)] */
  logic [1:0] es_14_6MyFalse_6QNode_Int_emitted;
  logic [1:0] es_14_6MyFalse_6QNode_Int_done;
  assign es_14_6MyFalse_6QNode_Int_1_d = (es_14_6MyFalse_6QNode_Int_d[0] && (! es_14_6MyFalse_6QNode_Int_emitted[0]));
  assign es_14_6MyFalse_6QNode_Int_2_d = (es_14_6MyFalse_6QNode_Int_d[0] && (! es_14_6MyFalse_6QNode_Int_emitted[1]));
  assign es_14_6MyFalse_6QNode_Int_done = (es_14_6MyFalse_6QNode_Int_emitted | ({es_14_6MyFalse_6QNode_Int_2_d[0],
                                                                                 es_14_6MyFalse_6QNode_Int_1_d[0]} & {es_14_6MyFalse_6QNode_Int_2_r,
                                                                                                                      es_14_6MyFalse_6QNode_Int_1_r}));
  assign es_14_6MyFalse_6QNode_Int_r = (& es_14_6MyFalse_6QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_14_6MyFalse_6QNode_Int_emitted <= 2'd0;
    else
      es_14_6MyFalse_6QNode_Int_emitted <= (es_14_6MyFalse_6QNode_Int_r ? 2'd0 :
                                            es_14_6MyFalse_6QNode_Int_done);
  
  /* dcon (Ty QTree_Int,
      Dcon QError_Int) : [(es_14_6MyFalse_6QNode_Int_1,Go)] > (es_14_6MyFalse_6QNode_Int_1QError_Int,QTree_Int) */
  assign es_14_6MyFalse_6QNode_Int_1QError_Int_d = QError_Int_dc((& {es_14_6MyFalse_6QNode_Int_1_d[0]}), es_14_6MyFalse_6QNode_Int_1_d);
  assign {es_14_6MyFalse_6QNode_Int_1_r} = {1 {(es_14_6MyFalse_6QNode_Int_1QError_Int_r && es_14_6MyFalse_6QNode_Int_1QError_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (es_14_6MyFalse_6QNode_Int_1QError_Int,QTree_Int) > (lizzieLet39_1_1_argbuf,QTree_Int) */
  QTree_Int_t es_14_6MyFalse_6QNode_Int_1QError_Int_bufchan_d;
  logic es_14_6MyFalse_6QNode_Int_1QError_Int_bufchan_r;
  assign es_14_6MyFalse_6QNode_Int_1QError_Int_r = ((! es_14_6MyFalse_6QNode_Int_1QError_Int_bufchan_d[0]) || es_14_6MyFalse_6QNode_Int_1QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_14_6MyFalse_6QNode_Int_1QError_Int_bufchan_d <= {66'd0, 1'd0};
    else
      if (es_14_6MyFalse_6QNode_Int_1QError_Int_r)
        es_14_6MyFalse_6QNode_Int_1QError_Int_bufchan_d <= es_14_6MyFalse_6QNode_Int_1QError_Int_d;
  QTree_Int_t es_14_6MyFalse_6QNode_Int_1QError_Int_bufchan_buf;
  assign es_14_6MyFalse_6QNode_Int_1QError_Int_bufchan_r = (! es_14_6MyFalse_6QNode_Int_1QError_Int_bufchan_buf[0]);
  assign lizzieLet39_1_1_argbuf_d = (es_14_6MyFalse_6QNode_Int_1QError_Int_bufchan_buf[0] ? es_14_6MyFalse_6QNode_Int_1QError_Int_bufchan_buf :
                                     es_14_6MyFalse_6QNode_Int_1QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_14_6MyFalse_6QNode_Int_1QError_Int_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((lizzieLet39_1_1_argbuf_r && es_14_6MyFalse_6QNode_Int_1QError_Int_bufchan_buf[0]))
        es_14_6MyFalse_6QNode_Int_1QError_Int_bufchan_buf <= {66'd0, 1'd0};
      else if (((! lizzieLet39_1_1_argbuf_r) && (! es_14_6MyFalse_6QNode_Int_1QError_Int_bufchan_buf[0])))
        es_14_6MyFalse_6QNode_Int_1QError_Int_bufchan_buf <= es_14_6MyFalse_6QNode_Int_1QError_Int_bufchan_d;
  
  /* buf (Ty Go) : (es_14_6MyFalse_6QNode_Int_2,Go) > (es_14_6MyFalse_6QNode_Int_2_argbuf,Go) */
  Go_t es_14_6MyFalse_6QNode_Int_2_bufchan_d;
  logic es_14_6MyFalse_6QNode_Int_2_bufchan_r;
  assign es_14_6MyFalse_6QNode_Int_2_r = ((! es_14_6MyFalse_6QNode_Int_2_bufchan_d[0]) || es_14_6MyFalse_6QNode_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_14_6MyFalse_6QNode_Int_2_bufchan_d <= 1'd0;
    else
      if (es_14_6MyFalse_6QNode_Int_2_r)
        es_14_6MyFalse_6QNode_Int_2_bufchan_d <= es_14_6MyFalse_6QNode_Int_2_d;
  Go_t es_14_6MyFalse_6QNode_Int_2_bufchan_buf;
  assign es_14_6MyFalse_6QNode_Int_2_bufchan_r = (! es_14_6MyFalse_6QNode_Int_2_bufchan_buf[0]);
  assign es_14_6MyFalse_6QNode_Int_2_argbuf_d = (es_14_6MyFalse_6QNode_Int_2_bufchan_buf[0] ? es_14_6MyFalse_6QNode_Int_2_bufchan_buf :
                                                 es_14_6MyFalse_6QNode_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_14_6MyFalse_6QNode_Int_2_bufchan_buf <= 1'd0;
    else
      if ((es_14_6MyFalse_6QNode_Int_2_argbuf_r && es_14_6MyFalse_6QNode_Int_2_bufchan_buf[0]))
        es_14_6MyFalse_6QNode_Int_2_bufchan_buf <= 1'd0;
      else if (((! es_14_6MyFalse_6QNode_Int_2_argbuf_r) && (! es_14_6MyFalse_6QNode_Int_2_bufchan_buf[0])))
        es_14_6MyFalse_6QNode_Int_2_bufchan_buf <= es_14_6MyFalse_6QNode_Int_2_bufchan_d;
  
  /* buf (Ty Go) : (es_14_6MyFalse_6QNone_Int,Go) > (es_14_6MyFalse_6QNone_Int_1_argbuf,Go) */
  Go_t es_14_6MyFalse_6QNone_Int_bufchan_d;
  logic es_14_6MyFalse_6QNone_Int_bufchan_r;
  assign es_14_6MyFalse_6QNone_Int_r = ((! es_14_6MyFalse_6QNone_Int_bufchan_d[0]) || es_14_6MyFalse_6QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_14_6MyFalse_6QNone_Int_bufchan_d <= 1'd0;
    else
      if (es_14_6MyFalse_6QNone_Int_r)
        es_14_6MyFalse_6QNone_Int_bufchan_d <= es_14_6MyFalse_6QNone_Int_d;
  Go_t es_14_6MyFalse_6QNone_Int_bufchan_buf;
  assign es_14_6MyFalse_6QNone_Int_bufchan_r = (! es_14_6MyFalse_6QNone_Int_bufchan_buf[0]);
  assign es_14_6MyFalse_6QNone_Int_1_argbuf_d = (es_14_6MyFalse_6QNone_Int_bufchan_buf[0] ? es_14_6MyFalse_6QNone_Int_bufchan_buf :
                                                 es_14_6MyFalse_6QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_14_6MyFalse_6QNone_Int_bufchan_buf <= 1'd0;
    else
      if ((es_14_6MyFalse_6QNone_Int_1_argbuf_r && es_14_6MyFalse_6QNone_Int_bufchan_buf[0]))
        es_14_6MyFalse_6QNone_Int_bufchan_buf <= 1'd0;
      else if (((! es_14_6MyFalse_6QNone_Int_1_argbuf_r) && (! es_14_6MyFalse_6QNone_Int_bufchan_buf[0])))
        es_14_6MyFalse_6QNone_Int_bufchan_buf <= es_14_6MyFalse_6QNone_Int_bufchan_d;
  
  /* fork (Ty Go) : (es_14_6MyFalse_6QVal_Int,Go) > [(es_14_6MyFalse_6QVal_Int_1,Go),
                                                (es_14_6MyFalse_6QVal_Int_2,Go)] */
  logic [1:0] es_14_6MyFalse_6QVal_Int_emitted;
  logic [1:0] es_14_6MyFalse_6QVal_Int_done;
  assign es_14_6MyFalse_6QVal_Int_1_d = (es_14_6MyFalse_6QVal_Int_d[0] && (! es_14_6MyFalse_6QVal_Int_emitted[0]));
  assign es_14_6MyFalse_6QVal_Int_2_d = (es_14_6MyFalse_6QVal_Int_d[0] && (! es_14_6MyFalse_6QVal_Int_emitted[1]));
  assign es_14_6MyFalse_6QVal_Int_done = (es_14_6MyFalse_6QVal_Int_emitted | ({es_14_6MyFalse_6QVal_Int_2_d[0],
                                                                               es_14_6MyFalse_6QVal_Int_1_d[0]} & {es_14_6MyFalse_6QVal_Int_2_r,
                                                                                                                   es_14_6MyFalse_6QVal_Int_1_r}));
  assign es_14_6MyFalse_6QVal_Int_r = (& es_14_6MyFalse_6QVal_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_14_6MyFalse_6QVal_Int_emitted <= 2'd0;
    else
      es_14_6MyFalse_6QVal_Int_emitted <= (es_14_6MyFalse_6QVal_Int_r ? 2'd0 :
                                           es_14_6MyFalse_6QVal_Int_done);
  
  /* buf (Ty Go) : (es_14_6MyFalse_6QVal_Int_1,Go) > (es_14_6MyFalse_6QVal_Int_1_argbuf,Go) */
  Go_t es_14_6MyFalse_6QVal_Int_1_bufchan_d;
  logic es_14_6MyFalse_6QVal_Int_1_bufchan_r;
  assign es_14_6MyFalse_6QVal_Int_1_r = ((! es_14_6MyFalse_6QVal_Int_1_bufchan_d[0]) || es_14_6MyFalse_6QVal_Int_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_14_6MyFalse_6QVal_Int_1_bufchan_d <= 1'd0;
    else
      if (es_14_6MyFalse_6QVal_Int_1_r)
        es_14_6MyFalse_6QVal_Int_1_bufchan_d <= es_14_6MyFalse_6QVal_Int_1_d;
  Go_t es_14_6MyFalse_6QVal_Int_1_bufchan_buf;
  assign es_14_6MyFalse_6QVal_Int_1_bufchan_r = (! es_14_6MyFalse_6QVal_Int_1_bufchan_buf[0]);
  assign es_14_6MyFalse_6QVal_Int_1_argbuf_d = (es_14_6MyFalse_6QVal_Int_1_bufchan_buf[0] ? es_14_6MyFalse_6QVal_Int_1_bufchan_buf :
                                                es_14_6MyFalse_6QVal_Int_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_14_6MyFalse_6QVal_Int_1_bufchan_buf <= 1'd0;
    else
      if ((es_14_6MyFalse_6QVal_Int_1_argbuf_r && es_14_6MyFalse_6QVal_Int_1_bufchan_buf[0]))
        es_14_6MyFalse_6QVal_Int_1_bufchan_buf <= 1'd0;
      else if (((! es_14_6MyFalse_6QVal_Int_1_argbuf_r) && (! es_14_6MyFalse_6QVal_Int_1_bufchan_buf[0])))
        es_14_6MyFalse_6QVal_Int_1_bufchan_buf <= es_14_6MyFalse_6QVal_Int_1_bufchan_d;
  
  /* dcon (Ty TupGo___MyDTInt_Bool___Int,
      Dcon TupGo___MyDTInt_Bool___Int) : [(es_14_6MyFalse_6QVal_Int_1_argbuf,Go),
                                          (es_14_6MyFalse_7QVal_Int_1_argbuf,MyDTInt_Bool),
                                          (es_17_1_argbuf,Int)] > (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int5,TupGo___MyDTInt_Bool___Int) */
  assign applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int5_d = TupGo___MyDTInt_Bool___Int_dc((& {es_14_6MyFalse_6QVal_Int_1_argbuf_d[0],
                                                                                            es_14_6MyFalse_7QVal_Int_1_argbuf_d[0],
                                                                                            es_17_1_argbuf_d[0]}), es_14_6MyFalse_6QVal_Int_1_argbuf_d, es_14_6MyFalse_7QVal_Int_1_argbuf_d, es_17_1_argbuf_d);
  assign {es_14_6MyFalse_6QVal_Int_1_argbuf_r,
          es_14_6MyFalse_7QVal_Int_1_argbuf_r,
          es_17_1_argbuf_r} = {3 {(applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int5_r && applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int5_d[0])}};
  
  /* demux (Ty QTree_Int,
       Ty MyDTInt_Bool) : (es_14_6MyFalse_7,QTree_Int) (es_14_5MyFalse,MyDTInt_Bool) > [(_241,MyDTInt_Bool),
                                                                                        (es_14_6MyFalse_7QVal_Int,MyDTInt_Bool),
                                                                                        (_240,MyDTInt_Bool),
                                                                                        (_239,MyDTInt_Bool)] */
  logic [3:0] es_14_5MyFalse_onehotd;
  always_comb
    if ((es_14_6MyFalse_7_d[0] && es_14_5MyFalse_d[0]))
      unique case (es_14_6MyFalse_7_d[2:1])
        2'd0: es_14_5MyFalse_onehotd = 4'd1;
        2'd1: es_14_5MyFalse_onehotd = 4'd2;
        2'd2: es_14_5MyFalse_onehotd = 4'd4;
        2'd3: es_14_5MyFalse_onehotd = 4'd8;
        default: es_14_5MyFalse_onehotd = 4'd0;
      endcase
    else es_14_5MyFalse_onehotd = 4'd0;
  assign _241_d = es_14_5MyFalse_onehotd[0];
  assign es_14_6MyFalse_7QVal_Int_d = es_14_5MyFalse_onehotd[1];
  assign _240_d = es_14_5MyFalse_onehotd[2];
  assign _239_d = es_14_5MyFalse_onehotd[3];
  assign es_14_5MyFalse_r = (| (es_14_5MyFalse_onehotd & {_239_r,
                                                          _240_r,
                                                          es_14_6MyFalse_7QVal_Int_r,
                                                          _241_r}));
  assign es_14_6MyFalse_7_r = es_14_5MyFalse_r;
  
  /* buf (Ty MyDTInt_Bool) : (es_14_6MyFalse_7QVal_Int,MyDTInt_Bool) > (es_14_6MyFalse_7QVal_Int_1_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t es_14_6MyFalse_7QVal_Int_bufchan_d;
  logic es_14_6MyFalse_7QVal_Int_bufchan_r;
  assign es_14_6MyFalse_7QVal_Int_r = ((! es_14_6MyFalse_7QVal_Int_bufchan_d[0]) || es_14_6MyFalse_7QVal_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_14_6MyFalse_7QVal_Int_bufchan_d <= 1'd0;
    else
      if (es_14_6MyFalse_7QVal_Int_r)
        es_14_6MyFalse_7QVal_Int_bufchan_d <= es_14_6MyFalse_7QVal_Int_d;
  MyDTInt_Bool_t es_14_6MyFalse_7QVal_Int_bufchan_buf;
  assign es_14_6MyFalse_7QVal_Int_bufchan_r = (! es_14_6MyFalse_7QVal_Int_bufchan_buf[0]);
  assign es_14_6MyFalse_7QVal_Int_1_argbuf_d = (es_14_6MyFalse_7QVal_Int_bufchan_buf[0] ? es_14_6MyFalse_7QVal_Int_bufchan_buf :
                                                es_14_6MyFalse_7QVal_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_14_6MyFalse_7QVal_Int_bufchan_buf <= 1'd0;
    else
      if ((es_14_6MyFalse_7QVal_Int_1_argbuf_r && es_14_6MyFalse_7QVal_Int_bufchan_buf[0]))
        es_14_6MyFalse_7QVal_Int_bufchan_buf <= 1'd0;
      else if (((! es_14_6MyFalse_7QVal_Int_1_argbuf_r) && (! es_14_6MyFalse_7QVal_Int_bufchan_buf[0])))
        es_14_6MyFalse_7QVal_Int_bufchan_buf <= es_14_6MyFalse_7QVal_Int_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Int) : (es_14_6MyFalse_8,QTree_Int) (es_14_8MyFalse,Int) > [(es_14_6MyFalse_8QNone_Int,Int),
                                                                      (es_14_6MyFalse_8QVal_Int,Int),
                                                                      (_238,Int),
                                                                      (_237,Int)] */
  logic [3:0] es_14_8MyFalse_onehotd;
  always_comb
    if ((es_14_6MyFalse_8_d[0] && es_14_8MyFalse_d[0]))
      unique case (es_14_6MyFalse_8_d[2:1])
        2'd0: es_14_8MyFalse_onehotd = 4'd1;
        2'd1: es_14_8MyFalse_onehotd = 4'd2;
        2'd2: es_14_8MyFalse_onehotd = 4'd4;
        2'd3: es_14_8MyFalse_onehotd = 4'd8;
        default: es_14_8MyFalse_onehotd = 4'd0;
      endcase
    else es_14_8MyFalse_onehotd = 4'd0;
  assign es_14_6MyFalse_8QNone_Int_d = {es_14_8MyFalse_d[32:1],
                                        es_14_8MyFalse_onehotd[0]};
  assign es_14_6MyFalse_8QVal_Int_d = {es_14_8MyFalse_d[32:1],
                                       es_14_8MyFalse_onehotd[1]};
  assign _238_d = {es_14_8MyFalse_d[32:1],
                   es_14_8MyFalse_onehotd[2]};
  assign _237_d = {es_14_8MyFalse_d[32:1],
                   es_14_8MyFalse_onehotd[3]};
  assign es_14_8MyFalse_r = (| (es_14_8MyFalse_onehotd & {_237_r,
                                                          _238_r,
                                                          es_14_6MyFalse_8QVal_Int_r,
                                                          es_14_6MyFalse_8QNone_Int_r}));
  assign es_14_6MyFalse_8_r = es_14_8MyFalse_r;
  
  /* buf (Ty Int) : (es_14_6MyFalse_8QNone_Int,Int) > (es_14_6MyFalse_8QNone_Int_1_argbuf,Int) */
  Int_t es_14_6MyFalse_8QNone_Int_bufchan_d;
  logic es_14_6MyFalse_8QNone_Int_bufchan_r;
  assign es_14_6MyFalse_8QNone_Int_r = ((! es_14_6MyFalse_8QNone_Int_bufchan_d[0]) || es_14_6MyFalse_8QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_14_6MyFalse_8QNone_Int_bufchan_d <= {32'd0, 1'd0};
    else
      if (es_14_6MyFalse_8QNone_Int_r)
        es_14_6MyFalse_8QNone_Int_bufchan_d <= es_14_6MyFalse_8QNone_Int_d;
  Int_t es_14_6MyFalse_8QNone_Int_bufchan_buf;
  assign es_14_6MyFalse_8QNone_Int_bufchan_r = (! es_14_6MyFalse_8QNone_Int_bufchan_buf[0]);
  assign es_14_6MyFalse_8QNone_Int_1_argbuf_d = (es_14_6MyFalse_8QNone_Int_bufchan_buf[0] ? es_14_6MyFalse_8QNone_Int_bufchan_buf :
                                                 es_14_6MyFalse_8QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_14_6MyFalse_8QNone_Int_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((es_14_6MyFalse_8QNone_Int_1_argbuf_r && es_14_6MyFalse_8QNone_Int_bufchan_buf[0]))
        es_14_6MyFalse_8QNone_Int_bufchan_buf <= {32'd0, 1'd0};
      else if (((! es_14_6MyFalse_8QNone_Int_1_argbuf_r) && (! es_14_6MyFalse_8QNone_Int_bufchan_buf[0])))
        es_14_6MyFalse_8QNone_Int_bufchan_buf <= es_14_6MyFalse_8QNone_Int_bufchan_d;
  
  /* fork (Ty Int) : (es_14_6MyFalse_8QVal_Int,Int) > [(es_14_6MyFalse_8QVal_Int_1,Int),
                                                  (es_14_6MyFalse_8QVal_Int_2,Int)] */
  logic [1:0] es_14_6MyFalse_8QVal_Int_emitted;
  logic [1:0] es_14_6MyFalse_8QVal_Int_done;
  assign es_14_6MyFalse_8QVal_Int_1_d = {es_14_6MyFalse_8QVal_Int_d[32:1],
                                         (es_14_6MyFalse_8QVal_Int_d[0] && (! es_14_6MyFalse_8QVal_Int_emitted[0]))};
  assign es_14_6MyFalse_8QVal_Int_2_d = {es_14_6MyFalse_8QVal_Int_d[32:1],
                                         (es_14_6MyFalse_8QVal_Int_d[0] && (! es_14_6MyFalse_8QVal_Int_emitted[1]))};
  assign es_14_6MyFalse_8QVal_Int_done = (es_14_6MyFalse_8QVal_Int_emitted | ({es_14_6MyFalse_8QVal_Int_2_d[0],
                                                                               es_14_6MyFalse_8QVal_Int_1_d[0]} & {es_14_6MyFalse_8QVal_Int_2_r,
                                                                                                                   es_14_6MyFalse_8QVal_Int_1_r}));
  assign es_14_6MyFalse_8QVal_Int_r = (& es_14_6MyFalse_8QVal_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_14_6MyFalse_8QVal_Int_emitted <= 2'd0;
    else
      es_14_6MyFalse_8QVal_Int_emitted <= (es_14_6MyFalse_8QVal_Int_r ? 2'd0 :
                                           es_14_6MyFalse_8QVal_Int_done);
  
  /* buf (Ty Int) : (es_14_6MyFalse_8QVal_Int_1,Int) > (es_14_6MyFalse_8QVal_Int_1_argbuf,Int) */
  Int_t es_14_6MyFalse_8QVal_Int_1_bufchan_d;
  logic es_14_6MyFalse_8QVal_Int_1_bufchan_r;
  assign es_14_6MyFalse_8QVal_Int_1_r = ((! es_14_6MyFalse_8QVal_Int_1_bufchan_d[0]) || es_14_6MyFalse_8QVal_Int_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_14_6MyFalse_8QVal_Int_1_bufchan_d <= {32'd0, 1'd0};
    else
      if (es_14_6MyFalse_8QVal_Int_1_r)
        es_14_6MyFalse_8QVal_Int_1_bufchan_d <= es_14_6MyFalse_8QVal_Int_1_d;
  Int_t es_14_6MyFalse_8QVal_Int_1_bufchan_buf;
  assign es_14_6MyFalse_8QVal_Int_1_bufchan_r = (! es_14_6MyFalse_8QVal_Int_1_bufchan_buf[0]);
  assign es_14_6MyFalse_8QVal_Int_1_argbuf_d = (es_14_6MyFalse_8QVal_Int_1_bufchan_buf[0] ? es_14_6MyFalse_8QVal_Int_1_bufchan_buf :
                                                es_14_6MyFalse_8QVal_Int_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_14_6MyFalse_8QVal_Int_1_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((es_14_6MyFalse_8QVal_Int_1_argbuf_r && es_14_6MyFalse_8QVal_Int_1_bufchan_buf[0]))
        es_14_6MyFalse_8QVal_Int_1_bufchan_buf <= {32'd0, 1'd0};
      else if (((! es_14_6MyFalse_8QVal_Int_1_argbuf_r) && (! es_14_6MyFalse_8QVal_Int_1_bufchan_buf[0])))
        es_14_6MyFalse_8QVal_Int_1_bufchan_buf <= es_14_6MyFalse_8QVal_Int_1_bufchan_d;
  
  /* demux (Ty MyBool,
       Ty Pointer_QTree_Int) : (es_14_7,MyBool) (lizzieLet17_5QVal_Int_9QVal_Int,Pointer_QTree_Int) > [(_236,Pointer_QTree_Int),
                                                                                                       (es_14_7MyTrue,Pointer_QTree_Int)] */
  logic [1:0] lizzieLet17_5QVal_Int_9QVal_Int_onehotd;
  always_comb
    if ((es_14_7_d[0] && lizzieLet17_5QVal_Int_9QVal_Int_d[0]))
      unique case (es_14_7_d[1:1])
        1'd0: lizzieLet17_5QVal_Int_9QVal_Int_onehotd = 2'd1;
        1'd1: lizzieLet17_5QVal_Int_9QVal_Int_onehotd = 2'd2;
        default: lizzieLet17_5QVal_Int_9QVal_Int_onehotd = 2'd0;
      endcase
    else lizzieLet17_5QVal_Int_9QVal_Int_onehotd = 2'd0;
  assign _236_d = {lizzieLet17_5QVal_Int_9QVal_Int_d[16:1],
                   lizzieLet17_5QVal_Int_9QVal_Int_onehotd[0]};
  assign es_14_7MyTrue_d = {lizzieLet17_5QVal_Int_9QVal_Int_d[16:1],
                            lizzieLet17_5QVal_Int_9QVal_Int_onehotd[1]};
  assign lizzieLet17_5QVal_Int_9QVal_Int_r = (| (lizzieLet17_5QVal_Int_9QVal_Int_onehotd & {es_14_7MyTrue_r,
                                                                                            _236_r}));
  assign es_14_7_r = lizzieLet17_5QVal_Int_9QVal_Int_r;
  
  /* buf (Ty Pointer_QTree_Int) : (es_14_7MyTrue,Pointer_QTree_Int) > (es_14_7MyTrue_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t es_14_7MyTrue_bufchan_d;
  logic es_14_7MyTrue_bufchan_r;
  assign es_14_7MyTrue_r = ((! es_14_7MyTrue_bufchan_d[0]) || es_14_7MyTrue_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_14_7MyTrue_bufchan_d <= {16'd0, 1'd0};
    else
      if (es_14_7MyTrue_r) es_14_7MyTrue_bufchan_d <= es_14_7MyTrue_d;
  Pointer_QTree_Int_t es_14_7MyTrue_bufchan_buf;
  assign es_14_7MyTrue_bufchan_r = (! es_14_7MyTrue_bufchan_buf[0]);
  assign es_14_7MyTrue_1_argbuf_d = (es_14_7MyTrue_bufchan_buf[0] ? es_14_7MyTrue_bufchan_buf :
                                     es_14_7MyTrue_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_14_7MyTrue_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((es_14_7MyTrue_1_argbuf_r && es_14_7MyTrue_bufchan_buf[0]))
        es_14_7MyTrue_bufchan_buf <= {16'd0, 1'd0};
      else if (((! es_14_7MyTrue_1_argbuf_r) && (! es_14_7MyTrue_bufchan_buf[0])))
        es_14_7MyTrue_bufchan_buf <= es_14_7MyTrue_bufchan_d;
  
  /* demux (Ty MyBool,
       Ty Int) : (es_14_8,MyBool) (vaeQ_2,Int) > [(es_14_8MyFalse,Int),
                                                  (_235,Int)] */
  logic [1:0] vaeQ_2_onehotd;
  always_comb
    if ((es_14_8_d[0] && vaeQ_2_d[0]))
      unique case (es_14_8_d[1:1])
        1'd0: vaeQ_2_onehotd = 2'd1;
        1'd1: vaeQ_2_onehotd = 2'd2;
        default: vaeQ_2_onehotd = 2'd0;
      endcase
    else vaeQ_2_onehotd = 2'd0;
  assign es_14_8MyFalse_d = {vaeQ_2_d[32:1], vaeQ_2_onehotd[0]};
  assign _235_d = {vaeQ_2_d[32:1], vaeQ_2_onehotd[1]};
  assign vaeQ_2_r = (| (vaeQ_2_onehotd & {_235_r,
                                          es_14_8MyFalse_r}));
  assign es_14_8_r = vaeQ_2_r;
  
  /* buf (Ty QTree_Int) : (es_15_1QVal_Int,QTree_Int) > (lizzieLet36_1_argbuf,QTree_Int) */
  QTree_Int_t es_15_1QVal_Int_bufchan_d;
  logic es_15_1QVal_Int_bufchan_r;
  assign es_15_1QVal_Int_r = ((! es_15_1QVal_Int_bufchan_d[0]) || es_15_1QVal_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_15_1QVal_Int_bufchan_d <= {66'd0, 1'd0};
    else
      if (es_15_1QVal_Int_r)
        es_15_1QVal_Int_bufchan_d <= es_15_1QVal_Int_d;
  QTree_Int_t es_15_1QVal_Int_bufchan_buf;
  assign es_15_1QVal_Int_bufchan_r = (! es_15_1QVal_Int_bufchan_buf[0]);
  assign lizzieLet36_1_argbuf_d = (es_15_1QVal_Int_bufchan_buf[0] ? es_15_1QVal_Int_bufchan_buf :
                                   es_15_1QVal_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_15_1QVal_Int_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((lizzieLet36_1_argbuf_r && es_15_1QVal_Int_bufchan_buf[0]))
        es_15_1QVal_Int_bufchan_buf <= {66'd0, 1'd0};
      else if (((! lizzieLet36_1_argbuf_r) && (! es_15_1QVal_Int_bufchan_buf[0])))
        es_15_1QVal_Int_bufchan_buf <= es_15_1QVal_Int_bufchan_d;
  
  /* demux (Ty MyBool,
       Ty Int) : (es_21_1,MyBool) (es_14_6MyFalse_3QVal_Int_2,Int) > [(es_21_1MyFalse,Int),
                                                                      (_234,Int)] */
  logic [1:0] es_14_6MyFalse_3QVal_Int_2_onehotd;
  always_comb
    if ((es_21_1_d[0] && es_14_6MyFalse_3QVal_Int_2_d[0]))
      unique case (es_21_1_d[1:1])
        1'd0: es_14_6MyFalse_3QVal_Int_2_onehotd = 2'd1;
        1'd1: es_14_6MyFalse_3QVal_Int_2_onehotd = 2'd2;
        default: es_14_6MyFalse_3QVal_Int_2_onehotd = 2'd0;
      endcase
    else es_14_6MyFalse_3QVal_Int_2_onehotd = 2'd0;
  assign es_21_1MyFalse_d = {es_14_6MyFalse_3QVal_Int_2_d[32:1],
                             es_14_6MyFalse_3QVal_Int_2_onehotd[0]};
  assign _234_d = {es_14_6MyFalse_3QVal_Int_2_d[32:1],
                   es_14_6MyFalse_3QVal_Int_2_onehotd[1]};
  assign es_14_6MyFalse_3QVal_Int_2_r = (| (es_14_6MyFalse_3QVal_Int_2_onehotd & {_234_r,
                                                                                  es_21_1MyFalse_r}));
  assign es_21_1_r = es_14_6MyFalse_3QVal_Int_2_r;
  
  /* buf (Ty Int) : (es_21_1MyFalse,Int) > (es_21_1MyFalse_1_argbuf,Int) */
  Int_t es_21_1MyFalse_bufchan_d;
  logic es_21_1MyFalse_bufchan_r;
  assign es_21_1MyFalse_r = ((! es_21_1MyFalse_bufchan_d[0]) || es_21_1MyFalse_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_21_1MyFalse_bufchan_d <= {32'd0, 1'd0};
    else
      if (es_21_1MyFalse_r) es_21_1MyFalse_bufchan_d <= es_21_1MyFalse_d;
  Int_t es_21_1MyFalse_bufchan_buf;
  assign es_21_1MyFalse_bufchan_r = (! es_21_1MyFalse_bufchan_buf[0]);
  assign es_21_1MyFalse_1_argbuf_d = (es_21_1MyFalse_bufchan_buf[0] ? es_21_1MyFalse_bufchan_buf :
                                      es_21_1MyFalse_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_21_1MyFalse_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((es_21_1MyFalse_1_argbuf_r && es_21_1MyFalse_bufchan_buf[0]))
        es_21_1MyFalse_bufchan_buf <= {32'd0, 1'd0};
      else if (((! es_21_1MyFalse_1_argbuf_r) && (! es_21_1MyFalse_bufchan_buf[0])))
        es_21_1MyFalse_bufchan_buf <= es_21_1MyFalse_bufchan_d;
  
  /* demux (Ty MyBool,
       Ty MyDTInt_Int_Int) : (es_21_2,MyBool) (es_14_6MyFalse_4QVal_Int_3,MyDTInt_Int_Int) > [(es_21_2MyFalse,MyDTInt_Int_Int),
                                                                                              (_233,MyDTInt_Int_Int)] */
  logic [1:0] es_14_6MyFalse_4QVal_Int_3_onehotd;
  always_comb
    if ((es_21_2_d[0] && es_14_6MyFalse_4QVal_Int_3_d[0]))
      unique case (es_21_2_d[1:1])
        1'd0: es_14_6MyFalse_4QVal_Int_3_onehotd = 2'd1;
        1'd1: es_14_6MyFalse_4QVal_Int_3_onehotd = 2'd2;
        default: es_14_6MyFalse_4QVal_Int_3_onehotd = 2'd0;
      endcase
    else es_14_6MyFalse_4QVal_Int_3_onehotd = 2'd0;
  assign es_21_2MyFalse_d = es_14_6MyFalse_4QVal_Int_3_onehotd[0];
  assign _233_d = es_14_6MyFalse_4QVal_Int_3_onehotd[1];
  assign es_14_6MyFalse_4QVal_Int_3_r = (| (es_14_6MyFalse_4QVal_Int_3_onehotd & {_233_r,
                                                                                  es_21_2MyFalse_r}));
  assign es_21_2_r = es_14_6MyFalse_4QVal_Int_3_r;
  
  /* fork (Ty MyDTInt_Int_Int) : (es_21_2MyFalse,MyDTInt_Int_Int) > [(es_21_2MyFalse_1,MyDTInt_Int_Int),
                                                                (es_21_2MyFalse_2,MyDTInt_Int_Int)] */
  logic [1:0] es_21_2MyFalse_emitted;
  logic [1:0] es_21_2MyFalse_done;
  assign es_21_2MyFalse_1_d = (es_21_2MyFalse_d[0] && (! es_21_2MyFalse_emitted[0]));
  assign es_21_2MyFalse_2_d = (es_21_2MyFalse_d[0] && (! es_21_2MyFalse_emitted[1]));
  assign es_21_2MyFalse_done = (es_21_2MyFalse_emitted | ({es_21_2MyFalse_2_d[0],
                                                           es_21_2MyFalse_1_d[0]} & {es_21_2MyFalse_2_r,
                                                                                     es_21_2MyFalse_1_r}));
  assign es_21_2MyFalse_r = (& es_21_2MyFalse_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_21_2MyFalse_emitted <= 2'd0;
    else
      es_21_2MyFalse_emitted <= (es_21_2MyFalse_r ? 2'd0 :
                                 es_21_2MyFalse_done);
  
  /* buf (Ty MyDTInt_Int_Int) : (es_21_2MyFalse_1,MyDTInt_Int_Int) > (es_21_2MyFalse_1_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t es_21_2MyFalse_1_bufchan_d;
  logic es_21_2MyFalse_1_bufchan_r;
  assign es_21_2MyFalse_1_r = ((! es_21_2MyFalse_1_bufchan_d[0]) || es_21_2MyFalse_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_21_2MyFalse_1_bufchan_d <= 1'd0;
    else
      if (es_21_2MyFalse_1_r)
        es_21_2MyFalse_1_bufchan_d <= es_21_2MyFalse_1_d;
  MyDTInt_Int_Int_t es_21_2MyFalse_1_bufchan_buf;
  assign es_21_2MyFalse_1_bufchan_r = (! es_21_2MyFalse_1_bufchan_buf[0]);
  assign es_21_2MyFalse_1_argbuf_d = (es_21_2MyFalse_1_bufchan_buf[0] ? es_21_2MyFalse_1_bufchan_buf :
                                      es_21_2MyFalse_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_21_2MyFalse_1_bufchan_buf <= 1'd0;
    else
      if ((es_21_2MyFalse_1_argbuf_r && es_21_2MyFalse_1_bufchan_buf[0]))
        es_21_2MyFalse_1_bufchan_buf <= 1'd0;
      else if (((! es_21_2MyFalse_1_argbuf_r) && (! es_21_2MyFalse_1_bufchan_buf[0])))
        es_21_2MyFalse_1_bufchan_buf <= es_21_2MyFalse_1_bufchan_d;
  
  /* dcon (Ty TupMyDTInt_Int_Int___Int___Int,
      Dcon TupMyDTInt_Int_Int___Int___Int) : [(es_21_2MyFalse_1_argbuf,MyDTInt_Int_Int),
                                              (es_21_1MyFalse_1_argbuf,Int),
                                              (es_21_5MyFalse_1_argbuf,Int)] > (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int11,TupMyDTInt_Int_Int___Int___Int) */
  assign applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int11_d = TupMyDTInt_Int_Int___Int___Int_dc((& {es_21_2MyFalse_1_argbuf_d[0],
                                                                                                        es_21_1MyFalse_1_argbuf_d[0],
                                                                                                        es_21_5MyFalse_1_argbuf_d[0]}), es_21_2MyFalse_1_argbuf_d, es_21_1MyFalse_1_argbuf_d, es_21_5MyFalse_1_argbuf_d);
  assign {es_21_2MyFalse_1_argbuf_r,
          es_21_1MyFalse_1_argbuf_r,
          es_21_5MyFalse_1_argbuf_r} = {3 {(applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int11_r && applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int11_d[0])}};
  
  /* buf (Ty MyDTInt_Int_Int) : (es_21_2MyFalse_2,MyDTInt_Int_Int) > (es_21_2MyFalse_2_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t es_21_2MyFalse_2_bufchan_d;
  logic es_21_2MyFalse_2_bufchan_r;
  assign es_21_2MyFalse_2_r = ((! es_21_2MyFalse_2_bufchan_d[0]) || es_21_2MyFalse_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_21_2MyFalse_2_bufchan_d <= 1'd0;
    else
      if (es_21_2MyFalse_2_r)
        es_21_2MyFalse_2_bufchan_d <= es_21_2MyFalse_2_d;
  MyDTInt_Int_Int_t es_21_2MyFalse_2_bufchan_buf;
  assign es_21_2MyFalse_2_bufchan_r = (! es_21_2MyFalse_2_bufchan_buf[0]);
  assign es_21_2MyFalse_2_argbuf_d = (es_21_2MyFalse_2_bufchan_buf[0] ? es_21_2MyFalse_2_bufchan_buf :
                                      es_21_2MyFalse_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_21_2MyFalse_2_bufchan_buf <= 1'd0;
    else
      if ((es_21_2MyFalse_2_argbuf_r && es_21_2MyFalse_2_bufchan_buf[0]))
        es_21_2MyFalse_2_bufchan_buf <= 1'd0;
      else if (((! es_21_2MyFalse_2_argbuf_r) && (! es_21_2MyFalse_2_bufchan_buf[0])))
        es_21_2MyFalse_2_bufchan_buf <= es_21_2MyFalse_2_bufchan_d;
  
  /* dcon (Ty TupMyDTInt_Int_Int___Int___Int,
      Dcon TupMyDTInt_Int_Int___Int___Int) : [(es_21_2MyFalse_2_argbuf,MyDTInt_Int_Int),
                                              (es_24_1_argbuf,Int),
                                              (es_21_6MyFalse_1_argbuf,Int)] > (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int12,TupMyDTInt_Int_Int___Int___Int) */
  assign applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int12_d = TupMyDTInt_Int_Int___Int___Int_dc((& {es_21_2MyFalse_2_argbuf_d[0],
                                                                                                        es_24_1_argbuf_d[0],
                                                                                                        es_21_6MyFalse_1_argbuf_d[0]}), es_21_2MyFalse_2_argbuf_d, es_24_1_argbuf_d, es_21_6MyFalse_1_argbuf_d);
  assign {es_21_2MyFalse_2_argbuf_r,
          es_24_1_argbuf_r,
          es_21_6MyFalse_1_argbuf_r} = {3 {(applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int12_r && applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int12_d[0])}};
  
  /* demux (Ty MyBool,
       Ty Pointer_CTf_f_Int) : (es_21_3,MyBool) (es_14_6MyFalse_5QVal_Int,Pointer_CTf_f_Int) > [(es_21_3MyFalse,Pointer_CTf_f_Int),
                                                                                                (es_21_3MyTrue,Pointer_CTf_f_Int)] */
  logic [1:0] es_14_6MyFalse_5QVal_Int_onehotd;
  always_comb
    if ((es_21_3_d[0] && es_14_6MyFalse_5QVal_Int_d[0]))
      unique case (es_21_3_d[1:1])
        1'd0: es_14_6MyFalse_5QVal_Int_onehotd = 2'd1;
        1'd1: es_14_6MyFalse_5QVal_Int_onehotd = 2'd2;
        default: es_14_6MyFalse_5QVal_Int_onehotd = 2'd0;
      endcase
    else es_14_6MyFalse_5QVal_Int_onehotd = 2'd0;
  assign es_21_3MyFalse_d = {es_14_6MyFalse_5QVal_Int_d[16:1],
                             es_14_6MyFalse_5QVal_Int_onehotd[0]};
  assign es_21_3MyTrue_d = {es_14_6MyFalse_5QVal_Int_d[16:1],
                            es_14_6MyFalse_5QVal_Int_onehotd[1]};
  assign es_14_6MyFalse_5QVal_Int_r = (| (es_14_6MyFalse_5QVal_Int_onehotd & {es_21_3MyTrue_r,
                                                                              es_21_3MyFalse_r}));
  assign es_21_3_r = es_14_6MyFalse_5QVal_Int_r;
  
  /* buf (Ty Pointer_CTf_f_Int) : (es_21_3MyFalse,Pointer_CTf_f_Int) > (es_21_3MyFalse_1_argbuf,Pointer_CTf_f_Int) */
  Pointer_CTf_f_Int_t es_21_3MyFalse_bufchan_d;
  logic es_21_3MyFalse_bufchan_r;
  assign es_21_3MyFalse_r = ((! es_21_3MyFalse_bufchan_d[0]) || es_21_3MyFalse_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_21_3MyFalse_bufchan_d <= {16'd0, 1'd0};
    else
      if (es_21_3MyFalse_r) es_21_3MyFalse_bufchan_d <= es_21_3MyFalse_d;
  Pointer_CTf_f_Int_t es_21_3MyFalse_bufchan_buf;
  assign es_21_3MyFalse_bufchan_r = (! es_21_3MyFalse_bufchan_buf[0]);
  assign es_21_3MyFalse_1_argbuf_d = (es_21_3MyFalse_bufchan_buf[0] ? es_21_3MyFalse_bufchan_buf :
                                      es_21_3MyFalse_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_21_3MyFalse_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((es_21_3MyFalse_1_argbuf_r && es_21_3MyFalse_bufchan_buf[0]))
        es_21_3MyFalse_bufchan_buf <= {16'd0, 1'd0};
      else if (((! es_21_3MyFalse_1_argbuf_r) && (! es_21_3MyFalse_bufchan_buf[0])))
        es_21_3MyFalse_bufchan_buf <= es_21_3MyFalse_bufchan_d;
  
  /* buf (Ty Pointer_CTf_f_Int) : (es_21_3MyTrue,Pointer_CTf_f_Int) > (es_21_3MyTrue_1_argbuf,Pointer_CTf_f_Int) */
  Pointer_CTf_f_Int_t es_21_3MyTrue_bufchan_d;
  logic es_21_3MyTrue_bufchan_r;
  assign es_21_3MyTrue_r = ((! es_21_3MyTrue_bufchan_d[0]) || es_21_3MyTrue_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_21_3MyTrue_bufchan_d <= {16'd0, 1'd0};
    else
      if (es_21_3MyTrue_r) es_21_3MyTrue_bufchan_d <= es_21_3MyTrue_d;
  Pointer_CTf_f_Int_t es_21_3MyTrue_bufchan_buf;
  assign es_21_3MyTrue_bufchan_r = (! es_21_3MyTrue_bufchan_buf[0]);
  assign es_21_3MyTrue_1_argbuf_d = (es_21_3MyTrue_bufchan_buf[0] ? es_21_3MyTrue_bufchan_buf :
                                     es_21_3MyTrue_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_21_3MyTrue_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((es_21_3MyTrue_1_argbuf_r && es_21_3MyTrue_bufchan_buf[0]))
        es_21_3MyTrue_bufchan_buf <= {16'd0, 1'd0};
      else if (((! es_21_3MyTrue_1_argbuf_r) && (! es_21_3MyTrue_bufchan_buf[0])))
        es_21_3MyTrue_bufchan_buf <= es_21_3MyTrue_bufchan_d;
  
  /* demux (Ty MyBool,
       Ty Go) : (es_21_4,MyBool) (es_14_6MyFalse_6QVal_Int_2,Go) > [(es_21_4MyFalse,Go),
                                                                    (es_21_4MyTrue,Go)] */
  logic [1:0] es_14_6MyFalse_6QVal_Int_2_onehotd;
  always_comb
    if ((es_21_4_d[0] && es_14_6MyFalse_6QVal_Int_2_d[0]))
      unique case (es_21_4_d[1:1])
        1'd0: es_14_6MyFalse_6QVal_Int_2_onehotd = 2'd1;
        1'd1: es_14_6MyFalse_6QVal_Int_2_onehotd = 2'd2;
        default: es_14_6MyFalse_6QVal_Int_2_onehotd = 2'd0;
      endcase
    else es_14_6MyFalse_6QVal_Int_2_onehotd = 2'd0;
  assign es_21_4MyFalse_d = es_14_6MyFalse_6QVal_Int_2_onehotd[0];
  assign es_21_4MyTrue_d = es_14_6MyFalse_6QVal_Int_2_onehotd[1];
  assign es_14_6MyFalse_6QVal_Int_2_r = (| (es_14_6MyFalse_6QVal_Int_2_onehotd & {es_21_4MyTrue_r,
                                                                                  es_21_4MyFalse_r}));
  assign es_21_4_r = es_14_6MyFalse_6QVal_Int_2_r;
  
  /* buf (Ty Go) : (es_21_4MyFalse,Go) > (es_21_4MyFalse_1_argbuf,Go) */
  Go_t es_21_4MyFalse_bufchan_d;
  logic es_21_4MyFalse_bufchan_r;
  assign es_21_4MyFalse_r = ((! es_21_4MyFalse_bufchan_d[0]) || es_21_4MyFalse_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_21_4MyFalse_bufchan_d <= 1'd0;
    else
      if (es_21_4MyFalse_r) es_21_4MyFalse_bufchan_d <= es_21_4MyFalse_d;
  Go_t es_21_4MyFalse_bufchan_buf;
  assign es_21_4MyFalse_bufchan_r = (! es_21_4MyFalse_bufchan_buf[0]);
  assign es_21_4MyFalse_1_argbuf_d = (es_21_4MyFalse_bufchan_buf[0] ? es_21_4MyFalse_bufchan_buf :
                                      es_21_4MyFalse_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_21_4MyFalse_bufchan_buf <= 1'd0;
    else
      if ((es_21_4MyFalse_1_argbuf_r && es_21_4MyFalse_bufchan_buf[0]))
        es_21_4MyFalse_bufchan_buf <= 1'd0;
      else if (((! es_21_4MyFalse_1_argbuf_r) && (! es_21_4MyFalse_bufchan_buf[0])))
        es_21_4MyFalse_bufchan_buf <= es_21_4MyFalse_bufchan_d;
  
  /* fork (Ty Go) : (es_21_4MyTrue,Go) > [(es_21_4MyTrue_1,Go),
                                     (es_21_4MyTrue_2,Go)] */
  logic [1:0] es_21_4MyTrue_emitted;
  logic [1:0] es_21_4MyTrue_done;
  assign es_21_4MyTrue_1_d = (es_21_4MyTrue_d[0] && (! es_21_4MyTrue_emitted[0]));
  assign es_21_4MyTrue_2_d = (es_21_4MyTrue_d[0] && (! es_21_4MyTrue_emitted[1]));
  assign es_21_4MyTrue_done = (es_21_4MyTrue_emitted | ({es_21_4MyTrue_2_d[0],
                                                         es_21_4MyTrue_1_d[0]} & {es_21_4MyTrue_2_r,
                                                                                  es_21_4MyTrue_1_r}));
  assign es_21_4MyTrue_r = (& es_21_4MyTrue_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_21_4MyTrue_emitted <= 2'd0;
    else
      es_21_4MyTrue_emitted <= (es_21_4MyTrue_r ? 2'd0 :
                                es_21_4MyTrue_done);
  
  /* dcon (Ty QTree_Int,
      Dcon QNone_Int) : [(es_21_4MyTrue_1,Go)] > (es_21_4MyTrue_1QNone_Int,QTree_Int) */
  assign es_21_4MyTrue_1QNone_Int_d = QNone_Int_dc((& {es_21_4MyTrue_1_d[0]}), es_21_4MyTrue_1_d);
  assign {es_21_4MyTrue_1_r} = {1 {(es_21_4MyTrue_1QNone_Int_r && es_21_4MyTrue_1QNone_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (es_21_4MyTrue_1QNone_Int,QTree_Int) > (lizzieLet38_1_1_argbuf,QTree_Int) */
  QTree_Int_t es_21_4MyTrue_1QNone_Int_bufchan_d;
  logic es_21_4MyTrue_1QNone_Int_bufchan_r;
  assign es_21_4MyTrue_1QNone_Int_r = ((! es_21_4MyTrue_1QNone_Int_bufchan_d[0]) || es_21_4MyTrue_1QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_21_4MyTrue_1QNone_Int_bufchan_d <= {66'd0, 1'd0};
    else
      if (es_21_4MyTrue_1QNone_Int_r)
        es_21_4MyTrue_1QNone_Int_bufchan_d <= es_21_4MyTrue_1QNone_Int_d;
  QTree_Int_t es_21_4MyTrue_1QNone_Int_bufchan_buf;
  assign es_21_4MyTrue_1QNone_Int_bufchan_r = (! es_21_4MyTrue_1QNone_Int_bufchan_buf[0]);
  assign lizzieLet38_1_1_argbuf_d = (es_21_4MyTrue_1QNone_Int_bufchan_buf[0] ? es_21_4MyTrue_1QNone_Int_bufchan_buf :
                                     es_21_4MyTrue_1QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_21_4MyTrue_1QNone_Int_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((lizzieLet38_1_1_argbuf_r && es_21_4MyTrue_1QNone_Int_bufchan_buf[0]))
        es_21_4MyTrue_1QNone_Int_bufchan_buf <= {66'd0, 1'd0};
      else if (((! lizzieLet38_1_1_argbuf_r) && (! es_21_4MyTrue_1QNone_Int_bufchan_buf[0])))
        es_21_4MyTrue_1QNone_Int_bufchan_buf <= es_21_4MyTrue_1QNone_Int_bufchan_d;
  
  /* buf (Ty Go) : (es_21_4MyTrue_2,Go) > (es_21_4MyTrue_2_argbuf,Go) */
  Go_t es_21_4MyTrue_2_bufchan_d;
  logic es_21_4MyTrue_2_bufchan_r;
  assign es_21_4MyTrue_2_r = ((! es_21_4MyTrue_2_bufchan_d[0]) || es_21_4MyTrue_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_21_4MyTrue_2_bufchan_d <= 1'd0;
    else
      if (es_21_4MyTrue_2_r)
        es_21_4MyTrue_2_bufchan_d <= es_21_4MyTrue_2_d;
  Go_t es_21_4MyTrue_2_bufchan_buf;
  assign es_21_4MyTrue_2_bufchan_r = (! es_21_4MyTrue_2_bufchan_buf[0]);
  assign es_21_4MyTrue_2_argbuf_d = (es_21_4MyTrue_2_bufchan_buf[0] ? es_21_4MyTrue_2_bufchan_buf :
                                     es_21_4MyTrue_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_21_4MyTrue_2_bufchan_buf <= 1'd0;
    else
      if ((es_21_4MyTrue_2_argbuf_r && es_21_4MyTrue_2_bufchan_buf[0]))
        es_21_4MyTrue_2_bufchan_buf <= 1'd0;
      else if (((! es_21_4MyTrue_2_argbuf_r) && (! es_21_4MyTrue_2_bufchan_buf[0])))
        es_21_4MyTrue_2_bufchan_buf <= es_21_4MyTrue_2_bufchan_d;
  
  /* demux (Ty MyBool,
       Ty Int) : (es_21_5,MyBool) (es_14_6MyFalse_8QVal_Int_2,Int) > [(es_21_5MyFalse,Int),
                                                                      (_232,Int)] */
  logic [1:0] es_14_6MyFalse_8QVal_Int_2_onehotd;
  always_comb
    if ((es_21_5_d[0] && es_14_6MyFalse_8QVal_Int_2_d[0]))
      unique case (es_21_5_d[1:1])
        1'd0: es_14_6MyFalse_8QVal_Int_2_onehotd = 2'd1;
        1'd1: es_14_6MyFalse_8QVal_Int_2_onehotd = 2'd2;
        default: es_14_6MyFalse_8QVal_Int_2_onehotd = 2'd0;
      endcase
    else es_14_6MyFalse_8QVal_Int_2_onehotd = 2'd0;
  assign es_21_5MyFalse_d = {es_14_6MyFalse_8QVal_Int_2_d[32:1],
                             es_14_6MyFalse_8QVal_Int_2_onehotd[0]};
  assign _232_d = {es_14_6MyFalse_8QVal_Int_2_d[32:1],
                   es_14_6MyFalse_8QVal_Int_2_onehotd[1]};
  assign es_14_6MyFalse_8QVal_Int_2_r = (| (es_14_6MyFalse_8QVal_Int_2_onehotd & {_232_r,
                                                                                  es_21_5MyFalse_r}));
  assign es_21_5_r = es_14_6MyFalse_8QVal_Int_2_r;
  
  /* buf (Ty Int) : (es_21_5MyFalse,Int) > (es_21_5MyFalse_1_argbuf,Int) */
  Int_t es_21_5MyFalse_bufchan_d;
  logic es_21_5MyFalse_bufchan_r;
  assign es_21_5MyFalse_r = ((! es_21_5MyFalse_bufchan_d[0]) || es_21_5MyFalse_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_21_5MyFalse_bufchan_d <= {32'd0, 1'd0};
    else
      if (es_21_5MyFalse_r) es_21_5MyFalse_bufchan_d <= es_21_5MyFalse_d;
  Int_t es_21_5MyFalse_bufchan_buf;
  assign es_21_5MyFalse_bufchan_r = (! es_21_5MyFalse_bufchan_buf[0]);
  assign es_21_5MyFalse_1_argbuf_d = (es_21_5MyFalse_bufchan_buf[0] ? es_21_5MyFalse_bufchan_buf :
                                      es_21_5MyFalse_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_21_5MyFalse_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((es_21_5MyFalse_1_argbuf_r && es_21_5MyFalse_bufchan_buf[0]))
        es_21_5MyFalse_bufchan_buf <= {32'd0, 1'd0};
      else if (((! es_21_5MyFalse_1_argbuf_r) && (! es_21_5MyFalse_bufchan_buf[0])))
        es_21_5MyFalse_bufchan_buf <= es_21_5MyFalse_bufchan_d;
  
  /* demux (Ty MyBool,
       Ty Int) : (es_21_6,MyBool) (v'aeR_2,Int) > [(es_21_6MyFalse,Int),
                                                   (_231,Int)] */
  logic [1:0] \v'aeR_2_onehotd ;
  always_comb
    if ((es_21_6_d[0] && \v'aeR_2_d [0]))
      unique case (es_21_6_d[1:1])
        1'd0: \v'aeR_2_onehotd  = 2'd1;
        1'd1: \v'aeR_2_onehotd  = 2'd2;
        default: \v'aeR_2_onehotd  = 2'd0;
      endcase
    else \v'aeR_2_onehotd  = 2'd0;
  assign es_21_6MyFalse_d = {\v'aeR_2_d [32:1],
                             \v'aeR_2_onehotd [0]};
  assign _231_d = {\v'aeR_2_d [32:1], \v'aeR_2_onehotd [1]};
  assign \v'aeR_2_r  = (| (\v'aeR_2_onehotd  & {_231_r,
                                                es_21_6MyFalse_r}));
  assign es_21_6_r = \v'aeR_2_r ;
  
  /* buf (Ty Int) : (es_21_6MyFalse,Int) > (es_21_6MyFalse_1_argbuf,Int) */
  Int_t es_21_6MyFalse_bufchan_d;
  logic es_21_6MyFalse_bufchan_r;
  assign es_21_6MyFalse_r = ((! es_21_6MyFalse_bufchan_d[0]) || es_21_6MyFalse_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_21_6MyFalse_bufchan_d <= {32'd0, 1'd0};
    else
      if (es_21_6MyFalse_r) es_21_6MyFalse_bufchan_d <= es_21_6MyFalse_d;
  Int_t es_21_6MyFalse_bufchan_buf;
  assign es_21_6MyFalse_bufchan_r = (! es_21_6MyFalse_bufchan_buf[0]);
  assign es_21_6MyFalse_1_argbuf_d = (es_21_6MyFalse_bufchan_buf[0] ? es_21_6MyFalse_bufchan_buf :
                                      es_21_6MyFalse_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_21_6MyFalse_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((es_21_6MyFalse_1_argbuf_r && es_21_6MyFalse_bufchan_buf[0]))
        es_21_6MyFalse_bufchan_buf <= {32'd0, 1'd0};
      else if (((! es_21_6MyFalse_1_argbuf_r) && (! es_21_6MyFalse_bufchan_buf[0])))
        es_21_6MyFalse_bufchan_buf <= es_21_6MyFalse_bufchan_d;
  
  /* buf (Ty QTree_Int) : (es_22_1QVal_Int,QTree_Int) > (lizzieLet37_2_1_argbuf,QTree_Int) */
  QTree_Int_t es_22_1QVal_Int_bufchan_d;
  logic es_22_1QVal_Int_bufchan_r;
  assign es_22_1QVal_Int_r = ((! es_22_1QVal_Int_bufchan_d[0]) || es_22_1QVal_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_22_1QVal_Int_bufchan_d <= {66'd0, 1'd0};
    else
      if (es_22_1QVal_Int_r)
        es_22_1QVal_Int_bufchan_d <= es_22_1QVal_Int_d;
  QTree_Int_t es_22_1QVal_Int_bufchan_buf;
  assign es_22_1QVal_Int_bufchan_r = (! es_22_1QVal_Int_bufchan_buf[0]);
  assign lizzieLet37_2_1_argbuf_d = (es_22_1QVal_Int_bufchan_buf[0] ? es_22_1QVal_Int_bufchan_buf :
                                     es_22_1QVal_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_22_1QVal_Int_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((lizzieLet37_2_1_argbuf_r && es_22_1QVal_Int_bufchan_buf[0]))
        es_22_1QVal_Int_bufchan_buf <= {66'd0, 1'd0};
      else if (((! lizzieLet37_2_1_argbuf_r) && (! es_22_1QVal_Int_bufchan_buf[0])))
        es_22_1QVal_Int_bufchan_buf <= es_22_1QVal_Int_bufchan_d;
  
  /* buf (Ty QTree_Int) : (es_26_1es_27_1es_28_1es_29_1QNode_Int,QTree_Int) > (lizzieLet46_1_argbuf,QTree_Int) */
  QTree_Int_t es_26_1es_27_1es_28_1es_29_1QNode_Int_bufchan_d;
  logic es_26_1es_27_1es_28_1es_29_1QNode_Int_bufchan_r;
  assign es_26_1es_27_1es_28_1es_29_1QNode_Int_r = ((! es_26_1es_27_1es_28_1es_29_1QNode_Int_bufchan_d[0]) || es_26_1es_27_1es_28_1es_29_1QNode_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_26_1es_27_1es_28_1es_29_1QNode_Int_bufchan_d <= {66'd0, 1'd0};
    else
      if (es_26_1es_27_1es_28_1es_29_1QNode_Int_r)
        es_26_1es_27_1es_28_1es_29_1QNode_Int_bufchan_d <= es_26_1es_27_1es_28_1es_29_1QNode_Int_d;
  QTree_Int_t es_26_1es_27_1es_28_1es_29_1QNode_Int_bufchan_buf;
  assign es_26_1es_27_1es_28_1es_29_1QNode_Int_bufchan_r = (! es_26_1es_27_1es_28_1es_29_1QNode_Int_bufchan_buf[0]);
  assign lizzieLet46_1_argbuf_d = (es_26_1es_27_1es_28_1es_29_1QNode_Int_bufchan_buf[0] ? es_26_1es_27_1es_28_1es_29_1QNode_Int_bufchan_buf :
                                   es_26_1es_27_1es_28_1es_29_1QNode_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_26_1es_27_1es_28_1es_29_1QNode_Int_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((lizzieLet46_1_argbuf_r && es_26_1es_27_1es_28_1es_29_1QNode_Int_bufchan_buf[0]))
        es_26_1es_27_1es_28_1es_29_1QNode_Int_bufchan_buf <= {66'd0, 1'd0};
      else if (((! lizzieLet46_1_argbuf_r) && (! es_26_1es_27_1es_28_1es_29_1QNode_Int_bufchan_buf[0])))
        es_26_1es_27_1es_28_1es_29_1QNode_Int_bufchan_buf <= es_26_1es_27_1es_28_1es_29_1QNode_Int_bufchan_d;
  
  /* demux (Ty MyBool,
       Ty Go) : (es_2_1,MyBool) (lizzieLet6_5QVal_Int_3QVal_Int_2,Go) > [(es_2_1MyFalse,Go),
                                                                         (es_2_1MyTrue,Go)] */
  logic [1:0] lizzieLet6_5QVal_Int_3QVal_Int_2_onehotd;
  always_comb
    if ((es_2_1_d[0] && lizzieLet6_5QVal_Int_3QVal_Int_2_d[0]))
      unique case (es_2_1_d[1:1])
        1'd0: lizzieLet6_5QVal_Int_3QVal_Int_2_onehotd = 2'd1;
        1'd1: lizzieLet6_5QVal_Int_3QVal_Int_2_onehotd = 2'd2;
        default: lizzieLet6_5QVal_Int_3QVal_Int_2_onehotd = 2'd0;
      endcase
    else lizzieLet6_5QVal_Int_3QVal_Int_2_onehotd = 2'd0;
  assign es_2_1MyFalse_d = lizzieLet6_5QVal_Int_3QVal_Int_2_onehotd[0];
  assign es_2_1MyTrue_d = lizzieLet6_5QVal_Int_3QVal_Int_2_onehotd[1];
  assign lizzieLet6_5QVal_Int_3QVal_Int_2_r = (| (lizzieLet6_5QVal_Int_3QVal_Int_2_onehotd & {es_2_1MyTrue_r,
                                                                                              es_2_1MyFalse_r}));
  assign es_2_1_r = lizzieLet6_5QVal_Int_3QVal_Int_2_r;
  
  /* buf (Ty Go) : (es_2_1MyFalse,Go) > (es_2_1MyFalse_1_argbuf,Go) */
  Go_t es_2_1MyFalse_bufchan_d;
  logic es_2_1MyFalse_bufchan_r;
  assign es_2_1MyFalse_r = ((! es_2_1MyFalse_bufchan_d[0]) || es_2_1MyFalse_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_2_1MyFalse_bufchan_d <= 1'd0;
    else
      if (es_2_1MyFalse_r) es_2_1MyFalse_bufchan_d <= es_2_1MyFalse_d;
  Go_t es_2_1MyFalse_bufchan_buf;
  assign es_2_1MyFalse_bufchan_r = (! es_2_1MyFalse_bufchan_buf[0]);
  assign es_2_1MyFalse_1_argbuf_d = (es_2_1MyFalse_bufchan_buf[0] ? es_2_1MyFalse_bufchan_buf :
                                     es_2_1MyFalse_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_2_1MyFalse_bufchan_buf <= 1'd0;
    else
      if ((es_2_1MyFalse_1_argbuf_r && es_2_1MyFalse_bufchan_buf[0]))
        es_2_1MyFalse_bufchan_buf <= 1'd0;
      else if (((! es_2_1MyFalse_1_argbuf_r) && (! es_2_1MyFalse_bufchan_buf[0])))
        es_2_1MyFalse_bufchan_buf <= es_2_1MyFalse_bufchan_d;
  
  /* fork (Ty Go) : (es_2_1MyTrue,Go) > [(es_2_1MyTrue_1,Go),
                                    (es_2_1MyTrue_2,Go)] */
  logic [1:0] es_2_1MyTrue_emitted;
  logic [1:0] es_2_1MyTrue_done;
  assign es_2_1MyTrue_1_d = (es_2_1MyTrue_d[0] && (! es_2_1MyTrue_emitted[0]));
  assign es_2_1MyTrue_2_d = (es_2_1MyTrue_d[0] && (! es_2_1MyTrue_emitted[1]));
  assign es_2_1MyTrue_done = (es_2_1MyTrue_emitted | ({es_2_1MyTrue_2_d[0],
                                                       es_2_1MyTrue_1_d[0]} & {es_2_1MyTrue_2_r,
                                                                               es_2_1MyTrue_1_r}));
  assign es_2_1MyTrue_r = (& es_2_1MyTrue_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_2_1MyTrue_emitted <= 2'd0;
    else
      es_2_1MyTrue_emitted <= (es_2_1MyTrue_r ? 2'd0 :
                               es_2_1MyTrue_done);
  
  /* dcon (Ty QTree_Int,
      Dcon QNone_Int) : [(es_2_1MyTrue_1,Go)] > (es_2_1MyTrue_1QNone_Int,QTree_Int) */
  assign es_2_1MyTrue_1QNone_Int_d = QNone_Int_dc((& {es_2_1MyTrue_1_d[0]}), es_2_1MyTrue_1_d);
  assign {es_2_1MyTrue_1_r} = {1 {(es_2_1MyTrue_1QNone_Int_r && es_2_1MyTrue_1QNone_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (es_2_1MyTrue_1QNone_Int,QTree_Int) > (lizzieLet9_1_argbuf,QTree_Int) */
  QTree_Int_t es_2_1MyTrue_1QNone_Int_bufchan_d;
  logic es_2_1MyTrue_1QNone_Int_bufchan_r;
  assign es_2_1MyTrue_1QNone_Int_r = ((! es_2_1MyTrue_1QNone_Int_bufchan_d[0]) || es_2_1MyTrue_1QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_2_1MyTrue_1QNone_Int_bufchan_d <= {66'd0, 1'd0};
    else
      if (es_2_1MyTrue_1QNone_Int_r)
        es_2_1MyTrue_1QNone_Int_bufchan_d <= es_2_1MyTrue_1QNone_Int_d;
  QTree_Int_t es_2_1MyTrue_1QNone_Int_bufchan_buf;
  assign es_2_1MyTrue_1QNone_Int_bufchan_r = (! es_2_1MyTrue_1QNone_Int_bufchan_buf[0]);
  assign lizzieLet9_1_argbuf_d = (es_2_1MyTrue_1QNone_Int_bufchan_buf[0] ? es_2_1MyTrue_1QNone_Int_bufchan_buf :
                                  es_2_1MyTrue_1QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_2_1MyTrue_1QNone_Int_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((lizzieLet9_1_argbuf_r && es_2_1MyTrue_1QNone_Int_bufchan_buf[0]))
        es_2_1MyTrue_1QNone_Int_bufchan_buf <= {66'd0, 1'd0};
      else if (((! lizzieLet9_1_argbuf_r) && (! es_2_1MyTrue_1QNone_Int_bufchan_buf[0])))
        es_2_1MyTrue_1QNone_Int_bufchan_buf <= es_2_1MyTrue_1QNone_Int_bufchan_d;
  
  /* buf (Ty Go) : (es_2_1MyTrue_2,Go) > (es_2_1MyTrue_2_argbuf,Go) */
  Go_t es_2_1MyTrue_2_bufchan_d;
  logic es_2_1MyTrue_2_bufchan_r;
  assign es_2_1MyTrue_2_r = ((! es_2_1MyTrue_2_bufchan_d[0]) || es_2_1MyTrue_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_2_1MyTrue_2_bufchan_d <= 1'd0;
    else
      if (es_2_1MyTrue_2_r) es_2_1MyTrue_2_bufchan_d <= es_2_1MyTrue_2_d;
  Go_t es_2_1MyTrue_2_bufchan_buf;
  assign es_2_1MyTrue_2_bufchan_r = (! es_2_1MyTrue_2_bufchan_buf[0]);
  assign es_2_1MyTrue_2_argbuf_d = (es_2_1MyTrue_2_bufchan_buf[0] ? es_2_1MyTrue_2_bufchan_buf :
                                    es_2_1MyTrue_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_2_1MyTrue_2_bufchan_buf <= 1'd0;
    else
      if ((es_2_1MyTrue_2_argbuf_r && es_2_1MyTrue_2_bufchan_buf[0]))
        es_2_1MyTrue_2_bufchan_buf <= 1'd0;
      else if (((! es_2_1MyTrue_2_argbuf_r) && (! es_2_1MyTrue_2_bufchan_buf[0])))
        es_2_1MyTrue_2_bufchan_buf <= es_2_1MyTrue_2_bufchan_d;
  
  /* demux (Ty MyBool,
       Ty MyDTInt_Int_Int) : (es_2_1_1,MyBool) (lizzieLet17_5QNone_Int_7QVal_Int_3QVal_Int_2,MyDTInt_Int_Int) > [(es_2_1_1MyFalse,MyDTInt_Int_Int),
                                                                                                                 (_230,MyDTInt_Int_Int)] */
  logic [1:0] lizzieLet17_5QNone_Int_7QVal_Int_3QVal_Int_2_onehotd;
  always_comb
    if ((es_2_1_1_d[0] && lizzieLet17_5QNone_Int_7QVal_Int_3QVal_Int_2_d[0]))
      unique case (es_2_1_1_d[1:1])
        1'd0: lizzieLet17_5QNone_Int_7QVal_Int_3QVal_Int_2_onehotd = 2'd1;
        1'd1: lizzieLet17_5QNone_Int_7QVal_Int_3QVal_Int_2_onehotd = 2'd2;
        default:
          lizzieLet17_5QNone_Int_7QVal_Int_3QVal_Int_2_onehotd = 2'd0;
      endcase
    else lizzieLet17_5QNone_Int_7QVal_Int_3QVal_Int_2_onehotd = 2'd0;
  assign es_2_1_1MyFalse_d = lizzieLet17_5QNone_Int_7QVal_Int_3QVal_Int_2_onehotd[0];
  assign _230_d = lizzieLet17_5QNone_Int_7QVal_Int_3QVal_Int_2_onehotd[1];
  assign lizzieLet17_5QNone_Int_7QVal_Int_3QVal_Int_2_r = (| (lizzieLet17_5QNone_Int_7QVal_Int_3QVal_Int_2_onehotd & {_230_r,
                                                                                                                      es_2_1_1MyFalse_r}));
  assign es_2_1_1_r = lizzieLet17_5QNone_Int_7QVal_Int_3QVal_Int_2_r;
  
  /* buf (Ty MyDTInt_Int_Int) : (es_2_1_1MyFalse,MyDTInt_Int_Int) > (es_2_1_1MyFalse_1_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t es_2_1_1MyFalse_bufchan_d;
  logic es_2_1_1MyFalse_bufchan_r;
  assign es_2_1_1MyFalse_r = ((! es_2_1_1MyFalse_bufchan_d[0]) || es_2_1_1MyFalse_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_2_1_1MyFalse_bufchan_d <= 1'd0;
    else
      if (es_2_1_1MyFalse_r)
        es_2_1_1MyFalse_bufchan_d <= es_2_1_1MyFalse_d;
  MyDTInt_Int_Int_t es_2_1_1MyFalse_bufchan_buf;
  assign es_2_1_1MyFalse_bufchan_r = (! es_2_1_1MyFalse_bufchan_buf[0]);
  assign es_2_1_1MyFalse_1_argbuf_d = (es_2_1_1MyFalse_bufchan_buf[0] ? es_2_1_1MyFalse_bufchan_buf :
                                       es_2_1_1MyFalse_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_2_1_1MyFalse_bufchan_buf <= 1'd0;
    else
      if ((es_2_1_1MyFalse_1_argbuf_r && es_2_1_1MyFalse_bufchan_buf[0]))
        es_2_1_1MyFalse_bufchan_buf <= 1'd0;
      else if (((! es_2_1_1MyFalse_1_argbuf_r) && (! es_2_1_1MyFalse_bufchan_buf[0])))
        es_2_1_1MyFalse_bufchan_buf <= es_2_1_1MyFalse_bufchan_d;
  
  /* dcon (Ty TupMyDTInt_Int_Int___Int___Int,
      Dcon TupMyDTInt_Int_Int___Int___Int) : [(es_2_1_1MyFalse_1_argbuf,MyDTInt_Int_Int),
                                              (es_2_1_4MyFalse_1_argbuf,Int),
                                              (es_2_1_5MyFalse_1_argbuf,Int)] > (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int2,TupMyDTInt_Int_Int___Int___Int) */
  assign applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int2_d = TupMyDTInt_Int_Int___Int___Int_dc((& {es_2_1_1MyFalse_1_argbuf_d[0],
                                                                                                       es_2_1_4MyFalse_1_argbuf_d[0],
                                                                                                       es_2_1_5MyFalse_1_argbuf_d[0]}), es_2_1_1MyFalse_1_argbuf_d, es_2_1_4MyFalse_1_argbuf_d, es_2_1_5MyFalse_1_argbuf_d);
  assign {es_2_1_1MyFalse_1_argbuf_r,
          es_2_1_4MyFalse_1_argbuf_r,
          es_2_1_5MyFalse_1_argbuf_r} = {3 {(applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int2_r && applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int2_d[0])}};
  
  /* demux (Ty MyBool,
       Ty Pointer_CTf_f_Int) : (es_2_1_2,MyBool) (lizzieLet17_5QNone_Int_7QVal_Int_4QVal_Int,Pointer_CTf_f_Int) > [(es_2_1_2MyFalse,Pointer_CTf_f_Int),
                                                                                                                   (es_2_1_2MyTrue,Pointer_CTf_f_Int)] */
  logic [1:0] lizzieLet17_5QNone_Int_7QVal_Int_4QVal_Int_onehotd;
  always_comb
    if ((es_2_1_2_d[0] && lizzieLet17_5QNone_Int_7QVal_Int_4QVal_Int_d[0]))
      unique case (es_2_1_2_d[1:1])
        1'd0: lizzieLet17_5QNone_Int_7QVal_Int_4QVal_Int_onehotd = 2'd1;
        1'd1: lizzieLet17_5QNone_Int_7QVal_Int_4QVal_Int_onehotd = 2'd2;
        default: lizzieLet17_5QNone_Int_7QVal_Int_4QVal_Int_onehotd = 2'd0;
      endcase
    else lizzieLet17_5QNone_Int_7QVal_Int_4QVal_Int_onehotd = 2'd0;
  assign es_2_1_2MyFalse_d = {lizzieLet17_5QNone_Int_7QVal_Int_4QVal_Int_d[16:1],
                              lizzieLet17_5QNone_Int_7QVal_Int_4QVal_Int_onehotd[0]};
  assign es_2_1_2MyTrue_d = {lizzieLet17_5QNone_Int_7QVal_Int_4QVal_Int_d[16:1],
                             lizzieLet17_5QNone_Int_7QVal_Int_4QVal_Int_onehotd[1]};
  assign lizzieLet17_5QNone_Int_7QVal_Int_4QVal_Int_r = (| (lizzieLet17_5QNone_Int_7QVal_Int_4QVal_Int_onehotd & {es_2_1_2MyTrue_r,
                                                                                                                  es_2_1_2MyFalse_r}));
  assign es_2_1_2_r = lizzieLet17_5QNone_Int_7QVal_Int_4QVal_Int_r;
  
  /* buf (Ty Pointer_CTf_f_Int) : (es_2_1_2MyFalse,Pointer_CTf_f_Int) > (es_2_1_2MyFalse_1_argbuf,Pointer_CTf_f_Int) */
  Pointer_CTf_f_Int_t es_2_1_2MyFalse_bufchan_d;
  logic es_2_1_2MyFalse_bufchan_r;
  assign es_2_1_2MyFalse_r = ((! es_2_1_2MyFalse_bufchan_d[0]) || es_2_1_2MyFalse_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_2_1_2MyFalse_bufchan_d <= {16'd0, 1'd0};
    else
      if (es_2_1_2MyFalse_r)
        es_2_1_2MyFalse_bufchan_d <= es_2_1_2MyFalse_d;
  Pointer_CTf_f_Int_t es_2_1_2MyFalse_bufchan_buf;
  assign es_2_1_2MyFalse_bufchan_r = (! es_2_1_2MyFalse_bufchan_buf[0]);
  assign es_2_1_2MyFalse_1_argbuf_d = (es_2_1_2MyFalse_bufchan_buf[0] ? es_2_1_2MyFalse_bufchan_buf :
                                       es_2_1_2MyFalse_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_2_1_2MyFalse_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((es_2_1_2MyFalse_1_argbuf_r && es_2_1_2MyFalse_bufchan_buf[0]))
        es_2_1_2MyFalse_bufchan_buf <= {16'd0, 1'd0};
      else if (((! es_2_1_2MyFalse_1_argbuf_r) && (! es_2_1_2MyFalse_bufchan_buf[0])))
        es_2_1_2MyFalse_bufchan_buf <= es_2_1_2MyFalse_bufchan_d;
  
  /* buf (Ty Pointer_CTf_f_Int) : (es_2_1_2MyTrue,Pointer_CTf_f_Int) > (es_2_1_2MyTrue_1_argbuf,Pointer_CTf_f_Int) */
  Pointer_CTf_f_Int_t es_2_1_2MyTrue_bufchan_d;
  logic es_2_1_2MyTrue_bufchan_r;
  assign es_2_1_2MyTrue_r = ((! es_2_1_2MyTrue_bufchan_d[0]) || es_2_1_2MyTrue_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_2_1_2MyTrue_bufchan_d <= {16'd0, 1'd0};
    else
      if (es_2_1_2MyTrue_r) es_2_1_2MyTrue_bufchan_d <= es_2_1_2MyTrue_d;
  Pointer_CTf_f_Int_t es_2_1_2MyTrue_bufchan_buf;
  assign es_2_1_2MyTrue_bufchan_r = (! es_2_1_2MyTrue_bufchan_buf[0]);
  assign es_2_1_2MyTrue_1_argbuf_d = (es_2_1_2MyTrue_bufchan_buf[0] ? es_2_1_2MyTrue_bufchan_buf :
                                      es_2_1_2MyTrue_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_2_1_2MyTrue_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((es_2_1_2MyTrue_1_argbuf_r && es_2_1_2MyTrue_bufchan_buf[0]))
        es_2_1_2MyTrue_bufchan_buf <= {16'd0, 1'd0};
      else if (((! es_2_1_2MyTrue_1_argbuf_r) && (! es_2_1_2MyTrue_bufchan_buf[0])))
        es_2_1_2MyTrue_bufchan_buf <= es_2_1_2MyTrue_bufchan_d;
  
  /* demux (Ty MyBool,
       Ty Go) : (es_2_1_3,MyBool) (lizzieLet17_5QNone_Int_7QVal_Int_5QVal_Int_2,Go) > [(es_2_1_3MyFalse,Go),
                                                                                       (es_2_1_3MyTrue,Go)] */
  logic [1:0] lizzieLet17_5QNone_Int_7QVal_Int_5QVal_Int_2_onehotd;
  always_comb
    if ((es_2_1_3_d[0] && lizzieLet17_5QNone_Int_7QVal_Int_5QVal_Int_2_d[0]))
      unique case (es_2_1_3_d[1:1])
        1'd0: lizzieLet17_5QNone_Int_7QVal_Int_5QVal_Int_2_onehotd = 2'd1;
        1'd1: lizzieLet17_5QNone_Int_7QVal_Int_5QVal_Int_2_onehotd = 2'd2;
        default:
          lizzieLet17_5QNone_Int_7QVal_Int_5QVal_Int_2_onehotd = 2'd0;
      endcase
    else lizzieLet17_5QNone_Int_7QVal_Int_5QVal_Int_2_onehotd = 2'd0;
  assign es_2_1_3MyFalse_d = lizzieLet17_5QNone_Int_7QVal_Int_5QVal_Int_2_onehotd[0];
  assign es_2_1_3MyTrue_d = lizzieLet17_5QNone_Int_7QVal_Int_5QVal_Int_2_onehotd[1];
  assign lizzieLet17_5QNone_Int_7QVal_Int_5QVal_Int_2_r = (| (lizzieLet17_5QNone_Int_7QVal_Int_5QVal_Int_2_onehotd & {es_2_1_3MyTrue_r,
                                                                                                                      es_2_1_3MyFalse_r}));
  assign es_2_1_3_r = lizzieLet17_5QNone_Int_7QVal_Int_5QVal_Int_2_r;
  
  /* buf (Ty Go) : (es_2_1_3MyFalse,Go) > (es_2_1_3MyFalse_1_argbuf,Go) */
  Go_t es_2_1_3MyFalse_bufchan_d;
  logic es_2_1_3MyFalse_bufchan_r;
  assign es_2_1_3MyFalse_r = ((! es_2_1_3MyFalse_bufchan_d[0]) || es_2_1_3MyFalse_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_2_1_3MyFalse_bufchan_d <= 1'd0;
    else
      if (es_2_1_3MyFalse_r)
        es_2_1_3MyFalse_bufchan_d <= es_2_1_3MyFalse_d;
  Go_t es_2_1_3MyFalse_bufchan_buf;
  assign es_2_1_3MyFalse_bufchan_r = (! es_2_1_3MyFalse_bufchan_buf[0]);
  assign es_2_1_3MyFalse_1_argbuf_d = (es_2_1_3MyFalse_bufchan_buf[0] ? es_2_1_3MyFalse_bufchan_buf :
                                       es_2_1_3MyFalse_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_2_1_3MyFalse_bufchan_buf <= 1'd0;
    else
      if ((es_2_1_3MyFalse_1_argbuf_r && es_2_1_3MyFalse_bufchan_buf[0]))
        es_2_1_3MyFalse_bufchan_buf <= 1'd0;
      else if (((! es_2_1_3MyFalse_1_argbuf_r) && (! es_2_1_3MyFalse_bufchan_buf[0])))
        es_2_1_3MyFalse_bufchan_buf <= es_2_1_3MyFalse_bufchan_d;
  
  /* fork (Ty Go) : (es_2_1_3MyTrue,Go) > [(es_2_1_3MyTrue_1,Go),
                                      (es_2_1_3MyTrue_2,Go)] */
  logic [1:0] es_2_1_3MyTrue_emitted;
  logic [1:0] es_2_1_3MyTrue_done;
  assign es_2_1_3MyTrue_1_d = (es_2_1_3MyTrue_d[0] && (! es_2_1_3MyTrue_emitted[0]));
  assign es_2_1_3MyTrue_2_d = (es_2_1_3MyTrue_d[0] && (! es_2_1_3MyTrue_emitted[1]));
  assign es_2_1_3MyTrue_done = (es_2_1_3MyTrue_emitted | ({es_2_1_3MyTrue_2_d[0],
                                                           es_2_1_3MyTrue_1_d[0]} & {es_2_1_3MyTrue_2_r,
                                                                                     es_2_1_3MyTrue_1_r}));
  assign es_2_1_3MyTrue_r = (& es_2_1_3MyTrue_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_2_1_3MyTrue_emitted <= 2'd0;
    else
      es_2_1_3MyTrue_emitted <= (es_2_1_3MyTrue_r ? 2'd0 :
                                 es_2_1_3MyTrue_done);
  
  /* dcon (Ty QTree_Int,
      Dcon QNone_Int) : [(es_2_1_3MyTrue_1,Go)] > (es_2_1_3MyTrue_1QNone_Int,QTree_Int) */
  assign es_2_1_3MyTrue_1QNone_Int_d = QNone_Int_dc((& {es_2_1_3MyTrue_1_d[0]}), es_2_1_3MyTrue_1_d);
  assign {es_2_1_3MyTrue_1_r} = {1 {(es_2_1_3MyTrue_1QNone_Int_r && es_2_1_3MyTrue_1QNone_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (es_2_1_3MyTrue_1QNone_Int,QTree_Int) > (lizzieLet21_1_argbuf,QTree_Int) */
  QTree_Int_t es_2_1_3MyTrue_1QNone_Int_bufchan_d;
  logic es_2_1_3MyTrue_1QNone_Int_bufchan_r;
  assign es_2_1_3MyTrue_1QNone_Int_r = ((! es_2_1_3MyTrue_1QNone_Int_bufchan_d[0]) || es_2_1_3MyTrue_1QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_2_1_3MyTrue_1QNone_Int_bufchan_d <= {66'd0, 1'd0};
    else
      if (es_2_1_3MyTrue_1QNone_Int_r)
        es_2_1_3MyTrue_1QNone_Int_bufchan_d <= es_2_1_3MyTrue_1QNone_Int_d;
  QTree_Int_t es_2_1_3MyTrue_1QNone_Int_bufchan_buf;
  assign es_2_1_3MyTrue_1QNone_Int_bufchan_r = (! es_2_1_3MyTrue_1QNone_Int_bufchan_buf[0]);
  assign lizzieLet21_1_argbuf_d = (es_2_1_3MyTrue_1QNone_Int_bufchan_buf[0] ? es_2_1_3MyTrue_1QNone_Int_bufchan_buf :
                                   es_2_1_3MyTrue_1QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_2_1_3MyTrue_1QNone_Int_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((lizzieLet21_1_argbuf_r && es_2_1_3MyTrue_1QNone_Int_bufchan_buf[0]))
        es_2_1_3MyTrue_1QNone_Int_bufchan_buf <= {66'd0, 1'd0};
      else if (((! lizzieLet21_1_argbuf_r) && (! es_2_1_3MyTrue_1QNone_Int_bufchan_buf[0])))
        es_2_1_3MyTrue_1QNone_Int_bufchan_buf <= es_2_1_3MyTrue_1QNone_Int_bufchan_d;
  
  /* buf (Ty Go) : (es_2_1_3MyTrue_2,Go) > (es_2_1_3MyTrue_2_argbuf,Go) */
  Go_t es_2_1_3MyTrue_2_bufchan_d;
  logic es_2_1_3MyTrue_2_bufchan_r;
  assign es_2_1_3MyTrue_2_r = ((! es_2_1_3MyTrue_2_bufchan_d[0]) || es_2_1_3MyTrue_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_2_1_3MyTrue_2_bufchan_d <= 1'd0;
    else
      if (es_2_1_3MyTrue_2_r)
        es_2_1_3MyTrue_2_bufchan_d <= es_2_1_3MyTrue_2_d;
  Go_t es_2_1_3MyTrue_2_bufchan_buf;
  assign es_2_1_3MyTrue_2_bufchan_r = (! es_2_1_3MyTrue_2_bufchan_buf[0]);
  assign es_2_1_3MyTrue_2_argbuf_d = (es_2_1_3MyTrue_2_bufchan_buf[0] ? es_2_1_3MyTrue_2_bufchan_buf :
                                      es_2_1_3MyTrue_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_2_1_3MyTrue_2_bufchan_buf <= 1'd0;
    else
      if ((es_2_1_3MyTrue_2_argbuf_r && es_2_1_3MyTrue_2_bufchan_buf[0]))
        es_2_1_3MyTrue_2_bufchan_buf <= 1'd0;
      else if (((! es_2_1_3MyTrue_2_argbuf_r) && (! es_2_1_3MyTrue_2_bufchan_buf[0])))
        es_2_1_3MyTrue_2_bufchan_buf <= es_2_1_3MyTrue_2_bufchan_d;
  
  /* demux (Ty MyBool,
       Ty Int) : (es_2_1_4,MyBool) (lizzieLet17_5QNone_Int_7QVal_Int_8QVal_Int_2,Int) > [(es_2_1_4MyFalse,Int),
                                                                                         (_229,Int)] */
  logic [1:0] lizzieLet17_5QNone_Int_7QVal_Int_8QVal_Int_2_onehotd;
  always_comb
    if ((es_2_1_4_d[0] && lizzieLet17_5QNone_Int_7QVal_Int_8QVal_Int_2_d[0]))
      unique case (es_2_1_4_d[1:1])
        1'd0: lizzieLet17_5QNone_Int_7QVal_Int_8QVal_Int_2_onehotd = 2'd1;
        1'd1: lizzieLet17_5QNone_Int_7QVal_Int_8QVal_Int_2_onehotd = 2'd2;
        default:
          lizzieLet17_5QNone_Int_7QVal_Int_8QVal_Int_2_onehotd = 2'd0;
      endcase
    else lizzieLet17_5QNone_Int_7QVal_Int_8QVal_Int_2_onehotd = 2'd0;
  assign es_2_1_4MyFalse_d = {lizzieLet17_5QNone_Int_7QVal_Int_8QVal_Int_2_d[32:1],
                              lizzieLet17_5QNone_Int_7QVal_Int_8QVal_Int_2_onehotd[0]};
  assign _229_d = {lizzieLet17_5QNone_Int_7QVal_Int_8QVal_Int_2_d[32:1],
                   lizzieLet17_5QNone_Int_7QVal_Int_8QVal_Int_2_onehotd[1]};
  assign lizzieLet17_5QNone_Int_7QVal_Int_8QVal_Int_2_r = (| (lizzieLet17_5QNone_Int_7QVal_Int_8QVal_Int_2_onehotd & {_229_r,
                                                                                                                      es_2_1_4MyFalse_r}));
  assign es_2_1_4_r = lizzieLet17_5QNone_Int_7QVal_Int_8QVal_Int_2_r;
  
  /* buf (Ty Int) : (es_2_1_4MyFalse,Int) > (es_2_1_4MyFalse_1_argbuf,Int) */
  Int_t es_2_1_4MyFalse_bufchan_d;
  logic es_2_1_4MyFalse_bufchan_r;
  assign es_2_1_4MyFalse_r = ((! es_2_1_4MyFalse_bufchan_d[0]) || es_2_1_4MyFalse_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_2_1_4MyFalse_bufchan_d <= {32'd0, 1'd0};
    else
      if (es_2_1_4MyFalse_r)
        es_2_1_4MyFalse_bufchan_d <= es_2_1_4MyFalse_d;
  Int_t es_2_1_4MyFalse_bufchan_buf;
  assign es_2_1_4MyFalse_bufchan_r = (! es_2_1_4MyFalse_bufchan_buf[0]);
  assign es_2_1_4MyFalse_1_argbuf_d = (es_2_1_4MyFalse_bufchan_buf[0] ? es_2_1_4MyFalse_bufchan_buf :
                                       es_2_1_4MyFalse_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_2_1_4MyFalse_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((es_2_1_4MyFalse_1_argbuf_r && es_2_1_4MyFalse_bufchan_buf[0]))
        es_2_1_4MyFalse_bufchan_buf <= {32'd0, 1'd0};
      else if (((! es_2_1_4MyFalse_1_argbuf_r) && (! es_2_1_4MyFalse_bufchan_buf[0])))
        es_2_1_4MyFalse_bufchan_buf <= es_2_1_4MyFalse_bufchan_d;
  
  /* demux (Ty MyBool,
       Ty Int) : (es_2_1_5,MyBool) (vaew_2,Int) > [(es_2_1_5MyFalse,Int),
                                                   (_228,Int)] */
  logic [1:0] vaew_2_onehotd;
  always_comb
    if ((es_2_1_5_d[0] && vaew_2_d[0]))
      unique case (es_2_1_5_d[1:1])
        1'd0: vaew_2_onehotd = 2'd1;
        1'd1: vaew_2_onehotd = 2'd2;
        default: vaew_2_onehotd = 2'd0;
      endcase
    else vaew_2_onehotd = 2'd0;
  assign es_2_1_5MyFalse_d = {vaew_2_d[32:1], vaew_2_onehotd[0]};
  assign _228_d = {vaew_2_d[32:1], vaew_2_onehotd[1]};
  assign vaew_2_r = (| (vaew_2_onehotd & {_228_r,
                                          es_2_1_5MyFalse_r}));
  assign es_2_1_5_r = vaew_2_r;
  
  /* buf (Ty Int) : (es_2_1_5MyFalse,Int) > (es_2_1_5MyFalse_1_argbuf,Int) */
  Int_t es_2_1_5MyFalse_bufchan_d;
  logic es_2_1_5MyFalse_bufchan_r;
  assign es_2_1_5MyFalse_r = ((! es_2_1_5MyFalse_bufchan_d[0]) || es_2_1_5MyFalse_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_2_1_5MyFalse_bufchan_d <= {32'd0, 1'd0};
    else
      if (es_2_1_5MyFalse_r)
        es_2_1_5MyFalse_bufchan_d <= es_2_1_5MyFalse_d;
  Int_t es_2_1_5MyFalse_bufchan_buf;
  assign es_2_1_5MyFalse_bufchan_r = (! es_2_1_5MyFalse_bufchan_buf[0]);
  assign es_2_1_5MyFalse_1_argbuf_d = (es_2_1_5MyFalse_bufchan_buf[0] ? es_2_1_5MyFalse_bufchan_buf :
                                       es_2_1_5MyFalse_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_2_1_5MyFalse_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((es_2_1_5MyFalse_1_argbuf_r && es_2_1_5MyFalse_bufchan_buf[0]))
        es_2_1_5MyFalse_bufchan_buf <= {32'd0, 1'd0};
      else if (((! es_2_1_5MyFalse_1_argbuf_r) && (! es_2_1_5MyFalse_bufchan_buf[0])))
        es_2_1_5MyFalse_bufchan_buf <= es_2_1_5MyFalse_bufchan_d;
  
  /* demux (Ty MyBool,
       Ty MyDTInt_Int_Int) : (es_2_2,MyBool) (lizzieLet6_5QVal_Int_5QVal_Int_2,MyDTInt_Int_Int) > [(es_2_2MyFalse,MyDTInt_Int_Int),
                                                                                                   (_227,MyDTInt_Int_Int)] */
  logic [1:0] lizzieLet6_5QVal_Int_5QVal_Int_2_onehotd;
  always_comb
    if ((es_2_2_d[0] && lizzieLet6_5QVal_Int_5QVal_Int_2_d[0]))
      unique case (es_2_2_d[1:1])
        1'd0: lizzieLet6_5QVal_Int_5QVal_Int_2_onehotd = 2'd1;
        1'd1: lizzieLet6_5QVal_Int_5QVal_Int_2_onehotd = 2'd2;
        default: lizzieLet6_5QVal_Int_5QVal_Int_2_onehotd = 2'd0;
      endcase
    else lizzieLet6_5QVal_Int_5QVal_Int_2_onehotd = 2'd0;
  assign es_2_2MyFalse_d = lizzieLet6_5QVal_Int_5QVal_Int_2_onehotd[0];
  assign _227_d = lizzieLet6_5QVal_Int_5QVal_Int_2_onehotd[1];
  assign lizzieLet6_5QVal_Int_5QVal_Int_2_r = (| (lizzieLet6_5QVal_Int_5QVal_Int_2_onehotd & {_227_r,
                                                                                              es_2_2MyFalse_r}));
  assign es_2_2_r = lizzieLet6_5QVal_Int_5QVal_Int_2_r;
  
  /* buf (Ty MyDTInt_Int_Int) : (es_2_2MyFalse,MyDTInt_Int_Int) > (es_2_2MyFalse_1_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t es_2_2MyFalse_bufchan_d;
  logic es_2_2MyFalse_bufchan_r;
  assign es_2_2MyFalse_r = ((! es_2_2MyFalse_bufchan_d[0]) || es_2_2MyFalse_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_2_2MyFalse_bufchan_d <= 1'd0;
    else
      if (es_2_2MyFalse_r) es_2_2MyFalse_bufchan_d <= es_2_2MyFalse_d;
  MyDTInt_Int_Int_t es_2_2MyFalse_bufchan_buf;
  assign es_2_2MyFalse_bufchan_r = (! es_2_2MyFalse_bufchan_buf[0]);
  assign es_2_2MyFalse_1_argbuf_d = (es_2_2MyFalse_bufchan_buf[0] ? es_2_2MyFalse_bufchan_buf :
                                     es_2_2MyFalse_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_2_2MyFalse_bufchan_buf <= 1'd0;
    else
      if ((es_2_2MyFalse_1_argbuf_r && es_2_2MyFalse_bufchan_buf[0]))
        es_2_2MyFalse_bufchan_buf <= 1'd0;
      else if (((! es_2_2MyFalse_1_argbuf_r) && (! es_2_2MyFalse_bufchan_buf[0])))
        es_2_2MyFalse_bufchan_buf <= es_2_2MyFalse_bufchan_d;
  
  /* dcon (Ty TupMyDTInt_Int_Int___Int___Int,
      Dcon TupMyDTInt_Int_Int___Int___Int) : [(es_2_2MyFalse_1_argbuf,MyDTInt_Int_Int),
                                              (es_2_4MyFalse_1_argbuf,Int),
                                              (es_2_5MyFalse_1_argbuf,Int)] > (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int4,TupMyDTInt_Int_Int___Int___Int) */
  assign applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int4_d = TupMyDTInt_Int_Int___Int___Int_dc((& {es_2_2MyFalse_1_argbuf_d[0],
                                                                                                       es_2_4MyFalse_1_argbuf_d[0],
                                                                                                       es_2_5MyFalse_1_argbuf_d[0]}), es_2_2MyFalse_1_argbuf_d, es_2_4MyFalse_1_argbuf_d, es_2_5MyFalse_1_argbuf_d);
  assign {es_2_2MyFalse_1_argbuf_r,
          es_2_4MyFalse_1_argbuf_r,
          es_2_5MyFalse_1_argbuf_r} = {3 {(applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int4_r && applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int4_d[0])}};
  
  /* demux (Ty MyBool,
       Ty Pointer_CTf''''''''''''_f''''''''''''_Int) : (es_2_3,MyBool) (lizzieLet6_5QVal_Int_7QVal_Int,Pointer_CTf''''''''''''_f''''''''''''_Int) > [(es_2_3MyFalse,Pointer_CTf''''''''''''_f''''''''''''_Int),
                                                                                                                                                     (es_2_3MyTrue,Pointer_CTf''''''''''''_f''''''''''''_Int)] */
  logic [1:0] lizzieLet6_5QVal_Int_7QVal_Int_onehotd;
  always_comb
    if ((es_2_3_d[0] && lizzieLet6_5QVal_Int_7QVal_Int_d[0]))
      unique case (es_2_3_d[1:1])
        1'd0: lizzieLet6_5QVal_Int_7QVal_Int_onehotd = 2'd1;
        1'd1: lizzieLet6_5QVal_Int_7QVal_Int_onehotd = 2'd2;
        default: lizzieLet6_5QVal_Int_7QVal_Int_onehotd = 2'd0;
      endcase
    else lizzieLet6_5QVal_Int_7QVal_Int_onehotd = 2'd0;
  assign es_2_3MyFalse_d = {lizzieLet6_5QVal_Int_7QVal_Int_d[16:1],
                            lizzieLet6_5QVal_Int_7QVal_Int_onehotd[0]};
  assign es_2_3MyTrue_d = {lizzieLet6_5QVal_Int_7QVal_Int_d[16:1],
                           lizzieLet6_5QVal_Int_7QVal_Int_onehotd[1]};
  assign lizzieLet6_5QVal_Int_7QVal_Int_r = (| (lizzieLet6_5QVal_Int_7QVal_Int_onehotd & {es_2_3MyTrue_r,
                                                                                          es_2_3MyFalse_r}));
  assign es_2_3_r = lizzieLet6_5QVal_Int_7QVal_Int_r;
  
  /* buf (Ty Pointer_CTf''''''''''''_f''''''''''''_Int) : (es_2_3MyFalse,Pointer_CTf''''''''''''_f''''''''''''_Int) > (es_2_3MyFalse_1_argbuf,Pointer_CTf''''''''''''_f''''''''''''_Int) */
  \Pointer_CTf''''''''''''_f''''''''''''_Int_t  es_2_3MyFalse_bufchan_d;
  logic es_2_3MyFalse_bufchan_r;
  assign es_2_3MyFalse_r = ((! es_2_3MyFalse_bufchan_d[0]) || es_2_3MyFalse_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_2_3MyFalse_bufchan_d <= {16'd0, 1'd0};
    else
      if (es_2_3MyFalse_r) es_2_3MyFalse_bufchan_d <= es_2_3MyFalse_d;
  \Pointer_CTf''''''''''''_f''''''''''''_Int_t  es_2_3MyFalse_bufchan_buf;
  assign es_2_3MyFalse_bufchan_r = (! es_2_3MyFalse_bufchan_buf[0]);
  assign es_2_3MyFalse_1_argbuf_d = (es_2_3MyFalse_bufchan_buf[0] ? es_2_3MyFalse_bufchan_buf :
                                     es_2_3MyFalse_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_2_3MyFalse_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((es_2_3MyFalse_1_argbuf_r && es_2_3MyFalse_bufchan_buf[0]))
        es_2_3MyFalse_bufchan_buf <= {16'd0, 1'd0};
      else if (((! es_2_3MyFalse_1_argbuf_r) && (! es_2_3MyFalse_bufchan_buf[0])))
        es_2_3MyFalse_bufchan_buf <= es_2_3MyFalse_bufchan_d;
  
  /* buf (Ty Pointer_CTf''''''''''''_f''''''''''''_Int) : (es_2_3MyTrue,Pointer_CTf''''''''''''_f''''''''''''_Int) > (es_2_3MyTrue_1_argbuf,Pointer_CTf''''''''''''_f''''''''''''_Int) */
  \Pointer_CTf''''''''''''_f''''''''''''_Int_t  es_2_3MyTrue_bufchan_d;
  logic es_2_3MyTrue_bufchan_r;
  assign es_2_3MyTrue_r = ((! es_2_3MyTrue_bufchan_d[0]) || es_2_3MyTrue_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_2_3MyTrue_bufchan_d <= {16'd0, 1'd0};
    else if (es_2_3MyTrue_r) es_2_3MyTrue_bufchan_d <= es_2_3MyTrue_d;
  \Pointer_CTf''''''''''''_f''''''''''''_Int_t  es_2_3MyTrue_bufchan_buf;
  assign es_2_3MyTrue_bufchan_r = (! es_2_3MyTrue_bufchan_buf[0]);
  assign es_2_3MyTrue_1_argbuf_d = (es_2_3MyTrue_bufchan_buf[0] ? es_2_3MyTrue_bufchan_buf :
                                    es_2_3MyTrue_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_2_3MyTrue_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((es_2_3MyTrue_1_argbuf_r && es_2_3MyTrue_bufchan_buf[0]))
        es_2_3MyTrue_bufchan_buf <= {16'd0, 1'd0};
      else if (((! es_2_3MyTrue_1_argbuf_r) && (! es_2_3MyTrue_bufchan_buf[0])))
        es_2_3MyTrue_bufchan_buf <= es_2_3MyTrue_bufchan_d;
  
  /* demux (Ty MyBool,
       Ty Int) : (es_2_4,MyBool) (lizzieLet6_5QVal_Int_8QVal_Int_2,Int) > [(es_2_4MyFalse,Int),
                                                                           (_226,Int)] */
  logic [1:0] lizzieLet6_5QVal_Int_8QVal_Int_2_onehotd;
  always_comb
    if ((es_2_4_d[0] && lizzieLet6_5QVal_Int_8QVal_Int_2_d[0]))
      unique case (es_2_4_d[1:1])
        1'd0: lizzieLet6_5QVal_Int_8QVal_Int_2_onehotd = 2'd1;
        1'd1: lizzieLet6_5QVal_Int_8QVal_Int_2_onehotd = 2'd2;
        default: lizzieLet6_5QVal_Int_8QVal_Int_2_onehotd = 2'd0;
      endcase
    else lizzieLet6_5QVal_Int_8QVal_Int_2_onehotd = 2'd0;
  assign es_2_4MyFalse_d = {lizzieLet6_5QVal_Int_8QVal_Int_2_d[32:1],
                            lizzieLet6_5QVal_Int_8QVal_Int_2_onehotd[0]};
  assign _226_d = {lizzieLet6_5QVal_Int_8QVal_Int_2_d[32:1],
                   lizzieLet6_5QVal_Int_8QVal_Int_2_onehotd[1]};
  assign lizzieLet6_5QVal_Int_8QVal_Int_2_r = (| (lizzieLet6_5QVal_Int_8QVal_Int_2_onehotd & {_226_r,
                                                                                              es_2_4MyFalse_r}));
  assign es_2_4_r = lizzieLet6_5QVal_Int_8QVal_Int_2_r;
  
  /* buf (Ty Int) : (es_2_4MyFalse,Int) > (es_2_4MyFalse_1_argbuf,Int) */
  Int_t es_2_4MyFalse_bufchan_d;
  logic es_2_4MyFalse_bufchan_r;
  assign es_2_4MyFalse_r = ((! es_2_4MyFalse_bufchan_d[0]) || es_2_4MyFalse_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_2_4MyFalse_bufchan_d <= {32'd0, 1'd0};
    else
      if (es_2_4MyFalse_r) es_2_4MyFalse_bufchan_d <= es_2_4MyFalse_d;
  Int_t es_2_4MyFalse_bufchan_buf;
  assign es_2_4MyFalse_bufchan_r = (! es_2_4MyFalse_bufchan_buf[0]);
  assign es_2_4MyFalse_1_argbuf_d = (es_2_4MyFalse_bufchan_buf[0] ? es_2_4MyFalse_bufchan_buf :
                                     es_2_4MyFalse_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_2_4MyFalse_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((es_2_4MyFalse_1_argbuf_r && es_2_4MyFalse_bufchan_buf[0]))
        es_2_4MyFalse_bufchan_buf <= {32'd0, 1'd0};
      else if (((! es_2_4MyFalse_1_argbuf_r) && (! es_2_4MyFalse_bufchan_buf[0])))
        es_2_4MyFalse_bufchan_buf <= es_2_4MyFalse_bufchan_d;
  
  /* demux (Ty MyBool,
       Ty Int) : (es_2_5,MyBool) (vafo_2,Int) > [(es_2_5MyFalse,Int),
                                                 (_225,Int)] */
  logic [1:0] vafo_2_onehotd;
  always_comb
    if ((es_2_5_d[0] && vafo_2_d[0]))
      unique case (es_2_5_d[1:1])
        1'd0: vafo_2_onehotd = 2'd1;
        1'd1: vafo_2_onehotd = 2'd2;
        default: vafo_2_onehotd = 2'd0;
      endcase
    else vafo_2_onehotd = 2'd0;
  assign es_2_5MyFalse_d = {vafo_2_d[32:1], vafo_2_onehotd[0]};
  assign _225_d = {vafo_2_d[32:1], vafo_2_onehotd[1]};
  assign vafo_2_r = (| (vafo_2_onehotd & {_225_r, es_2_5MyFalse_r}));
  assign es_2_5_r = vafo_2_r;
  
  /* buf (Ty Int) : (es_2_5MyFalse,Int) > (es_2_5MyFalse_1_argbuf,Int) */
  Int_t es_2_5MyFalse_bufchan_d;
  logic es_2_5MyFalse_bufchan_r;
  assign es_2_5MyFalse_r = ((! es_2_5MyFalse_bufchan_d[0]) || es_2_5MyFalse_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_2_5MyFalse_bufchan_d <= {32'd0, 1'd0};
    else
      if (es_2_5MyFalse_r) es_2_5MyFalse_bufchan_d <= es_2_5MyFalse_d;
  Int_t es_2_5MyFalse_bufchan_buf;
  assign es_2_5MyFalse_bufchan_r = (! es_2_5MyFalse_bufchan_buf[0]);
  assign es_2_5MyFalse_1_argbuf_d = (es_2_5MyFalse_bufchan_buf[0] ? es_2_5MyFalse_bufchan_buf :
                                     es_2_5MyFalse_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_2_5MyFalse_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((es_2_5MyFalse_1_argbuf_r && es_2_5MyFalse_bufchan_buf[0]))
        es_2_5MyFalse_bufchan_buf <= {32'd0, 1'd0};
      else if (((! es_2_5MyFalse_1_argbuf_r) && (! es_2_5MyFalse_bufchan_buf[0])))
        es_2_5MyFalse_bufchan_buf <= es_2_5MyFalse_bufchan_d;
  
  /* buf (Ty QTree_Int) : (es_30_1es_31_1es_32_1es_33_1QNode_Int,QTree_Int) > (lizzieLet50_1_argbuf,QTree_Int) */
  QTree_Int_t es_30_1es_31_1es_32_1es_33_1QNode_Int_bufchan_d;
  logic es_30_1es_31_1es_32_1es_33_1QNode_Int_bufchan_r;
  assign es_30_1es_31_1es_32_1es_33_1QNode_Int_r = ((! es_30_1es_31_1es_32_1es_33_1QNode_Int_bufchan_d[0]) || es_30_1es_31_1es_32_1es_33_1QNode_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_30_1es_31_1es_32_1es_33_1QNode_Int_bufchan_d <= {66'd0, 1'd0};
    else
      if (es_30_1es_31_1es_32_1es_33_1QNode_Int_r)
        es_30_1es_31_1es_32_1es_33_1QNode_Int_bufchan_d <= es_30_1es_31_1es_32_1es_33_1QNode_Int_d;
  QTree_Int_t es_30_1es_31_1es_32_1es_33_1QNode_Int_bufchan_buf;
  assign es_30_1es_31_1es_32_1es_33_1QNode_Int_bufchan_r = (! es_30_1es_31_1es_32_1es_33_1QNode_Int_bufchan_buf[0]);
  assign lizzieLet50_1_argbuf_d = (es_30_1es_31_1es_32_1es_33_1QNode_Int_bufchan_buf[0] ? es_30_1es_31_1es_32_1es_33_1QNode_Int_bufchan_buf :
                                   es_30_1es_31_1es_32_1es_33_1QNode_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_30_1es_31_1es_32_1es_33_1QNode_Int_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((lizzieLet50_1_argbuf_r && es_30_1es_31_1es_32_1es_33_1QNode_Int_bufchan_buf[0]))
        es_30_1es_31_1es_32_1es_33_1QNode_Int_bufchan_buf <= {66'd0, 1'd0};
      else if (((! lizzieLet50_1_argbuf_r) && (! es_30_1es_31_1es_32_1es_33_1QNode_Int_bufchan_buf[0])))
        es_30_1es_31_1es_32_1es_33_1QNode_Int_bufchan_buf <= es_30_1es_31_1es_32_1es_33_1QNode_Int_bufchan_d;
  
  /* buf (Ty QTree_Int) : (es_3_1QVal_Int,QTree_Int) > (lizzieLet8_1_argbuf,QTree_Int) */
  QTree_Int_t es_3_1QVal_Int_bufchan_d;
  logic es_3_1QVal_Int_bufchan_r;
  assign es_3_1QVal_Int_r = ((! es_3_1QVal_Int_bufchan_d[0]) || es_3_1QVal_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_3_1QVal_Int_bufchan_d <= {66'd0, 1'd0};
    else
      if (es_3_1QVal_Int_r) es_3_1QVal_Int_bufchan_d <= es_3_1QVal_Int_d;
  QTree_Int_t es_3_1QVal_Int_bufchan_buf;
  assign es_3_1QVal_Int_bufchan_r = (! es_3_1QVal_Int_bufchan_buf[0]);
  assign lizzieLet8_1_argbuf_d = (es_3_1QVal_Int_bufchan_buf[0] ? es_3_1QVal_Int_bufchan_buf :
                                  es_3_1QVal_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_3_1QVal_Int_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((lizzieLet8_1_argbuf_r && es_3_1QVal_Int_bufchan_buf[0]))
        es_3_1QVal_Int_bufchan_buf <= {66'd0, 1'd0};
      else if (((! lizzieLet8_1_argbuf_r) && (! es_3_1QVal_Int_bufchan_buf[0])))
        es_3_1QVal_Int_bufchan_buf <= es_3_1QVal_Int_bufchan_d;
  
  /* buf (Ty QTree_Int) : (es_3_1_1QVal_Int,QTree_Int) > (lizzieLet20_1_argbuf,QTree_Int) */
  QTree_Int_t es_3_1_1QVal_Int_bufchan_d;
  logic es_3_1_1QVal_Int_bufchan_r;
  assign es_3_1_1QVal_Int_r = ((! es_3_1_1QVal_Int_bufchan_d[0]) || es_3_1_1QVal_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_3_1_1QVal_Int_bufchan_d <= {66'd0, 1'd0};
    else
      if (es_3_1_1QVal_Int_r)
        es_3_1_1QVal_Int_bufchan_d <= es_3_1_1QVal_Int_d;
  QTree_Int_t es_3_1_1QVal_Int_bufchan_buf;
  assign es_3_1_1QVal_Int_bufchan_r = (! es_3_1_1QVal_Int_bufchan_buf[0]);
  assign lizzieLet20_1_argbuf_d = (es_3_1_1QVal_Int_bufchan_buf[0] ? es_3_1_1QVal_Int_bufchan_buf :
                                   es_3_1_1QVal_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_3_1_1QVal_Int_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((lizzieLet20_1_argbuf_r && es_3_1_1QVal_Int_bufchan_buf[0]))
        es_3_1_1QVal_Int_bufchan_buf <= {66'd0, 1'd0};
      else if (((! lizzieLet20_1_argbuf_r) && (! es_3_1_1QVal_Int_bufchan_buf[0])))
        es_3_1_1QVal_Int_bufchan_buf <= es_3_1_1QVal_Int_bufchan_d;
  
  /* buf (Ty QTree_Int) : (es_4_1_1es_5_1_1es_6_1_1es_7_1QNode_Int,QTree_Int) > (lizzieLet26_1_argbuf,QTree_Int) */
  QTree_Int_t es_4_1_1es_5_1_1es_6_1_1es_7_1QNode_Int_bufchan_d;
  logic es_4_1_1es_5_1_1es_6_1_1es_7_1QNode_Int_bufchan_r;
  assign es_4_1_1es_5_1_1es_6_1_1es_7_1QNode_Int_r = ((! es_4_1_1es_5_1_1es_6_1_1es_7_1QNode_Int_bufchan_d[0]) || es_4_1_1es_5_1_1es_6_1_1es_7_1QNode_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_4_1_1es_5_1_1es_6_1_1es_7_1QNode_Int_bufchan_d <= {66'd0, 1'd0};
    else
      if (es_4_1_1es_5_1_1es_6_1_1es_7_1QNode_Int_r)
        es_4_1_1es_5_1_1es_6_1_1es_7_1QNode_Int_bufchan_d <= es_4_1_1es_5_1_1es_6_1_1es_7_1QNode_Int_d;
  QTree_Int_t es_4_1_1es_5_1_1es_6_1_1es_7_1QNode_Int_bufchan_buf;
  assign es_4_1_1es_5_1_1es_6_1_1es_7_1QNode_Int_bufchan_r = (! es_4_1_1es_5_1_1es_6_1_1es_7_1QNode_Int_bufchan_buf[0]);
  assign lizzieLet26_1_argbuf_d = (es_4_1_1es_5_1_1es_6_1_1es_7_1QNode_Int_bufchan_buf[0] ? es_4_1_1es_5_1_1es_6_1_1es_7_1QNode_Int_bufchan_buf :
                                   es_4_1_1es_5_1_1es_6_1_1es_7_1QNode_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_4_1_1es_5_1_1es_6_1_1es_7_1QNode_Int_bufchan_buf <= {66'd0,
                                                              1'd0};
    else
      if ((lizzieLet26_1_argbuf_r && es_4_1_1es_5_1_1es_6_1_1es_7_1QNode_Int_bufchan_buf[0]))
        es_4_1_1es_5_1_1es_6_1_1es_7_1QNode_Int_bufchan_buf <= {66'd0,
                                                                1'd0};
      else if (((! lizzieLet26_1_argbuf_r) && (! es_4_1_1es_5_1_1es_6_1_1es_7_1QNode_Int_bufchan_buf[0])))
        es_4_1_1es_5_1_1es_6_1_1es_7_1QNode_Int_bufchan_buf <= es_4_1_1es_5_1_1es_6_1_1es_7_1QNode_Int_bufchan_d;
  
  /* buf (Ty Int#) : (es_4_2_1lizzieLet58_4Lcall_$wnnz0_1_Add32,Int#) > (contRet_0_1_argbuf,Int#) */
  \Int#_t  es_4_2_1lizzieLet58_4Lcall_$wnnz0_1_Add32_bufchan_d;
  logic es_4_2_1lizzieLet58_4Lcall_$wnnz0_1_Add32_bufchan_r;
  assign es_4_2_1lizzieLet58_4Lcall_$wnnz0_1_Add32_r = ((! es_4_2_1lizzieLet58_4Lcall_$wnnz0_1_Add32_bufchan_d[0]) || es_4_2_1lizzieLet58_4Lcall_$wnnz0_1_Add32_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_4_2_1lizzieLet58_4Lcall_$wnnz0_1_Add32_bufchan_d <= {32'd0,
                                                              1'd0};
    else
      if (es_4_2_1lizzieLet58_4Lcall_$wnnz0_1_Add32_r)
        es_4_2_1lizzieLet58_4Lcall_$wnnz0_1_Add32_bufchan_d <= es_4_2_1lizzieLet58_4Lcall_$wnnz0_1_Add32_d;
  \Int#_t  es_4_2_1lizzieLet58_4Lcall_$wnnz0_1_Add32_bufchan_buf;
  assign es_4_2_1lizzieLet58_4Lcall_$wnnz0_1_Add32_bufchan_r = (! es_4_2_1lizzieLet58_4Lcall_$wnnz0_1_Add32_bufchan_buf[0]);
  assign contRet_0_1_argbuf_d = (es_4_2_1lizzieLet58_4Lcall_$wnnz0_1_Add32_bufchan_buf[0] ? es_4_2_1lizzieLet58_4Lcall_$wnnz0_1_Add32_bufchan_buf :
                                 es_4_2_1lizzieLet58_4Lcall_$wnnz0_1_Add32_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_4_2_1lizzieLet58_4Lcall_$wnnz0_1_Add32_bufchan_buf <= {32'd0,
                                                                1'd0};
    else
      if ((contRet_0_1_argbuf_r && es_4_2_1lizzieLet58_4Lcall_$wnnz0_1_Add32_bufchan_buf[0]))
        es_4_2_1lizzieLet58_4Lcall_$wnnz0_1_Add32_bufchan_buf <= {32'd0,
                                                                  1'd0};
      else if (((! contRet_0_1_argbuf_r) && (! es_4_2_1lizzieLet58_4Lcall_$wnnz0_1_Add32_bufchan_buf[0])))
        es_4_2_1lizzieLet58_4Lcall_$wnnz0_1_Add32_bufchan_buf <= es_4_2_1lizzieLet58_4Lcall_$wnnz0_1_Add32_bufchan_d;
  
  /* sink (Ty Int) : (es_6_1I#,Int) > */
  assign {\es_6_1I#_r , \es_6_1I#_dout } = {\es_6_1I#_rout ,
                                            \es_6_1I#_d };
  
  /* op_add (Ty Int#) : (es_6_2_1ww2XmZ_1_1_Add32,Int#) (lizzieLet58_4Lcall_$wnnz0,Int#) > (es_4_2_1lizzieLet58_4Lcall_$wnnz0_1_Add32,Int#) */
  assign es_4_2_1lizzieLet58_4Lcall_$wnnz0_1_Add32_d = {(es_6_2_1ww2XmZ_1_1_Add32_d[32:1] + lizzieLet58_4Lcall_$wnnz0_d[32:1]),
                                                        (es_6_2_1ww2XmZ_1_1_Add32_d[0] && lizzieLet58_4Lcall_$wnnz0_d[0])};
  assign {es_6_2_1ww2XmZ_1_1_Add32_r,
          lizzieLet58_4Lcall_$wnnz0_r} = {2 {(es_4_2_1lizzieLet58_4Lcall_$wnnz0_1_Add32_r && es_4_2_1lizzieLet58_4Lcall_$wnnz0_1_Add32_d[0])}};
  
  /* mergectrl (Ty C12,
           Ty TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int) : [(f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1,TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int),
                                                                                                 (f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int2,TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int),
                                                                                                 (f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int3,TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int),
                                                                                                 (f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int4,TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int),
                                                                                                 (f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int5,TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int),
                                                                                                 (f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int6,TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int),
                                                                                                 (f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int7,TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int),
                                                                                                 (f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int8,TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int),
                                                                                                 (f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int9,TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int),
                                                                                                 (f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int10,TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int),
                                                                                                 (f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int11,TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int),
                                                                                                 (f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int12,TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int)] > (f''''''''''''_f''''''''''''_Int_choice,C12) (f''''''''''''_f''''''''''''_Int_data,TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int) */
  logic [11:0] \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_select_d ;
  assign \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_select_d  = ((| \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_select_q ) ? \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_select_q  :
                                                                                                                                       (\f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_d [0] ? 12'd1 :
                                                                                                                                        (\f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int2_d [0] ? 12'd2 :
                                                                                                                                         (\f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int3_d [0] ? 12'd4 :
                                                                                                                                          (\f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int4_d [0] ? 12'd8 :
                                                                                                                                           (\f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int5_d [0] ? 12'd16 :
                                                                                                                                            (\f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int6_d [0] ? 12'd32 :
                                                                                                                                             (\f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int7_d [0] ? 12'd64 :
                                                                                                                                              (\f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int8_d [0] ? 12'd128 :
                                                                                                                                               (\f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int9_d [0] ? 12'd256 :
                                                                                                                                                (\f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int10_d [0] ? 12'd512 :
                                                                                                                                                 (\f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int11_d [0] ? 12'd1024 :
                                                                                                                                                  (\f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int12_d [0] ? 12'd2048 :
                                                                                                                                                   12'd0)))))))))))));
  logic [11:0] \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_select_q ;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_select_q  <= 12'd0;
    else
      \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_select_q  <= (\f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_done  ? 12'd0 :
                                                                                                                                     \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_select_d );
  logic [1:0] \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_emit_q ;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_emit_q  <= 2'd0;
    else
      \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_emit_q  <= (\f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_done  ? 2'd0 :
                                                                                                                                   \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_emit_d );
  logic [1:0] \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_emit_d ;
  assign \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_emit_d  = (\f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_emit_q  | ({\f''''''''''''_f''''''''''''_Int_choice_d [0],
                                                                                                                                                                                                                                                                  \f''''''''''''_f''''''''''''_Int_data_d [0]} & {\f''''''''''''_f''''''''''''_Int_choice_r ,
                                                                                                                                                                                                                                                                                                                  \f''''''''''''_f''''''''''''_Int_data_r }));
  logic \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_done ;
  assign \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_done  = (& \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_emit_d );
  assign {\f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int12_r ,
          \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int11_r ,
          \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int10_r ,
          \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int9_r ,
          \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int8_r ,
          \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int7_r ,
          \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int6_r ,
          \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int5_r ,
          \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int4_r ,
          \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int3_r ,
          \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int2_r ,
          \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_r } = (\f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_done  ? \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_select_d  :
                                                                                                                                  12'd0);
  assign \f''''''''''''_f''''''''''''_Int_data_d  = ((\f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_select_d [0] && (! \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_emit_q [0])) ? \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_d  :
                                                     ((\f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_select_d [1] && (! \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_emit_q [0])) ? \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int2_d  :
                                                      ((\f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_select_d [2] && (! \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_emit_q [0])) ? \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int3_d  :
                                                       ((\f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_select_d [3] && (! \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_emit_q [0])) ? \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int4_d  :
                                                        ((\f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_select_d [4] && (! \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_emit_q [0])) ? \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int5_d  :
                                                         ((\f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_select_d [5] && (! \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_emit_q [0])) ? \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int6_d  :
                                                          ((\f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_select_d [6] && (! \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_emit_q [0])) ? \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int7_d  :
                                                           ((\f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_select_d [7] && (! \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_emit_q [0])) ? \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int8_d  :
                                                            ((\f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_select_d [8] && (! \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_emit_q [0])) ? \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int9_d  :
                                                             ((\f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_select_d [9] && (! \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_emit_q [0])) ? \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int10_d  :
                                                              ((\f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_select_d [10] && (! \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_emit_q [0])) ? \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int11_d  :
                                                               ((\f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_select_d [11] && (! \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_emit_q [0])) ? \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int12_d  :
                                                                {32'd0, 1'd0}))))))))))));
  assign \f''''''''''''_f''''''''''''_Int_choice_d  = ((\f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_select_d [0] && (! \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_emit_q [1])) ? C1_12_dc(1'd1) :
                                                       ((\f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_select_d [1] && (! \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_emit_q [1])) ? C2_12_dc(1'd1) :
                                                        ((\f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_select_d [2] && (! \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_emit_q [1])) ? C3_12_dc(1'd1) :
                                                         ((\f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_select_d [3] && (! \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_emit_q [1])) ? C4_12_dc(1'd1) :
                                                          ((\f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_select_d [4] && (! \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_emit_q [1])) ? C5_12_dc(1'd1) :
                                                           ((\f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_select_d [5] && (! \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_emit_q [1])) ? C6_12_dc(1'd1) :
                                                            ((\f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_select_d [6] && (! \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_emit_q [1])) ? C7_12_dc(1'd1) :
                                                             ((\f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_select_d [7] && (! \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_emit_q [1])) ? C8_12_dc(1'd1) :
                                                              ((\f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_select_d [8] && (! \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_emit_q [1])) ? C9_12_dc(1'd1) :
                                                               ((\f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_select_d [9] && (! \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_emit_q [1])) ? C10_12_dc(1'd1) :
                                                                ((\f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_select_d [10] && (! \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_emit_q [1])) ? C11_12_dc(1'd1) :
                                                                 ((\f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_select_d [11] && (! \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_emit_q [1])) ? C12_12_dc(1'd1) :
                                                                  {4'd0, 1'd0}))))))))))));
  
  /* fork (Ty Go) : (f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intgo_11,Go) > [(go_11_1,Go),
                                                                                                                                          (go_11_2,Go)] */
  logic [1:0] \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intgo_11_emitted ;
  logic [1:0] \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intgo_11_done ;
  assign go_11_1_d = (\f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intgo_11_d [0] && (! \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intgo_11_emitted [0]));
  assign go_11_2_d = (\f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intgo_11_d [0] && (! \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intgo_11_emitted [1]));
  assign \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intgo_11_done  = (\f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intgo_11_emitted  | ({go_11_2_d[0],
                                                                                                                                                                                                                                                                       go_11_1_d[0]} & {go_11_2_r,
                                                                                                                                                                                                                                                                                        go_11_1_r}));
  assign \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intgo_11_r  = (& \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intgo_11_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intgo_11_emitted  <= 2'd0;
    else
      \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intgo_11_emitted  <= (\f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intgo_11_r  ? 2'd0 :
                                                                                                                                       \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intgo_11_done );
  
  /* buf (Ty MyDTInt_Bool) : (f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zafl_1,MyDTInt_Bool) > (is_zafl_1_1_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zafl_1_bufchan_d ;
  logic \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zafl_1_bufchan_r ;
  assign \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zafl_1_r  = ((! \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zafl_1_bufchan_d [0]) || \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zafl_1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zafl_1_bufchan_d  <= 1'd0;
    else
      if (\f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zafl_1_r )
        \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zafl_1_bufchan_d  <= \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zafl_1_d ;
  MyDTInt_Bool_t \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zafl_1_bufchan_buf ;
  assign \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zafl_1_bufchan_r  = (! \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zafl_1_bufchan_buf [0]);
  assign is_zafl_1_1_argbuf_d = (\f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zafl_1_bufchan_buf [0] ? \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zafl_1_bufchan_buf  :
                                 \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zafl_1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zafl_1_bufchan_buf  <= 1'd0;
    else
      if ((is_zafl_1_1_argbuf_r && \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zafl_1_bufchan_buf [0]))
        \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zafl_1_bufchan_buf  <= 1'd0;
      else if (((! is_zafl_1_1_argbuf_r) && (! \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zafl_1_bufchan_buf [0])))
        \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zafl_1_bufchan_buf  <= \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zafl_1_bufchan_d ;
  
  /* buf (Ty MyDTInt_Int_Int) : (f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addafm_1,MyDTInt_Int_Int) > (op_addafm_1_1_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addafm_1_bufchan_d ;
  logic \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addafm_1_bufchan_r ;
  assign \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addafm_1_r  = ((! \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addafm_1_bufchan_d [0]) || \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addafm_1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addafm_1_bufchan_d  <= 1'd0;
    else
      if (\f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addafm_1_r )
        \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addafm_1_bufchan_d  <= \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addafm_1_d ;
  MyDTInt_Int_Int_t \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addafm_1_bufchan_buf ;
  assign \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addafm_1_bufchan_r  = (! \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addafm_1_bufchan_buf [0]);
  assign op_addafm_1_1_argbuf_d = (\f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addafm_1_bufchan_buf [0] ? \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addafm_1_bufchan_buf  :
                                   \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addafm_1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addafm_1_bufchan_buf  <= 1'd0;
    else
      if ((op_addafm_1_1_argbuf_r && \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addafm_1_bufchan_buf [0]))
        \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addafm_1_bufchan_buf  <= 1'd0;
      else if (((! op_addafm_1_1_argbuf_r) && (! \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addafm_1_bufchan_buf [0])))
        \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addafm_1_bufchan_buf  <= \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addafm_1_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Int) : (f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intq4afj_1,Pointer_QTree_Int) > (q4afj_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intq4afj_1_bufchan_d ;
  logic \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intq4afj_1_bufchan_r ;
  assign \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intq4afj_1_r  = ((! \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intq4afj_1_bufchan_d [0]) || \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intq4afj_1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intq4afj_1_bufchan_d  <= {16'd0,
                                                                                                                                           1'd0};
    else
      if (\f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intq4afj_1_r )
        \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intq4afj_1_bufchan_d  <= \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intq4afj_1_d ;
  Pointer_QTree_Int_t \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intq4afj_1_bufchan_buf ;
  assign \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intq4afj_1_bufchan_r  = (! \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intq4afj_1_bufchan_buf [0]);
  assign q4afj_1_1_argbuf_d = (\f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intq4afj_1_bufchan_buf [0] ? \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intq4afj_1_bufchan_buf  :
                               \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intq4afj_1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intq4afj_1_bufchan_buf  <= {16'd0,
                                                                                                                                             1'd0};
    else
      if ((q4afj_1_1_argbuf_r && \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intq4afj_1_bufchan_buf [0]))
        \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intq4afj_1_bufchan_buf  <= {16'd0,
                                                                                                                                               1'd0};
      else if (((! q4afj_1_1_argbuf_r) && (! \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intq4afj_1_bufchan_buf [0])))
        \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intq4afj_1_bufchan_buf  <= \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intq4afj_1_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Int) : (f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intt4afk_1,Pointer_QTree_Int) > (t4afk_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intt4afk_1_bufchan_d ;
  logic \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intt4afk_1_bufchan_r ;
  assign \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intt4afk_1_r  = ((! \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intt4afk_1_bufchan_d [0]) || \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intt4afk_1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intt4afk_1_bufchan_d  <= {16'd0,
                                                                                                                                           1'd0};
    else
      if (\f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intt4afk_1_r )
        \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intt4afk_1_bufchan_d  <= \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intt4afk_1_d ;
  Pointer_QTree_Int_t \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intt4afk_1_bufchan_buf ;
  assign \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intt4afk_1_bufchan_r  = (! \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intt4afk_1_bufchan_buf [0]);
  assign t4afk_1_1_argbuf_d = (\f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intt4afk_1_bufchan_buf [0] ? \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intt4afk_1_bufchan_buf  :
                               \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intt4afk_1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intt4afk_1_bufchan_buf  <= {16'd0,
                                                                                                                                             1'd0};
    else
      if ((t4afk_1_1_argbuf_r && \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intt4afk_1_bufchan_buf [0]))
        \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intt4afk_1_bufchan_buf  <= {16'd0,
                                                                                                                                               1'd0};
      else if (((! t4afk_1_1_argbuf_r) && (! \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intt4afk_1_bufchan_buf [0])))
        \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intt4afk_1_bufchan_buf  <= \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intt4afk_1_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Int) : (f''''''''''''_f''''''''''''_Int_1,Pointer_QTree_Int) > (f''''''''''''_f''''''''''''_Int_resbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t \f''''''''''''_f''''''''''''_Int_1_bufchan_d ;
  logic \f''''''''''''_f''''''''''''_Int_1_bufchan_r ;
  assign \f''''''''''''_f''''''''''''_Int_1_r  = ((! \f''''''''''''_f''''''''''''_Int_1_bufchan_d [0]) || \f''''''''''''_f''''''''''''_Int_1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''''''_f''''''''''''_Int_1_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\f''''''''''''_f''''''''''''_Int_1_r )
        \f''''''''''''_f''''''''''''_Int_1_bufchan_d  <= \f''''''''''''_f''''''''''''_Int_1_d ;
  Pointer_QTree_Int_t \f''''''''''''_f''''''''''''_Int_1_bufchan_buf ;
  assign \f''''''''''''_f''''''''''''_Int_1_bufchan_r  = (! \f''''''''''''_f''''''''''''_Int_1_bufchan_buf [0]);
  assign \f''''''''''''_f''''''''''''_Int_resbuf_d  = (\f''''''''''''_f''''''''''''_Int_1_bufchan_buf [0] ? \f''''''''''''_f''''''''''''_Int_1_bufchan_buf  :
                                                       \f''''''''''''_f''''''''''''_Int_1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''''''_f''''''''''''_Int_1_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((\f''''''''''''_f''''''''''''_Int_resbuf_r  && \f''''''''''''_f''''''''''''_Int_1_bufchan_buf [0]))
        \f''''''''''''_f''''''''''''_Int_1_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! \f''''''''''''_f''''''''''''_Int_resbuf_r ) && (! \f''''''''''''_f''''''''''''_Int_1_bufchan_buf [0])))
        \f''''''''''''_f''''''''''''_Int_1_bufchan_buf  <= \f''''''''''''_f''''''''''''_Int_1_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Int) : (f''''''''''''_f''''''''''''_Int_10,Pointer_QTree_Int) > (f''''''''''''_f''''''''''''_Int_10_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t \f''''''''''''_f''''''''''''_Int_10_bufchan_d ;
  logic \f''''''''''''_f''''''''''''_Int_10_bufchan_r ;
  assign \f''''''''''''_f''''''''''''_Int_10_r  = ((! \f''''''''''''_f''''''''''''_Int_10_bufchan_d [0]) || \f''''''''''''_f''''''''''''_Int_10_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''''''_f''''''''''''_Int_10_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\f''''''''''''_f''''''''''''_Int_10_r )
        \f''''''''''''_f''''''''''''_Int_10_bufchan_d  <= \f''''''''''''_f''''''''''''_Int_10_d ;
  Pointer_QTree_Int_t \f''''''''''''_f''''''''''''_Int_10_bufchan_buf ;
  assign \f''''''''''''_f''''''''''''_Int_10_bufchan_r  = (! \f''''''''''''_f''''''''''''_Int_10_bufchan_buf [0]);
  assign \f''''''''''''_f''''''''''''_Int_10_argbuf_d  = (\f''''''''''''_f''''''''''''_Int_10_bufchan_buf [0] ? \f''''''''''''_f''''''''''''_Int_10_bufchan_buf  :
                                                          \f''''''''''''_f''''''''''''_Int_10_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''''''_f''''''''''''_Int_10_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((\f''''''''''''_f''''''''''''_Int_10_argbuf_r  && \f''''''''''''_f''''''''''''_Int_10_bufchan_buf [0]))
        \f''''''''''''_f''''''''''''_Int_10_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! \f''''''''''''_f''''''''''''_Int_10_argbuf_r ) && (! \f''''''''''''_f''''''''''''_Int_10_bufchan_buf [0])))
        \f''''''''''''_f''''''''''''_Int_10_bufchan_buf  <= \f''''''''''''_f''''''''''''_Int_10_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Int) : (f''''''''''''_f''''''''''''_Int_11,Pointer_QTree_Int) > (f''''''''''''_f''''''''''''_Int_11_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t \f''''''''''''_f''''''''''''_Int_11_bufchan_d ;
  logic \f''''''''''''_f''''''''''''_Int_11_bufchan_r ;
  assign \f''''''''''''_f''''''''''''_Int_11_r  = ((! \f''''''''''''_f''''''''''''_Int_11_bufchan_d [0]) || \f''''''''''''_f''''''''''''_Int_11_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''''''_f''''''''''''_Int_11_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\f''''''''''''_f''''''''''''_Int_11_r )
        \f''''''''''''_f''''''''''''_Int_11_bufchan_d  <= \f''''''''''''_f''''''''''''_Int_11_d ;
  Pointer_QTree_Int_t \f''''''''''''_f''''''''''''_Int_11_bufchan_buf ;
  assign \f''''''''''''_f''''''''''''_Int_11_bufchan_r  = (! \f''''''''''''_f''''''''''''_Int_11_bufchan_buf [0]);
  assign \f''''''''''''_f''''''''''''_Int_11_argbuf_d  = (\f''''''''''''_f''''''''''''_Int_11_bufchan_buf [0] ? \f''''''''''''_f''''''''''''_Int_11_bufchan_buf  :
                                                          \f''''''''''''_f''''''''''''_Int_11_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''''''_f''''''''''''_Int_11_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((\f''''''''''''_f''''''''''''_Int_11_argbuf_r  && \f''''''''''''_f''''''''''''_Int_11_bufchan_buf [0]))
        \f''''''''''''_f''''''''''''_Int_11_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! \f''''''''''''_f''''''''''''_Int_11_argbuf_r ) && (! \f''''''''''''_f''''''''''''_Int_11_bufchan_buf [0])))
        \f''''''''''''_f''''''''''''_Int_11_bufchan_buf  <= \f''''''''''''_f''''''''''''_Int_11_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Int) : (f''''''''''''_f''''''''''''_Int_12,Pointer_QTree_Int) > (f''''''''''''_f''''''''''''_Int_12_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t \f''''''''''''_f''''''''''''_Int_12_bufchan_d ;
  logic \f''''''''''''_f''''''''''''_Int_12_bufchan_r ;
  assign \f''''''''''''_f''''''''''''_Int_12_r  = ((! \f''''''''''''_f''''''''''''_Int_12_bufchan_d [0]) || \f''''''''''''_f''''''''''''_Int_12_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''''''_f''''''''''''_Int_12_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\f''''''''''''_f''''''''''''_Int_12_r )
        \f''''''''''''_f''''''''''''_Int_12_bufchan_d  <= \f''''''''''''_f''''''''''''_Int_12_d ;
  Pointer_QTree_Int_t \f''''''''''''_f''''''''''''_Int_12_bufchan_buf ;
  assign \f''''''''''''_f''''''''''''_Int_12_bufchan_r  = (! \f''''''''''''_f''''''''''''_Int_12_bufchan_buf [0]);
  assign \f''''''''''''_f''''''''''''_Int_12_argbuf_d  = (\f''''''''''''_f''''''''''''_Int_12_bufchan_buf [0] ? \f''''''''''''_f''''''''''''_Int_12_bufchan_buf  :
                                                          \f''''''''''''_f''''''''''''_Int_12_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''''''_f''''''''''''_Int_12_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((\f''''''''''''_f''''''''''''_Int_12_argbuf_r  && \f''''''''''''_f''''''''''''_Int_12_bufchan_buf [0]))
        \f''''''''''''_f''''''''''''_Int_12_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! \f''''''''''''_f''''''''''''_Int_12_argbuf_r ) && (! \f''''''''''''_f''''''''''''_Int_12_bufchan_buf [0])))
        \f''''''''''''_f''''''''''''_Int_12_bufchan_buf  <= \f''''''''''''_f''''''''''''_Int_12_bufchan_d ;
  
  /* dcon (Ty QTree_Int,
      Dcon QNode_Int) : [(f''''''''''''_f''''''''''''_Int_12_argbuf,Pointer_QTree_Int),
                         (f''''''''''''_f''''''''''''_Int_11_argbuf,Pointer_QTree_Int),
                         (f''''''''''''_f''''''''''''_Int_10_argbuf,Pointer_QTree_Int),
                         (f''''''''''''_f''''''''''''_Int_9_argbuf,Pointer_QTree_Int)] > (es_30_1es_31_1es_32_1es_33_1QNode_Int,QTree_Int) */
  assign es_30_1es_31_1es_32_1es_33_1QNode_Int_d = QNode_Int_dc((& {\f''''''''''''_f''''''''''''_Int_12_argbuf_d [0],
                                                                    \f''''''''''''_f''''''''''''_Int_11_argbuf_d [0],
                                                                    \f''''''''''''_f''''''''''''_Int_10_argbuf_d [0],
                                                                    \f''''''''''''_f''''''''''''_Int_9_argbuf_d [0]}), \f''''''''''''_f''''''''''''_Int_12_argbuf_d , \f''''''''''''_f''''''''''''_Int_11_argbuf_d , \f''''''''''''_f''''''''''''_Int_10_argbuf_d , \f''''''''''''_f''''''''''''_Int_9_argbuf_d );
  assign {\f''''''''''''_f''''''''''''_Int_12_argbuf_r ,
          \f''''''''''''_f''''''''''''_Int_11_argbuf_r ,
          \f''''''''''''_f''''''''''''_Int_10_argbuf_r ,
          \f''''''''''''_f''''''''''''_Int_9_argbuf_r } = {4 {(es_30_1es_31_1es_32_1es_33_1QNode_Int_r && es_30_1es_31_1es_32_1es_33_1QNode_Int_d[0])}};
  
  /* buf (Ty Pointer_QTree_Int) : (f''''''''''''_f''''''''''''_Int_2,Pointer_QTree_Int) > (f''''''''''''_f''''''''''''_Int_2_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t \f''''''''''''_f''''''''''''_Int_2_bufchan_d ;
  logic \f''''''''''''_f''''''''''''_Int_2_bufchan_r ;
  assign \f''''''''''''_f''''''''''''_Int_2_r  = ((! \f''''''''''''_f''''''''''''_Int_2_bufchan_d [0]) || \f''''''''''''_f''''''''''''_Int_2_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''''''_f''''''''''''_Int_2_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\f''''''''''''_f''''''''''''_Int_2_r )
        \f''''''''''''_f''''''''''''_Int_2_bufchan_d  <= \f''''''''''''_f''''''''''''_Int_2_d ;
  Pointer_QTree_Int_t \f''''''''''''_f''''''''''''_Int_2_bufchan_buf ;
  assign \f''''''''''''_f''''''''''''_Int_2_bufchan_r  = (! \f''''''''''''_f''''''''''''_Int_2_bufchan_buf [0]);
  assign \f''''''''''''_f''''''''''''_Int_2_argbuf_d  = (\f''''''''''''_f''''''''''''_Int_2_bufchan_buf [0] ? \f''''''''''''_f''''''''''''_Int_2_bufchan_buf  :
                                                         \f''''''''''''_f''''''''''''_Int_2_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''''''_f''''''''''''_Int_2_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((\f''''''''''''_f''''''''''''_Int_2_argbuf_r  && \f''''''''''''_f''''''''''''_Int_2_bufchan_buf [0]))
        \f''''''''''''_f''''''''''''_Int_2_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! \f''''''''''''_f''''''''''''_Int_2_argbuf_r ) && (! \f''''''''''''_f''''''''''''_Int_2_bufchan_buf [0])))
        \f''''''''''''_f''''''''''''_Int_2_bufchan_buf  <= \f''''''''''''_f''''''''''''_Int_2_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Int) : (f''''''''''''_f''''''''''''_Int_3,Pointer_QTree_Int) > (f''''''''''''_f''''''''''''_Int_3_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t \f''''''''''''_f''''''''''''_Int_3_bufchan_d ;
  logic \f''''''''''''_f''''''''''''_Int_3_bufchan_r ;
  assign \f''''''''''''_f''''''''''''_Int_3_r  = ((! \f''''''''''''_f''''''''''''_Int_3_bufchan_d [0]) || \f''''''''''''_f''''''''''''_Int_3_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''''''_f''''''''''''_Int_3_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\f''''''''''''_f''''''''''''_Int_3_r )
        \f''''''''''''_f''''''''''''_Int_3_bufchan_d  <= \f''''''''''''_f''''''''''''_Int_3_d ;
  Pointer_QTree_Int_t \f''''''''''''_f''''''''''''_Int_3_bufchan_buf ;
  assign \f''''''''''''_f''''''''''''_Int_3_bufchan_r  = (! \f''''''''''''_f''''''''''''_Int_3_bufchan_buf [0]);
  assign \f''''''''''''_f''''''''''''_Int_3_argbuf_d  = (\f''''''''''''_f''''''''''''_Int_3_bufchan_buf [0] ? \f''''''''''''_f''''''''''''_Int_3_bufchan_buf  :
                                                         \f''''''''''''_f''''''''''''_Int_3_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''''''_f''''''''''''_Int_3_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((\f''''''''''''_f''''''''''''_Int_3_argbuf_r  && \f''''''''''''_f''''''''''''_Int_3_bufchan_buf [0]))
        \f''''''''''''_f''''''''''''_Int_3_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! \f''''''''''''_f''''''''''''_Int_3_argbuf_r ) && (! \f''''''''''''_f''''''''''''_Int_3_bufchan_buf [0])))
        \f''''''''''''_f''''''''''''_Int_3_bufchan_buf  <= \f''''''''''''_f''''''''''''_Int_3_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Int) : (f''''''''''''_f''''''''''''_Int_4,Pointer_QTree_Int) > (f''''''''''''_f''''''''''''_Int_4_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t \f''''''''''''_f''''''''''''_Int_4_bufchan_d ;
  logic \f''''''''''''_f''''''''''''_Int_4_bufchan_r ;
  assign \f''''''''''''_f''''''''''''_Int_4_r  = ((! \f''''''''''''_f''''''''''''_Int_4_bufchan_d [0]) || \f''''''''''''_f''''''''''''_Int_4_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''''''_f''''''''''''_Int_4_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\f''''''''''''_f''''''''''''_Int_4_r )
        \f''''''''''''_f''''''''''''_Int_4_bufchan_d  <= \f''''''''''''_f''''''''''''_Int_4_d ;
  Pointer_QTree_Int_t \f''''''''''''_f''''''''''''_Int_4_bufchan_buf ;
  assign \f''''''''''''_f''''''''''''_Int_4_bufchan_r  = (! \f''''''''''''_f''''''''''''_Int_4_bufchan_buf [0]);
  assign \f''''''''''''_f''''''''''''_Int_4_argbuf_d  = (\f''''''''''''_f''''''''''''_Int_4_bufchan_buf [0] ? \f''''''''''''_f''''''''''''_Int_4_bufchan_buf  :
                                                         \f''''''''''''_f''''''''''''_Int_4_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''''''_f''''''''''''_Int_4_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((\f''''''''''''_f''''''''''''_Int_4_argbuf_r  && \f''''''''''''_f''''''''''''_Int_4_bufchan_buf [0]))
        \f''''''''''''_f''''''''''''_Int_4_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! \f''''''''''''_f''''''''''''_Int_4_argbuf_r ) && (! \f''''''''''''_f''''''''''''_Int_4_bufchan_buf [0])))
        \f''''''''''''_f''''''''''''_Int_4_bufchan_buf  <= \f''''''''''''_f''''''''''''_Int_4_bufchan_d ;
  
  /* dcon (Ty QTree_Int,
      Dcon QNode_Int) : [(f''''''''''''_f''''''''''''_Int_4_argbuf,Pointer_QTree_Int),
                         (f''''''''''''_f''''''''''''_Int_3_argbuf,Pointer_QTree_Int),
                         (f''''''''''''_f''''''''''''_Int_2_argbuf,Pointer_QTree_Int),
                         (f''''''''''''_f''''''''''''_Int_resbuf,Pointer_QTree_Int)] > (es_4_1_1es_5_1_1es_6_1_1es_7_1QNode_Int,QTree_Int) */
  assign es_4_1_1es_5_1_1es_6_1_1es_7_1QNode_Int_d = QNode_Int_dc((& {\f''''''''''''_f''''''''''''_Int_4_argbuf_d [0],
                                                                      \f''''''''''''_f''''''''''''_Int_3_argbuf_d [0],
                                                                      \f''''''''''''_f''''''''''''_Int_2_argbuf_d [0],
                                                                      \f''''''''''''_f''''''''''''_Int_resbuf_d [0]}), \f''''''''''''_f''''''''''''_Int_4_argbuf_d , \f''''''''''''_f''''''''''''_Int_3_argbuf_d , \f''''''''''''_f''''''''''''_Int_2_argbuf_d , \f''''''''''''_f''''''''''''_Int_resbuf_d );
  assign {\f''''''''''''_f''''''''''''_Int_4_argbuf_r ,
          \f''''''''''''_f''''''''''''_Int_3_argbuf_r ,
          \f''''''''''''_f''''''''''''_Int_2_argbuf_r ,
          \f''''''''''''_f''''''''''''_Int_resbuf_r } = {4 {(es_4_1_1es_5_1_1es_6_1_1es_7_1QNode_Int_r && es_4_1_1es_5_1_1es_6_1_1es_7_1QNode_Int_d[0])}};
  
  /* buf (Ty Pointer_QTree_Int) : (f''''''''''''_f''''''''''''_Int_5,Pointer_QTree_Int) > (f''''''''''''_f''''''''''''_Int_5_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t \f''''''''''''_f''''''''''''_Int_5_bufchan_d ;
  logic \f''''''''''''_f''''''''''''_Int_5_bufchan_r ;
  assign \f''''''''''''_f''''''''''''_Int_5_r  = ((! \f''''''''''''_f''''''''''''_Int_5_bufchan_d [0]) || \f''''''''''''_f''''''''''''_Int_5_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''''''_f''''''''''''_Int_5_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\f''''''''''''_f''''''''''''_Int_5_r )
        \f''''''''''''_f''''''''''''_Int_5_bufchan_d  <= \f''''''''''''_f''''''''''''_Int_5_d ;
  Pointer_QTree_Int_t \f''''''''''''_f''''''''''''_Int_5_bufchan_buf ;
  assign \f''''''''''''_f''''''''''''_Int_5_bufchan_r  = (! \f''''''''''''_f''''''''''''_Int_5_bufchan_buf [0]);
  assign \f''''''''''''_f''''''''''''_Int_5_argbuf_d  = (\f''''''''''''_f''''''''''''_Int_5_bufchan_buf [0] ? \f''''''''''''_f''''''''''''_Int_5_bufchan_buf  :
                                                         \f''''''''''''_f''''''''''''_Int_5_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''''''_f''''''''''''_Int_5_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((\f''''''''''''_f''''''''''''_Int_5_argbuf_r  && \f''''''''''''_f''''''''''''_Int_5_bufchan_buf [0]))
        \f''''''''''''_f''''''''''''_Int_5_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! \f''''''''''''_f''''''''''''_Int_5_argbuf_r ) && (! \f''''''''''''_f''''''''''''_Int_5_bufchan_buf [0])))
        \f''''''''''''_f''''''''''''_Int_5_bufchan_buf  <= \f''''''''''''_f''''''''''''_Int_5_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Int) : (f''''''''''''_f''''''''''''_Int_6,Pointer_QTree_Int) > (f''''''''''''_f''''''''''''_Int_6_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t \f''''''''''''_f''''''''''''_Int_6_bufchan_d ;
  logic \f''''''''''''_f''''''''''''_Int_6_bufchan_r ;
  assign \f''''''''''''_f''''''''''''_Int_6_r  = ((! \f''''''''''''_f''''''''''''_Int_6_bufchan_d [0]) || \f''''''''''''_f''''''''''''_Int_6_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''''''_f''''''''''''_Int_6_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\f''''''''''''_f''''''''''''_Int_6_r )
        \f''''''''''''_f''''''''''''_Int_6_bufchan_d  <= \f''''''''''''_f''''''''''''_Int_6_d ;
  Pointer_QTree_Int_t \f''''''''''''_f''''''''''''_Int_6_bufchan_buf ;
  assign \f''''''''''''_f''''''''''''_Int_6_bufchan_r  = (! \f''''''''''''_f''''''''''''_Int_6_bufchan_buf [0]);
  assign \f''''''''''''_f''''''''''''_Int_6_argbuf_d  = (\f''''''''''''_f''''''''''''_Int_6_bufchan_buf [0] ? \f''''''''''''_f''''''''''''_Int_6_bufchan_buf  :
                                                         \f''''''''''''_f''''''''''''_Int_6_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''''''_f''''''''''''_Int_6_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((\f''''''''''''_f''''''''''''_Int_6_argbuf_r  && \f''''''''''''_f''''''''''''_Int_6_bufchan_buf [0]))
        \f''''''''''''_f''''''''''''_Int_6_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! \f''''''''''''_f''''''''''''_Int_6_argbuf_r ) && (! \f''''''''''''_f''''''''''''_Int_6_bufchan_buf [0])))
        \f''''''''''''_f''''''''''''_Int_6_bufchan_buf  <= \f''''''''''''_f''''''''''''_Int_6_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Int) : (f''''''''''''_f''''''''''''_Int_7,Pointer_QTree_Int) > (f''''''''''''_f''''''''''''_Int_7_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t \f''''''''''''_f''''''''''''_Int_7_bufchan_d ;
  logic \f''''''''''''_f''''''''''''_Int_7_bufchan_r ;
  assign \f''''''''''''_f''''''''''''_Int_7_r  = ((! \f''''''''''''_f''''''''''''_Int_7_bufchan_d [0]) || \f''''''''''''_f''''''''''''_Int_7_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''''''_f''''''''''''_Int_7_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\f''''''''''''_f''''''''''''_Int_7_r )
        \f''''''''''''_f''''''''''''_Int_7_bufchan_d  <= \f''''''''''''_f''''''''''''_Int_7_d ;
  Pointer_QTree_Int_t \f''''''''''''_f''''''''''''_Int_7_bufchan_buf ;
  assign \f''''''''''''_f''''''''''''_Int_7_bufchan_r  = (! \f''''''''''''_f''''''''''''_Int_7_bufchan_buf [0]);
  assign \f''''''''''''_f''''''''''''_Int_7_argbuf_d  = (\f''''''''''''_f''''''''''''_Int_7_bufchan_buf [0] ? \f''''''''''''_f''''''''''''_Int_7_bufchan_buf  :
                                                         \f''''''''''''_f''''''''''''_Int_7_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''''''_f''''''''''''_Int_7_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((\f''''''''''''_f''''''''''''_Int_7_argbuf_r  && \f''''''''''''_f''''''''''''_Int_7_bufchan_buf [0]))
        \f''''''''''''_f''''''''''''_Int_7_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! \f''''''''''''_f''''''''''''_Int_7_argbuf_r ) && (! \f''''''''''''_f''''''''''''_Int_7_bufchan_buf [0])))
        \f''''''''''''_f''''''''''''_Int_7_bufchan_buf  <= \f''''''''''''_f''''''''''''_Int_7_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Int) : (f''''''''''''_f''''''''''''_Int_8,Pointer_QTree_Int) > (f''''''''''''_f''''''''''''_Int_8_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t \f''''''''''''_f''''''''''''_Int_8_bufchan_d ;
  logic \f''''''''''''_f''''''''''''_Int_8_bufchan_r ;
  assign \f''''''''''''_f''''''''''''_Int_8_r  = ((! \f''''''''''''_f''''''''''''_Int_8_bufchan_d [0]) || \f''''''''''''_f''''''''''''_Int_8_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''''''_f''''''''''''_Int_8_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\f''''''''''''_f''''''''''''_Int_8_r )
        \f''''''''''''_f''''''''''''_Int_8_bufchan_d  <= \f''''''''''''_f''''''''''''_Int_8_d ;
  Pointer_QTree_Int_t \f''''''''''''_f''''''''''''_Int_8_bufchan_buf ;
  assign \f''''''''''''_f''''''''''''_Int_8_bufchan_r  = (! \f''''''''''''_f''''''''''''_Int_8_bufchan_buf [0]);
  assign \f''''''''''''_f''''''''''''_Int_8_argbuf_d  = (\f''''''''''''_f''''''''''''_Int_8_bufchan_buf [0] ? \f''''''''''''_f''''''''''''_Int_8_bufchan_buf  :
                                                         \f''''''''''''_f''''''''''''_Int_8_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''''''_f''''''''''''_Int_8_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((\f''''''''''''_f''''''''''''_Int_8_argbuf_r  && \f''''''''''''_f''''''''''''_Int_8_bufchan_buf [0]))
        \f''''''''''''_f''''''''''''_Int_8_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! \f''''''''''''_f''''''''''''_Int_8_argbuf_r ) && (! \f''''''''''''_f''''''''''''_Int_8_bufchan_buf [0])))
        \f''''''''''''_f''''''''''''_Int_8_bufchan_buf  <= \f''''''''''''_f''''''''''''_Int_8_bufchan_d ;
  
  /* dcon (Ty QTree_Int,
      Dcon QNode_Int) : [(f''''''''''''_f''''''''''''_Int_8_argbuf,Pointer_QTree_Int),
                         (f''''''''''''_f''''''''''''_Int_7_argbuf,Pointer_QTree_Int),
                         (f''''''''''''_f''''''''''''_Int_6_argbuf,Pointer_QTree_Int),
                         (f''''''''''''_f''''''''''''_Int_5_argbuf,Pointer_QTree_Int)] > (es_26_1es_27_1es_28_1es_29_1QNode_Int,QTree_Int) */
  assign es_26_1es_27_1es_28_1es_29_1QNode_Int_d = QNode_Int_dc((& {\f''''''''''''_f''''''''''''_Int_8_argbuf_d [0],
                                                                    \f''''''''''''_f''''''''''''_Int_7_argbuf_d [0],
                                                                    \f''''''''''''_f''''''''''''_Int_6_argbuf_d [0],
                                                                    \f''''''''''''_f''''''''''''_Int_5_argbuf_d [0]}), \f''''''''''''_f''''''''''''_Int_8_argbuf_d , \f''''''''''''_f''''''''''''_Int_7_argbuf_d , \f''''''''''''_f''''''''''''_Int_6_argbuf_d , \f''''''''''''_f''''''''''''_Int_5_argbuf_d );
  assign {\f''''''''''''_f''''''''''''_Int_8_argbuf_r ,
          \f''''''''''''_f''''''''''''_Int_7_argbuf_r ,
          \f''''''''''''_f''''''''''''_Int_6_argbuf_r ,
          \f''''''''''''_f''''''''''''_Int_5_argbuf_r } = {4 {(es_26_1es_27_1es_28_1es_29_1QNode_Int_r && es_26_1es_27_1es_28_1es_29_1QNode_Int_d[0])}};
  
  /* buf (Ty Pointer_QTree_Int) : (f''''''''''''_f''''''''''''_Int_9,Pointer_QTree_Int) > (f''''''''''''_f''''''''''''_Int_9_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t \f''''''''''''_f''''''''''''_Int_9_bufchan_d ;
  logic \f''''''''''''_f''''''''''''_Int_9_bufchan_r ;
  assign \f''''''''''''_f''''''''''''_Int_9_r  = ((! \f''''''''''''_f''''''''''''_Int_9_bufchan_d [0]) || \f''''''''''''_f''''''''''''_Int_9_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''''''_f''''''''''''_Int_9_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\f''''''''''''_f''''''''''''_Int_9_r )
        \f''''''''''''_f''''''''''''_Int_9_bufchan_d  <= \f''''''''''''_f''''''''''''_Int_9_d ;
  Pointer_QTree_Int_t \f''''''''''''_f''''''''''''_Int_9_bufchan_buf ;
  assign \f''''''''''''_f''''''''''''_Int_9_bufchan_r  = (! \f''''''''''''_f''''''''''''_Int_9_bufchan_buf [0]);
  assign \f''''''''''''_f''''''''''''_Int_9_argbuf_d  = (\f''''''''''''_f''''''''''''_Int_9_bufchan_buf [0] ? \f''''''''''''_f''''''''''''_Int_9_bufchan_buf  :
                                                         \f''''''''''''_f''''''''''''_Int_9_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''''''_f''''''''''''_Int_9_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((\f''''''''''''_f''''''''''''_Int_9_argbuf_r  && \f''''''''''''_f''''''''''''_Int_9_bufchan_buf [0]))
        \f''''''''''''_f''''''''''''_Int_9_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! \f''''''''''''_f''''''''''''_Int_9_argbuf_r ) && (! \f''''''''''''_f''''''''''''_Int_9_bufchan_buf [0])))
        \f''''''''''''_f''''''''''''_Int_9_bufchan_buf  <= \f''''''''''''_f''''''''''''_Int_9_bufchan_d ;
  
  /* demux (Ty C12,
       Ty Pointer_QTree_Int) : (f''''''''''''_f''''''''''''_Int_choice,C12) (lizzieLet62_4Lf''''''''''''_f''''''''''''_Intsbos_1_merge_merge_fork_2,Pointer_QTree_Int) > [(f''''''''''''_f''''''''''''_Int_1,Pointer_QTree_Int),
                                                                                                                                                                          (f''''''''''''_f''''''''''''_Int_2,Pointer_QTree_Int),
                                                                                                                                                                          (f''''''''''''_f''''''''''''_Int_3,Pointer_QTree_Int),
                                                                                                                                                                          (f''''''''''''_f''''''''''''_Int_4,Pointer_QTree_Int),
                                                                                                                                                                          (f''''''''''''_f''''''''''''_Int_5,Pointer_QTree_Int),
                                                                                                                                                                          (f''''''''''''_f''''''''''''_Int_6,Pointer_QTree_Int),
                                                                                                                                                                          (f''''''''''''_f''''''''''''_Int_7,Pointer_QTree_Int),
                                                                                                                                                                          (f''''''''''''_f''''''''''''_Int_8,Pointer_QTree_Int),
                                                                                                                                                                          (f''''''''''''_f''''''''''''_Int_9,Pointer_QTree_Int),
                                                                                                                                                                          (f''''''''''''_f''''''''''''_Int_10,Pointer_QTree_Int),
                                                                                                                                                                          (f''''''''''''_f''''''''''''_Int_11,Pointer_QTree_Int),
                                                                                                                                                                          (f''''''''''''_f''''''''''''_Int_12,Pointer_QTree_Int)] */
  logic [11:0] \lizzieLet62_4Lf''''''''''''_f''''''''''''_Intsbos_1_merge_merge_fork_2_onehotd ;
  always_comb
    if ((\f''''''''''''_f''''''''''''_Int_choice_d [0] && \lizzieLet62_4Lf''''''''''''_f''''''''''''_Intsbos_1_merge_merge_fork_2_d [0]))
      unique case (\f''''''''''''_f''''''''''''_Int_choice_d [4:1])
        4'd0:
          \lizzieLet62_4Lf''''''''''''_f''''''''''''_Intsbos_1_merge_merge_fork_2_onehotd  = 12'd1;
        4'd1:
          \lizzieLet62_4Lf''''''''''''_f''''''''''''_Intsbos_1_merge_merge_fork_2_onehotd  = 12'd2;
        4'd2:
          \lizzieLet62_4Lf''''''''''''_f''''''''''''_Intsbos_1_merge_merge_fork_2_onehotd  = 12'd4;
        4'd3:
          \lizzieLet62_4Lf''''''''''''_f''''''''''''_Intsbos_1_merge_merge_fork_2_onehotd  = 12'd8;
        4'd4:
          \lizzieLet62_4Lf''''''''''''_f''''''''''''_Intsbos_1_merge_merge_fork_2_onehotd  = 12'd16;
        4'd5:
          \lizzieLet62_4Lf''''''''''''_f''''''''''''_Intsbos_1_merge_merge_fork_2_onehotd  = 12'd32;
        4'd6:
          \lizzieLet62_4Lf''''''''''''_f''''''''''''_Intsbos_1_merge_merge_fork_2_onehotd  = 12'd64;
        4'd7:
          \lizzieLet62_4Lf''''''''''''_f''''''''''''_Intsbos_1_merge_merge_fork_2_onehotd  = 12'd128;
        4'd8:
          \lizzieLet62_4Lf''''''''''''_f''''''''''''_Intsbos_1_merge_merge_fork_2_onehotd  = 12'd256;
        4'd9:
          \lizzieLet62_4Lf''''''''''''_f''''''''''''_Intsbos_1_merge_merge_fork_2_onehotd  = 12'd512;
        4'd10:
          \lizzieLet62_4Lf''''''''''''_f''''''''''''_Intsbos_1_merge_merge_fork_2_onehotd  = 12'd1024;
        4'd11:
          \lizzieLet62_4Lf''''''''''''_f''''''''''''_Intsbos_1_merge_merge_fork_2_onehotd  = 12'd2048;
        default:
          \lizzieLet62_4Lf''''''''''''_f''''''''''''_Intsbos_1_merge_merge_fork_2_onehotd  = 12'd0;
      endcase
    else
      \lizzieLet62_4Lf''''''''''''_f''''''''''''_Intsbos_1_merge_merge_fork_2_onehotd  = 12'd0;
  assign \f''''''''''''_f''''''''''''_Int_1_d  = {\lizzieLet62_4Lf''''''''''''_f''''''''''''_Intsbos_1_merge_merge_fork_2_d [16:1],
                                                  \lizzieLet62_4Lf''''''''''''_f''''''''''''_Intsbos_1_merge_merge_fork_2_onehotd [0]};
  assign \f''''''''''''_f''''''''''''_Int_2_d  = {\lizzieLet62_4Lf''''''''''''_f''''''''''''_Intsbos_1_merge_merge_fork_2_d [16:1],
                                                  \lizzieLet62_4Lf''''''''''''_f''''''''''''_Intsbos_1_merge_merge_fork_2_onehotd [1]};
  assign \f''''''''''''_f''''''''''''_Int_3_d  = {\lizzieLet62_4Lf''''''''''''_f''''''''''''_Intsbos_1_merge_merge_fork_2_d [16:1],
                                                  \lizzieLet62_4Lf''''''''''''_f''''''''''''_Intsbos_1_merge_merge_fork_2_onehotd [2]};
  assign \f''''''''''''_f''''''''''''_Int_4_d  = {\lizzieLet62_4Lf''''''''''''_f''''''''''''_Intsbos_1_merge_merge_fork_2_d [16:1],
                                                  \lizzieLet62_4Lf''''''''''''_f''''''''''''_Intsbos_1_merge_merge_fork_2_onehotd [3]};
  assign \f''''''''''''_f''''''''''''_Int_5_d  = {\lizzieLet62_4Lf''''''''''''_f''''''''''''_Intsbos_1_merge_merge_fork_2_d [16:1],
                                                  \lizzieLet62_4Lf''''''''''''_f''''''''''''_Intsbos_1_merge_merge_fork_2_onehotd [4]};
  assign \f''''''''''''_f''''''''''''_Int_6_d  = {\lizzieLet62_4Lf''''''''''''_f''''''''''''_Intsbos_1_merge_merge_fork_2_d [16:1],
                                                  \lizzieLet62_4Lf''''''''''''_f''''''''''''_Intsbos_1_merge_merge_fork_2_onehotd [5]};
  assign \f''''''''''''_f''''''''''''_Int_7_d  = {\lizzieLet62_4Lf''''''''''''_f''''''''''''_Intsbos_1_merge_merge_fork_2_d [16:1],
                                                  \lizzieLet62_4Lf''''''''''''_f''''''''''''_Intsbos_1_merge_merge_fork_2_onehotd [6]};
  assign \f''''''''''''_f''''''''''''_Int_8_d  = {\lizzieLet62_4Lf''''''''''''_f''''''''''''_Intsbos_1_merge_merge_fork_2_d [16:1],
                                                  \lizzieLet62_4Lf''''''''''''_f''''''''''''_Intsbos_1_merge_merge_fork_2_onehotd [7]};
  assign \f''''''''''''_f''''''''''''_Int_9_d  = {\lizzieLet62_4Lf''''''''''''_f''''''''''''_Intsbos_1_merge_merge_fork_2_d [16:1],
                                                  \lizzieLet62_4Lf''''''''''''_f''''''''''''_Intsbos_1_merge_merge_fork_2_onehotd [8]};
  assign \f''''''''''''_f''''''''''''_Int_10_d  = {\lizzieLet62_4Lf''''''''''''_f''''''''''''_Intsbos_1_merge_merge_fork_2_d [16:1],
                                                   \lizzieLet62_4Lf''''''''''''_f''''''''''''_Intsbos_1_merge_merge_fork_2_onehotd [9]};
  assign \f''''''''''''_f''''''''''''_Int_11_d  = {\lizzieLet62_4Lf''''''''''''_f''''''''''''_Intsbos_1_merge_merge_fork_2_d [16:1],
                                                   \lizzieLet62_4Lf''''''''''''_f''''''''''''_Intsbos_1_merge_merge_fork_2_onehotd [10]};
  assign \f''''''''''''_f''''''''''''_Int_12_d  = {\lizzieLet62_4Lf''''''''''''_f''''''''''''_Intsbos_1_merge_merge_fork_2_d [16:1],
                                                   \lizzieLet62_4Lf''''''''''''_f''''''''''''_Intsbos_1_merge_merge_fork_2_onehotd [11]};
  assign \lizzieLet62_4Lf''''''''''''_f''''''''''''_Intsbos_1_merge_merge_fork_2_r  = (| (\lizzieLet62_4Lf''''''''''''_f''''''''''''_Intsbos_1_merge_merge_fork_2_onehotd  & {\f''''''''''''_f''''''''''''_Int_12_r ,
                                                                                                                                                                              \f''''''''''''_f''''''''''''_Int_11_r ,
                                                                                                                                                                              \f''''''''''''_f''''''''''''_Int_10_r ,
                                                                                                                                                                              \f''''''''''''_f''''''''''''_Int_9_r ,
                                                                                                                                                                              \f''''''''''''_f''''''''''''_Int_8_r ,
                                                                                                                                                                              \f''''''''''''_f''''''''''''_Int_7_r ,
                                                                                                                                                                              \f''''''''''''_f''''''''''''_Int_6_r ,
                                                                                                                                                                              \f''''''''''''_f''''''''''''_Int_5_r ,
                                                                                                                                                                              \f''''''''''''_f''''''''''''_Int_4_r ,
                                                                                                                                                                              \f''''''''''''_f''''''''''''_Int_3_r ,
                                                                                                                                                                              \f''''''''''''_f''''''''''''_Int_2_r ,
                                                                                                                                                                              \f''''''''''''_f''''''''''''_Int_1_r }));
  assign \f''''''''''''_f''''''''''''_Int_choice_r  = \lizzieLet62_4Lf''''''''''''_f''''''''''''_Intsbos_1_merge_merge_fork_2_r ;
  
  /* destruct (Ty TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int,
          Dcon TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int) : (f''''''''''''_f''''''''''''_Int_data,TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int) > [(f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intgo_11,Go),
                                                                                                                                                                                                                          (f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intq4afj_1,Pointer_QTree_Int),
                                                                                                                                                                                                                          (f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intt4afk_1,Pointer_QTree_Int),
                                                                                                                                                                                                                          (f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zafl_1,MyDTInt_Bool),
                                                                                                                                                                                                                          (f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addafm_1,MyDTInt_Int_Int)] */
  logic [4:0] \f''''''''''''_f''''''''''''_Int_data_emitted ;
  logic [4:0] \f''''''''''''_f''''''''''''_Int_data_done ;
  assign \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intgo_11_d  = (\f''''''''''''_f''''''''''''_Int_data_d [0] && (! \f''''''''''''_f''''''''''''_Int_data_emitted [0]));
  assign \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intq4afj_1_d  = {\f''''''''''''_f''''''''''''_Int_data_d [16:1],
                                                                                                                                     (\f''''''''''''_f''''''''''''_Int_data_d [0] && (! \f''''''''''''_f''''''''''''_Int_data_emitted [1]))};
  assign \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intt4afk_1_d  = {\f''''''''''''_f''''''''''''_Int_data_d [32:17],
                                                                                                                                     (\f''''''''''''_f''''''''''''_Int_data_d [0] && (! \f''''''''''''_f''''''''''''_Int_data_emitted [2]))};
  assign \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zafl_1_d  = (\f''''''''''''_f''''''''''''_Int_data_d [0] && (! \f''''''''''''_f''''''''''''_Int_data_emitted [3]));
  assign \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addafm_1_d  = (\f''''''''''''_f''''''''''''_Int_data_d [0] && (! \f''''''''''''_f''''''''''''_Int_data_emitted [4]));
  assign \f''''''''''''_f''''''''''''_Int_data_done  = (\f''''''''''''_f''''''''''''_Int_data_emitted  | ({\f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addafm_1_d [0],
                                                                                                           \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zafl_1_d [0],
                                                                                                           \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intt4afk_1_d [0],
                                                                                                           \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intq4afj_1_d [0],
                                                                                                           \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intgo_11_d [0]} & {\f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addafm_1_r ,
                                                                                                                                                                                                                                         \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zafl_1_r ,
                                                                                                                                                                                                                                         \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intt4afk_1_r ,
                                                                                                                                                                                                                                         \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intq4afj_1_r ,
                                                                                                                                                                                                                                         \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intgo_11_r }));
  assign \f''''''''''''_f''''''''''''_Int_data_r  = (& \f''''''''''''_f''''''''''''_Int_data_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''''''_f''''''''''''_Int_data_emitted  <= 5'd0;
    else
      \f''''''''''''_f''''''''''''_Int_data_emitted  <= (\f''''''''''''_f''''''''''''_Int_data_r  ? 5'd0 :
                                                         \f''''''''''''_f''''''''''''_Int_data_done );
  
  /* destruct (Ty TupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int,
          Dcon TupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int) : (f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1,TupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int) > [(f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intgo_12,Go),
                                                                                                                                                                                                                                                                                                                                         (f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm1aeq_1,Pointer_QTree_Int),
                                                                                                                                                                                                                                                                                                                                         (f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm2aer_1,Pointer_QTree_Int),
                                                                                                                                                                                                                                                                                                                                         (f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm3aes_1,Pointer_QTree_Int),
                                                                                                                                                                                                                                                                                                                                         (f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zaet_1,MyDTInt_Bool),
                                                                                                                                                                                                                                                                                                                                         (f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addaeu_1,MyDTInt_Int_Int)] */
  logic [5:0] f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_emitted;
  logic [5:0] f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_done;
  assign f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intgo_12_d = (f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_d[0] && (! f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_emitted[0]));
  assign f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm1aeq_1_d = {f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_d[16:1],
                                                                                                                               (f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_d[0] && (! f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_emitted[1]))};
  assign f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm2aer_1_d = {f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_d[32:17],
                                                                                                                               (f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_d[0] && (! f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_emitted[2]))};
  assign f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm3aes_1_d = {f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_d[48:33],
                                                                                                                               (f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_d[0] && (! f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_emitted[3]))};
  assign f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zaet_1_d = (f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_d[0] && (! f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_emitted[4]));
  assign f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addaeu_1_d = (f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_d[0] && (! f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_emitted[5]));
  assign f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_done = (f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_emitted | ({f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addaeu_1_d[0],
                                                                                                                                                                                                                                                     f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zaet_1_d[0],
                                                                                                                                                                                                                                                     f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm3aes_1_d[0],
                                                                                                                                                                                                                                                     f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm2aer_1_d[0],
                                                                                                                                                                                                                                                     f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm1aeq_1_d[0],
                                                                                                                                                                                                                                                     f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intgo_12_d[0]} & {f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addaeu_1_r,
                                                                                                                                                                                                                                                                                                                                                                             f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zaet_1_r,
                                                                                                                                                                                                                                                                                                                                                                             f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm3aes_1_r,
                                                                                                                                                                                                                                                                                                                                                                             f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm2aer_1_r,
                                                                                                                                                                                                                                                                                                                                                                             f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm1aeq_1_r,
                                                                                                                                                                                                                                                                                                                                                                             f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intgo_12_r}));
  assign f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_r = (& f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_emitted <= 6'd0;
    else
      f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_emitted <= (f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_r ? 6'd0 :
                                                                                                                              f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_done);
  
  /* fork (Ty Go) : (f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intgo_12,Go) > [(go_12_1,Go),
                                                                                                                                      (go_12_2,Go)] */
  logic [1:0] f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intgo_12_emitted;
  logic [1:0] f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intgo_12_done;
  assign go_12_1_d = (f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intgo_12_d[0] && (! f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intgo_12_emitted[0]));
  assign go_12_2_d = (f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intgo_12_d[0] && (! f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intgo_12_emitted[1]));
  assign f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intgo_12_done = (f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intgo_12_emitted | ({go_12_2_d[0],
                                                                                                                                                                                                                                                           go_12_1_d[0]} & {go_12_2_r,
                                                                                                                                                                                                                                                                            go_12_1_r}));
  assign f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intgo_12_r = (& f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intgo_12_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intgo_12_emitted <= 2'd0;
    else
      f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intgo_12_emitted <= (f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intgo_12_r ? 2'd0 :
                                                                                                                                 f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intgo_12_done);
  
  /* buf (Ty MyDTInt_Bool) : (f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zaet_1,MyDTInt_Bool) > (is_zaet_1_1_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zaet_1_bufchan_d;
  logic f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zaet_1_bufchan_r;
  assign f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zaet_1_r = ((! f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zaet_1_bufchan_d[0]) || f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zaet_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zaet_1_bufchan_d <= 1'd0;
    else
      if (f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zaet_1_r)
        f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zaet_1_bufchan_d <= f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zaet_1_d;
  MyDTInt_Bool_t f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zaet_1_bufchan_buf;
  assign f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zaet_1_bufchan_r = (! f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zaet_1_bufchan_buf[0]);
  assign is_zaet_1_1_argbuf_d = (f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zaet_1_bufchan_buf[0] ? f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zaet_1_bufchan_buf :
                                 f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zaet_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zaet_1_bufchan_buf <= 1'd0;
    else
      if ((is_zaet_1_1_argbuf_r && f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zaet_1_bufchan_buf[0]))
        f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zaet_1_bufchan_buf <= 1'd0;
      else if (((! is_zaet_1_1_argbuf_r) && (! f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zaet_1_bufchan_buf[0])))
        f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zaet_1_bufchan_buf <= f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zaet_1_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm1aeq_1,Pointer_QTree_Int) > (m1aeq_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm1aeq_1_bufchan_d;
  logic f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm1aeq_1_bufchan_r;
  assign f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm1aeq_1_r = ((! f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm1aeq_1_bufchan_d[0]) || f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm1aeq_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm1aeq_1_bufchan_d <= {16'd0,
                                                                                                                                     1'd0};
    else
      if (f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm1aeq_1_r)
        f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm1aeq_1_bufchan_d <= f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm1aeq_1_d;
  Pointer_QTree_Int_t f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm1aeq_1_bufchan_buf;
  assign f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm1aeq_1_bufchan_r = (! f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm1aeq_1_bufchan_buf[0]);
  assign m1aeq_1_1_argbuf_d = (f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm1aeq_1_bufchan_buf[0] ? f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm1aeq_1_bufchan_buf :
                               f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm1aeq_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm1aeq_1_bufchan_buf <= {16'd0,
                                                                                                                                       1'd0};
    else
      if ((m1aeq_1_1_argbuf_r && f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm1aeq_1_bufchan_buf[0]))
        f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm1aeq_1_bufchan_buf <= {16'd0,
                                                                                                                                         1'd0};
      else if (((! m1aeq_1_1_argbuf_r) && (! f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm1aeq_1_bufchan_buf[0])))
        f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm1aeq_1_bufchan_buf <= f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm1aeq_1_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm2aer_1,Pointer_QTree_Int) > (m2aer_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm2aer_1_bufchan_d;
  logic f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm2aer_1_bufchan_r;
  assign f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm2aer_1_r = ((! f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm2aer_1_bufchan_d[0]) || f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm2aer_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm2aer_1_bufchan_d <= {16'd0,
                                                                                                                                     1'd0};
    else
      if (f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm2aer_1_r)
        f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm2aer_1_bufchan_d <= f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm2aer_1_d;
  Pointer_QTree_Int_t f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm2aer_1_bufchan_buf;
  assign f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm2aer_1_bufchan_r = (! f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm2aer_1_bufchan_buf[0]);
  assign m2aer_1_1_argbuf_d = (f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm2aer_1_bufchan_buf[0] ? f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm2aer_1_bufchan_buf :
                               f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm2aer_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm2aer_1_bufchan_buf <= {16'd0,
                                                                                                                                       1'd0};
    else
      if ((m2aer_1_1_argbuf_r && f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm2aer_1_bufchan_buf[0]))
        f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm2aer_1_bufchan_buf <= {16'd0,
                                                                                                                                         1'd0};
      else if (((! m2aer_1_1_argbuf_r) && (! f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm2aer_1_bufchan_buf[0])))
        f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm2aer_1_bufchan_buf <= f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm2aer_1_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm3aes_1,Pointer_QTree_Int) > (m3aes_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm3aes_1_bufchan_d;
  logic f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm3aes_1_bufchan_r;
  assign f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm3aes_1_r = ((! f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm3aes_1_bufchan_d[0]) || f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm3aes_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm3aes_1_bufchan_d <= {16'd0,
                                                                                                                                     1'd0};
    else
      if (f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm3aes_1_r)
        f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm3aes_1_bufchan_d <= f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm3aes_1_d;
  Pointer_QTree_Int_t f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm3aes_1_bufchan_buf;
  assign f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm3aes_1_bufchan_r = (! f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm3aes_1_bufchan_buf[0]);
  assign m3aes_1_1_argbuf_d = (f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm3aes_1_bufchan_buf[0] ? f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm3aes_1_bufchan_buf :
                               f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm3aes_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm3aes_1_bufchan_buf <= {16'd0,
                                                                                                                                       1'd0};
    else
      if ((m3aes_1_1_argbuf_r && f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm3aes_1_bufchan_buf[0]))
        f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm3aes_1_bufchan_buf <= {16'd0,
                                                                                                                                         1'd0};
      else if (((! m3aes_1_1_argbuf_r) && (! f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm3aes_1_bufchan_buf[0])))
        f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm3aes_1_bufchan_buf <= f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm3aes_1_bufchan_d;
  
  /* buf (Ty MyDTInt_Int_Int) : (f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addaeu_1,MyDTInt_Int_Int) > (op_addaeu_1_1_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addaeu_1_bufchan_d;
  logic f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addaeu_1_bufchan_r;
  assign f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addaeu_1_r = ((! f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addaeu_1_bufchan_d[0]) || f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addaeu_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addaeu_1_bufchan_d <= 1'd0;
    else
      if (f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addaeu_1_r)
        f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addaeu_1_bufchan_d <= f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addaeu_1_d;
  MyDTInt_Int_Int_t f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addaeu_1_bufchan_buf;
  assign f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addaeu_1_bufchan_r = (! f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addaeu_1_bufchan_buf[0]);
  assign op_addaeu_1_1_argbuf_d = (f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addaeu_1_bufchan_buf[0] ? f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addaeu_1_bufchan_buf :
                                   f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addaeu_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addaeu_1_bufchan_buf <= 1'd0;
    else
      if ((op_addaeu_1_1_argbuf_r && f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addaeu_1_bufchan_buf[0]))
        f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addaeu_1_bufchan_buf <= 1'd0;
      else if (((! op_addaeu_1_1_argbuf_r) && (! f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addaeu_1_bufchan_buf[0])))
        f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addaeu_1_bufchan_buf <= f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addaeu_1_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (f_f_Int_resbuf,Pointer_QTree_Int) > (es_0_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t f_f_Int_resbuf_bufchan_d;
  logic f_f_Int_resbuf_bufchan_r;
  assign f_f_Int_resbuf_r = ((! f_f_Int_resbuf_bufchan_d[0]) || f_f_Int_resbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) f_f_Int_resbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (f_f_Int_resbuf_r) f_f_Int_resbuf_bufchan_d <= f_f_Int_resbuf_d;
  Pointer_QTree_Int_t f_f_Int_resbuf_bufchan_buf;
  assign f_f_Int_resbuf_bufchan_r = (! f_f_Int_resbuf_bufchan_buf[0]);
  assign es_0_1_argbuf_d = (f_f_Int_resbuf_bufchan_buf[0] ? f_f_Int_resbuf_bufchan_buf :
                            f_f_Int_resbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) f_f_Int_resbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((es_0_1_argbuf_r && f_f_Int_resbuf_bufchan_buf[0]))
        f_f_Int_resbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! es_0_1_argbuf_r) && (! f_f_Int_resbuf_bufchan_buf[0])))
        f_f_Int_resbuf_bufchan_buf <= f_f_Int_resbuf_bufchan_d;
  
  /* dcon (Ty MyDTInt_Int_Int,
      Dcon Dcon_$fNumInt_$c+) : [(go_1,Go)] > (go_1Dcon_$fNumInt_$c+,MyDTInt_Int_Int) */
  assign \go_1Dcon_$fNumInt_$c+_d  = \Dcon_$fNumInt_$c+_dc ((& {go_1_d[0]}), go_1_d);
  assign {go_1_r} = {1 {(\go_1Dcon_$fNumInt_$c+_r  && \go_1Dcon_$fNumInt_$c+_d [0])}};
  
  /* fork (Ty C5) : (go_10_goMux_choice,C5) > [(go_10_goMux_choice_1,C5),
                                          (go_10_goMux_choice_2,C5),
                                          (go_10_goMux_choice_3,C5),
                                          (go_10_goMux_choice_4,C5),
                                          (go_10_goMux_choice_5,C5),
                                          (go_10_goMux_choice_6,C5)] */
  logic [5:0] go_10_goMux_choice_emitted;
  logic [5:0] go_10_goMux_choice_done;
  assign go_10_goMux_choice_1_d = {go_10_goMux_choice_d[3:1],
                                   (go_10_goMux_choice_d[0] && (! go_10_goMux_choice_emitted[0]))};
  assign go_10_goMux_choice_2_d = {go_10_goMux_choice_d[3:1],
                                   (go_10_goMux_choice_d[0] && (! go_10_goMux_choice_emitted[1]))};
  assign go_10_goMux_choice_3_d = {go_10_goMux_choice_d[3:1],
                                   (go_10_goMux_choice_d[0] && (! go_10_goMux_choice_emitted[2]))};
  assign go_10_goMux_choice_4_d = {go_10_goMux_choice_d[3:1],
                                   (go_10_goMux_choice_d[0] && (! go_10_goMux_choice_emitted[3]))};
  assign go_10_goMux_choice_5_d = {go_10_goMux_choice_d[3:1],
                                   (go_10_goMux_choice_d[0] && (! go_10_goMux_choice_emitted[4]))};
  assign go_10_goMux_choice_6_d = {go_10_goMux_choice_d[3:1],
                                   (go_10_goMux_choice_d[0] && (! go_10_goMux_choice_emitted[5]))};
  assign go_10_goMux_choice_done = (go_10_goMux_choice_emitted | ({go_10_goMux_choice_6_d[0],
                                                                   go_10_goMux_choice_5_d[0],
                                                                   go_10_goMux_choice_4_d[0],
                                                                   go_10_goMux_choice_3_d[0],
                                                                   go_10_goMux_choice_2_d[0],
                                                                   go_10_goMux_choice_1_d[0]} & {go_10_goMux_choice_6_r,
                                                                                                 go_10_goMux_choice_5_r,
                                                                                                 go_10_goMux_choice_4_r,
                                                                                                 go_10_goMux_choice_3_r,
                                                                                                 go_10_goMux_choice_2_r,
                                                                                                 go_10_goMux_choice_1_r}));
  assign go_10_goMux_choice_r = (& go_10_goMux_choice_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_10_goMux_choice_emitted <= 6'd0;
    else
      go_10_goMux_choice_emitted <= (go_10_goMux_choice_r ? 6'd0 :
                                     go_10_goMux_choice_done);
  
  /* mux (Ty C5,
     Ty Pointer_QTree_Int) : (go_10_goMux_choice_1,C5) [(call_f_f_Int_goMux2,Pointer_QTree_Int),
                                                        (q3af2_1_1_argbuf,Pointer_QTree_Int),
                                                        (q2af1_2_1_argbuf,Pointer_QTree_Int),
                                                        (q1af0_3_1_argbuf,Pointer_QTree_Int),
                                                        (lizzieLet17_5QNode_Int_7QNode_Int_5QNode_Int_1_argbuf,Pointer_QTree_Int)] > (m1aeq_goMux_mux,Pointer_QTree_Int) */
  logic [16:0] m1aeq_goMux_mux_mux;
  logic [4:0] m1aeq_goMux_mux_onehot;
  always_comb
    unique case (go_10_goMux_choice_1_d[3:1])
      3'd0:
        {m1aeq_goMux_mux_onehot, m1aeq_goMux_mux_mux} = {5'd1,
                                                         call_f_f_Int_goMux2_d};
      3'd1:
        {m1aeq_goMux_mux_onehot, m1aeq_goMux_mux_mux} = {5'd2,
                                                         q3af2_1_1_argbuf_d};
      3'd2:
        {m1aeq_goMux_mux_onehot, m1aeq_goMux_mux_mux} = {5'd4,
                                                         q2af1_2_1_argbuf_d};
      3'd3:
        {m1aeq_goMux_mux_onehot, m1aeq_goMux_mux_mux} = {5'd8,
                                                         q1af0_3_1_argbuf_d};
      3'd4:
        {m1aeq_goMux_mux_onehot, m1aeq_goMux_mux_mux} = {5'd16,
                                                         lizzieLet17_5QNode_Int_7QNode_Int_5QNode_Int_1_argbuf_d};
      default:
        {m1aeq_goMux_mux_onehot, m1aeq_goMux_mux_mux} = {5'd0,
                                                         {16'd0, 1'd0}};
    endcase
  assign m1aeq_goMux_mux_d = {m1aeq_goMux_mux_mux[16:1],
                              (m1aeq_goMux_mux_mux[0] && go_10_goMux_choice_1_d[0])};
  assign go_10_goMux_choice_1_r = (m1aeq_goMux_mux_d[0] && m1aeq_goMux_mux_r);
  assign {lizzieLet17_5QNode_Int_7QNode_Int_5QNode_Int_1_argbuf_r,
          q1af0_3_1_argbuf_r,
          q2af1_2_1_argbuf_r,
          q3af2_1_1_argbuf_r,
          call_f_f_Int_goMux2_r} = (go_10_goMux_choice_1_r ? m1aeq_goMux_mux_onehot :
                                    5'd0);
  
  /* mux (Ty C5,
     Ty Pointer_QTree_Int) : (go_10_goMux_choice_2,C5) [(call_f_f_Int_goMux3,Pointer_QTree_Int),
                                                        (t3afc_1_1_argbuf,Pointer_QTree_Int),
                                                        (t2afb_2_1_argbuf,Pointer_QTree_Int),
                                                        (t1afa_3_1_argbuf,Pointer_QTree_Int),
                                                        (lizzieLet17_5QNode_Int_7QNode_Int_14QNode_Int_1_argbuf,Pointer_QTree_Int)] > (m2aer_goMux_mux,Pointer_QTree_Int) */
  logic [16:0] m2aer_goMux_mux_mux;
  logic [4:0] m2aer_goMux_mux_onehot;
  always_comb
    unique case (go_10_goMux_choice_2_d[3:1])
      3'd0:
        {m2aer_goMux_mux_onehot, m2aer_goMux_mux_mux} = {5'd1,
                                                         call_f_f_Int_goMux3_d};
      3'd1:
        {m2aer_goMux_mux_onehot, m2aer_goMux_mux_mux} = {5'd2,
                                                         t3afc_1_1_argbuf_d};
      3'd2:
        {m2aer_goMux_mux_onehot, m2aer_goMux_mux_mux} = {5'd4,
                                                         t2afb_2_1_argbuf_d};
      3'd3:
        {m2aer_goMux_mux_onehot, m2aer_goMux_mux_mux} = {5'd8,
                                                         t1afa_3_1_argbuf_d};
      3'd4:
        {m2aer_goMux_mux_onehot, m2aer_goMux_mux_mux} = {5'd16,
                                                         lizzieLet17_5QNode_Int_7QNode_Int_14QNode_Int_1_argbuf_d};
      default:
        {m2aer_goMux_mux_onehot, m2aer_goMux_mux_mux} = {5'd0,
                                                         {16'd0, 1'd0}};
    endcase
  assign m2aer_goMux_mux_d = {m2aer_goMux_mux_mux[16:1],
                              (m2aer_goMux_mux_mux[0] && go_10_goMux_choice_2_d[0])};
  assign go_10_goMux_choice_2_r = (m2aer_goMux_mux_d[0] && m2aer_goMux_mux_r);
  assign {lizzieLet17_5QNode_Int_7QNode_Int_14QNode_Int_1_argbuf_r,
          t1afa_3_1_argbuf_r,
          t2afb_2_1_argbuf_r,
          t3afc_1_1_argbuf_r,
          call_f_f_Int_goMux3_r} = (go_10_goMux_choice_2_r ? m2aer_goMux_mux_onehot :
                                    5'd0);
  
  /* mux (Ty C5,
     Ty Pointer_QTree_Int) : (go_10_goMux_choice_3,C5) [(call_f_f_Int_goMux4,Pointer_QTree_Int),
                                                        (t3'afh_1_1_argbuf,Pointer_QTree_Int),
                                                        (t2'afg_2_1_argbuf,Pointer_QTree_Int),
                                                        (t1'aff_3_1_argbuf,Pointer_QTree_Int),
                                                        (t4'afi_1_argbuf,Pointer_QTree_Int)] > (m3aes_goMux_mux,Pointer_QTree_Int) */
  logic [16:0] m3aes_goMux_mux_mux;
  logic [4:0] m3aes_goMux_mux_onehot;
  always_comb
    unique case (go_10_goMux_choice_3_d[3:1])
      3'd0:
        {m3aes_goMux_mux_onehot, m3aes_goMux_mux_mux} = {5'd1,
                                                         call_f_f_Int_goMux4_d};
      3'd1:
        {m3aes_goMux_mux_onehot, m3aes_goMux_mux_mux} = {5'd2,
                                                         \t3'afh_1_1_argbuf_d };
      3'd2:
        {m3aes_goMux_mux_onehot, m3aes_goMux_mux_mux} = {5'd4,
                                                         \t2'afg_2_1_argbuf_d };
      3'd3:
        {m3aes_goMux_mux_onehot, m3aes_goMux_mux_mux} = {5'd8,
                                                         \t1'aff_3_1_argbuf_d };
      3'd4:
        {m3aes_goMux_mux_onehot, m3aes_goMux_mux_mux} = {5'd16,
                                                         \t4'afi_1_argbuf_d };
      default:
        {m3aes_goMux_mux_onehot, m3aes_goMux_mux_mux} = {5'd0,
                                                         {16'd0, 1'd0}};
    endcase
  assign m3aes_goMux_mux_d = {m3aes_goMux_mux_mux[16:1],
                              (m3aes_goMux_mux_mux[0] && go_10_goMux_choice_3_d[0])};
  assign go_10_goMux_choice_3_r = (m3aes_goMux_mux_d[0] && m3aes_goMux_mux_r);
  assign {\t4'afi_1_argbuf_r ,
          \t1'aff_3_1_argbuf_r ,
          \t2'afg_2_1_argbuf_r ,
          \t3'afh_1_1_argbuf_r ,
          call_f_f_Int_goMux4_r} = (go_10_goMux_choice_3_r ? m3aes_goMux_mux_onehot :
                                    5'd0);
  
  /* mux (Ty C5,
     Ty MyDTInt_Bool) : (go_10_goMux_choice_4,C5) [(call_f_f_Int_goMux5,MyDTInt_Bool),
                                                   (is_zaet_2_2_argbuf,MyDTInt_Bool),
                                                   (is_zaet_3_2_argbuf,MyDTInt_Bool),
                                                   (is_zaet_4_1_argbuf,MyDTInt_Bool),
                                                   (lizzieLet17_5QNode_Int_7QNode_Int_9QNode_Int_2_argbuf,MyDTInt_Bool)] > (is_zaet_goMux_mux,MyDTInt_Bool) */
  logic [0:0] is_zaet_goMux_mux_mux;
  logic [4:0] is_zaet_goMux_mux_onehot;
  always_comb
    unique case (go_10_goMux_choice_4_d[3:1])
      3'd0:
        {is_zaet_goMux_mux_onehot, is_zaet_goMux_mux_mux} = {5'd1,
                                                             call_f_f_Int_goMux5_d};
      3'd1:
        {is_zaet_goMux_mux_onehot, is_zaet_goMux_mux_mux} = {5'd2,
                                                             is_zaet_2_2_argbuf_d};
      3'd2:
        {is_zaet_goMux_mux_onehot, is_zaet_goMux_mux_mux} = {5'd4,
                                                             is_zaet_3_2_argbuf_d};
      3'd3:
        {is_zaet_goMux_mux_onehot, is_zaet_goMux_mux_mux} = {5'd8,
                                                             is_zaet_4_1_argbuf_d};
      3'd4:
        {is_zaet_goMux_mux_onehot, is_zaet_goMux_mux_mux} = {5'd16,
                                                             lizzieLet17_5QNode_Int_7QNode_Int_9QNode_Int_2_argbuf_d};
      default:
        {is_zaet_goMux_mux_onehot, is_zaet_goMux_mux_mux} = {5'd0, 1'd0};
    endcase
  assign is_zaet_goMux_mux_d = (is_zaet_goMux_mux_mux[0] && go_10_goMux_choice_4_d[0]);
  assign go_10_goMux_choice_4_r = (is_zaet_goMux_mux_d[0] && is_zaet_goMux_mux_r);
  assign {lizzieLet17_5QNode_Int_7QNode_Int_9QNode_Int_2_argbuf_r,
          is_zaet_4_1_argbuf_r,
          is_zaet_3_2_argbuf_r,
          is_zaet_2_2_argbuf_r,
          call_f_f_Int_goMux5_r} = (go_10_goMux_choice_4_r ? is_zaet_goMux_mux_onehot :
                                    5'd0);
  
  /* mux (Ty C5,
     Ty MyDTInt_Int_Int) : (go_10_goMux_choice_5,C5) [(call_f_f_Int_goMux6,MyDTInt_Int_Int),
                                                      (op_addaeu_2_2_argbuf,MyDTInt_Int_Int),
                                                      (op_addaeu_3_2_argbuf,MyDTInt_Int_Int),
                                                      (op_addaeu_4_1_argbuf,MyDTInt_Int_Int),
                                                      (lizzieLet17_5QNode_Int_7QNode_Int_6QNode_Int_2_argbuf,MyDTInt_Int_Int)] > (op_addaeu_goMux_mux,MyDTInt_Int_Int) */
  logic [0:0] op_addaeu_goMux_mux_mux;
  logic [4:0] op_addaeu_goMux_mux_onehot;
  always_comb
    unique case (go_10_goMux_choice_5_d[3:1])
      3'd0:
        {op_addaeu_goMux_mux_onehot, op_addaeu_goMux_mux_mux} = {5'd1,
                                                                 call_f_f_Int_goMux6_d};
      3'd1:
        {op_addaeu_goMux_mux_onehot, op_addaeu_goMux_mux_mux} = {5'd2,
                                                                 op_addaeu_2_2_argbuf_d};
      3'd2:
        {op_addaeu_goMux_mux_onehot, op_addaeu_goMux_mux_mux} = {5'd4,
                                                                 op_addaeu_3_2_argbuf_d};
      3'd3:
        {op_addaeu_goMux_mux_onehot, op_addaeu_goMux_mux_mux} = {5'd8,
                                                                 op_addaeu_4_1_argbuf_d};
      3'd4:
        {op_addaeu_goMux_mux_onehot, op_addaeu_goMux_mux_mux} = {5'd16,
                                                                 lizzieLet17_5QNode_Int_7QNode_Int_6QNode_Int_2_argbuf_d};
      default:
        {op_addaeu_goMux_mux_onehot, op_addaeu_goMux_mux_mux} = {5'd0,
                                                                 1'd0};
    endcase
  assign op_addaeu_goMux_mux_d = (op_addaeu_goMux_mux_mux[0] && go_10_goMux_choice_5_d[0]);
  assign go_10_goMux_choice_5_r = (op_addaeu_goMux_mux_d[0] && op_addaeu_goMux_mux_r);
  assign {lizzieLet17_5QNode_Int_7QNode_Int_6QNode_Int_2_argbuf_r,
          op_addaeu_4_1_argbuf_r,
          op_addaeu_3_2_argbuf_r,
          op_addaeu_2_2_argbuf_r,
          call_f_f_Int_goMux6_r} = (go_10_goMux_choice_5_r ? op_addaeu_goMux_mux_onehot :
                                    5'd0);
  
  /* mux (Ty C5,
     Ty Pointer_CTf_f_Int) : (go_10_goMux_choice_6,C5) [(call_f_f_Int_goMux7,Pointer_CTf_f_Int),
                                                        (sca2_2_1_argbuf,Pointer_CTf_f_Int),
                                                        (sca1_2_1_argbuf,Pointer_CTf_f_Int),
                                                        (sca0_2_1_argbuf,Pointer_CTf_f_Int),
                                                        (sca3_2_1_argbuf,Pointer_CTf_f_Int)] > (sc_0_2_goMux_mux,Pointer_CTf_f_Int) */
  logic [16:0] sc_0_2_goMux_mux_mux;
  logic [4:0] sc_0_2_goMux_mux_onehot;
  always_comb
    unique case (go_10_goMux_choice_6_d[3:1])
      3'd0:
        {sc_0_2_goMux_mux_onehot, sc_0_2_goMux_mux_mux} = {5'd1,
                                                           call_f_f_Int_goMux7_d};
      3'd1:
        {sc_0_2_goMux_mux_onehot, sc_0_2_goMux_mux_mux} = {5'd2,
                                                           sca2_2_1_argbuf_d};
      3'd2:
        {sc_0_2_goMux_mux_onehot, sc_0_2_goMux_mux_mux} = {5'd4,
                                                           sca1_2_1_argbuf_d};
      3'd3:
        {sc_0_2_goMux_mux_onehot, sc_0_2_goMux_mux_mux} = {5'd8,
                                                           sca0_2_1_argbuf_d};
      3'd4:
        {sc_0_2_goMux_mux_onehot, sc_0_2_goMux_mux_mux} = {5'd16,
                                                           sca3_2_1_argbuf_d};
      default:
        {sc_0_2_goMux_mux_onehot, sc_0_2_goMux_mux_mux} = {5'd0,
                                                           {16'd0, 1'd0}};
    endcase
  assign sc_0_2_goMux_mux_d = {sc_0_2_goMux_mux_mux[16:1],
                               (sc_0_2_goMux_mux_mux[0] && go_10_goMux_choice_6_d[0])};
  assign go_10_goMux_choice_6_r = (sc_0_2_goMux_mux_d[0] && sc_0_2_goMux_mux_r);
  assign {sca3_2_1_argbuf_r,
          sca0_2_1_argbuf_r,
          sca1_2_1_argbuf_r,
          sca2_2_1_argbuf_r,
          call_f_f_Int_goMux7_r} = (go_10_goMux_choice_6_r ? sc_0_2_goMux_mux_onehot :
                                    5'd0);
  
  /* dcon (Ty CTf''''''''''''_f''''''''''''_Int,
      Dcon Lf''''''''''''_f''''''''''''_Intsbos) : [(go_11_1,Go)] > (go_11_1Lf''''''''''''_f''''''''''''_Intsbos,CTf''''''''''''_f''''''''''''_Int) */
  assign \go_11_1Lf''''''''''''_f''''''''''''_Intsbos_d  = \Lf''''''''''''_f''''''''''''_Intsbos_dc ((& {go_11_1_d[0]}), go_11_1_d);
  assign {go_11_1_r} = {1 {(\go_11_1Lf''''''''''''_f''''''''''''_Intsbos_r  && \go_11_1Lf''''''''''''_f''''''''''''_Intsbos_d [0])}};
  
  /* buf (Ty CTf''''''''''''_f''''''''''''_Int) : (go_11_1Lf''''''''''''_f''''''''''''_Intsbos,CTf''''''''''''_f''''''''''''_Int) > (lizzieLet56_1_argbuf,CTf''''''''''''_f''''''''''''_Int) */
  \CTf''''''''''''_f''''''''''''_Int_t  \go_11_1Lf''''''''''''_f''''''''''''_Intsbos_bufchan_d ;
  logic \go_11_1Lf''''''''''''_f''''''''''''_Intsbos_bufchan_r ;
  assign \go_11_1Lf''''''''''''_f''''''''''''_Intsbos_r  = ((! \go_11_1Lf''''''''''''_f''''''''''''_Intsbos_bufchan_d [0]) || \go_11_1Lf''''''''''''_f''''''''''''_Intsbos_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \go_11_1Lf''''''''''''_f''''''''''''_Intsbos_bufchan_d  <= {115'd0,
                                                                  1'd0};
    else
      if (\go_11_1Lf''''''''''''_f''''''''''''_Intsbos_r )
        \go_11_1Lf''''''''''''_f''''''''''''_Intsbos_bufchan_d  <= \go_11_1Lf''''''''''''_f''''''''''''_Intsbos_d ;
  \CTf''''''''''''_f''''''''''''_Int_t  \go_11_1Lf''''''''''''_f''''''''''''_Intsbos_bufchan_buf ;
  assign \go_11_1Lf''''''''''''_f''''''''''''_Intsbos_bufchan_r  = (! \go_11_1Lf''''''''''''_f''''''''''''_Intsbos_bufchan_buf [0]);
  assign lizzieLet56_1_argbuf_d = (\go_11_1Lf''''''''''''_f''''''''''''_Intsbos_bufchan_buf [0] ? \go_11_1Lf''''''''''''_f''''''''''''_Intsbos_bufchan_buf  :
                                   \go_11_1Lf''''''''''''_f''''''''''''_Intsbos_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \go_11_1Lf''''''''''''_f''''''''''''_Intsbos_bufchan_buf  <= {115'd0,
                                                                    1'd0};
    else
      if ((lizzieLet56_1_argbuf_r && \go_11_1Lf''''''''''''_f''''''''''''_Intsbos_bufchan_buf [0]))
        \go_11_1Lf''''''''''''_f''''''''''''_Intsbos_bufchan_buf  <= {115'd0,
                                                                      1'd0};
      else if (((! lizzieLet56_1_argbuf_r) && (! \go_11_1Lf''''''''''''_f''''''''''''_Intsbos_bufchan_buf [0])))
        \go_11_1Lf''''''''''''_f''''''''''''_Intsbos_bufchan_buf  <= \go_11_1Lf''''''''''''_f''''''''''''_Intsbos_bufchan_d ;
  
  /* buf (Ty Go) : (go_11_2,Go) > (go_11_2_argbuf,Go) */
  Go_t go_11_2_bufchan_d;
  logic go_11_2_bufchan_r;
  assign go_11_2_r = ((! go_11_2_bufchan_d[0]) || go_11_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_11_2_bufchan_d <= 1'd0;
    else if (go_11_2_r) go_11_2_bufchan_d <= go_11_2_d;
  Go_t go_11_2_bufchan_buf;
  assign go_11_2_bufchan_r = (! go_11_2_bufchan_buf[0]);
  assign go_11_2_argbuf_d = (go_11_2_bufchan_buf[0] ? go_11_2_bufchan_buf :
                             go_11_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_11_2_bufchan_buf <= 1'd0;
    else
      if ((go_11_2_argbuf_r && go_11_2_bufchan_buf[0]))
        go_11_2_bufchan_buf <= 1'd0;
      else if (((! go_11_2_argbuf_r) && (! go_11_2_bufchan_buf[0])))
        go_11_2_bufchan_buf <= go_11_2_bufchan_d;
  
  /* dcon (Ty TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf''''''''''''_f''''''''''''_Int,
      Dcon TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf''''''''''''_f''''''''''''_Int) : [(go_11_2_argbuf,Go),
                                                                                                                                          (q4afj_1_1_argbuf,Pointer_QTree_Int),
                                                                                                                                          (t4afk_1_1_argbuf,Pointer_QTree_Int),
                                                                                                                                          (is_zafl_1_1_argbuf,MyDTInt_Bool),
                                                                                                                                          (op_addafm_1_1_argbuf,MyDTInt_Int_Int),
                                                                                                                                          (lizzieLet7_1_1_argbuf,Pointer_CTf''''''''''''_f''''''''''''_Int)] > (call_f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf''''''''''''_f''''''''''''_Int_1,TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf''''''''''''_f''''''''''''_Int) */
  assign \call_f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf''''''''''''_f''''''''''''_Int_1_d  = \TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf''''''''''''_f''''''''''''_Int_dc ((& {go_11_2_argbuf_d[0],
                                                                                                                                                                                                                                                                                                                    q4afj_1_1_argbuf_d[0],
                                                                                                                                                                                                                                                                                                                    t4afk_1_1_argbuf_d[0],
                                                                                                                                                                                                                                                                                                                    is_zafl_1_1_argbuf_d[0],
                                                                                                                                                                                                                                                                                                                    op_addafm_1_1_argbuf_d[0],
                                                                                                                                                                                                                                                                                                                    lizzieLet7_1_1_argbuf_d[0]}), go_11_2_argbuf_d, q4afj_1_1_argbuf_d, t4afk_1_1_argbuf_d, is_zafl_1_1_argbuf_d, op_addafm_1_1_argbuf_d, lizzieLet7_1_1_argbuf_d);
  assign {go_11_2_argbuf_r,
          q4afj_1_1_argbuf_r,
          t4afk_1_1_argbuf_r,
          is_zafl_1_1_argbuf_r,
          op_addafm_1_1_argbuf_r,
          lizzieLet7_1_1_argbuf_r} = {6 {(\call_f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf''''''''''''_f''''''''''''_Int_1_r  && \call_f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf''''''''''''_f''''''''''''_Int_1_d [0])}};
  
  /* dcon (Ty CTf_f_Int,
      Dcon Lf_f_Intsbos) : [(go_12_1,Go)] > (go_12_1Lf_f_Intsbos,CTf_f_Int) */
  assign go_12_1Lf_f_Intsbos_d = Lf_f_Intsbos_dc((& {go_12_1_d[0]}), go_12_1_d);
  assign {go_12_1_r} = {1 {(go_12_1Lf_f_Intsbos_r && go_12_1Lf_f_Intsbos_d[0])}};
  
  /* buf (Ty CTf_f_Int) : (go_12_1Lf_f_Intsbos,CTf_f_Int) > (lizzieLet57_1_argbuf,CTf_f_Int) */
  CTf_f_Int_t go_12_1Lf_f_Intsbos_bufchan_d;
  logic go_12_1Lf_f_Intsbos_bufchan_r;
  assign go_12_1Lf_f_Intsbos_r = ((! go_12_1Lf_f_Intsbos_bufchan_d[0]) || go_12_1Lf_f_Intsbos_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      go_12_1Lf_f_Intsbos_bufchan_d <= {163'd0, 1'd0};
    else
      if (go_12_1Lf_f_Intsbos_r)
        go_12_1Lf_f_Intsbos_bufchan_d <= go_12_1Lf_f_Intsbos_d;
  CTf_f_Int_t go_12_1Lf_f_Intsbos_bufchan_buf;
  assign go_12_1Lf_f_Intsbos_bufchan_r = (! go_12_1Lf_f_Intsbos_bufchan_buf[0]);
  assign lizzieLet57_1_argbuf_d = (go_12_1Lf_f_Intsbos_bufchan_buf[0] ? go_12_1Lf_f_Intsbos_bufchan_buf :
                                   go_12_1Lf_f_Intsbos_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      go_12_1Lf_f_Intsbos_bufchan_buf <= {163'd0, 1'd0};
    else
      if ((lizzieLet57_1_argbuf_r && go_12_1Lf_f_Intsbos_bufchan_buf[0]))
        go_12_1Lf_f_Intsbos_bufchan_buf <= {163'd0, 1'd0};
      else if (((! lizzieLet57_1_argbuf_r) && (! go_12_1Lf_f_Intsbos_bufchan_buf[0])))
        go_12_1Lf_f_Intsbos_bufchan_buf <= go_12_1Lf_f_Intsbos_bufchan_d;
  
  /* buf (Ty Go) : (go_12_2,Go) > (go_12_2_argbuf,Go) */
  Go_t go_12_2_bufchan_d;
  logic go_12_2_bufchan_r;
  assign go_12_2_r = ((! go_12_2_bufchan_d[0]) || go_12_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_12_2_bufchan_d <= 1'd0;
    else if (go_12_2_r) go_12_2_bufchan_d <= go_12_2_d;
  Go_t go_12_2_bufchan_buf;
  assign go_12_2_bufchan_r = (! go_12_2_bufchan_buf[0]);
  assign go_12_2_argbuf_d = (go_12_2_bufchan_buf[0] ? go_12_2_bufchan_buf :
                             go_12_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_12_2_bufchan_buf <= 1'd0;
    else
      if ((go_12_2_argbuf_r && go_12_2_bufchan_buf[0]))
        go_12_2_bufchan_buf <= 1'd0;
      else if (((! go_12_2_argbuf_r) && (! go_12_2_bufchan_buf[0])))
        go_12_2_bufchan_buf <= go_12_2_bufchan_d;
  
  /* dcon (Ty TupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int,
      Dcon TupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int) : [(go_12_2_argbuf,Go),
                                                                                                                                      (m1aeq_1_1_argbuf,Pointer_QTree_Int),
                                                                                                                                      (m2aer_1_1_argbuf,Pointer_QTree_Int),
                                                                                                                                      (m3aes_1_1_argbuf,Pointer_QTree_Int),
                                                                                                                                      (is_zaet_1_1_argbuf,MyDTInt_Bool),
                                                                                                                                      (op_addaeu_1_1_argbuf,MyDTInt_Int_Int),
                                                                                                                                      (lizzieLet36_1_1_argbuf,Pointer_CTf_f_Int)] > (call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_1,TupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int) */
  assign call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_1_d = TupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_dc((& {go_12_2_argbuf_d[0],
                                                                                                                                                                                                                                                                                m1aeq_1_1_argbuf_d[0],
                                                                                                                                                                                                                                                                                m2aer_1_1_argbuf_d[0],
                                                                                                                                                                                                                                                                                m3aes_1_1_argbuf_d[0],
                                                                                                                                                                                                                                                                                is_zaet_1_1_argbuf_d[0],
                                                                                                                                                                                                                                                                                op_addaeu_1_1_argbuf_d[0],
                                                                                                                                                                                                                                                                                lizzieLet36_1_1_argbuf_d[0]}), go_12_2_argbuf_d, m1aeq_1_1_argbuf_d, m2aer_1_1_argbuf_d, m3aes_1_1_argbuf_d, is_zaet_1_1_argbuf_d, op_addaeu_1_1_argbuf_d, lizzieLet36_1_1_argbuf_d);
  assign {go_12_2_argbuf_r,
          m1aeq_1_1_argbuf_r,
          m2aer_1_1_argbuf_r,
          m3aes_1_1_argbuf_r,
          is_zaet_1_1_argbuf_r,
          op_addaeu_1_1_argbuf_r,
          lizzieLet36_1_1_argbuf_r} = {7 {(call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_1_r && call_f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_1_d[0])}};
  
  /* fork (Ty C4) : (go_13_goMux_choice,C4) > [(go_13_goMux_choice_1,C4),
                                          (go_13_goMux_choice_2,C4)] */
  logic [1:0] go_13_goMux_choice_emitted;
  logic [1:0] go_13_goMux_choice_done;
  assign go_13_goMux_choice_1_d = {go_13_goMux_choice_d[2:1],
                                   (go_13_goMux_choice_d[0] && (! go_13_goMux_choice_emitted[0]))};
  assign go_13_goMux_choice_2_d = {go_13_goMux_choice_d[2:1],
                                   (go_13_goMux_choice_d[0] && (! go_13_goMux_choice_emitted[1]))};
  assign go_13_goMux_choice_done = (go_13_goMux_choice_emitted | ({go_13_goMux_choice_2_d[0],
                                                                   go_13_goMux_choice_1_d[0]} & {go_13_goMux_choice_2_r,
                                                                                                 go_13_goMux_choice_1_r}));
  assign go_13_goMux_choice_r = (& go_13_goMux_choice_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_13_goMux_choice_emitted <= 2'd0;
    else
      go_13_goMux_choice_emitted <= (go_13_goMux_choice_r ? 2'd0 :
                                     go_13_goMux_choice_done);
  
  /* mux (Ty C4,
     Ty Int#) : (go_13_goMux_choice_1,C4) [(lizzieLet37_1_argbuf,Int#),
                                           (contRet_0_1_argbuf,Int#),
                                           (lizzieLet38_1_argbuf,Int#),
                                           (lizzieLet37_1_1_argbuf,Int#)] > (srtarg_0_goMux_mux,Int#) */
  logic [32:0] srtarg_0_goMux_mux_mux;
  logic [3:0] srtarg_0_goMux_mux_onehot;
  always_comb
    unique case (go_13_goMux_choice_1_d[2:1])
      2'd0:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {4'd1,
                                                               lizzieLet37_1_argbuf_d};
      2'd1:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {4'd2,
                                                               contRet_0_1_argbuf_d};
      2'd2:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {4'd4,
                                                               lizzieLet38_1_argbuf_d};
      2'd3:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {4'd8,
                                                               lizzieLet37_1_1_argbuf_d};
      default:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {4'd0,
                                                               {32'd0, 1'd0}};
    endcase
  assign srtarg_0_goMux_mux_d = {srtarg_0_goMux_mux_mux[32:1],
                                 (srtarg_0_goMux_mux_mux[0] && go_13_goMux_choice_1_d[0])};
  assign go_13_goMux_choice_1_r = (srtarg_0_goMux_mux_d[0] && srtarg_0_goMux_mux_r);
  assign {lizzieLet37_1_1_argbuf_r,
          lizzieLet38_1_argbuf_r,
          contRet_0_1_argbuf_r,
          lizzieLet37_1_argbuf_r} = (go_13_goMux_choice_1_r ? srtarg_0_goMux_mux_onehot :
                                     4'd0);
  
  /* mux (Ty C4,
     Ty Pointer_CT$wnnz) : (go_13_goMux_choice_2,C4) [(lizzieLet4_4QNone_Int_1_argbuf,Pointer_CT$wnnz),
                                                      (sc_0_6_1_argbuf,Pointer_CT$wnnz),
                                                      (lizzieLet4_4QVal_Int_1_argbuf,Pointer_CT$wnnz),
                                                      (lizzieLet4_4QError_Int_1_argbuf,Pointer_CT$wnnz)] > (scfarg_0_goMux_mux,Pointer_CT$wnnz) */
  logic [16:0] scfarg_0_goMux_mux_mux;
  logic [3:0] scfarg_0_goMux_mux_onehot;
  always_comb
    unique case (go_13_goMux_choice_2_d[2:1])
      2'd0:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {4'd1,
                                                               lizzieLet4_4QNone_Int_1_argbuf_d};
      2'd1:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {4'd2,
                                                               sc_0_6_1_argbuf_d};
      2'd2:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {4'd4,
                                                               lizzieLet4_4QVal_Int_1_argbuf_d};
      2'd3:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {4'd8,
                                                               lizzieLet4_4QError_Int_1_argbuf_d};
      default:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {4'd0,
                                                               {16'd0, 1'd0}};
    endcase
  assign scfarg_0_goMux_mux_d = {scfarg_0_goMux_mux_mux[16:1],
                                 (scfarg_0_goMux_mux_mux[0] && go_13_goMux_choice_2_d[0])};
  assign go_13_goMux_choice_2_r = (scfarg_0_goMux_mux_d[0] && scfarg_0_goMux_mux_r);
  assign {lizzieLet4_4QError_Int_1_argbuf_r,
          lizzieLet4_4QVal_Int_1_argbuf_r,
          sc_0_6_1_argbuf_r,
          lizzieLet4_4QNone_Int_1_argbuf_r} = (go_13_goMux_choice_2_r ? scfarg_0_goMux_mux_onehot :
                                               4'd0);
  
  /* fork (Ty C11) : (go_14_goMux_choice,C11) > [(go_14_goMux_choice_1,C11),
                                            (go_14_goMux_choice_2,C11)] */
  logic [1:0] go_14_goMux_choice_emitted;
  logic [1:0] go_14_goMux_choice_done;
  assign go_14_goMux_choice_1_d = {go_14_goMux_choice_d[4:1],
                                   (go_14_goMux_choice_d[0] && (! go_14_goMux_choice_emitted[0]))};
  assign go_14_goMux_choice_2_d = {go_14_goMux_choice_d[4:1],
                                   (go_14_goMux_choice_d[0] && (! go_14_goMux_choice_emitted[1]))};
  assign go_14_goMux_choice_done = (go_14_goMux_choice_emitted | ({go_14_goMux_choice_2_d[0],
                                                                   go_14_goMux_choice_1_d[0]} & {go_14_goMux_choice_2_r,
                                                                                                 go_14_goMux_choice_1_r}));
  assign go_14_goMux_choice_r = (& go_14_goMux_choice_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_14_goMux_choice_emitted <= 2'd0;
    else
      go_14_goMux_choice_emitted <= (go_14_goMux_choice_r ? 2'd0 :
                                     go_14_goMux_choice_done);
  
  /* mux (Ty C11,
     Ty Pointer_QTree_Int) : (go_14_goMux_choice_1,C11) [(lizzieLet6_9QNone_Int_1_argbuf,Pointer_QTree_Int),
                                                         (contRet_0_1_1_argbuf,Pointer_QTree_Int),
                                                         (lizzieLet6_5QVal_Int_6QNone_Int_1_argbuf,Pointer_QTree_Int),
                                                         (lizzieLet0_1_1_argbuf,Pointer_QTree_Int),
                                                         (lizzieLet1_1_1_argbuf,Pointer_QTree_Int),
                                                         (lizzieLet2_1_1_argbuf,Pointer_QTree_Int),
                                                         (lizzieLet3_1_1_argbuf,Pointer_QTree_Int),
                                                         (lizzieLet6_5QNode_Int_6QNone_Int_1_argbuf,Pointer_QTree_Int),
                                                         (lizzieLet4_1_1_argbuf,Pointer_QTree_Int),
                                                         (lizzieLet5_1_1_argbuf,Pointer_QTree_Int),
                                                         (lizzieLet6_1_1_argbuf,Pointer_QTree_Int)] > (srtarg_0_1_goMux_mux,Pointer_QTree_Int) */
  logic [16:0] srtarg_0_1_goMux_mux_mux;
  logic [10:0] srtarg_0_1_goMux_mux_onehot;
  always_comb
    unique case (go_14_goMux_choice_1_d[4:1])
      4'd0:
        {srtarg_0_1_goMux_mux_onehot, srtarg_0_1_goMux_mux_mux} = {11'd1,
                                                                   lizzieLet6_9QNone_Int_1_argbuf_d};
      4'd1:
        {srtarg_0_1_goMux_mux_onehot, srtarg_0_1_goMux_mux_mux} = {11'd2,
                                                                   contRet_0_1_1_argbuf_d};
      4'd2:
        {srtarg_0_1_goMux_mux_onehot, srtarg_0_1_goMux_mux_mux} = {11'd4,
                                                                   lizzieLet6_5QVal_Int_6QNone_Int_1_argbuf_d};
      4'd3:
        {srtarg_0_1_goMux_mux_onehot, srtarg_0_1_goMux_mux_mux} = {11'd8,
                                                                   lizzieLet0_1_1_argbuf_d};
      4'd4:
        {srtarg_0_1_goMux_mux_onehot, srtarg_0_1_goMux_mux_mux} = {11'd16,
                                                                   lizzieLet1_1_1_argbuf_d};
      4'd5:
        {srtarg_0_1_goMux_mux_onehot, srtarg_0_1_goMux_mux_mux} = {11'd32,
                                                                   lizzieLet2_1_1_argbuf_d};
      4'd6:
        {srtarg_0_1_goMux_mux_onehot, srtarg_0_1_goMux_mux_mux} = {11'd64,
                                                                   lizzieLet3_1_1_argbuf_d};
      4'd7:
        {srtarg_0_1_goMux_mux_onehot, srtarg_0_1_goMux_mux_mux} = {11'd128,
                                                                   lizzieLet6_5QNode_Int_6QNone_Int_1_argbuf_d};
      4'd8:
        {srtarg_0_1_goMux_mux_onehot, srtarg_0_1_goMux_mux_mux} = {11'd256,
                                                                   lizzieLet4_1_1_argbuf_d};
      4'd9:
        {srtarg_0_1_goMux_mux_onehot, srtarg_0_1_goMux_mux_mux} = {11'd512,
                                                                   lizzieLet5_1_1_argbuf_d};
      4'd10:
        {srtarg_0_1_goMux_mux_onehot,
         srtarg_0_1_goMux_mux_mux} = {11'd1024, lizzieLet6_1_1_argbuf_d};
      default:
        {srtarg_0_1_goMux_mux_onehot, srtarg_0_1_goMux_mux_mux} = {11'd0,
                                                                   {16'd0, 1'd0}};
    endcase
  assign srtarg_0_1_goMux_mux_d = {srtarg_0_1_goMux_mux_mux[16:1],
                                   (srtarg_0_1_goMux_mux_mux[0] && go_14_goMux_choice_1_d[0])};
  assign go_14_goMux_choice_1_r = (srtarg_0_1_goMux_mux_d[0] && srtarg_0_1_goMux_mux_r);
  assign {lizzieLet6_1_1_argbuf_r,
          lizzieLet5_1_1_argbuf_r,
          lizzieLet4_1_1_argbuf_r,
          lizzieLet6_5QNode_Int_6QNone_Int_1_argbuf_r,
          lizzieLet3_1_1_argbuf_r,
          lizzieLet2_1_1_argbuf_r,
          lizzieLet1_1_1_argbuf_r,
          lizzieLet0_1_1_argbuf_r,
          lizzieLet6_5QVal_Int_6QNone_Int_1_argbuf_r,
          contRet_0_1_1_argbuf_r,
          lizzieLet6_9QNone_Int_1_argbuf_r} = (go_14_goMux_choice_1_r ? srtarg_0_1_goMux_mux_onehot :
                                               11'd0);
  
  /* mux (Ty C11,
     Ty Pointer_CTf''''''''''''_f''''''''''''_Int) : (go_14_goMux_choice_2,C11) [(lizzieLet6_8QNone_Int_1_argbuf,Pointer_CTf''''''''''''_f''''''''''''_Int),
                                                                                 (sc_0_10_1_argbuf,Pointer_CTf''''''''''''_f''''''''''''_Int),
                                                                                 (lizzieLet6_5QVal_Int_7QNone_Int_1_argbuf,Pointer_CTf''''''''''''_f''''''''''''_Int),
                                                                                 (es_2_3MyFalse_1_argbuf,Pointer_CTf''''''''''''_f''''''''''''_Int),
                                                                                 (es_2_3MyTrue_1_argbuf,Pointer_CTf''''''''''''_f''''''''''''_Int),
                                                                                 (lizzieLet6_5QVal_Int_7QNode_Int_1_argbuf,Pointer_CTf''''''''''''_f''''''''''''_Int),
                                                                                 (lizzieLet6_5QVal_Int_7QError_Int_1_argbuf,Pointer_CTf''''''''''''_f''''''''''''_Int),
                                                                                 (lizzieLet6_5QNode_Int_7QNone_Int_1_argbuf,Pointer_CTf''''''''''''_f''''''''''''_Int),
                                                                                 (lizzieLet6_5QNode_Int_7QVal_Int_1_argbuf,Pointer_CTf''''''''''''_f''''''''''''_Int),
                                                                                 (lizzieLet6_5QNode_Int_7QError_Int_1_argbuf,Pointer_CTf''''''''''''_f''''''''''''_Int),
                                                                                 (lizzieLet6_8QError_Int_1_argbuf,Pointer_CTf''''''''''''_f''''''''''''_Int)] > (scfarg_0_1_goMux_mux,Pointer_CTf''''''''''''_f''''''''''''_Int) */
  logic [16:0] scfarg_0_1_goMux_mux_mux;
  logic [10:0] scfarg_0_1_goMux_mux_onehot;
  always_comb
    unique case (go_14_goMux_choice_2_d[4:1])
      4'd0:
        {scfarg_0_1_goMux_mux_onehot, scfarg_0_1_goMux_mux_mux} = {11'd1,
                                                                   lizzieLet6_8QNone_Int_1_argbuf_d};
      4'd1:
        {scfarg_0_1_goMux_mux_onehot, scfarg_0_1_goMux_mux_mux} = {11'd2,
                                                                   sc_0_10_1_argbuf_d};
      4'd2:
        {scfarg_0_1_goMux_mux_onehot, scfarg_0_1_goMux_mux_mux} = {11'd4,
                                                                   lizzieLet6_5QVal_Int_7QNone_Int_1_argbuf_d};
      4'd3:
        {scfarg_0_1_goMux_mux_onehot, scfarg_0_1_goMux_mux_mux} = {11'd8,
                                                                   es_2_3MyFalse_1_argbuf_d};
      4'd4:
        {scfarg_0_1_goMux_mux_onehot, scfarg_0_1_goMux_mux_mux} = {11'd16,
                                                                   es_2_3MyTrue_1_argbuf_d};
      4'd5:
        {scfarg_0_1_goMux_mux_onehot, scfarg_0_1_goMux_mux_mux} = {11'd32,
                                                                   lizzieLet6_5QVal_Int_7QNode_Int_1_argbuf_d};
      4'd6:
        {scfarg_0_1_goMux_mux_onehot, scfarg_0_1_goMux_mux_mux} = {11'd64,
                                                                   lizzieLet6_5QVal_Int_7QError_Int_1_argbuf_d};
      4'd7:
        {scfarg_0_1_goMux_mux_onehot, scfarg_0_1_goMux_mux_mux} = {11'd128,
                                                                   lizzieLet6_5QNode_Int_7QNone_Int_1_argbuf_d};
      4'd8:
        {scfarg_0_1_goMux_mux_onehot, scfarg_0_1_goMux_mux_mux} = {11'd256,
                                                                   lizzieLet6_5QNode_Int_7QVal_Int_1_argbuf_d};
      4'd9:
        {scfarg_0_1_goMux_mux_onehot, scfarg_0_1_goMux_mux_mux} = {11'd512,
                                                                   lizzieLet6_5QNode_Int_7QError_Int_1_argbuf_d};
      4'd10:
        {scfarg_0_1_goMux_mux_onehot,
         scfarg_0_1_goMux_mux_mux} = {11'd1024,
                                      lizzieLet6_8QError_Int_1_argbuf_d};
      default:
        {scfarg_0_1_goMux_mux_onehot, scfarg_0_1_goMux_mux_mux} = {11'd0,
                                                                   {16'd0, 1'd0}};
    endcase
  assign scfarg_0_1_goMux_mux_d = {scfarg_0_1_goMux_mux_mux[16:1],
                                   (scfarg_0_1_goMux_mux_mux[0] && go_14_goMux_choice_2_d[0])};
  assign go_14_goMux_choice_2_r = (scfarg_0_1_goMux_mux_d[0] && scfarg_0_1_goMux_mux_r);
  assign {lizzieLet6_8QError_Int_1_argbuf_r,
          lizzieLet6_5QNode_Int_7QError_Int_1_argbuf_r,
          lizzieLet6_5QNode_Int_7QVal_Int_1_argbuf_r,
          lizzieLet6_5QNode_Int_7QNone_Int_1_argbuf_r,
          lizzieLet6_5QVal_Int_7QError_Int_1_argbuf_r,
          lizzieLet6_5QVal_Int_7QNode_Int_1_argbuf_r,
          es_2_3MyTrue_1_argbuf_r,
          es_2_3MyFalse_1_argbuf_r,
          lizzieLet6_5QVal_Int_7QNone_Int_1_argbuf_r,
          sc_0_10_1_argbuf_r,
          lizzieLet6_8QNone_Int_1_argbuf_r} = (go_14_goMux_choice_2_r ? scfarg_0_1_goMux_mux_onehot :
                                               11'd0);
  
  /* fork (Ty C35) : (go_15_goMux_choice,C35) > [(go_15_goMux_choice_1,C35),
                                            (go_15_goMux_choice_2,C35)] */
  logic [1:0] go_15_goMux_choice_emitted;
  logic [1:0] go_15_goMux_choice_done;
  assign go_15_goMux_choice_1_d = {go_15_goMux_choice_d[6:1],
                                   (go_15_goMux_choice_d[0] && (! go_15_goMux_choice_emitted[0]))};
  assign go_15_goMux_choice_2_d = {go_15_goMux_choice_d[6:1],
                                   (go_15_goMux_choice_d[0] && (! go_15_goMux_choice_emitted[1]))};
  assign go_15_goMux_choice_done = (go_15_goMux_choice_emitted | ({go_15_goMux_choice_2_d[0],
                                                                   go_15_goMux_choice_1_d[0]} & {go_15_goMux_choice_2_r,
                                                                                                 go_15_goMux_choice_1_r}));
  assign go_15_goMux_choice_r = (& go_15_goMux_choice_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_15_goMux_choice_emitted <= 2'd0;
    else
      go_15_goMux_choice_emitted <= (go_15_goMux_choice_r ? 2'd0 :
                                     go_15_goMux_choice_done);
  
  /* mux (Ty C35,
     Ty Pointer_QTree_Int) : (go_15_goMux_choice_1,C35) [(lizzieLet17_5QNone_Int_9QNone_Int_1_argbuf,Pointer_QTree_Int),
                                                         (contRet_0_2_1_argbuf,Pointer_QTree_Int),
                                                         (lizzieLet17_5QNone_Int_7QVal_Int_7QNone_Int_1_argbuf,Pointer_QTree_Int),
                                                         (lizzieLet8_1_1_argbuf,Pointer_QTree_Int),
                                                         (lizzieLet9_1_1_argbuf,Pointer_QTree_Int),
                                                         (lizzieLet10_1_1_argbuf,Pointer_QTree_Int),
                                                         (lizzieLet11_1_1_argbuf,Pointer_QTree_Int),
                                                         (lizzieLet17_5QNone_Int_7QNode_Int_7QNone_Int_1_argbuf,Pointer_QTree_Int),
                                                         (lizzieLet12_1_argbuf,Pointer_QTree_Int),
                                                         (lizzieLet13_1_1_argbuf,Pointer_QTree_Int),
                                                         (lizzieLet14_1_1_argbuf,Pointer_QTree_Int),
                                                         (lizzieLet15_1_1_argbuf,Pointer_QTree_Int),
                                                         (lizzieLet17_5QVal_Int_7QNone_Int_8QNone_Int_1_argbuf,Pointer_QTree_Int),
                                                         (lizzieLet16_1_1_argbuf,Pointer_QTree_Int),
                                                         (lizzieLet17_1_1_argbuf,Pointer_QTree_Int),
                                                         (lizzieLet18_1_1_argbuf,Pointer_QTree_Int),
                                                         (lizzieLet19_1_1_argbuf,Pointer_QTree_Int),
                                                         (lizzieLet20_1_1_argbuf,Pointer_QTree_Int),
                                                         (lizzieLet21_1_1_argbuf,Pointer_QTree_Int),
                                                         (lizzieLet22_1_1_argbuf,Pointer_QTree_Int),
                                                         (lizzieLet23_1_1_argbuf,Pointer_QTree_Int),
                                                         (lizzieLet24_1_argbuf,Pointer_QTree_Int),
                                                         (es_14_7MyTrue_1_argbuf,Pointer_QTree_Int),
                                                         (lizzieLet25_1_1_argbuf,Pointer_QTree_Int),
                                                         (lizzieLet26_1_1_argbuf,Pointer_QTree_Int),
                                                         (lizzieLet17_5QNode_Int_7QNone_Int_10QNone_Int_1_argbuf,Pointer_QTree_Int),
                                                         (lizzieLet27_1_1_argbuf,Pointer_QTree_Int),
                                                         (lizzieLet28_1_1_argbuf,Pointer_QTree_Int),
                                                         (lizzieLet29_1_argbuf,Pointer_QTree_Int),
                                                         (lizzieLet30_1_argbuf,Pointer_QTree_Int),
                                                         (lizzieLet31_1_1_argbuf,Pointer_QTree_Int),
                                                         (lizzieLet32_1_1_argbuf,Pointer_QTree_Int),
                                                         (lizzieLet33_1_1_argbuf,Pointer_QTree_Int),
                                                         (lizzieLet34_1_1_argbuf,Pointer_QTree_Int),
                                                         (lizzieLet35_1_argbuf,Pointer_QTree_Int)] > (srtarg_0_2_goMux_mux,Pointer_QTree_Int) */
  logic [16:0] srtarg_0_2_goMux_mux_mux;
  logic [34:0] srtarg_0_2_goMux_mux_onehot;
  always_comb
    unique case (go_15_goMux_choice_1_d[6:1])
      6'd0:
        {srtarg_0_2_goMux_mux_onehot, srtarg_0_2_goMux_mux_mux} = {35'd1,
                                                                   lizzieLet17_5QNone_Int_9QNone_Int_1_argbuf_d};
      6'd1:
        {srtarg_0_2_goMux_mux_onehot, srtarg_0_2_goMux_mux_mux} = {35'd2,
                                                                   contRet_0_2_1_argbuf_d};
      6'd2:
        {srtarg_0_2_goMux_mux_onehot, srtarg_0_2_goMux_mux_mux} = {35'd4,
                                                                   lizzieLet17_5QNone_Int_7QVal_Int_7QNone_Int_1_argbuf_d};
      6'd3:
        {srtarg_0_2_goMux_mux_onehot, srtarg_0_2_goMux_mux_mux} = {35'd8,
                                                                   lizzieLet8_1_1_argbuf_d};
      6'd4:
        {srtarg_0_2_goMux_mux_onehot, srtarg_0_2_goMux_mux_mux} = {35'd16,
                                                                   lizzieLet9_1_1_argbuf_d};
      6'd5:
        {srtarg_0_2_goMux_mux_onehot, srtarg_0_2_goMux_mux_mux} = {35'd32,
                                                                   lizzieLet10_1_1_argbuf_d};
      6'd6:
        {srtarg_0_2_goMux_mux_onehot, srtarg_0_2_goMux_mux_mux} = {35'd64,
                                                                   lizzieLet11_1_1_argbuf_d};
      6'd7:
        {srtarg_0_2_goMux_mux_onehot, srtarg_0_2_goMux_mux_mux} = {35'd128,
                                                                   lizzieLet17_5QNone_Int_7QNode_Int_7QNone_Int_1_argbuf_d};
      6'd8:
        {srtarg_0_2_goMux_mux_onehot, srtarg_0_2_goMux_mux_mux} = {35'd256,
                                                                   lizzieLet12_1_argbuf_d};
      6'd9:
        {srtarg_0_2_goMux_mux_onehot, srtarg_0_2_goMux_mux_mux} = {35'd512,
                                                                   lizzieLet13_1_1_argbuf_d};
      6'd10:
        {srtarg_0_2_goMux_mux_onehot,
         srtarg_0_2_goMux_mux_mux} = {35'd1024, lizzieLet14_1_1_argbuf_d};
      6'd11:
        {srtarg_0_2_goMux_mux_onehot,
         srtarg_0_2_goMux_mux_mux} = {35'd2048, lizzieLet15_1_1_argbuf_d};
      6'd12:
        {srtarg_0_2_goMux_mux_onehot,
         srtarg_0_2_goMux_mux_mux} = {35'd4096,
                                      lizzieLet17_5QVal_Int_7QNone_Int_8QNone_Int_1_argbuf_d};
      6'd13:
        {srtarg_0_2_goMux_mux_onehot,
         srtarg_0_2_goMux_mux_mux} = {35'd8192, lizzieLet16_1_1_argbuf_d};
      6'd14:
        {srtarg_0_2_goMux_mux_onehot,
         srtarg_0_2_goMux_mux_mux} = {35'd16384, lizzieLet17_1_1_argbuf_d};
      6'd15:
        {srtarg_0_2_goMux_mux_onehot,
         srtarg_0_2_goMux_mux_mux} = {35'd32768, lizzieLet18_1_1_argbuf_d};
      6'd16:
        {srtarg_0_2_goMux_mux_onehot,
         srtarg_0_2_goMux_mux_mux} = {35'd65536, lizzieLet19_1_1_argbuf_d};
      6'd17:
        {srtarg_0_2_goMux_mux_onehot,
         srtarg_0_2_goMux_mux_mux} = {35'd131072, lizzieLet20_1_1_argbuf_d};
      6'd18:
        {srtarg_0_2_goMux_mux_onehot,
         srtarg_0_2_goMux_mux_mux} = {35'd262144, lizzieLet21_1_1_argbuf_d};
      6'd19:
        {srtarg_0_2_goMux_mux_onehot,
         srtarg_0_2_goMux_mux_mux} = {35'd524288, lizzieLet22_1_1_argbuf_d};
      6'd20:
        {srtarg_0_2_goMux_mux_onehot,
         srtarg_0_2_goMux_mux_mux} = {35'd1048576,
                                      lizzieLet23_1_1_argbuf_d};
      6'd21:
        {srtarg_0_2_goMux_mux_onehot,
         srtarg_0_2_goMux_mux_mux} = {35'd2097152, lizzieLet24_1_argbuf_d};
      6'd22:
        {srtarg_0_2_goMux_mux_onehot,
         srtarg_0_2_goMux_mux_mux} = {35'd4194304,
                                      es_14_7MyTrue_1_argbuf_d};
      6'd23:
        {srtarg_0_2_goMux_mux_onehot,
         srtarg_0_2_goMux_mux_mux} = {35'd8388608,
                                      lizzieLet25_1_1_argbuf_d};
      6'd24:
        {srtarg_0_2_goMux_mux_onehot,
         srtarg_0_2_goMux_mux_mux} = {35'd16777216,
                                      lizzieLet26_1_1_argbuf_d};
      6'd25:
        {srtarg_0_2_goMux_mux_onehot,
         srtarg_0_2_goMux_mux_mux} = {35'd33554432,
                                      lizzieLet17_5QNode_Int_7QNone_Int_10QNone_Int_1_argbuf_d};
      6'd26:
        {srtarg_0_2_goMux_mux_onehot,
         srtarg_0_2_goMux_mux_mux} = {35'd67108864,
                                      lizzieLet27_1_1_argbuf_d};
      6'd27:
        {srtarg_0_2_goMux_mux_onehot,
         srtarg_0_2_goMux_mux_mux} = {35'd134217728,
                                      lizzieLet28_1_1_argbuf_d};
      6'd28:
        {srtarg_0_2_goMux_mux_onehot,
         srtarg_0_2_goMux_mux_mux} = {35'd268435456,
                                      lizzieLet29_1_argbuf_d};
      6'd29:
        {srtarg_0_2_goMux_mux_onehot,
         srtarg_0_2_goMux_mux_mux} = {35'd536870912,
                                      lizzieLet30_1_argbuf_d};
      6'd30:
        {srtarg_0_2_goMux_mux_onehot,
         srtarg_0_2_goMux_mux_mux} = {35'd1073741824,
                                      lizzieLet31_1_1_argbuf_d};
      6'd31:
        {srtarg_0_2_goMux_mux_onehot,
         srtarg_0_2_goMux_mux_mux} = {35'd2147483648,
                                      lizzieLet32_1_1_argbuf_d};
      6'd32:
        {srtarg_0_2_goMux_mux_onehot,
         srtarg_0_2_goMux_mux_mux} = {35'd4294967296,
                                      lizzieLet33_1_1_argbuf_d};
      6'd33:
        {srtarg_0_2_goMux_mux_onehot,
         srtarg_0_2_goMux_mux_mux} = {35'd8589934592,
                                      lizzieLet34_1_1_argbuf_d};
      6'd34:
        {srtarg_0_2_goMux_mux_onehot,
         srtarg_0_2_goMux_mux_mux} = {35'd17179869184,
                                      lizzieLet35_1_argbuf_d};
      default:
        {srtarg_0_2_goMux_mux_onehot, srtarg_0_2_goMux_mux_mux} = {35'd0,
                                                                   {16'd0, 1'd0}};
    endcase
  assign srtarg_0_2_goMux_mux_d = {srtarg_0_2_goMux_mux_mux[16:1],
                                   (srtarg_0_2_goMux_mux_mux[0] && go_15_goMux_choice_1_d[0])};
  assign go_15_goMux_choice_1_r = (srtarg_0_2_goMux_mux_d[0] && srtarg_0_2_goMux_mux_r);
  assign {lizzieLet35_1_argbuf_r,
          lizzieLet34_1_1_argbuf_r,
          lizzieLet33_1_1_argbuf_r,
          lizzieLet32_1_1_argbuf_r,
          lizzieLet31_1_1_argbuf_r,
          lizzieLet30_1_argbuf_r,
          lizzieLet29_1_argbuf_r,
          lizzieLet28_1_1_argbuf_r,
          lizzieLet27_1_1_argbuf_r,
          lizzieLet17_5QNode_Int_7QNone_Int_10QNone_Int_1_argbuf_r,
          lizzieLet26_1_1_argbuf_r,
          lizzieLet25_1_1_argbuf_r,
          es_14_7MyTrue_1_argbuf_r,
          lizzieLet24_1_argbuf_r,
          lizzieLet23_1_1_argbuf_r,
          lizzieLet22_1_1_argbuf_r,
          lizzieLet21_1_1_argbuf_r,
          lizzieLet20_1_1_argbuf_r,
          lizzieLet19_1_1_argbuf_r,
          lizzieLet18_1_1_argbuf_r,
          lizzieLet17_1_1_argbuf_r,
          lizzieLet16_1_1_argbuf_r,
          lizzieLet17_5QVal_Int_7QNone_Int_8QNone_Int_1_argbuf_r,
          lizzieLet15_1_1_argbuf_r,
          lizzieLet14_1_1_argbuf_r,
          lizzieLet13_1_1_argbuf_r,
          lizzieLet12_1_argbuf_r,
          lizzieLet17_5QNone_Int_7QNode_Int_7QNone_Int_1_argbuf_r,
          lizzieLet11_1_1_argbuf_r,
          lizzieLet10_1_1_argbuf_r,
          lizzieLet9_1_1_argbuf_r,
          lizzieLet8_1_1_argbuf_r,
          lizzieLet17_5QNone_Int_7QVal_Int_7QNone_Int_1_argbuf_r,
          contRet_0_2_1_argbuf_r,
          lizzieLet17_5QNone_Int_9QNone_Int_1_argbuf_r} = (go_15_goMux_choice_1_r ? srtarg_0_2_goMux_mux_onehot :
                                                           35'd0);
  
  /* mux (Ty C35,
     Ty Pointer_CTf_f_Int) : (go_15_goMux_choice_2,C35) [(lizzieLet17_5QNone_Int_4QNone_Int_1_argbuf,Pointer_CTf_f_Int),
                                                         (sc_0_14_1_argbuf,Pointer_CTf_f_Int),
                                                         (lizzieLet17_5QNone_Int_7QVal_Int_4QNone_Int_1_argbuf,Pointer_CTf_f_Int),
                                                         (es_2_1_2MyFalse_1_argbuf,Pointer_CTf_f_Int),
                                                         (es_2_1_2MyTrue_1_argbuf,Pointer_CTf_f_Int),
                                                         (lizzieLet17_5QNone_Int_7QVal_Int_4QNode_Int_1_argbuf,Pointer_CTf_f_Int),
                                                         (lizzieLet17_5QNone_Int_7QVal_Int_4QError_Int_1_argbuf,Pointer_CTf_f_Int),
                                                         (lizzieLet17_5QNone_Int_7QNode_Int_4QNone_Int_1_argbuf,Pointer_CTf_f_Int),
                                                         (lizzieLet17_5QNone_Int_7QNode_Int_4QVal_Int_1_argbuf,Pointer_CTf_f_Int),
                                                         (lizzieLet17_5QNone_Int_7QNode_Int_4QNode_Int_1_argbuf,Pointer_CTf_f_Int),
                                                         (lizzieLet17_5QNone_Int_7QNode_Int_4QError_Int_1_argbuf,Pointer_CTf_f_Int),
                                                         (lizzieLet17_5QNone_Int_4QError_Int_1_argbuf,Pointer_CTf_f_Int),
                                                         (lizzieLet17_5QVal_Int_7QNone_Int_5QNone_Int_1_argbuf,Pointer_CTf_f_Int),
                                                         (es_10_3MyFalse_1_argbuf,Pointer_CTf_f_Int),
                                                         (es_10_3MyTrue_1_argbuf,Pointer_CTf_f_Int),
                                                         (lizzieLet17_5QVal_Int_7QNone_Int_5QNode_Int_1_argbuf,Pointer_CTf_f_Int),
                                                         (lizzieLet17_5QVal_Int_7QNone_Int_5QError_Int_1_argbuf,Pointer_CTf_f_Int),
                                                         (es_14_6MyFalse_5QNone_Int_1_argbuf,Pointer_CTf_f_Int),
                                                         (es_21_3MyFalse_1_argbuf,Pointer_CTf_f_Int),
                                                         (es_21_3MyTrue_1_argbuf,Pointer_CTf_f_Int),
                                                         (es_14_6MyFalse_5QNode_Int_1_argbuf,Pointer_CTf_f_Int),
                                                         (es_14_6MyFalse_5QError_Int_1_argbuf,Pointer_CTf_f_Int),
                                                         (es_14_3MyTrue_1_argbuf,Pointer_CTf_f_Int),
                                                         (lizzieLet17_5QVal_Int_4QNode_Int_1_argbuf,Pointer_CTf_f_Int),
                                                         (lizzieLet17_5QVal_Int_4QError_Int_1_argbuf,Pointer_CTf_f_Int),
                                                         (lizzieLet17_5QNode_Int_7QNone_Int_7QNone_Int_1_argbuf,Pointer_CTf_f_Int),
                                                         (lizzieLet17_5QNode_Int_7QNone_Int_7QVal_Int_1_argbuf,Pointer_CTf_f_Int),
                                                         (lizzieLet17_5QNode_Int_7QNone_Int_7QNode_Int_1_argbuf,Pointer_CTf_f_Int),
                                                         (lizzieLet17_5QNode_Int_7QNone_Int_7QError_Int_1_argbuf,Pointer_CTf_f_Int),
                                                         (lizzieLet17_5QNode_Int_4QVal_Int_1_argbuf,Pointer_CTf_f_Int),
                                                         (lizzieLet17_5QNode_Int_7QNode_Int_7QNone_Int_1_argbuf,Pointer_CTf_f_Int),
                                                         (lizzieLet17_5QNode_Int_7QNode_Int_7QVal_Int_1_argbuf,Pointer_CTf_f_Int),
                                                         (lizzieLet17_5QNode_Int_7QNode_Int_7QError_Int_1_argbuf,Pointer_CTf_f_Int),
                                                         (lizzieLet17_5QNode_Int_4QError_Int_1_argbuf,Pointer_CTf_f_Int),
                                                         (lizzieLet17_11QError_Int_1_argbuf,Pointer_CTf_f_Int)] > (scfarg_0_2_goMux_mux,Pointer_CTf_f_Int) */
  logic [16:0] scfarg_0_2_goMux_mux_mux;
  logic [34:0] scfarg_0_2_goMux_mux_onehot;
  always_comb
    unique case (go_15_goMux_choice_2_d[6:1])
      6'd0:
        {scfarg_0_2_goMux_mux_onehot, scfarg_0_2_goMux_mux_mux} = {35'd1,
                                                                   lizzieLet17_5QNone_Int_4QNone_Int_1_argbuf_d};
      6'd1:
        {scfarg_0_2_goMux_mux_onehot, scfarg_0_2_goMux_mux_mux} = {35'd2,
                                                                   sc_0_14_1_argbuf_d};
      6'd2:
        {scfarg_0_2_goMux_mux_onehot, scfarg_0_2_goMux_mux_mux} = {35'd4,
                                                                   lizzieLet17_5QNone_Int_7QVal_Int_4QNone_Int_1_argbuf_d};
      6'd3:
        {scfarg_0_2_goMux_mux_onehot, scfarg_0_2_goMux_mux_mux} = {35'd8,
                                                                   es_2_1_2MyFalse_1_argbuf_d};
      6'd4:
        {scfarg_0_2_goMux_mux_onehot, scfarg_0_2_goMux_mux_mux} = {35'd16,
                                                                   es_2_1_2MyTrue_1_argbuf_d};
      6'd5:
        {scfarg_0_2_goMux_mux_onehot, scfarg_0_2_goMux_mux_mux} = {35'd32,
                                                                   lizzieLet17_5QNone_Int_7QVal_Int_4QNode_Int_1_argbuf_d};
      6'd6:
        {scfarg_0_2_goMux_mux_onehot, scfarg_0_2_goMux_mux_mux} = {35'd64,
                                                                   lizzieLet17_5QNone_Int_7QVal_Int_4QError_Int_1_argbuf_d};
      6'd7:
        {scfarg_0_2_goMux_mux_onehot, scfarg_0_2_goMux_mux_mux} = {35'd128,
                                                                   lizzieLet17_5QNone_Int_7QNode_Int_4QNone_Int_1_argbuf_d};
      6'd8:
        {scfarg_0_2_goMux_mux_onehot, scfarg_0_2_goMux_mux_mux} = {35'd256,
                                                                   lizzieLet17_5QNone_Int_7QNode_Int_4QVal_Int_1_argbuf_d};
      6'd9:
        {scfarg_0_2_goMux_mux_onehot, scfarg_0_2_goMux_mux_mux} = {35'd512,
                                                                   lizzieLet17_5QNone_Int_7QNode_Int_4QNode_Int_1_argbuf_d};
      6'd10:
        {scfarg_0_2_goMux_mux_onehot,
         scfarg_0_2_goMux_mux_mux} = {35'd1024,
                                      lizzieLet17_5QNone_Int_7QNode_Int_4QError_Int_1_argbuf_d};
      6'd11:
        {scfarg_0_2_goMux_mux_onehot,
         scfarg_0_2_goMux_mux_mux} = {35'd2048,
                                      lizzieLet17_5QNone_Int_4QError_Int_1_argbuf_d};
      6'd12:
        {scfarg_0_2_goMux_mux_onehot,
         scfarg_0_2_goMux_mux_mux} = {35'd4096,
                                      lizzieLet17_5QVal_Int_7QNone_Int_5QNone_Int_1_argbuf_d};
      6'd13:
        {scfarg_0_2_goMux_mux_onehot,
         scfarg_0_2_goMux_mux_mux} = {35'd8192, es_10_3MyFalse_1_argbuf_d};
      6'd14:
        {scfarg_0_2_goMux_mux_onehot,
         scfarg_0_2_goMux_mux_mux} = {35'd16384, es_10_3MyTrue_1_argbuf_d};
      6'd15:
        {scfarg_0_2_goMux_mux_onehot,
         scfarg_0_2_goMux_mux_mux} = {35'd32768,
                                      lizzieLet17_5QVal_Int_7QNone_Int_5QNode_Int_1_argbuf_d};
      6'd16:
        {scfarg_0_2_goMux_mux_onehot,
         scfarg_0_2_goMux_mux_mux} = {35'd65536,
                                      lizzieLet17_5QVal_Int_7QNone_Int_5QError_Int_1_argbuf_d};
      6'd17:
        {scfarg_0_2_goMux_mux_onehot,
         scfarg_0_2_goMux_mux_mux} = {35'd131072,
                                      es_14_6MyFalse_5QNone_Int_1_argbuf_d};
      6'd18:
        {scfarg_0_2_goMux_mux_onehot,
         scfarg_0_2_goMux_mux_mux} = {35'd262144,
                                      es_21_3MyFalse_1_argbuf_d};
      6'd19:
        {scfarg_0_2_goMux_mux_onehot,
         scfarg_0_2_goMux_mux_mux} = {35'd524288, es_21_3MyTrue_1_argbuf_d};
      6'd20:
        {scfarg_0_2_goMux_mux_onehot,
         scfarg_0_2_goMux_mux_mux} = {35'd1048576,
                                      es_14_6MyFalse_5QNode_Int_1_argbuf_d};
      6'd21:
        {scfarg_0_2_goMux_mux_onehot,
         scfarg_0_2_goMux_mux_mux} = {35'd2097152,
                                      es_14_6MyFalse_5QError_Int_1_argbuf_d};
      6'd22:
        {scfarg_0_2_goMux_mux_onehot,
         scfarg_0_2_goMux_mux_mux} = {35'd4194304,
                                      es_14_3MyTrue_1_argbuf_d};
      6'd23:
        {scfarg_0_2_goMux_mux_onehot,
         scfarg_0_2_goMux_mux_mux} = {35'd8388608,
                                      lizzieLet17_5QVal_Int_4QNode_Int_1_argbuf_d};
      6'd24:
        {scfarg_0_2_goMux_mux_onehot,
         scfarg_0_2_goMux_mux_mux} = {35'd16777216,
                                      lizzieLet17_5QVal_Int_4QError_Int_1_argbuf_d};
      6'd25:
        {scfarg_0_2_goMux_mux_onehot,
         scfarg_0_2_goMux_mux_mux} = {35'd33554432,
                                      lizzieLet17_5QNode_Int_7QNone_Int_7QNone_Int_1_argbuf_d};
      6'd26:
        {scfarg_0_2_goMux_mux_onehot,
         scfarg_0_2_goMux_mux_mux} = {35'd67108864,
                                      lizzieLet17_5QNode_Int_7QNone_Int_7QVal_Int_1_argbuf_d};
      6'd27:
        {scfarg_0_2_goMux_mux_onehot,
         scfarg_0_2_goMux_mux_mux} = {35'd134217728,
                                      lizzieLet17_5QNode_Int_7QNone_Int_7QNode_Int_1_argbuf_d};
      6'd28:
        {scfarg_0_2_goMux_mux_onehot,
         scfarg_0_2_goMux_mux_mux} = {35'd268435456,
                                      lizzieLet17_5QNode_Int_7QNone_Int_7QError_Int_1_argbuf_d};
      6'd29:
        {scfarg_0_2_goMux_mux_onehot,
         scfarg_0_2_goMux_mux_mux} = {35'd536870912,
                                      lizzieLet17_5QNode_Int_4QVal_Int_1_argbuf_d};
      6'd30:
        {scfarg_0_2_goMux_mux_onehot,
         scfarg_0_2_goMux_mux_mux} = {35'd1073741824,
                                      lizzieLet17_5QNode_Int_7QNode_Int_7QNone_Int_1_argbuf_d};
      6'd31:
        {scfarg_0_2_goMux_mux_onehot,
         scfarg_0_2_goMux_mux_mux} = {35'd2147483648,
                                      lizzieLet17_5QNode_Int_7QNode_Int_7QVal_Int_1_argbuf_d};
      6'd32:
        {scfarg_0_2_goMux_mux_onehot,
         scfarg_0_2_goMux_mux_mux} = {35'd4294967296,
                                      lizzieLet17_5QNode_Int_7QNode_Int_7QError_Int_1_argbuf_d};
      6'd33:
        {scfarg_0_2_goMux_mux_onehot,
         scfarg_0_2_goMux_mux_mux} = {35'd8589934592,
                                      lizzieLet17_5QNode_Int_4QError_Int_1_argbuf_d};
      6'd34:
        {scfarg_0_2_goMux_mux_onehot,
         scfarg_0_2_goMux_mux_mux} = {35'd17179869184,
                                      lizzieLet17_11QError_Int_1_argbuf_d};
      default:
        {scfarg_0_2_goMux_mux_onehot, scfarg_0_2_goMux_mux_mux} = {35'd0,
                                                                   {16'd0, 1'd0}};
    endcase
  assign scfarg_0_2_goMux_mux_d = {scfarg_0_2_goMux_mux_mux[16:1],
                                   (scfarg_0_2_goMux_mux_mux[0] && go_15_goMux_choice_2_d[0])};
  assign go_15_goMux_choice_2_r = (scfarg_0_2_goMux_mux_d[0] && scfarg_0_2_goMux_mux_r);
  assign {lizzieLet17_11QError_Int_1_argbuf_r,
          lizzieLet17_5QNode_Int_4QError_Int_1_argbuf_r,
          lizzieLet17_5QNode_Int_7QNode_Int_7QError_Int_1_argbuf_r,
          lizzieLet17_5QNode_Int_7QNode_Int_7QVal_Int_1_argbuf_r,
          lizzieLet17_5QNode_Int_7QNode_Int_7QNone_Int_1_argbuf_r,
          lizzieLet17_5QNode_Int_4QVal_Int_1_argbuf_r,
          lizzieLet17_5QNode_Int_7QNone_Int_7QError_Int_1_argbuf_r,
          lizzieLet17_5QNode_Int_7QNone_Int_7QNode_Int_1_argbuf_r,
          lizzieLet17_5QNode_Int_7QNone_Int_7QVal_Int_1_argbuf_r,
          lizzieLet17_5QNode_Int_7QNone_Int_7QNone_Int_1_argbuf_r,
          lizzieLet17_5QVal_Int_4QError_Int_1_argbuf_r,
          lizzieLet17_5QVal_Int_4QNode_Int_1_argbuf_r,
          es_14_3MyTrue_1_argbuf_r,
          es_14_6MyFalse_5QError_Int_1_argbuf_r,
          es_14_6MyFalse_5QNode_Int_1_argbuf_r,
          es_21_3MyTrue_1_argbuf_r,
          es_21_3MyFalse_1_argbuf_r,
          es_14_6MyFalse_5QNone_Int_1_argbuf_r,
          lizzieLet17_5QVal_Int_7QNone_Int_5QError_Int_1_argbuf_r,
          lizzieLet17_5QVal_Int_7QNone_Int_5QNode_Int_1_argbuf_r,
          es_10_3MyTrue_1_argbuf_r,
          es_10_3MyFalse_1_argbuf_r,
          lizzieLet17_5QVal_Int_7QNone_Int_5QNone_Int_1_argbuf_r,
          lizzieLet17_5QNone_Int_4QError_Int_1_argbuf_r,
          lizzieLet17_5QNone_Int_7QNode_Int_4QError_Int_1_argbuf_r,
          lizzieLet17_5QNone_Int_7QNode_Int_4QNode_Int_1_argbuf_r,
          lizzieLet17_5QNone_Int_7QNode_Int_4QVal_Int_1_argbuf_r,
          lizzieLet17_5QNone_Int_7QNode_Int_4QNone_Int_1_argbuf_r,
          lizzieLet17_5QNone_Int_7QVal_Int_4QError_Int_1_argbuf_r,
          lizzieLet17_5QNone_Int_7QVal_Int_4QNode_Int_1_argbuf_r,
          es_2_1_2MyTrue_1_argbuf_r,
          es_2_1_2MyFalse_1_argbuf_r,
          lizzieLet17_5QNone_Int_7QVal_Int_4QNone_Int_1_argbuf_r,
          sc_0_14_1_argbuf_r,
          lizzieLet17_5QNone_Int_4QNone_Int_1_argbuf_r} = (go_15_goMux_choice_2_r ? scfarg_0_2_goMux_mux_onehot :
                                                           35'd0);
  
  /* buf (Ty MyDTInt_Int_Int) : (go_1Dcon_$fNumInt_$c+,MyDTInt_Int_Int) > (es_5_1_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t \go_1Dcon_$fNumInt_$c+_bufchan_d ;
  logic \go_1Dcon_$fNumInt_$c+_bufchan_r ;
  assign \go_1Dcon_$fNumInt_$c+_r  = ((! \go_1Dcon_$fNumInt_$c+_bufchan_d [0]) || \go_1Dcon_$fNumInt_$c+_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \go_1Dcon_$fNumInt_$c+_bufchan_d  <= 1'd0;
    else
      if (\go_1Dcon_$fNumInt_$c+_r )
        \go_1Dcon_$fNumInt_$c+_bufchan_d  <= \go_1Dcon_$fNumInt_$c+_d ;
  MyDTInt_Int_Int_t \go_1Dcon_$fNumInt_$c+_bufchan_buf ;
  assign \go_1Dcon_$fNumInt_$c+_bufchan_r  = (! \go_1Dcon_$fNumInt_$c+_bufchan_buf [0]);
  assign es_5_1_argbuf_d = (\go_1Dcon_$fNumInt_$c+_bufchan_buf [0] ? \go_1Dcon_$fNumInt_$c+_bufchan_buf  :
                            \go_1Dcon_$fNumInt_$c+_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \go_1Dcon_$fNumInt_$c+_bufchan_buf  <= 1'd0;
    else
      if ((es_5_1_argbuf_r && \go_1Dcon_$fNumInt_$c+_bufchan_buf [0]))
        \go_1Dcon_$fNumInt_$c+_bufchan_buf  <= 1'd0;
      else if (((! es_5_1_argbuf_r) && (! \go_1Dcon_$fNumInt_$c+_bufchan_buf [0])))
        \go_1Dcon_$fNumInt_$c+_bufchan_buf  <= \go_1Dcon_$fNumInt_$c+_bufchan_d ;
  
  /* dcon (Ty MyDTInt_Bool,
      Dcon Dcon_isZ) : [(go_2,Go)] > (go_2Dcon_isZ,MyDTInt_Bool) */
  assign go_2Dcon_isZ_d = Dcon_isZ_dc((& {go_2_d[0]}), go_2_d);
  assign {go_2_r} = {1 {(go_2Dcon_isZ_r && go_2Dcon_isZ_d[0])}};
  
  /* buf (Ty MyDTInt_Bool) : (go_2Dcon_isZ,MyDTInt_Bool) > (es_4_1_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t go_2Dcon_isZ_bufchan_d;
  logic go_2Dcon_isZ_bufchan_r;
  assign go_2Dcon_isZ_r = ((! go_2Dcon_isZ_bufchan_d[0]) || go_2Dcon_isZ_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_2Dcon_isZ_bufchan_d <= 1'd0;
    else if (go_2Dcon_isZ_r) go_2Dcon_isZ_bufchan_d <= go_2Dcon_isZ_d;
  MyDTInt_Bool_t go_2Dcon_isZ_bufchan_buf;
  assign go_2Dcon_isZ_bufchan_r = (! go_2Dcon_isZ_bufchan_buf[0]);
  assign es_4_1_argbuf_d = (go_2Dcon_isZ_bufchan_buf[0] ? go_2Dcon_isZ_bufchan_buf :
                            go_2Dcon_isZ_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_2Dcon_isZ_bufchan_buf <= 1'd0;
    else
      if ((es_4_1_argbuf_r && go_2Dcon_isZ_bufchan_buf[0]))
        go_2Dcon_isZ_bufchan_buf <= 1'd0;
      else if (((! es_4_1_argbuf_r) && (! go_2Dcon_isZ_bufchan_buf[0])))
        go_2Dcon_isZ_bufchan_buf <= go_2Dcon_isZ_bufchan_d;
  
  /* buf (Ty Go) : (go_3,Go) > (go_3_argbuf,Go) */
  Go_t go_3_bufchan_d;
  logic go_3_bufchan_r;
  assign go_3_r = ((! go_3_bufchan_d[0]) || go_3_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_3_bufchan_d <= 1'd0;
    else if (go_3_r) go_3_bufchan_d <= go_3_d;
  Go_t go_3_bufchan_buf;
  assign go_3_bufchan_r = (! go_3_bufchan_buf[0]);
  assign go_3_argbuf_d = (go_3_bufchan_buf[0] ? go_3_bufchan_buf :
                          go_3_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_3_bufchan_buf <= 1'd0;
    else
      if ((go_3_argbuf_r && go_3_bufchan_buf[0]))
        go_3_bufchan_buf <= 1'd0;
      else if (((! go_3_argbuf_r) && (! go_3_bufchan_buf[0])))
        go_3_bufchan_buf <= go_3_bufchan_d;
  
  /* dcon (Ty TupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int,
      Dcon TupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int) : [(go_3_argbuf,Go),
                                                                                                                  (m1aen_0,Pointer_QTree_Int),
                                                                                                                  (m2aeo_1,Pointer_QTree_Int),
                                                                                                                  (m3aep_2,Pointer_QTree_Int),
                                                                                                                  (es_4_1_argbuf,MyDTInt_Bool),
                                                                                                                  (es_5_1_argbuf,MyDTInt_Int_Int)] > (f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1,TupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int) */
  assign f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_d = TupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_dc((& {go_3_argbuf_d[0],
                                                                                                                                                                                                                                   m1aen_0_d[0],
                                                                                                                                                                                                                                   m2aeo_1_d[0],
                                                                                                                                                                                                                                   m3aep_2_d[0],
                                                                                                                                                                                                                                   es_4_1_argbuf_d[0],
                                                                                                                                                                                                                                   es_5_1_argbuf_d[0]}), go_3_argbuf_d, m1aen_0_d, m2aeo_1_d, m3aep_2_d, es_4_1_argbuf_d, es_5_1_argbuf_d);
  assign {go_3_argbuf_r,
          m1aen_0_r,
          m2aeo_1_r,
          m3aep_2_r,
          es_4_1_argbuf_r,
          es_5_1_argbuf_r} = {6 {(f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_r && f_f_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_d[0])}};
  
  /* buf (Ty Go) : (go_4,Go) > (go_4_argbuf,Go) */
  Go_t go_4_bufchan_d;
  logic go_4_bufchan_r;
  assign go_4_r = ((! go_4_bufchan_d[0]) || go_4_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_4_bufchan_d <= 1'd0;
    else if (go_4_r) go_4_bufchan_d <= go_4_d;
  Go_t go_4_bufchan_buf;
  assign go_4_bufchan_r = (! go_4_bufchan_buf[0]);
  assign go_4_argbuf_d = (go_4_bufchan_buf[0] ? go_4_bufchan_buf :
                          go_4_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_4_bufchan_buf <= 1'd0;
    else
      if ((go_4_argbuf_r && go_4_bufchan_buf[0]))
        go_4_bufchan_buf <= 1'd0;
      else if (((! go_4_argbuf_r) && (! go_4_bufchan_buf[0])))
        go_4_bufchan_buf <= go_4_bufchan_d;
  
  /* dcon (Ty TupGo___Pointer_QTree_Int,
      Dcon TupGo___Pointer_QTree_Int) : [(go_4_argbuf,Go),
                                         (es_0_1_argbuf,Pointer_QTree_Int)] > ($wnnzTupGo___Pointer_QTree_Int_1,TupGo___Pointer_QTree_Int) */
  assign \$wnnzTupGo___Pointer_QTree_Int_1_d  = TupGo___Pointer_QTree_Int_dc((& {go_4_argbuf_d[0],
                                                                                 es_0_1_argbuf_d[0]}), go_4_argbuf_d, es_0_1_argbuf_d);
  assign {go_4_argbuf_r,
          es_0_1_argbuf_r} = {2 {(\$wnnzTupGo___Pointer_QTree_Int_1_r  && \$wnnzTupGo___Pointer_QTree_Int_1_d [0])}};
  
  /* dcon (Ty CT$wnnz,
      Dcon L$wnnzsbos) : [(go_6_1,Go)] > (go_6_1L$wnnzsbos,CT$wnnz) */
  assign go_6_1L$wnnzsbos_d = L$wnnzsbos_dc((& {go_6_1_d[0]}), go_6_1_d);
  assign {go_6_1_r} = {1 {(go_6_1L$wnnzsbos_r && go_6_1L$wnnzsbos_d[0])}};
  
  /* buf (Ty CT$wnnz) : (go_6_1L$wnnzsbos,CT$wnnz) > (lizzieLet0_1_argbuf,CT$wnnz) */
  CT$wnnz_t go_6_1L$wnnzsbos_bufchan_d;
  logic go_6_1L$wnnzsbos_bufchan_r;
  assign go_6_1L$wnnzsbos_r = ((! go_6_1L$wnnzsbos_bufchan_d[0]) || go_6_1L$wnnzsbos_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_6_1L$wnnzsbos_bufchan_d <= {115'd0, 1'd0};
    else
      if (go_6_1L$wnnzsbos_r)
        go_6_1L$wnnzsbos_bufchan_d <= go_6_1L$wnnzsbos_d;
  CT$wnnz_t go_6_1L$wnnzsbos_bufchan_buf;
  assign go_6_1L$wnnzsbos_bufchan_r = (! go_6_1L$wnnzsbos_bufchan_buf[0]);
  assign lizzieLet0_1_argbuf_d = (go_6_1L$wnnzsbos_bufchan_buf[0] ? go_6_1L$wnnzsbos_bufchan_buf :
                                  go_6_1L$wnnzsbos_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      go_6_1L$wnnzsbos_bufchan_buf <= {115'd0, 1'd0};
    else
      if ((lizzieLet0_1_argbuf_r && go_6_1L$wnnzsbos_bufchan_buf[0]))
        go_6_1L$wnnzsbos_bufchan_buf <= {115'd0, 1'd0};
      else if (((! lizzieLet0_1_argbuf_r) && (! go_6_1L$wnnzsbos_bufchan_buf[0])))
        go_6_1L$wnnzsbos_bufchan_buf <= go_6_1L$wnnzsbos_bufchan_d;
  
  /* buf (Ty Go) : (go_6_2,Go) > (go_6_2_argbuf,Go) */
  Go_t go_6_2_bufchan_d;
  logic go_6_2_bufchan_r;
  assign go_6_2_r = ((! go_6_2_bufchan_d[0]) || go_6_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_6_2_bufchan_d <= 1'd0;
    else if (go_6_2_r) go_6_2_bufchan_d <= go_6_2_d;
  Go_t go_6_2_bufchan_buf;
  assign go_6_2_bufchan_r = (! go_6_2_bufchan_buf[0]);
  assign go_6_2_argbuf_d = (go_6_2_bufchan_buf[0] ? go_6_2_bufchan_buf :
                            go_6_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_6_2_bufchan_buf <= 1'd0;
    else
      if ((go_6_2_argbuf_r && go_6_2_bufchan_buf[0]))
        go_6_2_bufchan_buf <= 1'd0;
      else if (((! go_6_2_argbuf_r) && (! go_6_2_bufchan_buf[0])))
        go_6_2_bufchan_buf <= go_6_2_bufchan_d;
  
  /* dcon (Ty TupGo___Pointer_QTree_Int___Pointer_CT$wnnz,
      Dcon TupGo___Pointer_QTree_Int___Pointer_CT$wnnz) : [(go_6_2_argbuf,Go),
                                                           (wsmk_1_argbuf,Pointer_QTree_Int),
                                                           (lizzieLet39_1_argbuf,Pointer_CT$wnnz)] > (call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_1,TupGo___Pointer_QTree_Int___Pointer_CT$wnnz) */
  assign call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_1_d = TupGo___Pointer_QTree_Int___Pointer_CT$wnnz_dc((& {go_6_2_argbuf_d[0],
                                                                                                                        wsmk_1_argbuf_d[0],
                                                                                                                        lizzieLet39_1_argbuf_d[0]}), go_6_2_argbuf_d, wsmk_1_argbuf_d, lizzieLet39_1_argbuf_d);
  assign {go_6_2_argbuf_r,
          wsmk_1_argbuf_r,
          lizzieLet39_1_argbuf_r} = {3 {(call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_1_r && call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_1_d[0])}};
  
  /* fork (Ty C5) : (go_8_goMux_choice,C5) > [(go_8_goMux_choice_1,C5),
                                         (go_8_goMux_choice_2,C5)] */
  logic [1:0] go_8_goMux_choice_emitted;
  logic [1:0] go_8_goMux_choice_done;
  assign go_8_goMux_choice_1_d = {go_8_goMux_choice_d[3:1],
                                  (go_8_goMux_choice_d[0] && (! go_8_goMux_choice_emitted[0]))};
  assign go_8_goMux_choice_2_d = {go_8_goMux_choice_d[3:1],
                                  (go_8_goMux_choice_d[0] && (! go_8_goMux_choice_emitted[1]))};
  assign go_8_goMux_choice_done = (go_8_goMux_choice_emitted | ({go_8_goMux_choice_2_d[0],
                                                                 go_8_goMux_choice_1_d[0]} & {go_8_goMux_choice_2_r,
                                                                                              go_8_goMux_choice_1_r}));
  assign go_8_goMux_choice_r = (& go_8_goMux_choice_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_8_goMux_choice_emitted <= 2'd0;
    else
      go_8_goMux_choice_emitted <= (go_8_goMux_choice_r ? 2'd0 :
                                    go_8_goMux_choice_done);
  
  /* mux (Ty C5,
     Ty Pointer_QTree_Int) : (go_8_goMux_choice_1,C5) [(call_$wnnz_goMux2,Pointer_QTree_Int),
                                                       (q2a8s_1_1_argbuf,Pointer_QTree_Int),
                                                       (q3a8t_2_1_argbuf,Pointer_QTree_Int),
                                                       (q4a8u_3_1_argbuf,Pointer_QTree_Int),
                                                       (q1a8r_1_argbuf,Pointer_QTree_Int)] > (wsmk_1_goMux_mux,Pointer_QTree_Int) */
  logic [16:0] wsmk_1_goMux_mux_mux;
  logic [4:0] wsmk_1_goMux_mux_onehot;
  always_comb
    unique case (go_8_goMux_choice_1_d[3:1])
      3'd0:
        {wsmk_1_goMux_mux_onehot, wsmk_1_goMux_mux_mux} = {5'd1,
                                                           call_$wnnz_goMux2_d};
      3'd1:
        {wsmk_1_goMux_mux_onehot, wsmk_1_goMux_mux_mux} = {5'd2,
                                                           q2a8s_1_1_argbuf_d};
      3'd2:
        {wsmk_1_goMux_mux_onehot, wsmk_1_goMux_mux_mux} = {5'd4,
                                                           q3a8t_2_1_argbuf_d};
      3'd3:
        {wsmk_1_goMux_mux_onehot, wsmk_1_goMux_mux_mux} = {5'd8,
                                                           q4a8u_3_1_argbuf_d};
      3'd4:
        {wsmk_1_goMux_mux_onehot, wsmk_1_goMux_mux_mux} = {5'd16,
                                                           q1a8r_1_argbuf_d};
      default:
        {wsmk_1_goMux_mux_onehot, wsmk_1_goMux_mux_mux} = {5'd0,
                                                           {16'd0, 1'd0}};
    endcase
  assign wsmk_1_goMux_mux_d = {wsmk_1_goMux_mux_mux[16:1],
                               (wsmk_1_goMux_mux_mux[0] && go_8_goMux_choice_1_d[0])};
  assign go_8_goMux_choice_1_r = (wsmk_1_goMux_mux_d[0] && wsmk_1_goMux_mux_r);
  assign {q1a8r_1_argbuf_r,
          q4a8u_3_1_argbuf_r,
          q3a8t_2_1_argbuf_r,
          q2a8s_1_1_argbuf_r,
          call_$wnnz_goMux2_r} = (go_8_goMux_choice_1_r ? wsmk_1_goMux_mux_onehot :
                                  5'd0);
  
  /* mux (Ty C5,
     Ty Pointer_CT$wnnz) : (go_8_goMux_choice_2,C5) [(call_$wnnz_goMux3,Pointer_CT$wnnz),
                                                     (sca2_1_argbuf,Pointer_CT$wnnz),
                                                     (sca1_1_argbuf,Pointer_CT$wnnz),
                                                     (sca0_1_argbuf,Pointer_CT$wnnz),
                                                     (sca3_1_argbuf,Pointer_CT$wnnz)] > (sc_0_goMux_mux,Pointer_CT$wnnz) */
  logic [16:0] sc_0_goMux_mux_mux;
  logic [4:0] sc_0_goMux_mux_onehot;
  always_comb
    unique case (go_8_goMux_choice_2_d[3:1])
      3'd0:
        {sc_0_goMux_mux_onehot, sc_0_goMux_mux_mux} = {5'd1,
                                                       call_$wnnz_goMux3_d};
      3'd1:
        {sc_0_goMux_mux_onehot, sc_0_goMux_mux_mux} = {5'd2,
                                                       sca2_1_argbuf_d};
      3'd2:
        {sc_0_goMux_mux_onehot, sc_0_goMux_mux_mux} = {5'd4,
                                                       sca1_1_argbuf_d};
      3'd3:
        {sc_0_goMux_mux_onehot, sc_0_goMux_mux_mux} = {5'd8,
                                                       sca0_1_argbuf_d};
      3'd4:
        {sc_0_goMux_mux_onehot, sc_0_goMux_mux_mux} = {5'd16,
                                                       sca3_1_argbuf_d};
      default:
        {sc_0_goMux_mux_onehot, sc_0_goMux_mux_mux} = {5'd0,
                                                       {16'd0, 1'd0}};
    endcase
  assign sc_0_goMux_mux_d = {sc_0_goMux_mux_mux[16:1],
                             (sc_0_goMux_mux_mux[0] && go_8_goMux_choice_2_d[0])};
  assign go_8_goMux_choice_2_r = (sc_0_goMux_mux_d[0] && sc_0_goMux_mux_r);
  assign {sca3_1_argbuf_r,
          sca0_1_argbuf_r,
          sca1_1_argbuf_r,
          sca2_1_argbuf_r,
          call_$wnnz_goMux3_r} = (go_8_goMux_choice_2_r ? sc_0_goMux_mux_onehot :
                                  5'd0);
  
  /* fork (Ty C5) : (go_9_goMux_choice,C5) > [(go_9_goMux_choice_1,C5),
                                         (go_9_goMux_choice_2,C5),
                                         (go_9_goMux_choice_3,C5),
                                         (go_9_goMux_choice_4,C5),
                                         (go_9_goMux_choice_5,C5)] */
  logic [4:0] go_9_goMux_choice_emitted;
  logic [4:0] go_9_goMux_choice_done;
  assign go_9_goMux_choice_1_d = {go_9_goMux_choice_d[3:1],
                                  (go_9_goMux_choice_d[0] && (! go_9_goMux_choice_emitted[0]))};
  assign go_9_goMux_choice_2_d = {go_9_goMux_choice_d[3:1],
                                  (go_9_goMux_choice_d[0] && (! go_9_goMux_choice_emitted[1]))};
  assign go_9_goMux_choice_3_d = {go_9_goMux_choice_d[3:1],
                                  (go_9_goMux_choice_d[0] && (! go_9_goMux_choice_emitted[2]))};
  assign go_9_goMux_choice_4_d = {go_9_goMux_choice_d[3:1],
                                  (go_9_goMux_choice_d[0] && (! go_9_goMux_choice_emitted[3]))};
  assign go_9_goMux_choice_5_d = {go_9_goMux_choice_d[3:1],
                                  (go_9_goMux_choice_d[0] && (! go_9_goMux_choice_emitted[4]))};
  assign go_9_goMux_choice_done = (go_9_goMux_choice_emitted | ({go_9_goMux_choice_5_d[0],
                                                                 go_9_goMux_choice_4_d[0],
                                                                 go_9_goMux_choice_3_d[0],
                                                                 go_9_goMux_choice_2_d[0],
                                                                 go_9_goMux_choice_1_d[0]} & {go_9_goMux_choice_5_r,
                                                                                              go_9_goMux_choice_4_r,
                                                                                              go_9_goMux_choice_3_r,
                                                                                              go_9_goMux_choice_2_r,
                                                                                              go_9_goMux_choice_1_r}));
  assign go_9_goMux_choice_r = (& go_9_goMux_choice_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_9_goMux_choice_emitted <= 5'd0;
    else
      go_9_goMux_choice_emitted <= (go_9_goMux_choice_r ? 5'd0 :
                                    go_9_goMux_choice_done);
  
  /* mux (Ty C5,
     Ty Pointer_QTree_Int) : (go_9_goMux_choice_1,C5) [(call_f''''''''''''_f''''''''''''_Int_goMux2,Pointer_QTree_Int),
                                                       (q3afv_1_1_argbuf,Pointer_QTree_Int),
                                                       (q2afu_2_1_argbuf,Pointer_QTree_Int),
                                                       (q1aft_3_1_argbuf,Pointer_QTree_Int),
                                                       (lizzieLet6_5QNode_Int_11QNode_Int_1_argbuf,Pointer_QTree_Int)] > (q4afj_goMux_mux,Pointer_QTree_Int) */
  logic [16:0] q4afj_goMux_mux_mux;
  logic [4:0] q4afj_goMux_mux_onehot;
  always_comb
    unique case (go_9_goMux_choice_1_d[3:1])
      3'd0:
        {q4afj_goMux_mux_onehot, q4afj_goMux_mux_mux} = {5'd1,
                                                         \call_f''''''''''''_f''''''''''''_Int_goMux2_d };
      3'd1:
        {q4afj_goMux_mux_onehot, q4afj_goMux_mux_mux} = {5'd2,
                                                         q3afv_1_1_argbuf_d};
      3'd2:
        {q4afj_goMux_mux_onehot, q4afj_goMux_mux_mux} = {5'd4,
                                                         q2afu_2_1_argbuf_d};
      3'd3:
        {q4afj_goMux_mux_onehot, q4afj_goMux_mux_mux} = {5'd8,
                                                         q1aft_3_1_argbuf_d};
      3'd4:
        {q4afj_goMux_mux_onehot, q4afj_goMux_mux_mux} = {5'd16,
                                                         lizzieLet6_5QNode_Int_11QNode_Int_1_argbuf_d};
      default:
        {q4afj_goMux_mux_onehot, q4afj_goMux_mux_mux} = {5'd0,
                                                         {16'd0, 1'd0}};
    endcase
  assign q4afj_goMux_mux_d = {q4afj_goMux_mux_mux[16:1],
                              (q4afj_goMux_mux_mux[0] && go_9_goMux_choice_1_d[0])};
  assign go_9_goMux_choice_1_r = (q4afj_goMux_mux_d[0] && q4afj_goMux_mux_r);
  assign {lizzieLet6_5QNode_Int_11QNode_Int_1_argbuf_r,
          q1aft_3_1_argbuf_r,
          q2afu_2_1_argbuf_r,
          q3afv_1_1_argbuf_r,
          \call_f''''''''''''_f''''''''''''_Int_goMux2_r } = (go_9_goMux_choice_1_r ? q4afj_goMux_mux_onehot :
                                                              5'd0);
  
  /* mux (Ty C5,
     Ty Pointer_QTree_Int) : (go_9_goMux_choice_2,C5) [(call_f''''''''''''_f''''''''''''_Int_goMux3,Pointer_QTree_Int),
                                                       (t3afA_1_1_argbuf,Pointer_QTree_Int),
                                                       (t2afz_2_1_argbuf,Pointer_QTree_Int),
                                                       (t1afy_3_1_argbuf,Pointer_QTree_Int),
                                                       (t5afB_1_argbuf,Pointer_QTree_Int)] > (t4afk_goMux_mux,Pointer_QTree_Int) */
  logic [16:0] t4afk_goMux_mux_mux;
  logic [4:0] t4afk_goMux_mux_onehot;
  always_comb
    unique case (go_9_goMux_choice_2_d[3:1])
      3'd0:
        {t4afk_goMux_mux_onehot, t4afk_goMux_mux_mux} = {5'd1,
                                                         \call_f''''''''''''_f''''''''''''_Int_goMux3_d };
      3'd1:
        {t4afk_goMux_mux_onehot, t4afk_goMux_mux_mux} = {5'd2,
                                                         t3afA_1_1_argbuf_d};
      3'd2:
        {t4afk_goMux_mux_onehot, t4afk_goMux_mux_mux} = {5'd4,
                                                         t2afz_2_1_argbuf_d};
      3'd3:
        {t4afk_goMux_mux_onehot, t4afk_goMux_mux_mux} = {5'd8,
                                                         t1afy_3_1_argbuf_d};
      3'd4:
        {t4afk_goMux_mux_onehot, t4afk_goMux_mux_mux} = {5'd16,
                                                         t5afB_1_argbuf_d};
      default:
        {t4afk_goMux_mux_onehot, t4afk_goMux_mux_mux} = {5'd0,
                                                         {16'd0, 1'd0}};
    endcase
  assign t4afk_goMux_mux_d = {t4afk_goMux_mux_mux[16:1],
                              (t4afk_goMux_mux_mux[0] && go_9_goMux_choice_2_d[0])};
  assign go_9_goMux_choice_2_r = (t4afk_goMux_mux_d[0] && t4afk_goMux_mux_r);
  assign {t5afB_1_argbuf_r,
          t1afy_3_1_argbuf_r,
          t2afz_2_1_argbuf_r,
          t3afA_1_1_argbuf_r,
          \call_f''''''''''''_f''''''''''''_Int_goMux3_r } = (go_9_goMux_choice_2_r ? t4afk_goMux_mux_onehot :
                                                              5'd0);
  
  /* mux (Ty C5,
     Ty MyDTInt_Bool) : (go_9_goMux_choice_3,C5) [(call_f''''''''''''_f''''''''''''_Int_goMux4,MyDTInt_Bool),
                                                  (is_zafl_2_2_argbuf,MyDTInt_Bool),
                                                  (is_zafl_3_2_argbuf,MyDTInt_Bool),
                                                  (is_zafl_4_1_argbuf,MyDTInt_Bool),
                                                  (lizzieLet6_5QNode_Int_4QNode_Int_2_argbuf,MyDTInt_Bool)] > (is_zafl_goMux_mux,MyDTInt_Bool) */
  logic [0:0] is_zafl_goMux_mux_mux;
  logic [4:0] is_zafl_goMux_mux_onehot;
  always_comb
    unique case (go_9_goMux_choice_3_d[3:1])
      3'd0:
        {is_zafl_goMux_mux_onehot, is_zafl_goMux_mux_mux} = {5'd1,
                                                             \call_f''''''''''''_f''''''''''''_Int_goMux4_d };
      3'd1:
        {is_zafl_goMux_mux_onehot, is_zafl_goMux_mux_mux} = {5'd2,
                                                             is_zafl_2_2_argbuf_d};
      3'd2:
        {is_zafl_goMux_mux_onehot, is_zafl_goMux_mux_mux} = {5'd4,
                                                             is_zafl_3_2_argbuf_d};
      3'd3:
        {is_zafl_goMux_mux_onehot, is_zafl_goMux_mux_mux} = {5'd8,
                                                             is_zafl_4_1_argbuf_d};
      3'd4:
        {is_zafl_goMux_mux_onehot, is_zafl_goMux_mux_mux} = {5'd16,
                                                             lizzieLet6_5QNode_Int_4QNode_Int_2_argbuf_d};
      default:
        {is_zafl_goMux_mux_onehot, is_zafl_goMux_mux_mux} = {5'd0, 1'd0};
    endcase
  assign is_zafl_goMux_mux_d = (is_zafl_goMux_mux_mux[0] && go_9_goMux_choice_3_d[0]);
  assign go_9_goMux_choice_3_r = (is_zafl_goMux_mux_d[0] && is_zafl_goMux_mux_r);
  assign {lizzieLet6_5QNode_Int_4QNode_Int_2_argbuf_r,
          is_zafl_4_1_argbuf_r,
          is_zafl_3_2_argbuf_r,
          is_zafl_2_2_argbuf_r,
          \call_f''''''''''''_f''''''''''''_Int_goMux4_r } = (go_9_goMux_choice_3_r ? is_zafl_goMux_mux_onehot :
                                                              5'd0);
  
  /* mux (Ty C5,
     Ty MyDTInt_Int_Int) : (go_9_goMux_choice_4,C5) [(call_f''''''''''''_f''''''''''''_Int_goMux5,MyDTInt_Int_Int),
                                                     (op_addafm_2_2_argbuf,MyDTInt_Int_Int),
                                                     (op_addafm_3_2_argbuf,MyDTInt_Int_Int),
                                                     (op_addafm_4_1_argbuf,MyDTInt_Int_Int),
                                                     (lizzieLet6_5QNode_Int_5QNode_Int_2_argbuf,MyDTInt_Int_Int)] > (op_addafm_goMux_mux,MyDTInt_Int_Int) */
  logic [0:0] op_addafm_goMux_mux_mux;
  logic [4:0] op_addafm_goMux_mux_onehot;
  always_comb
    unique case (go_9_goMux_choice_4_d[3:1])
      3'd0:
        {op_addafm_goMux_mux_onehot, op_addafm_goMux_mux_mux} = {5'd1,
                                                                 \call_f''''''''''''_f''''''''''''_Int_goMux5_d };
      3'd1:
        {op_addafm_goMux_mux_onehot, op_addafm_goMux_mux_mux} = {5'd2,
                                                                 op_addafm_2_2_argbuf_d};
      3'd2:
        {op_addafm_goMux_mux_onehot, op_addafm_goMux_mux_mux} = {5'd4,
                                                                 op_addafm_3_2_argbuf_d};
      3'd3:
        {op_addafm_goMux_mux_onehot, op_addafm_goMux_mux_mux} = {5'd8,
                                                                 op_addafm_4_1_argbuf_d};
      3'd4:
        {op_addafm_goMux_mux_onehot, op_addafm_goMux_mux_mux} = {5'd16,
                                                                 lizzieLet6_5QNode_Int_5QNode_Int_2_argbuf_d};
      default:
        {op_addafm_goMux_mux_onehot, op_addafm_goMux_mux_mux} = {5'd0,
                                                                 1'd0};
    endcase
  assign op_addafm_goMux_mux_d = (op_addafm_goMux_mux_mux[0] && go_9_goMux_choice_4_d[0]);
  assign go_9_goMux_choice_4_r = (op_addafm_goMux_mux_d[0] && op_addafm_goMux_mux_r);
  assign {lizzieLet6_5QNode_Int_5QNode_Int_2_argbuf_r,
          op_addafm_4_1_argbuf_r,
          op_addafm_3_2_argbuf_r,
          op_addafm_2_2_argbuf_r,
          \call_f''''''''''''_f''''''''''''_Int_goMux5_r } = (go_9_goMux_choice_4_r ? op_addafm_goMux_mux_onehot :
                                                              5'd0);
  
  /* mux (Ty C5,
     Ty Pointer_CTf''''''''''''_f''''''''''''_Int) : (go_9_goMux_choice_5,C5) [(call_f''''''''''''_f''''''''''''_Int_goMux6,Pointer_CTf''''''''''''_f''''''''''''_Int),
                                                                               (sca2_1_1_argbuf,Pointer_CTf''''''''''''_f''''''''''''_Int),
                                                                               (sca1_1_1_argbuf,Pointer_CTf''''''''''''_f''''''''''''_Int),
                                                                               (sca0_1_1_argbuf,Pointer_CTf''''''''''''_f''''''''''''_Int),
                                                                               (sca3_1_1_argbuf,Pointer_CTf''''''''''''_f''''''''''''_Int)] > (sc_0_1_goMux_mux,Pointer_CTf''''''''''''_f''''''''''''_Int) */
  logic [16:0] sc_0_1_goMux_mux_mux;
  logic [4:0] sc_0_1_goMux_mux_onehot;
  always_comb
    unique case (go_9_goMux_choice_5_d[3:1])
      3'd0:
        {sc_0_1_goMux_mux_onehot, sc_0_1_goMux_mux_mux} = {5'd1,
                                                           \call_f''''''''''''_f''''''''''''_Int_goMux6_d };
      3'd1:
        {sc_0_1_goMux_mux_onehot, sc_0_1_goMux_mux_mux} = {5'd2,
                                                           sca2_1_1_argbuf_d};
      3'd2:
        {sc_0_1_goMux_mux_onehot, sc_0_1_goMux_mux_mux} = {5'd4,
                                                           sca1_1_1_argbuf_d};
      3'd3:
        {sc_0_1_goMux_mux_onehot, sc_0_1_goMux_mux_mux} = {5'd8,
                                                           sca0_1_1_argbuf_d};
      3'd4:
        {sc_0_1_goMux_mux_onehot, sc_0_1_goMux_mux_mux} = {5'd16,
                                                           sca3_1_1_argbuf_d};
      default:
        {sc_0_1_goMux_mux_onehot, sc_0_1_goMux_mux_mux} = {5'd0,
                                                           {16'd0, 1'd0}};
    endcase
  assign sc_0_1_goMux_mux_d = {sc_0_1_goMux_mux_mux[16:1],
                               (sc_0_1_goMux_mux_mux[0] && go_9_goMux_choice_5_d[0])};
  assign go_9_goMux_choice_5_r = (sc_0_1_goMux_mux_d[0] && sc_0_1_goMux_mux_r);
  assign {sca3_1_1_argbuf_r,
          sca0_1_1_argbuf_r,
          sca1_1_1_argbuf_r,
          sca2_1_1_argbuf_r,
          \call_f''''''''''''_f''''''''''''_Int_goMux6_r } = (go_9_goMux_choice_5_r ? sc_0_1_goMux_mux_onehot :
                                                              5'd0);
  
  /* buf (Ty MyDTInt_Bool) : (is_zaet_2_2,MyDTInt_Bool) > (is_zaet_2_2_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t is_zaet_2_2_bufchan_d;
  logic is_zaet_2_2_bufchan_r;
  assign is_zaet_2_2_r = ((! is_zaet_2_2_bufchan_d[0]) || is_zaet_2_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) is_zaet_2_2_bufchan_d <= 1'd0;
    else if (is_zaet_2_2_r) is_zaet_2_2_bufchan_d <= is_zaet_2_2_d;
  MyDTInt_Bool_t is_zaet_2_2_bufchan_buf;
  assign is_zaet_2_2_bufchan_r = (! is_zaet_2_2_bufchan_buf[0]);
  assign is_zaet_2_2_argbuf_d = (is_zaet_2_2_bufchan_buf[0] ? is_zaet_2_2_bufchan_buf :
                                 is_zaet_2_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) is_zaet_2_2_bufchan_buf <= 1'd0;
    else
      if ((is_zaet_2_2_argbuf_r && is_zaet_2_2_bufchan_buf[0]))
        is_zaet_2_2_bufchan_buf <= 1'd0;
      else if (((! is_zaet_2_2_argbuf_r) && (! is_zaet_2_2_bufchan_buf[0])))
        is_zaet_2_2_bufchan_buf <= is_zaet_2_2_bufchan_d;
  
  /* fork (Ty MyDTInt_Bool) : (is_zaet_2_destruct,MyDTInt_Bool) > [(is_zaet_2_1,MyDTInt_Bool),
                                                              (is_zaet_2_2,MyDTInt_Bool)] */
  logic [1:0] is_zaet_2_destruct_emitted;
  logic [1:0] is_zaet_2_destruct_done;
  assign is_zaet_2_1_d = (is_zaet_2_destruct_d[0] && (! is_zaet_2_destruct_emitted[0]));
  assign is_zaet_2_2_d = (is_zaet_2_destruct_d[0] && (! is_zaet_2_destruct_emitted[1]));
  assign is_zaet_2_destruct_done = (is_zaet_2_destruct_emitted | ({is_zaet_2_2_d[0],
                                                                   is_zaet_2_1_d[0]} & {is_zaet_2_2_r,
                                                                                        is_zaet_2_1_r}));
  assign is_zaet_2_destruct_r = (& is_zaet_2_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) is_zaet_2_destruct_emitted <= 2'd0;
    else
      is_zaet_2_destruct_emitted <= (is_zaet_2_destruct_r ? 2'd0 :
                                     is_zaet_2_destruct_done);
  
  /* buf (Ty MyDTInt_Bool) : (is_zaet_3_2,MyDTInt_Bool) > (is_zaet_3_2_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t is_zaet_3_2_bufchan_d;
  logic is_zaet_3_2_bufchan_r;
  assign is_zaet_3_2_r = ((! is_zaet_3_2_bufchan_d[0]) || is_zaet_3_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) is_zaet_3_2_bufchan_d <= 1'd0;
    else if (is_zaet_3_2_r) is_zaet_3_2_bufchan_d <= is_zaet_3_2_d;
  MyDTInt_Bool_t is_zaet_3_2_bufchan_buf;
  assign is_zaet_3_2_bufchan_r = (! is_zaet_3_2_bufchan_buf[0]);
  assign is_zaet_3_2_argbuf_d = (is_zaet_3_2_bufchan_buf[0] ? is_zaet_3_2_bufchan_buf :
                                 is_zaet_3_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) is_zaet_3_2_bufchan_buf <= 1'd0;
    else
      if ((is_zaet_3_2_argbuf_r && is_zaet_3_2_bufchan_buf[0]))
        is_zaet_3_2_bufchan_buf <= 1'd0;
      else if (((! is_zaet_3_2_argbuf_r) && (! is_zaet_3_2_bufchan_buf[0])))
        is_zaet_3_2_bufchan_buf <= is_zaet_3_2_bufchan_d;
  
  /* fork (Ty MyDTInt_Bool) : (is_zaet_3_destruct,MyDTInt_Bool) > [(is_zaet_3_1,MyDTInt_Bool),
                                                              (is_zaet_3_2,MyDTInt_Bool)] */
  logic [1:0] is_zaet_3_destruct_emitted;
  logic [1:0] is_zaet_3_destruct_done;
  assign is_zaet_3_1_d = (is_zaet_3_destruct_d[0] && (! is_zaet_3_destruct_emitted[0]));
  assign is_zaet_3_2_d = (is_zaet_3_destruct_d[0] && (! is_zaet_3_destruct_emitted[1]));
  assign is_zaet_3_destruct_done = (is_zaet_3_destruct_emitted | ({is_zaet_3_2_d[0],
                                                                   is_zaet_3_1_d[0]} & {is_zaet_3_2_r,
                                                                                        is_zaet_3_1_r}));
  assign is_zaet_3_destruct_r = (& is_zaet_3_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) is_zaet_3_destruct_emitted <= 2'd0;
    else
      is_zaet_3_destruct_emitted <= (is_zaet_3_destruct_r ? 2'd0 :
                                     is_zaet_3_destruct_done);
  
  /* buf (Ty MyDTInt_Bool) : (is_zaet_4_destruct,MyDTInt_Bool) > (is_zaet_4_1_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t is_zaet_4_destruct_bufchan_d;
  logic is_zaet_4_destruct_bufchan_r;
  assign is_zaet_4_destruct_r = ((! is_zaet_4_destruct_bufchan_d[0]) || is_zaet_4_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) is_zaet_4_destruct_bufchan_d <= 1'd0;
    else
      if (is_zaet_4_destruct_r)
        is_zaet_4_destruct_bufchan_d <= is_zaet_4_destruct_d;
  MyDTInt_Bool_t is_zaet_4_destruct_bufchan_buf;
  assign is_zaet_4_destruct_bufchan_r = (! is_zaet_4_destruct_bufchan_buf[0]);
  assign is_zaet_4_1_argbuf_d = (is_zaet_4_destruct_bufchan_buf[0] ? is_zaet_4_destruct_bufchan_buf :
                                 is_zaet_4_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) is_zaet_4_destruct_bufchan_buf <= 1'd0;
    else
      if ((is_zaet_4_1_argbuf_r && is_zaet_4_destruct_bufchan_buf[0]))
        is_zaet_4_destruct_bufchan_buf <= 1'd0;
      else if (((! is_zaet_4_1_argbuf_r) && (! is_zaet_4_destruct_bufchan_buf[0])))
        is_zaet_4_destruct_bufchan_buf <= is_zaet_4_destruct_bufchan_d;
  
  /* buf (Ty MyDTInt_Bool) : (is_zafl_2_2,MyDTInt_Bool) > (is_zafl_2_2_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t is_zafl_2_2_bufchan_d;
  logic is_zafl_2_2_bufchan_r;
  assign is_zafl_2_2_r = ((! is_zafl_2_2_bufchan_d[0]) || is_zafl_2_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) is_zafl_2_2_bufchan_d <= 1'd0;
    else if (is_zafl_2_2_r) is_zafl_2_2_bufchan_d <= is_zafl_2_2_d;
  MyDTInt_Bool_t is_zafl_2_2_bufchan_buf;
  assign is_zafl_2_2_bufchan_r = (! is_zafl_2_2_bufchan_buf[0]);
  assign is_zafl_2_2_argbuf_d = (is_zafl_2_2_bufchan_buf[0] ? is_zafl_2_2_bufchan_buf :
                                 is_zafl_2_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) is_zafl_2_2_bufchan_buf <= 1'd0;
    else
      if ((is_zafl_2_2_argbuf_r && is_zafl_2_2_bufchan_buf[0]))
        is_zafl_2_2_bufchan_buf <= 1'd0;
      else if (((! is_zafl_2_2_argbuf_r) && (! is_zafl_2_2_bufchan_buf[0])))
        is_zafl_2_2_bufchan_buf <= is_zafl_2_2_bufchan_d;
  
  /* fork (Ty MyDTInt_Bool) : (is_zafl_2_destruct,MyDTInt_Bool) > [(is_zafl_2_1,MyDTInt_Bool),
                                                              (is_zafl_2_2,MyDTInt_Bool)] */
  logic [1:0] is_zafl_2_destruct_emitted;
  logic [1:0] is_zafl_2_destruct_done;
  assign is_zafl_2_1_d = (is_zafl_2_destruct_d[0] && (! is_zafl_2_destruct_emitted[0]));
  assign is_zafl_2_2_d = (is_zafl_2_destruct_d[0] && (! is_zafl_2_destruct_emitted[1]));
  assign is_zafl_2_destruct_done = (is_zafl_2_destruct_emitted | ({is_zafl_2_2_d[0],
                                                                   is_zafl_2_1_d[0]} & {is_zafl_2_2_r,
                                                                                        is_zafl_2_1_r}));
  assign is_zafl_2_destruct_r = (& is_zafl_2_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) is_zafl_2_destruct_emitted <= 2'd0;
    else
      is_zafl_2_destruct_emitted <= (is_zafl_2_destruct_r ? 2'd0 :
                                     is_zafl_2_destruct_done);
  
  /* buf (Ty MyDTInt_Bool) : (is_zafl_3_2,MyDTInt_Bool) > (is_zafl_3_2_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t is_zafl_3_2_bufchan_d;
  logic is_zafl_3_2_bufchan_r;
  assign is_zafl_3_2_r = ((! is_zafl_3_2_bufchan_d[0]) || is_zafl_3_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) is_zafl_3_2_bufchan_d <= 1'd0;
    else if (is_zafl_3_2_r) is_zafl_3_2_bufchan_d <= is_zafl_3_2_d;
  MyDTInt_Bool_t is_zafl_3_2_bufchan_buf;
  assign is_zafl_3_2_bufchan_r = (! is_zafl_3_2_bufchan_buf[0]);
  assign is_zafl_3_2_argbuf_d = (is_zafl_3_2_bufchan_buf[0] ? is_zafl_3_2_bufchan_buf :
                                 is_zafl_3_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) is_zafl_3_2_bufchan_buf <= 1'd0;
    else
      if ((is_zafl_3_2_argbuf_r && is_zafl_3_2_bufchan_buf[0]))
        is_zafl_3_2_bufchan_buf <= 1'd0;
      else if (((! is_zafl_3_2_argbuf_r) && (! is_zafl_3_2_bufchan_buf[0])))
        is_zafl_3_2_bufchan_buf <= is_zafl_3_2_bufchan_d;
  
  /* fork (Ty MyDTInt_Bool) : (is_zafl_3_destruct,MyDTInt_Bool) > [(is_zafl_3_1,MyDTInt_Bool),
                                                              (is_zafl_3_2,MyDTInt_Bool)] */
  logic [1:0] is_zafl_3_destruct_emitted;
  logic [1:0] is_zafl_3_destruct_done;
  assign is_zafl_3_1_d = (is_zafl_3_destruct_d[0] && (! is_zafl_3_destruct_emitted[0]));
  assign is_zafl_3_2_d = (is_zafl_3_destruct_d[0] && (! is_zafl_3_destruct_emitted[1]));
  assign is_zafl_3_destruct_done = (is_zafl_3_destruct_emitted | ({is_zafl_3_2_d[0],
                                                                   is_zafl_3_1_d[0]} & {is_zafl_3_2_r,
                                                                                        is_zafl_3_1_r}));
  assign is_zafl_3_destruct_r = (& is_zafl_3_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) is_zafl_3_destruct_emitted <= 2'd0;
    else
      is_zafl_3_destruct_emitted <= (is_zafl_3_destruct_r ? 2'd0 :
                                     is_zafl_3_destruct_done);
  
  /* buf (Ty MyDTInt_Bool) : (is_zafl_4_destruct,MyDTInt_Bool) > (is_zafl_4_1_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t is_zafl_4_destruct_bufchan_d;
  logic is_zafl_4_destruct_bufchan_r;
  assign is_zafl_4_destruct_r = ((! is_zafl_4_destruct_bufchan_d[0]) || is_zafl_4_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) is_zafl_4_destruct_bufchan_d <= 1'd0;
    else
      if (is_zafl_4_destruct_r)
        is_zafl_4_destruct_bufchan_d <= is_zafl_4_destruct_d;
  MyDTInt_Bool_t is_zafl_4_destruct_bufchan_buf;
  assign is_zafl_4_destruct_bufchan_r = (! is_zafl_4_destruct_bufchan_buf[0]);
  assign is_zafl_4_1_argbuf_d = (is_zafl_4_destruct_bufchan_buf[0] ? is_zafl_4_destruct_bufchan_buf :
                                 is_zafl_4_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) is_zafl_4_destruct_bufchan_buf <= 1'd0;
    else
      if ((is_zafl_4_1_argbuf_r && is_zafl_4_destruct_bufchan_buf[0]))
        is_zafl_4_destruct_bufchan_buf <= 1'd0;
      else if (((! is_zafl_4_1_argbuf_r) && (! is_zafl_4_destruct_bufchan_buf[0])))
        is_zafl_4_destruct_bufchan_buf <= is_zafl_4_destruct_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty MyDTInt_Int_Int) : (lizzieLet17_10,QTree_Int) (op_addaeu_goMux_mux,MyDTInt_Int_Int) > [(lizzieLet17_10QNone_Int,MyDTInt_Int_Int),
                                                                                                 (lizzieLet17_10QVal_Int,MyDTInt_Int_Int),
                                                                                                 (lizzieLet17_10QNode_Int,MyDTInt_Int_Int),
                                                                                                 (_224,MyDTInt_Int_Int)] */
  logic [3:0] op_addaeu_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet17_10_d[0] && op_addaeu_goMux_mux_d[0]))
      unique case (lizzieLet17_10_d[2:1])
        2'd0: op_addaeu_goMux_mux_onehotd = 4'd1;
        2'd1: op_addaeu_goMux_mux_onehotd = 4'd2;
        2'd2: op_addaeu_goMux_mux_onehotd = 4'd4;
        2'd3: op_addaeu_goMux_mux_onehotd = 4'd8;
        default: op_addaeu_goMux_mux_onehotd = 4'd0;
      endcase
    else op_addaeu_goMux_mux_onehotd = 4'd0;
  assign lizzieLet17_10QNone_Int_d = op_addaeu_goMux_mux_onehotd[0];
  assign lizzieLet17_10QVal_Int_d = op_addaeu_goMux_mux_onehotd[1];
  assign lizzieLet17_10QNode_Int_d = op_addaeu_goMux_mux_onehotd[2];
  assign _224_d = op_addaeu_goMux_mux_onehotd[3];
  assign op_addaeu_goMux_mux_r = (| (op_addaeu_goMux_mux_onehotd & {_224_r,
                                                                    lizzieLet17_10QNode_Int_r,
                                                                    lizzieLet17_10QVal_Int_r,
                                                                    lizzieLet17_10QNone_Int_r}));
  assign lizzieLet17_10_r = op_addaeu_goMux_mux_r;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_CTf_f_Int) : (lizzieLet17_11,QTree_Int) (sc_0_2_goMux_mux,Pointer_CTf_f_Int) > [(lizzieLet17_11QNone_Int,Pointer_CTf_f_Int),
                                                                                                  (lizzieLet17_11QVal_Int,Pointer_CTf_f_Int),
                                                                                                  (lizzieLet17_11QNode_Int,Pointer_CTf_f_Int),
                                                                                                  (lizzieLet17_11QError_Int,Pointer_CTf_f_Int)] */
  logic [3:0] sc_0_2_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet17_11_d[0] && sc_0_2_goMux_mux_d[0]))
      unique case (lizzieLet17_11_d[2:1])
        2'd0: sc_0_2_goMux_mux_onehotd = 4'd1;
        2'd1: sc_0_2_goMux_mux_onehotd = 4'd2;
        2'd2: sc_0_2_goMux_mux_onehotd = 4'd4;
        2'd3: sc_0_2_goMux_mux_onehotd = 4'd8;
        default: sc_0_2_goMux_mux_onehotd = 4'd0;
      endcase
    else sc_0_2_goMux_mux_onehotd = 4'd0;
  assign lizzieLet17_11QNone_Int_d = {sc_0_2_goMux_mux_d[16:1],
                                      sc_0_2_goMux_mux_onehotd[0]};
  assign lizzieLet17_11QVal_Int_d = {sc_0_2_goMux_mux_d[16:1],
                                     sc_0_2_goMux_mux_onehotd[1]};
  assign lizzieLet17_11QNode_Int_d = {sc_0_2_goMux_mux_d[16:1],
                                      sc_0_2_goMux_mux_onehotd[2]};
  assign lizzieLet17_11QError_Int_d = {sc_0_2_goMux_mux_d[16:1],
                                       sc_0_2_goMux_mux_onehotd[3]};
  assign sc_0_2_goMux_mux_r = (| (sc_0_2_goMux_mux_onehotd & {lizzieLet17_11QError_Int_r,
                                                              lizzieLet17_11QNode_Int_r,
                                                              lizzieLet17_11QVal_Int_r,
                                                              lizzieLet17_11QNone_Int_r}));
  assign lizzieLet17_11_r = sc_0_2_goMux_mux_r;
  
  /* buf (Ty Pointer_CTf_f_Int) : (lizzieLet17_11QError_Int,Pointer_CTf_f_Int) > (lizzieLet17_11QError_Int_1_argbuf,Pointer_CTf_f_Int) */
  Pointer_CTf_f_Int_t lizzieLet17_11QError_Int_bufchan_d;
  logic lizzieLet17_11QError_Int_bufchan_r;
  assign lizzieLet17_11QError_Int_r = ((! lizzieLet17_11QError_Int_bufchan_d[0]) || lizzieLet17_11QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_11QError_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet17_11QError_Int_r)
        lizzieLet17_11QError_Int_bufchan_d <= lizzieLet17_11QError_Int_d;
  Pointer_CTf_f_Int_t lizzieLet17_11QError_Int_bufchan_buf;
  assign lizzieLet17_11QError_Int_bufchan_r = (! lizzieLet17_11QError_Int_bufchan_buf[0]);
  assign lizzieLet17_11QError_Int_1_argbuf_d = (lizzieLet17_11QError_Int_bufchan_buf[0] ? lizzieLet17_11QError_Int_bufchan_buf :
                                                lizzieLet17_11QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_11QError_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet17_11QError_Int_1_argbuf_r && lizzieLet17_11QError_Int_bufchan_buf[0]))
        lizzieLet17_11QError_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet17_11QError_Int_1_argbuf_r) && (! lizzieLet17_11QError_Int_bufchan_buf[0])))
        lizzieLet17_11QError_Int_bufchan_buf <= lizzieLet17_11QError_Int_bufchan_d;
  
  /* destruct (Ty QTree_Int,
          Dcon QNode_Int) : (lizzieLet17_1QNode_Int,QTree_Int) > [(q1af0_destruct,Pointer_QTree_Int),
                                                                  (q2af1_destruct,Pointer_QTree_Int),
                                                                  (q3af2_destruct,Pointer_QTree_Int),
                                                                  (q4af3_destruct,Pointer_QTree_Int)] */
  logic [3:0] lizzieLet17_1QNode_Int_emitted;
  logic [3:0] lizzieLet17_1QNode_Int_done;
  assign q1af0_destruct_d = {lizzieLet17_1QNode_Int_d[18:3],
                             (lizzieLet17_1QNode_Int_d[0] && (! lizzieLet17_1QNode_Int_emitted[0]))};
  assign q2af1_destruct_d = {lizzieLet17_1QNode_Int_d[34:19],
                             (lizzieLet17_1QNode_Int_d[0] && (! lizzieLet17_1QNode_Int_emitted[1]))};
  assign q3af2_destruct_d = {lizzieLet17_1QNode_Int_d[50:35],
                             (lizzieLet17_1QNode_Int_d[0] && (! lizzieLet17_1QNode_Int_emitted[2]))};
  assign q4af3_destruct_d = {lizzieLet17_1QNode_Int_d[66:51],
                             (lizzieLet17_1QNode_Int_d[0] && (! lizzieLet17_1QNode_Int_emitted[3]))};
  assign lizzieLet17_1QNode_Int_done = (lizzieLet17_1QNode_Int_emitted | ({q4af3_destruct_d[0],
                                                                           q3af2_destruct_d[0],
                                                                           q2af1_destruct_d[0],
                                                                           q1af0_destruct_d[0]} & {q4af3_destruct_r,
                                                                                                   q3af2_destruct_r,
                                                                                                   q2af1_destruct_r,
                                                                                                   q1af0_destruct_r}));
  assign lizzieLet17_1QNode_Int_r = (& lizzieLet17_1QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet17_1QNode_Int_emitted <= 4'd0;
    else
      lizzieLet17_1QNode_Int_emitted <= (lizzieLet17_1QNode_Int_r ? 4'd0 :
                                         lizzieLet17_1QNode_Int_done);
  
  /* destruct (Ty QTree_Int,
          Dcon QVal_Int) : (lizzieLet17_1QVal_Int,QTree_Int) > [(v1aeK_destruct,Int)] */
  assign v1aeK_destruct_d = {lizzieLet17_1QVal_Int_d[34:3],
                             lizzieLet17_1QVal_Int_d[0]};
  assign lizzieLet17_1QVal_Int_r = v1aeK_destruct_r;
  
  /* demux (Ty QTree_Int,
       Ty QTree_Int) : (lizzieLet17_2,QTree_Int) (lizzieLet17_1,QTree_Int) > [(_223,QTree_Int),
                                                                              (lizzieLet17_1QVal_Int,QTree_Int),
                                                                              (lizzieLet17_1QNode_Int,QTree_Int),
                                                                              (_222,QTree_Int)] */
  logic [3:0] lizzieLet17_1_onehotd;
  always_comb
    if ((lizzieLet17_2_d[0] && lizzieLet17_1_d[0]))
      unique case (lizzieLet17_2_d[2:1])
        2'd0: lizzieLet17_1_onehotd = 4'd1;
        2'd1: lizzieLet17_1_onehotd = 4'd2;
        2'd2: lizzieLet17_1_onehotd = 4'd4;
        2'd3: lizzieLet17_1_onehotd = 4'd8;
        default: lizzieLet17_1_onehotd = 4'd0;
      endcase
    else lizzieLet17_1_onehotd = 4'd0;
  assign _223_d = {lizzieLet17_1_d[66:1], lizzieLet17_1_onehotd[0]};
  assign lizzieLet17_1QVal_Int_d = {lizzieLet17_1_d[66:1],
                                    lizzieLet17_1_onehotd[1]};
  assign lizzieLet17_1QNode_Int_d = {lizzieLet17_1_d[66:1],
                                     lizzieLet17_1_onehotd[2]};
  assign _222_d = {lizzieLet17_1_d[66:1], lizzieLet17_1_onehotd[3]};
  assign lizzieLet17_1_r = (| (lizzieLet17_1_onehotd & {_222_r,
                                                        lizzieLet17_1QNode_Int_r,
                                                        lizzieLet17_1QVal_Int_r,
                                                        _223_r}));
  assign lizzieLet17_2_r = lizzieLet17_1_r;
  
  /* demux (Ty QTree_Int,
       Ty Go) : (lizzieLet17_3,QTree_Int) (go_10_goMux_data,Go) > [(lizzieLet17_3QNone_Int,Go),
                                                                   (lizzieLet17_3QVal_Int,Go),
                                                                   (lizzieLet17_3QNode_Int,Go),
                                                                   (lizzieLet17_3QError_Int,Go)] */
  logic [3:0] go_10_goMux_data_onehotd;
  always_comb
    if ((lizzieLet17_3_d[0] && go_10_goMux_data_d[0]))
      unique case (lizzieLet17_3_d[2:1])
        2'd0: go_10_goMux_data_onehotd = 4'd1;
        2'd1: go_10_goMux_data_onehotd = 4'd2;
        2'd2: go_10_goMux_data_onehotd = 4'd4;
        2'd3: go_10_goMux_data_onehotd = 4'd8;
        default: go_10_goMux_data_onehotd = 4'd0;
      endcase
    else go_10_goMux_data_onehotd = 4'd0;
  assign lizzieLet17_3QNone_Int_d = go_10_goMux_data_onehotd[0];
  assign lizzieLet17_3QVal_Int_d = go_10_goMux_data_onehotd[1];
  assign lizzieLet17_3QNode_Int_d = go_10_goMux_data_onehotd[2];
  assign lizzieLet17_3QError_Int_d = go_10_goMux_data_onehotd[3];
  assign go_10_goMux_data_r = (| (go_10_goMux_data_onehotd & {lizzieLet17_3QError_Int_r,
                                                              lizzieLet17_3QNode_Int_r,
                                                              lizzieLet17_3QVal_Int_r,
                                                              lizzieLet17_3QNone_Int_r}));
  assign lizzieLet17_3_r = go_10_goMux_data_r;
  
  /* fork (Ty Go) : (lizzieLet17_3QError_Int,Go) > [(lizzieLet17_3QError_Int_1,Go),
                                               (lizzieLet17_3QError_Int_2,Go)] */
  logic [1:0] lizzieLet17_3QError_Int_emitted;
  logic [1:0] lizzieLet17_3QError_Int_done;
  assign lizzieLet17_3QError_Int_1_d = (lizzieLet17_3QError_Int_d[0] && (! lizzieLet17_3QError_Int_emitted[0]));
  assign lizzieLet17_3QError_Int_2_d = (lizzieLet17_3QError_Int_d[0] && (! lizzieLet17_3QError_Int_emitted[1]));
  assign lizzieLet17_3QError_Int_done = (lizzieLet17_3QError_Int_emitted | ({lizzieLet17_3QError_Int_2_d[0],
                                                                             lizzieLet17_3QError_Int_1_d[0]} & {lizzieLet17_3QError_Int_2_r,
                                                                                                                lizzieLet17_3QError_Int_1_r}));
  assign lizzieLet17_3QError_Int_r = (& lizzieLet17_3QError_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet17_3QError_Int_emitted <= 2'd0;
    else
      lizzieLet17_3QError_Int_emitted <= (lizzieLet17_3QError_Int_r ? 2'd0 :
                                          lizzieLet17_3QError_Int_done);
  
  /* dcon (Ty QTree_Int,
      Dcon QError_Int) : [(lizzieLet17_3QError_Int_1,Go)] > (lizzieLet17_3QError_Int_1QError_Int,QTree_Int) */
  assign lizzieLet17_3QError_Int_1QError_Int_d = QError_Int_dc((& {lizzieLet17_3QError_Int_1_d[0]}), lizzieLet17_3QError_Int_1_d);
  assign {lizzieLet17_3QError_Int_1_r} = {1 {(lizzieLet17_3QError_Int_1QError_Int_r && lizzieLet17_3QError_Int_1QError_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (lizzieLet17_3QError_Int_1QError_Int,QTree_Int) > (lizzieLet55_1_argbuf,QTree_Int) */
  QTree_Int_t lizzieLet17_3QError_Int_1QError_Int_bufchan_d;
  logic lizzieLet17_3QError_Int_1QError_Int_bufchan_r;
  assign lizzieLet17_3QError_Int_1QError_Int_r = ((! lizzieLet17_3QError_Int_1QError_Int_bufchan_d[0]) || lizzieLet17_3QError_Int_1QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_3QError_Int_1QError_Int_bufchan_d <= {66'd0, 1'd0};
    else
      if (lizzieLet17_3QError_Int_1QError_Int_r)
        lizzieLet17_3QError_Int_1QError_Int_bufchan_d <= lizzieLet17_3QError_Int_1QError_Int_d;
  QTree_Int_t lizzieLet17_3QError_Int_1QError_Int_bufchan_buf;
  assign lizzieLet17_3QError_Int_1QError_Int_bufchan_r = (! lizzieLet17_3QError_Int_1QError_Int_bufchan_buf[0]);
  assign lizzieLet55_1_argbuf_d = (lizzieLet17_3QError_Int_1QError_Int_bufchan_buf[0] ? lizzieLet17_3QError_Int_1QError_Int_bufchan_buf :
                                   lizzieLet17_3QError_Int_1QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_3QError_Int_1QError_Int_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((lizzieLet55_1_argbuf_r && lizzieLet17_3QError_Int_1QError_Int_bufchan_buf[0]))
        lizzieLet17_3QError_Int_1QError_Int_bufchan_buf <= {66'd0, 1'd0};
      else if (((! lizzieLet55_1_argbuf_r) && (! lizzieLet17_3QError_Int_1QError_Int_bufchan_buf[0])))
        lizzieLet17_3QError_Int_1QError_Int_bufchan_buf <= lizzieLet17_3QError_Int_1QError_Int_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet17_3QError_Int_2,Go) > (lizzieLet17_3QError_Int_2_argbuf,Go) */
  Go_t lizzieLet17_3QError_Int_2_bufchan_d;
  logic lizzieLet17_3QError_Int_2_bufchan_r;
  assign lizzieLet17_3QError_Int_2_r = ((! lizzieLet17_3QError_Int_2_bufchan_d[0]) || lizzieLet17_3QError_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet17_3QError_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet17_3QError_Int_2_r)
        lizzieLet17_3QError_Int_2_bufchan_d <= lizzieLet17_3QError_Int_2_d;
  Go_t lizzieLet17_3QError_Int_2_bufchan_buf;
  assign lizzieLet17_3QError_Int_2_bufchan_r = (! lizzieLet17_3QError_Int_2_bufchan_buf[0]);
  assign lizzieLet17_3QError_Int_2_argbuf_d = (lizzieLet17_3QError_Int_2_bufchan_buf[0] ? lizzieLet17_3QError_Int_2_bufchan_buf :
                                               lizzieLet17_3QError_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet17_3QError_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet17_3QError_Int_2_argbuf_r && lizzieLet17_3QError_Int_2_bufchan_buf[0]))
        lizzieLet17_3QError_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet17_3QError_Int_2_argbuf_r) && (! lizzieLet17_3QError_Int_2_bufchan_buf[0])))
        lizzieLet17_3QError_Int_2_bufchan_buf <= lizzieLet17_3QError_Int_2_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty MyDTInt_Bool) : (lizzieLet17_4,QTree_Int) (is_zaet_goMux_mux,MyDTInt_Bool) > [(lizzieLet17_4QNone_Int,MyDTInt_Bool),
                                                                                        (lizzieLet17_4QVal_Int,MyDTInt_Bool),
                                                                                        (lizzieLet17_4QNode_Int,MyDTInt_Bool),
                                                                                        (_221,MyDTInt_Bool)] */
  logic [3:0] is_zaet_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet17_4_d[0] && is_zaet_goMux_mux_d[0]))
      unique case (lizzieLet17_4_d[2:1])
        2'd0: is_zaet_goMux_mux_onehotd = 4'd1;
        2'd1: is_zaet_goMux_mux_onehotd = 4'd2;
        2'd2: is_zaet_goMux_mux_onehotd = 4'd4;
        2'd3: is_zaet_goMux_mux_onehotd = 4'd8;
        default: is_zaet_goMux_mux_onehotd = 4'd0;
      endcase
    else is_zaet_goMux_mux_onehotd = 4'd0;
  assign lizzieLet17_4QNone_Int_d = is_zaet_goMux_mux_onehotd[0];
  assign lizzieLet17_4QVal_Int_d = is_zaet_goMux_mux_onehotd[1];
  assign lizzieLet17_4QNode_Int_d = is_zaet_goMux_mux_onehotd[2];
  assign _221_d = is_zaet_goMux_mux_onehotd[3];
  assign is_zaet_goMux_mux_r = (| (is_zaet_goMux_mux_onehotd & {_221_r,
                                                                lizzieLet17_4QNode_Int_r,
                                                                lizzieLet17_4QVal_Int_r,
                                                                lizzieLet17_4QNone_Int_r}));
  assign lizzieLet17_4_r = is_zaet_goMux_mux_r;
  
  /* demux (Ty QTree_Int,
       Ty QTree_Int) : (lizzieLet17_5,QTree_Int) (readPointer_QTree_Intm2aer_1_argbuf_rwb,QTree_Int) > [(lizzieLet17_5QNone_Int,QTree_Int),
                                                                                                        (lizzieLet17_5QVal_Int,QTree_Int),
                                                                                                        (lizzieLet17_5QNode_Int,QTree_Int),
                                                                                                        (_220,QTree_Int)] */
  logic [3:0] readPointer_QTree_Intm2aer_1_argbuf_rwb_onehotd;
  always_comb
    if ((lizzieLet17_5_d[0] && readPointer_QTree_Intm2aer_1_argbuf_rwb_d[0]))
      unique case (lizzieLet17_5_d[2:1])
        2'd0: readPointer_QTree_Intm2aer_1_argbuf_rwb_onehotd = 4'd1;
        2'd1: readPointer_QTree_Intm2aer_1_argbuf_rwb_onehotd = 4'd2;
        2'd2: readPointer_QTree_Intm2aer_1_argbuf_rwb_onehotd = 4'd4;
        2'd3: readPointer_QTree_Intm2aer_1_argbuf_rwb_onehotd = 4'd8;
        default: readPointer_QTree_Intm2aer_1_argbuf_rwb_onehotd = 4'd0;
      endcase
    else readPointer_QTree_Intm2aer_1_argbuf_rwb_onehotd = 4'd0;
  assign lizzieLet17_5QNone_Int_d = {readPointer_QTree_Intm2aer_1_argbuf_rwb_d[66:1],
                                     readPointer_QTree_Intm2aer_1_argbuf_rwb_onehotd[0]};
  assign lizzieLet17_5QVal_Int_d = {readPointer_QTree_Intm2aer_1_argbuf_rwb_d[66:1],
                                    readPointer_QTree_Intm2aer_1_argbuf_rwb_onehotd[1]};
  assign lizzieLet17_5QNode_Int_d = {readPointer_QTree_Intm2aer_1_argbuf_rwb_d[66:1],
                                     readPointer_QTree_Intm2aer_1_argbuf_rwb_onehotd[2]};
  assign _220_d = {readPointer_QTree_Intm2aer_1_argbuf_rwb_d[66:1],
                   readPointer_QTree_Intm2aer_1_argbuf_rwb_onehotd[3]};
  assign readPointer_QTree_Intm2aer_1_argbuf_rwb_r = (| (readPointer_QTree_Intm2aer_1_argbuf_rwb_onehotd & {_220_r,
                                                                                                            lizzieLet17_5QNode_Int_r,
                                                                                                            lizzieLet17_5QVal_Int_r,
                                                                                                            lizzieLet17_5QNone_Int_r}));
  assign lizzieLet17_5_r = readPointer_QTree_Intm2aer_1_argbuf_rwb_r;
  
  /* fork (Ty QTree_Int) : (lizzieLet17_5QNode_Int,QTree_Int) > [(lizzieLet17_5QNode_Int_1,QTree_Int),
                                                            (lizzieLet17_5QNode_Int_2,QTree_Int),
                                                            (lizzieLet17_5QNode_Int_3,QTree_Int),
                                                            (lizzieLet17_5QNode_Int_4,QTree_Int),
                                                            (lizzieLet17_5QNode_Int_5,QTree_Int),
                                                            (lizzieLet17_5QNode_Int_6,QTree_Int),
                                                            (lizzieLet17_5QNode_Int_7,QTree_Int),
                                                            (lizzieLet17_5QNode_Int_8,QTree_Int),
                                                            (lizzieLet17_5QNode_Int_9,QTree_Int),
                                                            (lizzieLet17_5QNode_Int_10,QTree_Int),
                                                            (lizzieLet17_5QNode_Int_11,QTree_Int),
                                                            (lizzieLet17_5QNode_Int_12,QTree_Int)] */
  logic [11:0] lizzieLet17_5QNode_Int_emitted;
  logic [11:0] lizzieLet17_5QNode_Int_done;
  assign lizzieLet17_5QNode_Int_1_d = {lizzieLet17_5QNode_Int_d[66:1],
                                       (lizzieLet17_5QNode_Int_d[0] && (! lizzieLet17_5QNode_Int_emitted[0]))};
  assign lizzieLet17_5QNode_Int_2_d = {lizzieLet17_5QNode_Int_d[66:1],
                                       (lizzieLet17_5QNode_Int_d[0] && (! lizzieLet17_5QNode_Int_emitted[1]))};
  assign lizzieLet17_5QNode_Int_3_d = {lizzieLet17_5QNode_Int_d[66:1],
                                       (lizzieLet17_5QNode_Int_d[0] && (! lizzieLet17_5QNode_Int_emitted[2]))};
  assign lizzieLet17_5QNode_Int_4_d = {lizzieLet17_5QNode_Int_d[66:1],
                                       (lizzieLet17_5QNode_Int_d[0] && (! lizzieLet17_5QNode_Int_emitted[3]))};
  assign lizzieLet17_5QNode_Int_5_d = {lizzieLet17_5QNode_Int_d[66:1],
                                       (lizzieLet17_5QNode_Int_d[0] && (! lizzieLet17_5QNode_Int_emitted[4]))};
  assign lizzieLet17_5QNode_Int_6_d = {lizzieLet17_5QNode_Int_d[66:1],
                                       (lizzieLet17_5QNode_Int_d[0] && (! lizzieLet17_5QNode_Int_emitted[5]))};
  assign lizzieLet17_5QNode_Int_7_d = {lizzieLet17_5QNode_Int_d[66:1],
                                       (lizzieLet17_5QNode_Int_d[0] && (! lizzieLet17_5QNode_Int_emitted[6]))};
  assign lizzieLet17_5QNode_Int_8_d = {lizzieLet17_5QNode_Int_d[66:1],
                                       (lizzieLet17_5QNode_Int_d[0] && (! lizzieLet17_5QNode_Int_emitted[7]))};
  assign lizzieLet17_5QNode_Int_9_d = {lizzieLet17_5QNode_Int_d[66:1],
                                       (lizzieLet17_5QNode_Int_d[0] && (! lizzieLet17_5QNode_Int_emitted[8]))};
  assign lizzieLet17_5QNode_Int_10_d = {lizzieLet17_5QNode_Int_d[66:1],
                                        (lizzieLet17_5QNode_Int_d[0] && (! lizzieLet17_5QNode_Int_emitted[9]))};
  assign lizzieLet17_5QNode_Int_11_d = {lizzieLet17_5QNode_Int_d[66:1],
                                        (lizzieLet17_5QNode_Int_d[0] && (! lizzieLet17_5QNode_Int_emitted[10]))};
  assign lizzieLet17_5QNode_Int_12_d = {lizzieLet17_5QNode_Int_d[66:1],
                                        (lizzieLet17_5QNode_Int_d[0] && (! lizzieLet17_5QNode_Int_emitted[11]))};
  assign lizzieLet17_5QNode_Int_done = (lizzieLet17_5QNode_Int_emitted | ({lizzieLet17_5QNode_Int_12_d[0],
                                                                           lizzieLet17_5QNode_Int_11_d[0],
                                                                           lizzieLet17_5QNode_Int_10_d[0],
                                                                           lizzieLet17_5QNode_Int_9_d[0],
                                                                           lizzieLet17_5QNode_Int_8_d[0],
                                                                           lizzieLet17_5QNode_Int_7_d[0],
                                                                           lizzieLet17_5QNode_Int_6_d[0],
                                                                           lizzieLet17_5QNode_Int_5_d[0],
                                                                           lizzieLet17_5QNode_Int_4_d[0],
                                                                           lizzieLet17_5QNode_Int_3_d[0],
                                                                           lizzieLet17_5QNode_Int_2_d[0],
                                                                           lizzieLet17_5QNode_Int_1_d[0]} & {lizzieLet17_5QNode_Int_12_r,
                                                                                                             lizzieLet17_5QNode_Int_11_r,
                                                                                                             lizzieLet17_5QNode_Int_10_r,
                                                                                                             lizzieLet17_5QNode_Int_9_r,
                                                                                                             lizzieLet17_5QNode_Int_8_r,
                                                                                                             lizzieLet17_5QNode_Int_7_r,
                                                                                                             lizzieLet17_5QNode_Int_6_r,
                                                                                                             lizzieLet17_5QNode_Int_5_r,
                                                                                                             lizzieLet17_5QNode_Int_4_r,
                                                                                                             lizzieLet17_5QNode_Int_3_r,
                                                                                                             lizzieLet17_5QNode_Int_2_r,
                                                                                                             lizzieLet17_5QNode_Int_1_r}));
  assign lizzieLet17_5QNode_Int_r = (& lizzieLet17_5QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet17_5QNode_Int_emitted <= 12'd0;
    else
      lizzieLet17_5QNode_Int_emitted <= (lizzieLet17_5QNode_Int_r ? 12'd0 :
                                         lizzieLet17_5QNode_Int_done);
  
  /* demux (Ty QTree_Int,
       Ty Pointer_QTree_Int) : (lizzieLet17_5QNode_Int_10,QTree_Int) (q2af1_destruct,Pointer_QTree_Int) > [(lizzieLet17_5QNode_Int_10QNone_Int,Pointer_QTree_Int),
                                                                                                           (_219,Pointer_QTree_Int),
                                                                                                           (lizzieLet17_5QNode_Int_10QNode_Int,Pointer_QTree_Int),
                                                                                                           (_218,Pointer_QTree_Int)] */
  logic [3:0] q2af1_destruct_onehotd;
  always_comb
    if ((lizzieLet17_5QNode_Int_10_d[0] && q2af1_destruct_d[0]))
      unique case (lizzieLet17_5QNode_Int_10_d[2:1])
        2'd0: q2af1_destruct_onehotd = 4'd1;
        2'd1: q2af1_destruct_onehotd = 4'd2;
        2'd2: q2af1_destruct_onehotd = 4'd4;
        2'd3: q2af1_destruct_onehotd = 4'd8;
        default: q2af1_destruct_onehotd = 4'd0;
      endcase
    else q2af1_destruct_onehotd = 4'd0;
  assign lizzieLet17_5QNode_Int_10QNone_Int_d = {q2af1_destruct_d[16:1],
                                                 q2af1_destruct_onehotd[0]};
  assign _219_d = {q2af1_destruct_d[16:1],
                   q2af1_destruct_onehotd[1]};
  assign lizzieLet17_5QNode_Int_10QNode_Int_d = {q2af1_destruct_d[16:1],
                                                 q2af1_destruct_onehotd[2]};
  assign _218_d = {q2af1_destruct_d[16:1],
                   q2af1_destruct_onehotd[3]};
  assign q2af1_destruct_r = (| (q2af1_destruct_onehotd & {_218_r,
                                                          lizzieLet17_5QNode_Int_10QNode_Int_r,
                                                          _219_r,
                                                          lizzieLet17_5QNode_Int_10QNone_Int_r}));
  assign lizzieLet17_5QNode_Int_10_r = q2af1_destruct_r;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_QTree_Int) : (lizzieLet17_5QNode_Int_11,QTree_Int) (q3af2_destruct,Pointer_QTree_Int) > [(lizzieLet17_5QNode_Int_11QNone_Int,Pointer_QTree_Int),
                                                                                                           (_217,Pointer_QTree_Int),
                                                                                                           (lizzieLet17_5QNode_Int_11QNode_Int,Pointer_QTree_Int),
                                                                                                           (_216,Pointer_QTree_Int)] */
  logic [3:0] q3af2_destruct_onehotd;
  always_comb
    if ((lizzieLet17_5QNode_Int_11_d[0] && q3af2_destruct_d[0]))
      unique case (lizzieLet17_5QNode_Int_11_d[2:1])
        2'd0: q3af2_destruct_onehotd = 4'd1;
        2'd1: q3af2_destruct_onehotd = 4'd2;
        2'd2: q3af2_destruct_onehotd = 4'd4;
        2'd3: q3af2_destruct_onehotd = 4'd8;
        default: q3af2_destruct_onehotd = 4'd0;
      endcase
    else q3af2_destruct_onehotd = 4'd0;
  assign lizzieLet17_5QNode_Int_11QNone_Int_d = {q3af2_destruct_d[16:1],
                                                 q3af2_destruct_onehotd[0]};
  assign _217_d = {q3af2_destruct_d[16:1],
                   q3af2_destruct_onehotd[1]};
  assign lizzieLet17_5QNode_Int_11QNode_Int_d = {q3af2_destruct_d[16:1],
                                                 q3af2_destruct_onehotd[2]};
  assign _216_d = {q3af2_destruct_d[16:1],
                   q3af2_destruct_onehotd[3]};
  assign q3af2_destruct_r = (| (q3af2_destruct_onehotd & {_216_r,
                                                          lizzieLet17_5QNode_Int_11QNode_Int_r,
                                                          _217_r,
                                                          lizzieLet17_5QNode_Int_11QNone_Int_r}));
  assign lizzieLet17_5QNode_Int_11_r = q3af2_destruct_r;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_QTree_Int) : (lizzieLet17_5QNode_Int_12,QTree_Int) (q4af3_destruct,Pointer_QTree_Int) > [(lizzieLet17_5QNode_Int_12QNone_Int,Pointer_QTree_Int),
                                                                                                           (_215,Pointer_QTree_Int),
                                                                                                           (lizzieLet17_5QNode_Int_12QNode_Int,Pointer_QTree_Int),
                                                                                                           (_214,Pointer_QTree_Int)] */
  logic [3:0] q4af3_destruct_onehotd;
  always_comb
    if ((lizzieLet17_5QNode_Int_12_d[0] && q4af3_destruct_d[0]))
      unique case (lizzieLet17_5QNode_Int_12_d[2:1])
        2'd0: q4af3_destruct_onehotd = 4'd1;
        2'd1: q4af3_destruct_onehotd = 4'd2;
        2'd2: q4af3_destruct_onehotd = 4'd4;
        2'd3: q4af3_destruct_onehotd = 4'd8;
        default: q4af3_destruct_onehotd = 4'd0;
      endcase
    else q4af3_destruct_onehotd = 4'd0;
  assign lizzieLet17_5QNode_Int_12QNone_Int_d = {q4af3_destruct_d[16:1],
                                                 q4af3_destruct_onehotd[0]};
  assign _215_d = {q4af3_destruct_d[16:1],
                   q4af3_destruct_onehotd[1]};
  assign lizzieLet17_5QNode_Int_12QNode_Int_d = {q4af3_destruct_d[16:1],
                                                 q4af3_destruct_onehotd[2]};
  assign _214_d = {q4af3_destruct_d[16:1],
                   q4af3_destruct_onehotd[3]};
  assign q4af3_destruct_r = (| (q4af3_destruct_onehotd & {_214_r,
                                                          lizzieLet17_5QNode_Int_12QNode_Int_r,
                                                          _215_r,
                                                          lizzieLet17_5QNode_Int_12QNone_Int_r}));
  assign lizzieLet17_5QNode_Int_12_r = q4af3_destruct_r;
  
  /* destruct (Ty QTree_Int,
          Dcon QNode_Int) : (lizzieLet17_5QNode_Int_1QNode_Int,QTree_Int) > [(t1afa_destruct,Pointer_QTree_Int),
                                                                             (t2afb_destruct,Pointer_QTree_Int),
                                                                             (t3afc_destruct,Pointer_QTree_Int),
                                                                             (t4afd_destruct,Pointer_QTree_Int)] */
  logic [3:0] lizzieLet17_5QNode_Int_1QNode_Int_emitted;
  logic [3:0] lizzieLet17_5QNode_Int_1QNode_Int_done;
  assign t1afa_destruct_d = {lizzieLet17_5QNode_Int_1QNode_Int_d[18:3],
                             (lizzieLet17_5QNode_Int_1QNode_Int_d[0] && (! lizzieLet17_5QNode_Int_1QNode_Int_emitted[0]))};
  assign t2afb_destruct_d = {lizzieLet17_5QNode_Int_1QNode_Int_d[34:19],
                             (lizzieLet17_5QNode_Int_1QNode_Int_d[0] && (! lizzieLet17_5QNode_Int_1QNode_Int_emitted[1]))};
  assign t3afc_destruct_d = {lizzieLet17_5QNode_Int_1QNode_Int_d[50:35],
                             (lizzieLet17_5QNode_Int_1QNode_Int_d[0] && (! lizzieLet17_5QNode_Int_1QNode_Int_emitted[2]))};
  assign t4afd_destruct_d = {lizzieLet17_5QNode_Int_1QNode_Int_d[66:51],
                             (lizzieLet17_5QNode_Int_1QNode_Int_d[0] && (! lizzieLet17_5QNode_Int_1QNode_Int_emitted[3]))};
  assign lizzieLet17_5QNode_Int_1QNode_Int_done = (lizzieLet17_5QNode_Int_1QNode_Int_emitted | ({t4afd_destruct_d[0],
                                                                                                 t3afc_destruct_d[0],
                                                                                                 t2afb_destruct_d[0],
                                                                                                 t1afa_destruct_d[0]} & {t4afd_destruct_r,
                                                                                                                         t3afc_destruct_r,
                                                                                                                         t2afb_destruct_r,
                                                                                                                         t1afa_destruct_r}));
  assign lizzieLet17_5QNode_Int_1QNode_Int_r = (& lizzieLet17_5QNode_Int_1QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_1QNode_Int_emitted <= 4'd0;
    else
      lizzieLet17_5QNode_Int_1QNode_Int_emitted <= (lizzieLet17_5QNode_Int_1QNode_Int_r ? 4'd0 :
                                                    lizzieLet17_5QNode_Int_1QNode_Int_done);
  
  /* demux (Ty QTree_Int,
       Ty QTree_Int) : (lizzieLet17_5QNode_Int_2,QTree_Int) (lizzieLet17_5QNode_Int_1,QTree_Int) > [(_213,QTree_Int),
                                                                                                    (_212,QTree_Int),
                                                                                                    (lizzieLet17_5QNode_Int_1QNode_Int,QTree_Int),
                                                                                                    (_211,QTree_Int)] */
  logic [3:0] lizzieLet17_5QNode_Int_1_onehotd;
  always_comb
    if ((lizzieLet17_5QNode_Int_2_d[0] && lizzieLet17_5QNode_Int_1_d[0]))
      unique case (lizzieLet17_5QNode_Int_2_d[2:1])
        2'd0: lizzieLet17_5QNode_Int_1_onehotd = 4'd1;
        2'd1: lizzieLet17_5QNode_Int_1_onehotd = 4'd2;
        2'd2: lizzieLet17_5QNode_Int_1_onehotd = 4'd4;
        2'd3: lizzieLet17_5QNode_Int_1_onehotd = 4'd8;
        default: lizzieLet17_5QNode_Int_1_onehotd = 4'd0;
      endcase
    else lizzieLet17_5QNode_Int_1_onehotd = 4'd0;
  assign _213_d = {lizzieLet17_5QNode_Int_1_d[66:1],
                   lizzieLet17_5QNode_Int_1_onehotd[0]};
  assign _212_d = {lizzieLet17_5QNode_Int_1_d[66:1],
                   lizzieLet17_5QNode_Int_1_onehotd[1]};
  assign lizzieLet17_5QNode_Int_1QNode_Int_d = {lizzieLet17_5QNode_Int_1_d[66:1],
                                                lizzieLet17_5QNode_Int_1_onehotd[2]};
  assign _211_d = {lizzieLet17_5QNode_Int_1_d[66:1],
                   lizzieLet17_5QNode_Int_1_onehotd[3]};
  assign lizzieLet17_5QNode_Int_1_r = (| (lizzieLet17_5QNode_Int_1_onehotd & {_211_r,
                                                                              lizzieLet17_5QNode_Int_1QNode_Int_r,
                                                                              _212_r,
                                                                              _213_r}));
  assign lizzieLet17_5QNode_Int_2_r = lizzieLet17_5QNode_Int_1_r;
  
  /* demux (Ty QTree_Int,
       Ty MyDTInt_Int_Int) : (lizzieLet17_5QNode_Int_3,QTree_Int) (lizzieLet17_10QNode_Int,MyDTInt_Int_Int) > [(lizzieLet17_5QNode_Int_3QNone_Int,MyDTInt_Int_Int),
                                                                                                               (_210,MyDTInt_Int_Int),
                                                                                                               (lizzieLet17_5QNode_Int_3QNode_Int,MyDTInt_Int_Int),
                                                                                                               (_209,MyDTInt_Int_Int)] */
  logic [3:0] lizzieLet17_10QNode_Int_onehotd;
  always_comb
    if ((lizzieLet17_5QNode_Int_3_d[0] && lizzieLet17_10QNode_Int_d[0]))
      unique case (lizzieLet17_5QNode_Int_3_d[2:1])
        2'd0: lizzieLet17_10QNode_Int_onehotd = 4'd1;
        2'd1: lizzieLet17_10QNode_Int_onehotd = 4'd2;
        2'd2: lizzieLet17_10QNode_Int_onehotd = 4'd4;
        2'd3: lizzieLet17_10QNode_Int_onehotd = 4'd8;
        default: lizzieLet17_10QNode_Int_onehotd = 4'd0;
      endcase
    else lizzieLet17_10QNode_Int_onehotd = 4'd0;
  assign lizzieLet17_5QNode_Int_3QNone_Int_d = lizzieLet17_10QNode_Int_onehotd[0];
  assign _210_d = lizzieLet17_10QNode_Int_onehotd[1];
  assign lizzieLet17_5QNode_Int_3QNode_Int_d = lizzieLet17_10QNode_Int_onehotd[2];
  assign _209_d = lizzieLet17_10QNode_Int_onehotd[3];
  assign lizzieLet17_10QNode_Int_r = (| (lizzieLet17_10QNode_Int_onehotd & {_209_r,
                                                                            lizzieLet17_5QNode_Int_3QNode_Int_r,
                                                                            _210_r,
                                                                            lizzieLet17_5QNode_Int_3QNone_Int_r}));
  assign lizzieLet17_5QNode_Int_3_r = lizzieLet17_10QNode_Int_r;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_CTf_f_Int) : (lizzieLet17_5QNode_Int_4,QTree_Int) (lizzieLet17_11QNode_Int,Pointer_CTf_f_Int) > [(lizzieLet17_5QNode_Int_4QNone_Int,Pointer_CTf_f_Int),
                                                                                                                   (lizzieLet17_5QNode_Int_4QVal_Int,Pointer_CTf_f_Int),
                                                                                                                   (lizzieLet17_5QNode_Int_4QNode_Int,Pointer_CTf_f_Int),
                                                                                                                   (lizzieLet17_5QNode_Int_4QError_Int,Pointer_CTf_f_Int)] */
  logic [3:0] lizzieLet17_11QNode_Int_onehotd;
  always_comb
    if ((lizzieLet17_5QNode_Int_4_d[0] && lizzieLet17_11QNode_Int_d[0]))
      unique case (lizzieLet17_5QNode_Int_4_d[2:1])
        2'd0: lizzieLet17_11QNode_Int_onehotd = 4'd1;
        2'd1: lizzieLet17_11QNode_Int_onehotd = 4'd2;
        2'd2: lizzieLet17_11QNode_Int_onehotd = 4'd4;
        2'd3: lizzieLet17_11QNode_Int_onehotd = 4'd8;
        default: lizzieLet17_11QNode_Int_onehotd = 4'd0;
      endcase
    else lizzieLet17_11QNode_Int_onehotd = 4'd0;
  assign lizzieLet17_5QNode_Int_4QNone_Int_d = {lizzieLet17_11QNode_Int_d[16:1],
                                                lizzieLet17_11QNode_Int_onehotd[0]};
  assign lizzieLet17_5QNode_Int_4QVal_Int_d = {lizzieLet17_11QNode_Int_d[16:1],
                                               lizzieLet17_11QNode_Int_onehotd[1]};
  assign lizzieLet17_5QNode_Int_4QNode_Int_d = {lizzieLet17_11QNode_Int_d[16:1],
                                                lizzieLet17_11QNode_Int_onehotd[2]};
  assign lizzieLet17_5QNode_Int_4QError_Int_d = {lizzieLet17_11QNode_Int_d[16:1],
                                                 lizzieLet17_11QNode_Int_onehotd[3]};
  assign lizzieLet17_11QNode_Int_r = (| (lizzieLet17_11QNode_Int_onehotd & {lizzieLet17_5QNode_Int_4QError_Int_r,
                                                                            lizzieLet17_5QNode_Int_4QNode_Int_r,
                                                                            lizzieLet17_5QNode_Int_4QVal_Int_r,
                                                                            lizzieLet17_5QNode_Int_4QNone_Int_r}));
  assign lizzieLet17_5QNode_Int_4_r = lizzieLet17_11QNode_Int_r;
  
  /* buf (Ty Pointer_CTf_f_Int) : (lizzieLet17_5QNode_Int_4QError_Int,Pointer_CTf_f_Int) > (lizzieLet17_5QNode_Int_4QError_Int_1_argbuf,Pointer_CTf_f_Int) */
  Pointer_CTf_f_Int_t lizzieLet17_5QNode_Int_4QError_Int_bufchan_d;
  logic lizzieLet17_5QNode_Int_4QError_Int_bufchan_r;
  assign lizzieLet17_5QNode_Int_4QError_Int_r = ((! lizzieLet17_5QNode_Int_4QError_Int_bufchan_d[0]) || lizzieLet17_5QNode_Int_4QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_4QError_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet17_5QNode_Int_4QError_Int_r)
        lizzieLet17_5QNode_Int_4QError_Int_bufchan_d <= lizzieLet17_5QNode_Int_4QError_Int_d;
  Pointer_CTf_f_Int_t lizzieLet17_5QNode_Int_4QError_Int_bufchan_buf;
  assign lizzieLet17_5QNode_Int_4QError_Int_bufchan_r = (! lizzieLet17_5QNode_Int_4QError_Int_bufchan_buf[0]);
  assign lizzieLet17_5QNode_Int_4QError_Int_1_argbuf_d = (lizzieLet17_5QNode_Int_4QError_Int_bufchan_buf[0] ? lizzieLet17_5QNode_Int_4QError_Int_bufchan_buf :
                                                          lizzieLet17_5QNode_Int_4QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_4QError_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet17_5QNode_Int_4QError_Int_1_argbuf_r && lizzieLet17_5QNode_Int_4QError_Int_bufchan_buf[0]))
        lizzieLet17_5QNode_Int_4QError_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet17_5QNode_Int_4QError_Int_1_argbuf_r) && (! lizzieLet17_5QNode_Int_4QError_Int_bufchan_buf[0])))
        lizzieLet17_5QNode_Int_4QError_Int_bufchan_buf <= lizzieLet17_5QNode_Int_4QError_Int_bufchan_d;
  
  /* buf (Ty Pointer_CTf_f_Int) : (lizzieLet17_5QNode_Int_4QVal_Int,Pointer_CTf_f_Int) > (lizzieLet17_5QNode_Int_4QVal_Int_1_argbuf,Pointer_CTf_f_Int) */
  Pointer_CTf_f_Int_t lizzieLet17_5QNode_Int_4QVal_Int_bufchan_d;
  logic lizzieLet17_5QNode_Int_4QVal_Int_bufchan_r;
  assign lizzieLet17_5QNode_Int_4QVal_Int_r = ((! lizzieLet17_5QNode_Int_4QVal_Int_bufchan_d[0]) || lizzieLet17_5QNode_Int_4QVal_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_4QVal_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet17_5QNode_Int_4QVal_Int_r)
        lizzieLet17_5QNode_Int_4QVal_Int_bufchan_d <= lizzieLet17_5QNode_Int_4QVal_Int_d;
  Pointer_CTf_f_Int_t lizzieLet17_5QNode_Int_4QVal_Int_bufchan_buf;
  assign lizzieLet17_5QNode_Int_4QVal_Int_bufchan_r = (! lizzieLet17_5QNode_Int_4QVal_Int_bufchan_buf[0]);
  assign lizzieLet17_5QNode_Int_4QVal_Int_1_argbuf_d = (lizzieLet17_5QNode_Int_4QVal_Int_bufchan_buf[0] ? lizzieLet17_5QNode_Int_4QVal_Int_bufchan_buf :
                                                        lizzieLet17_5QNode_Int_4QVal_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_4QVal_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet17_5QNode_Int_4QVal_Int_1_argbuf_r && lizzieLet17_5QNode_Int_4QVal_Int_bufchan_buf[0]))
        lizzieLet17_5QNode_Int_4QVal_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet17_5QNode_Int_4QVal_Int_1_argbuf_r) && (! lizzieLet17_5QNode_Int_4QVal_Int_bufchan_buf[0])))
        lizzieLet17_5QNode_Int_4QVal_Int_bufchan_buf <= lizzieLet17_5QNode_Int_4QVal_Int_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Go) : (lizzieLet17_5QNode_Int_5,QTree_Int) (lizzieLet17_3QNode_Int,Go) > [(lizzieLet17_5QNode_Int_5QNone_Int,Go),
                                                                                    (lizzieLet17_5QNode_Int_5QVal_Int,Go),
                                                                                    (lizzieLet17_5QNode_Int_5QNode_Int,Go),
                                                                                    (lizzieLet17_5QNode_Int_5QError_Int,Go)] */
  logic [3:0] lizzieLet17_3QNode_Int_onehotd;
  always_comb
    if ((lizzieLet17_5QNode_Int_5_d[0] && lizzieLet17_3QNode_Int_d[0]))
      unique case (lizzieLet17_5QNode_Int_5_d[2:1])
        2'd0: lizzieLet17_3QNode_Int_onehotd = 4'd1;
        2'd1: lizzieLet17_3QNode_Int_onehotd = 4'd2;
        2'd2: lizzieLet17_3QNode_Int_onehotd = 4'd4;
        2'd3: lizzieLet17_3QNode_Int_onehotd = 4'd8;
        default: lizzieLet17_3QNode_Int_onehotd = 4'd0;
      endcase
    else lizzieLet17_3QNode_Int_onehotd = 4'd0;
  assign lizzieLet17_5QNode_Int_5QNone_Int_d = lizzieLet17_3QNode_Int_onehotd[0];
  assign lizzieLet17_5QNode_Int_5QVal_Int_d = lizzieLet17_3QNode_Int_onehotd[1];
  assign lizzieLet17_5QNode_Int_5QNode_Int_d = lizzieLet17_3QNode_Int_onehotd[2];
  assign lizzieLet17_5QNode_Int_5QError_Int_d = lizzieLet17_3QNode_Int_onehotd[3];
  assign lizzieLet17_3QNode_Int_r = (| (lizzieLet17_3QNode_Int_onehotd & {lizzieLet17_5QNode_Int_5QError_Int_r,
                                                                          lizzieLet17_5QNode_Int_5QNode_Int_r,
                                                                          lizzieLet17_5QNode_Int_5QVal_Int_r,
                                                                          lizzieLet17_5QNode_Int_5QNone_Int_r}));
  assign lizzieLet17_5QNode_Int_5_r = lizzieLet17_3QNode_Int_r;
  
  /* fork (Ty Go) : (lizzieLet17_5QNode_Int_5QError_Int,Go) > [(lizzieLet17_5QNode_Int_5QError_Int_1,Go),
                                                          (lizzieLet17_5QNode_Int_5QError_Int_2,Go)] */
  logic [1:0] lizzieLet17_5QNode_Int_5QError_Int_emitted;
  logic [1:0] lizzieLet17_5QNode_Int_5QError_Int_done;
  assign lizzieLet17_5QNode_Int_5QError_Int_1_d = (lizzieLet17_5QNode_Int_5QError_Int_d[0] && (! lizzieLet17_5QNode_Int_5QError_Int_emitted[0]));
  assign lizzieLet17_5QNode_Int_5QError_Int_2_d = (lizzieLet17_5QNode_Int_5QError_Int_d[0] && (! lizzieLet17_5QNode_Int_5QError_Int_emitted[1]));
  assign lizzieLet17_5QNode_Int_5QError_Int_done = (lizzieLet17_5QNode_Int_5QError_Int_emitted | ({lizzieLet17_5QNode_Int_5QError_Int_2_d[0],
                                                                                                   lizzieLet17_5QNode_Int_5QError_Int_1_d[0]} & {lizzieLet17_5QNode_Int_5QError_Int_2_r,
                                                                                                                                                 lizzieLet17_5QNode_Int_5QError_Int_1_r}));
  assign lizzieLet17_5QNode_Int_5QError_Int_r = (& lizzieLet17_5QNode_Int_5QError_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_5QError_Int_emitted <= 2'd0;
    else
      lizzieLet17_5QNode_Int_5QError_Int_emitted <= (lizzieLet17_5QNode_Int_5QError_Int_r ? 2'd0 :
                                                     lizzieLet17_5QNode_Int_5QError_Int_done);
  
  /* dcon (Ty QTree_Int,
      Dcon QError_Int) : [(lizzieLet17_5QNode_Int_5QError_Int_1,Go)] > (lizzieLet17_5QNode_Int_5QError_Int_1QError_Int,QTree_Int) */
  assign lizzieLet17_5QNode_Int_5QError_Int_1QError_Int_d = QError_Int_dc((& {lizzieLet17_5QNode_Int_5QError_Int_1_d[0]}), lizzieLet17_5QNode_Int_5QError_Int_1_d);
  assign {lizzieLet17_5QNode_Int_5QError_Int_1_r} = {1 {(lizzieLet17_5QNode_Int_5QError_Int_1QError_Int_r && lizzieLet17_5QNode_Int_5QError_Int_1QError_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (lizzieLet17_5QNode_Int_5QError_Int_1QError_Int,QTree_Int) > (lizzieLet54_1_argbuf,QTree_Int) */
  QTree_Int_t lizzieLet17_5QNode_Int_5QError_Int_1QError_Int_bufchan_d;
  logic lizzieLet17_5QNode_Int_5QError_Int_1QError_Int_bufchan_r;
  assign lizzieLet17_5QNode_Int_5QError_Int_1QError_Int_r = ((! lizzieLet17_5QNode_Int_5QError_Int_1QError_Int_bufchan_d[0]) || lizzieLet17_5QNode_Int_5QError_Int_1QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_5QError_Int_1QError_Int_bufchan_d <= {66'd0,
                                                                   1'd0};
    else
      if (lizzieLet17_5QNode_Int_5QError_Int_1QError_Int_r)
        lizzieLet17_5QNode_Int_5QError_Int_1QError_Int_bufchan_d <= lizzieLet17_5QNode_Int_5QError_Int_1QError_Int_d;
  QTree_Int_t lizzieLet17_5QNode_Int_5QError_Int_1QError_Int_bufchan_buf;
  assign lizzieLet17_5QNode_Int_5QError_Int_1QError_Int_bufchan_r = (! lizzieLet17_5QNode_Int_5QError_Int_1QError_Int_bufchan_buf[0]);
  assign lizzieLet54_1_argbuf_d = (lizzieLet17_5QNode_Int_5QError_Int_1QError_Int_bufchan_buf[0] ? lizzieLet17_5QNode_Int_5QError_Int_1QError_Int_bufchan_buf :
                                   lizzieLet17_5QNode_Int_5QError_Int_1QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_5QError_Int_1QError_Int_bufchan_buf <= {66'd0,
                                                                     1'd0};
    else
      if ((lizzieLet54_1_argbuf_r && lizzieLet17_5QNode_Int_5QError_Int_1QError_Int_bufchan_buf[0]))
        lizzieLet17_5QNode_Int_5QError_Int_1QError_Int_bufchan_buf <= {66'd0,
                                                                       1'd0};
      else if (((! lizzieLet54_1_argbuf_r) && (! lizzieLet17_5QNode_Int_5QError_Int_1QError_Int_bufchan_buf[0])))
        lizzieLet17_5QNode_Int_5QError_Int_1QError_Int_bufchan_buf <= lizzieLet17_5QNode_Int_5QError_Int_1QError_Int_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet17_5QNode_Int_5QError_Int_2,Go) > (lizzieLet17_5QNode_Int_5QError_Int_2_argbuf,Go) */
  Go_t lizzieLet17_5QNode_Int_5QError_Int_2_bufchan_d;
  logic lizzieLet17_5QNode_Int_5QError_Int_2_bufchan_r;
  assign lizzieLet17_5QNode_Int_5QError_Int_2_r = ((! lizzieLet17_5QNode_Int_5QError_Int_2_bufchan_d[0]) || lizzieLet17_5QNode_Int_5QError_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_5QError_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet17_5QNode_Int_5QError_Int_2_r)
        lizzieLet17_5QNode_Int_5QError_Int_2_bufchan_d <= lizzieLet17_5QNode_Int_5QError_Int_2_d;
  Go_t lizzieLet17_5QNode_Int_5QError_Int_2_bufchan_buf;
  assign lizzieLet17_5QNode_Int_5QError_Int_2_bufchan_r = (! lizzieLet17_5QNode_Int_5QError_Int_2_bufchan_buf[0]);
  assign lizzieLet17_5QNode_Int_5QError_Int_2_argbuf_d = (lizzieLet17_5QNode_Int_5QError_Int_2_bufchan_buf[0] ? lizzieLet17_5QNode_Int_5QError_Int_2_bufchan_buf :
                                                          lizzieLet17_5QNode_Int_5QError_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_5QError_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet17_5QNode_Int_5QError_Int_2_argbuf_r && lizzieLet17_5QNode_Int_5QError_Int_2_bufchan_buf[0]))
        lizzieLet17_5QNode_Int_5QError_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet17_5QNode_Int_5QError_Int_2_argbuf_r) && (! lizzieLet17_5QNode_Int_5QError_Int_2_bufchan_buf[0])))
        lizzieLet17_5QNode_Int_5QError_Int_2_bufchan_buf <= lizzieLet17_5QNode_Int_5QError_Int_2_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet17_5QNode_Int_5QVal_Int,Go) > [(lizzieLet17_5QNode_Int_5QVal_Int_1,Go),
                                                        (lizzieLet17_5QNode_Int_5QVal_Int_2,Go)] */
  logic [1:0] lizzieLet17_5QNode_Int_5QVal_Int_emitted;
  logic [1:0] lizzieLet17_5QNode_Int_5QVal_Int_done;
  assign lizzieLet17_5QNode_Int_5QVal_Int_1_d = (lizzieLet17_5QNode_Int_5QVal_Int_d[0] && (! lizzieLet17_5QNode_Int_5QVal_Int_emitted[0]));
  assign lizzieLet17_5QNode_Int_5QVal_Int_2_d = (lizzieLet17_5QNode_Int_5QVal_Int_d[0] && (! lizzieLet17_5QNode_Int_5QVal_Int_emitted[1]));
  assign lizzieLet17_5QNode_Int_5QVal_Int_done = (lizzieLet17_5QNode_Int_5QVal_Int_emitted | ({lizzieLet17_5QNode_Int_5QVal_Int_2_d[0],
                                                                                               lizzieLet17_5QNode_Int_5QVal_Int_1_d[0]} & {lizzieLet17_5QNode_Int_5QVal_Int_2_r,
                                                                                                                                           lizzieLet17_5QNode_Int_5QVal_Int_1_r}));
  assign lizzieLet17_5QNode_Int_5QVal_Int_r = (& lizzieLet17_5QNode_Int_5QVal_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_5QVal_Int_emitted <= 2'd0;
    else
      lizzieLet17_5QNode_Int_5QVal_Int_emitted <= (lizzieLet17_5QNode_Int_5QVal_Int_r ? 2'd0 :
                                                   lizzieLet17_5QNode_Int_5QVal_Int_done);
  
  /* dcon (Ty QTree_Int,
      Dcon QError_Int) : [(lizzieLet17_5QNode_Int_5QVal_Int_1,Go)] > (lizzieLet17_5QNode_Int_5QVal_Int_1QError_Int,QTree_Int) */
  assign lizzieLet17_5QNode_Int_5QVal_Int_1QError_Int_d = QError_Int_dc((& {lizzieLet17_5QNode_Int_5QVal_Int_1_d[0]}), lizzieLet17_5QNode_Int_5QVal_Int_1_d);
  assign {lizzieLet17_5QNode_Int_5QVal_Int_1_r} = {1 {(lizzieLet17_5QNode_Int_5QVal_Int_1QError_Int_r && lizzieLet17_5QNode_Int_5QVal_Int_1QError_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (lizzieLet17_5QNode_Int_5QVal_Int_1QError_Int,QTree_Int) > (lizzieLet48_1_argbuf,QTree_Int) */
  QTree_Int_t lizzieLet17_5QNode_Int_5QVal_Int_1QError_Int_bufchan_d;
  logic lizzieLet17_5QNode_Int_5QVal_Int_1QError_Int_bufchan_r;
  assign lizzieLet17_5QNode_Int_5QVal_Int_1QError_Int_r = ((! lizzieLet17_5QNode_Int_5QVal_Int_1QError_Int_bufchan_d[0]) || lizzieLet17_5QNode_Int_5QVal_Int_1QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_5QVal_Int_1QError_Int_bufchan_d <= {66'd0,
                                                                 1'd0};
    else
      if (lizzieLet17_5QNode_Int_5QVal_Int_1QError_Int_r)
        lizzieLet17_5QNode_Int_5QVal_Int_1QError_Int_bufchan_d <= lizzieLet17_5QNode_Int_5QVal_Int_1QError_Int_d;
  QTree_Int_t lizzieLet17_5QNode_Int_5QVal_Int_1QError_Int_bufchan_buf;
  assign lizzieLet17_5QNode_Int_5QVal_Int_1QError_Int_bufchan_r = (! lizzieLet17_5QNode_Int_5QVal_Int_1QError_Int_bufchan_buf[0]);
  assign lizzieLet48_1_argbuf_d = (lizzieLet17_5QNode_Int_5QVal_Int_1QError_Int_bufchan_buf[0] ? lizzieLet17_5QNode_Int_5QVal_Int_1QError_Int_bufchan_buf :
                                   lizzieLet17_5QNode_Int_5QVal_Int_1QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_5QVal_Int_1QError_Int_bufchan_buf <= {66'd0,
                                                                   1'd0};
    else
      if ((lizzieLet48_1_argbuf_r && lizzieLet17_5QNode_Int_5QVal_Int_1QError_Int_bufchan_buf[0]))
        lizzieLet17_5QNode_Int_5QVal_Int_1QError_Int_bufchan_buf <= {66'd0,
                                                                     1'd0};
      else if (((! lizzieLet48_1_argbuf_r) && (! lizzieLet17_5QNode_Int_5QVal_Int_1QError_Int_bufchan_buf[0])))
        lizzieLet17_5QNode_Int_5QVal_Int_1QError_Int_bufchan_buf <= lizzieLet17_5QNode_Int_5QVal_Int_1QError_Int_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet17_5QNode_Int_5QVal_Int_2,Go) > (lizzieLet17_5QNode_Int_5QVal_Int_2_argbuf,Go) */
  Go_t lizzieLet17_5QNode_Int_5QVal_Int_2_bufchan_d;
  logic lizzieLet17_5QNode_Int_5QVal_Int_2_bufchan_r;
  assign lizzieLet17_5QNode_Int_5QVal_Int_2_r = ((! lizzieLet17_5QNode_Int_5QVal_Int_2_bufchan_d[0]) || lizzieLet17_5QNode_Int_5QVal_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_5QVal_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet17_5QNode_Int_5QVal_Int_2_r)
        lizzieLet17_5QNode_Int_5QVal_Int_2_bufchan_d <= lizzieLet17_5QNode_Int_5QVal_Int_2_d;
  Go_t lizzieLet17_5QNode_Int_5QVal_Int_2_bufchan_buf;
  assign lizzieLet17_5QNode_Int_5QVal_Int_2_bufchan_r = (! lizzieLet17_5QNode_Int_5QVal_Int_2_bufchan_buf[0]);
  assign lizzieLet17_5QNode_Int_5QVal_Int_2_argbuf_d = (lizzieLet17_5QNode_Int_5QVal_Int_2_bufchan_buf[0] ? lizzieLet17_5QNode_Int_5QVal_Int_2_bufchan_buf :
                                                        lizzieLet17_5QNode_Int_5QVal_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_5QVal_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet17_5QNode_Int_5QVal_Int_2_argbuf_r && lizzieLet17_5QNode_Int_5QVal_Int_2_bufchan_buf[0]))
        lizzieLet17_5QNode_Int_5QVal_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet17_5QNode_Int_5QVal_Int_2_argbuf_r) && (! lizzieLet17_5QNode_Int_5QVal_Int_2_bufchan_buf[0])))
        lizzieLet17_5QNode_Int_5QVal_Int_2_bufchan_buf <= lizzieLet17_5QNode_Int_5QVal_Int_2_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty MyDTInt_Bool) : (lizzieLet17_5QNode_Int_6,QTree_Int) (lizzieLet17_4QNode_Int,MyDTInt_Bool) > [(lizzieLet17_5QNode_Int_6QNone_Int,MyDTInt_Bool),
                                                                                                        (_208,MyDTInt_Bool),
                                                                                                        (lizzieLet17_5QNode_Int_6QNode_Int,MyDTInt_Bool),
                                                                                                        (_207,MyDTInt_Bool)] */
  logic [3:0] lizzieLet17_4QNode_Int_onehotd;
  always_comb
    if ((lizzieLet17_5QNode_Int_6_d[0] && lizzieLet17_4QNode_Int_d[0]))
      unique case (lizzieLet17_5QNode_Int_6_d[2:1])
        2'd0: lizzieLet17_4QNode_Int_onehotd = 4'd1;
        2'd1: lizzieLet17_4QNode_Int_onehotd = 4'd2;
        2'd2: lizzieLet17_4QNode_Int_onehotd = 4'd4;
        2'd3: lizzieLet17_4QNode_Int_onehotd = 4'd8;
        default: lizzieLet17_4QNode_Int_onehotd = 4'd0;
      endcase
    else lizzieLet17_4QNode_Int_onehotd = 4'd0;
  assign lizzieLet17_5QNode_Int_6QNone_Int_d = lizzieLet17_4QNode_Int_onehotd[0];
  assign _208_d = lizzieLet17_4QNode_Int_onehotd[1];
  assign lizzieLet17_5QNode_Int_6QNode_Int_d = lizzieLet17_4QNode_Int_onehotd[2];
  assign _207_d = lizzieLet17_4QNode_Int_onehotd[3];
  assign lizzieLet17_4QNode_Int_r = (| (lizzieLet17_4QNode_Int_onehotd & {_207_r,
                                                                          lizzieLet17_5QNode_Int_6QNode_Int_r,
                                                                          _208_r,
                                                                          lizzieLet17_5QNode_Int_6QNone_Int_r}));
  assign lizzieLet17_5QNode_Int_6_r = lizzieLet17_4QNode_Int_r;
  
  /* demux (Ty QTree_Int,
       Ty QTree_Int) : (lizzieLet17_5QNode_Int_7,QTree_Int) (lizzieLet17_6QNode_Int,QTree_Int) > [(lizzieLet17_5QNode_Int_7QNone_Int,QTree_Int),
                                                                                                  (_206,QTree_Int),
                                                                                                  (lizzieLet17_5QNode_Int_7QNode_Int,QTree_Int),
                                                                                                  (_205,QTree_Int)] */
  logic [3:0] lizzieLet17_6QNode_Int_onehotd;
  always_comb
    if ((lizzieLet17_5QNode_Int_7_d[0] && lizzieLet17_6QNode_Int_d[0]))
      unique case (lizzieLet17_5QNode_Int_7_d[2:1])
        2'd0: lizzieLet17_6QNode_Int_onehotd = 4'd1;
        2'd1: lizzieLet17_6QNode_Int_onehotd = 4'd2;
        2'd2: lizzieLet17_6QNode_Int_onehotd = 4'd4;
        2'd3: lizzieLet17_6QNode_Int_onehotd = 4'd8;
        default: lizzieLet17_6QNode_Int_onehotd = 4'd0;
      endcase
    else lizzieLet17_6QNode_Int_onehotd = 4'd0;
  assign lizzieLet17_5QNode_Int_7QNone_Int_d = {lizzieLet17_6QNode_Int_d[66:1],
                                                lizzieLet17_6QNode_Int_onehotd[0]};
  assign _206_d = {lizzieLet17_6QNode_Int_d[66:1],
                   lizzieLet17_6QNode_Int_onehotd[1]};
  assign lizzieLet17_5QNode_Int_7QNode_Int_d = {lizzieLet17_6QNode_Int_d[66:1],
                                                lizzieLet17_6QNode_Int_onehotd[2]};
  assign _205_d = {lizzieLet17_6QNode_Int_d[66:1],
                   lizzieLet17_6QNode_Int_onehotd[3]};
  assign lizzieLet17_6QNode_Int_r = (| (lizzieLet17_6QNode_Int_onehotd & {_205_r,
                                                                          lizzieLet17_5QNode_Int_7QNode_Int_r,
                                                                          _206_r,
                                                                          lizzieLet17_5QNode_Int_7QNone_Int_r}));
  assign lizzieLet17_5QNode_Int_7_r = lizzieLet17_6QNode_Int_r;
  
  /* fork (Ty QTree_Int) : (lizzieLet17_5QNode_Int_7QNode_Int,QTree_Int) > [(lizzieLet17_5QNode_Int_7QNode_Int_1,QTree_Int),
                                                                       (lizzieLet17_5QNode_Int_7QNode_Int_2,QTree_Int),
                                                                       (lizzieLet17_5QNode_Int_7QNode_Int_3,QTree_Int),
                                                                       (lizzieLet17_5QNode_Int_7QNode_Int_4,QTree_Int),
                                                                       (lizzieLet17_5QNode_Int_7QNode_Int_5,QTree_Int),
                                                                       (lizzieLet17_5QNode_Int_7QNode_Int_6,QTree_Int),
                                                                       (lizzieLet17_5QNode_Int_7QNode_Int_7,QTree_Int),
                                                                       (lizzieLet17_5QNode_Int_7QNode_Int_8,QTree_Int),
                                                                       (lizzieLet17_5QNode_Int_7QNode_Int_9,QTree_Int),
                                                                       (lizzieLet17_5QNode_Int_7QNode_Int_10,QTree_Int),
                                                                       (lizzieLet17_5QNode_Int_7QNode_Int_11,QTree_Int),
                                                                       (lizzieLet17_5QNode_Int_7QNode_Int_12,QTree_Int),
                                                                       (lizzieLet17_5QNode_Int_7QNode_Int_13,QTree_Int),
                                                                       (lizzieLet17_5QNode_Int_7QNode_Int_14,QTree_Int)] */
  logic [13:0] lizzieLet17_5QNode_Int_7QNode_Int_emitted;
  logic [13:0] lizzieLet17_5QNode_Int_7QNode_Int_done;
  assign lizzieLet17_5QNode_Int_7QNode_Int_1_d = {lizzieLet17_5QNode_Int_7QNode_Int_d[66:1],
                                                  (lizzieLet17_5QNode_Int_7QNode_Int_d[0] && (! lizzieLet17_5QNode_Int_7QNode_Int_emitted[0]))};
  assign lizzieLet17_5QNode_Int_7QNode_Int_2_d = {lizzieLet17_5QNode_Int_7QNode_Int_d[66:1],
                                                  (lizzieLet17_5QNode_Int_7QNode_Int_d[0] && (! lizzieLet17_5QNode_Int_7QNode_Int_emitted[1]))};
  assign lizzieLet17_5QNode_Int_7QNode_Int_3_d = {lizzieLet17_5QNode_Int_7QNode_Int_d[66:1],
                                                  (lizzieLet17_5QNode_Int_7QNode_Int_d[0] && (! lizzieLet17_5QNode_Int_7QNode_Int_emitted[2]))};
  assign lizzieLet17_5QNode_Int_7QNode_Int_4_d = {lizzieLet17_5QNode_Int_7QNode_Int_d[66:1],
                                                  (lizzieLet17_5QNode_Int_7QNode_Int_d[0] && (! lizzieLet17_5QNode_Int_7QNode_Int_emitted[3]))};
  assign lizzieLet17_5QNode_Int_7QNode_Int_5_d = {lizzieLet17_5QNode_Int_7QNode_Int_d[66:1],
                                                  (lizzieLet17_5QNode_Int_7QNode_Int_d[0] && (! lizzieLet17_5QNode_Int_7QNode_Int_emitted[4]))};
  assign lizzieLet17_5QNode_Int_7QNode_Int_6_d = {lizzieLet17_5QNode_Int_7QNode_Int_d[66:1],
                                                  (lizzieLet17_5QNode_Int_7QNode_Int_d[0] && (! lizzieLet17_5QNode_Int_7QNode_Int_emitted[5]))};
  assign lizzieLet17_5QNode_Int_7QNode_Int_7_d = {lizzieLet17_5QNode_Int_7QNode_Int_d[66:1],
                                                  (lizzieLet17_5QNode_Int_7QNode_Int_d[0] && (! lizzieLet17_5QNode_Int_7QNode_Int_emitted[6]))};
  assign lizzieLet17_5QNode_Int_7QNode_Int_8_d = {lizzieLet17_5QNode_Int_7QNode_Int_d[66:1],
                                                  (lizzieLet17_5QNode_Int_7QNode_Int_d[0] && (! lizzieLet17_5QNode_Int_7QNode_Int_emitted[7]))};
  assign lizzieLet17_5QNode_Int_7QNode_Int_9_d = {lizzieLet17_5QNode_Int_7QNode_Int_d[66:1],
                                                  (lizzieLet17_5QNode_Int_7QNode_Int_d[0] && (! lizzieLet17_5QNode_Int_7QNode_Int_emitted[8]))};
  assign lizzieLet17_5QNode_Int_7QNode_Int_10_d = {lizzieLet17_5QNode_Int_7QNode_Int_d[66:1],
                                                   (lizzieLet17_5QNode_Int_7QNode_Int_d[0] && (! lizzieLet17_5QNode_Int_7QNode_Int_emitted[9]))};
  assign lizzieLet17_5QNode_Int_7QNode_Int_11_d = {lizzieLet17_5QNode_Int_7QNode_Int_d[66:1],
                                                   (lizzieLet17_5QNode_Int_7QNode_Int_d[0] && (! lizzieLet17_5QNode_Int_7QNode_Int_emitted[10]))};
  assign lizzieLet17_5QNode_Int_7QNode_Int_12_d = {lizzieLet17_5QNode_Int_7QNode_Int_d[66:1],
                                                   (lizzieLet17_5QNode_Int_7QNode_Int_d[0] && (! lizzieLet17_5QNode_Int_7QNode_Int_emitted[11]))};
  assign lizzieLet17_5QNode_Int_7QNode_Int_13_d = {lizzieLet17_5QNode_Int_7QNode_Int_d[66:1],
                                                   (lizzieLet17_5QNode_Int_7QNode_Int_d[0] && (! lizzieLet17_5QNode_Int_7QNode_Int_emitted[12]))};
  assign lizzieLet17_5QNode_Int_7QNode_Int_14_d = {lizzieLet17_5QNode_Int_7QNode_Int_d[66:1],
                                                   (lizzieLet17_5QNode_Int_7QNode_Int_d[0] && (! lizzieLet17_5QNode_Int_7QNode_Int_emitted[13]))};
  assign lizzieLet17_5QNode_Int_7QNode_Int_done = (lizzieLet17_5QNode_Int_7QNode_Int_emitted | ({lizzieLet17_5QNode_Int_7QNode_Int_14_d[0],
                                                                                                 lizzieLet17_5QNode_Int_7QNode_Int_13_d[0],
                                                                                                 lizzieLet17_5QNode_Int_7QNode_Int_12_d[0],
                                                                                                 lizzieLet17_5QNode_Int_7QNode_Int_11_d[0],
                                                                                                 lizzieLet17_5QNode_Int_7QNode_Int_10_d[0],
                                                                                                 lizzieLet17_5QNode_Int_7QNode_Int_9_d[0],
                                                                                                 lizzieLet17_5QNode_Int_7QNode_Int_8_d[0],
                                                                                                 lizzieLet17_5QNode_Int_7QNode_Int_7_d[0],
                                                                                                 lizzieLet17_5QNode_Int_7QNode_Int_6_d[0],
                                                                                                 lizzieLet17_5QNode_Int_7QNode_Int_5_d[0],
                                                                                                 lizzieLet17_5QNode_Int_7QNode_Int_4_d[0],
                                                                                                 lizzieLet17_5QNode_Int_7QNode_Int_3_d[0],
                                                                                                 lizzieLet17_5QNode_Int_7QNode_Int_2_d[0],
                                                                                                 lizzieLet17_5QNode_Int_7QNode_Int_1_d[0]} & {lizzieLet17_5QNode_Int_7QNode_Int_14_r,
                                                                                                                                              lizzieLet17_5QNode_Int_7QNode_Int_13_r,
                                                                                                                                              lizzieLet17_5QNode_Int_7QNode_Int_12_r,
                                                                                                                                              lizzieLet17_5QNode_Int_7QNode_Int_11_r,
                                                                                                                                              lizzieLet17_5QNode_Int_7QNode_Int_10_r,
                                                                                                                                              lizzieLet17_5QNode_Int_7QNode_Int_9_r,
                                                                                                                                              lizzieLet17_5QNode_Int_7QNode_Int_8_r,
                                                                                                                                              lizzieLet17_5QNode_Int_7QNode_Int_7_r,
                                                                                                                                              lizzieLet17_5QNode_Int_7QNode_Int_6_r,
                                                                                                                                              lizzieLet17_5QNode_Int_7QNode_Int_5_r,
                                                                                                                                              lizzieLet17_5QNode_Int_7QNode_Int_4_r,
                                                                                                                                              lizzieLet17_5QNode_Int_7QNode_Int_3_r,
                                                                                                                                              lizzieLet17_5QNode_Int_7QNode_Int_2_r,
                                                                                                                                              lizzieLet17_5QNode_Int_7QNode_Int_1_r}));
  assign lizzieLet17_5QNode_Int_7QNode_Int_r = (& lizzieLet17_5QNode_Int_7QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNode_Int_emitted <= 14'd0;
    else
      lizzieLet17_5QNode_Int_7QNode_Int_emitted <= (lizzieLet17_5QNode_Int_7QNode_Int_r ? 14'd0 :
                                                    lizzieLet17_5QNode_Int_7QNode_Int_done);
  
  /* demux (Ty QTree_Int,
       Ty Pointer_QTree_Int) : (lizzieLet17_5QNode_Int_7QNode_Int_10,QTree_Int) (lizzieLet17_5QNode_Int_9QNode_Int,Pointer_QTree_Int) > [(lizzieLet17_5QNode_Int_7QNode_Int_10QNone_Int,Pointer_QTree_Int),
                                                                                                                                         (_204,Pointer_QTree_Int),
                                                                                                                                         (lizzieLet17_5QNode_Int_7QNode_Int_10QNode_Int,Pointer_QTree_Int),
                                                                                                                                         (_203,Pointer_QTree_Int)] */
  logic [3:0] lizzieLet17_5QNode_Int_9QNode_Int_onehotd;
  always_comb
    if ((lizzieLet17_5QNode_Int_7QNode_Int_10_d[0] && lizzieLet17_5QNode_Int_9QNode_Int_d[0]))
      unique case (lizzieLet17_5QNode_Int_7QNode_Int_10_d[2:1])
        2'd0: lizzieLet17_5QNode_Int_9QNode_Int_onehotd = 4'd1;
        2'd1: lizzieLet17_5QNode_Int_9QNode_Int_onehotd = 4'd2;
        2'd2: lizzieLet17_5QNode_Int_9QNode_Int_onehotd = 4'd4;
        2'd3: lizzieLet17_5QNode_Int_9QNode_Int_onehotd = 4'd8;
        default: lizzieLet17_5QNode_Int_9QNode_Int_onehotd = 4'd0;
      endcase
    else lizzieLet17_5QNode_Int_9QNode_Int_onehotd = 4'd0;
  assign lizzieLet17_5QNode_Int_7QNode_Int_10QNone_Int_d = {lizzieLet17_5QNode_Int_9QNode_Int_d[16:1],
                                                            lizzieLet17_5QNode_Int_9QNode_Int_onehotd[0]};
  assign _204_d = {lizzieLet17_5QNode_Int_9QNode_Int_d[16:1],
                   lizzieLet17_5QNode_Int_9QNode_Int_onehotd[1]};
  assign lizzieLet17_5QNode_Int_7QNode_Int_10QNode_Int_d = {lizzieLet17_5QNode_Int_9QNode_Int_d[16:1],
                                                            lizzieLet17_5QNode_Int_9QNode_Int_onehotd[2]};
  assign _203_d = {lizzieLet17_5QNode_Int_9QNode_Int_d[16:1],
                   lizzieLet17_5QNode_Int_9QNode_Int_onehotd[3]};
  assign lizzieLet17_5QNode_Int_9QNode_Int_r = (| (lizzieLet17_5QNode_Int_9QNode_Int_onehotd & {_203_r,
                                                                                                lizzieLet17_5QNode_Int_7QNode_Int_10QNode_Int_r,
                                                                                                _204_r,
                                                                                                lizzieLet17_5QNode_Int_7QNode_Int_10QNone_Int_r}));
  assign lizzieLet17_5QNode_Int_7QNode_Int_10_r = lizzieLet17_5QNode_Int_9QNode_Int_r;
  
  /* buf (Ty Pointer_QTree_Int) : (lizzieLet17_5QNode_Int_7QNode_Int_10QNone_Int,Pointer_QTree_Int) > (lizzieLet17_5QNode_Int_7QNode_Int_10QNone_Int_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t lizzieLet17_5QNode_Int_7QNode_Int_10QNone_Int_bufchan_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_10QNone_Int_bufchan_r;
  assign lizzieLet17_5QNode_Int_7QNode_Int_10QNone_Int_r = ((! lizzieLet17_5QNode_Int_7QNode_Int_10QNone_Int_bufchan_d[0]) || lizzieLet17_5QNode_Int_7QNode_Int_10QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNode_Int_10QNone_Int_bufchan_d <= {16'd0,
                                                                  1'd0};
    else
      if (lizzieLet17_5QNode_Int_7QNode_Int_10QNone_Int_r)
        lizzieLet17_5QNode_Int_7QNode_Int_10QNone_Int_bufchan_d <= lizzieLet17_5QNode_Int_7QNode_Int_10QNone_Int_d;
  Pointer_QTree_Int_t lizzieLet17_5QNode_Int_7QNode_Int_10QNone_Int_bufchan_buf;
  assign lizzieLet17_5QNode_Int_7QNode_Int_10QNone_Int_bufchan_r = (! lizzieLet17_5QNode_Int_7QNode_Int_10QNone_Int_bufchan_buf[0]);
  assign lizzieLet17_5QNode_Int_7QNode_Int_10QNone_Int_1_argbuf_d = (lizzieLet17_5QNode_Int_7QNode_Int_10QNone_Int_bufchan_buf[0] ? lizzieLet17_5QNode_Int_7QNode_Int_10QNone_Int_bufchan_buf :
                                                                     lizzieLet17_5QNode_Int_7QNode_Int_10QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNode_Int_10QNone_Int_bufchan_buf <= {16'd0,
                                                                    1'd0};
    else
      if ((lizzieLet17_5QNode_Int_7QNode_Int_10QNone_Int_1_argbuf_r && lizzieLet17_5QNode_Int_7QNode_Int_10QNone_Int_bufchan_buf[0]))
        lizzieLet17_5QNode_Int_7QNode_Int_10QNone_Int_bufchan_buf <= {16'd0,
                                                                      1'd0};
      else if (((! lizzieLet17_5QNode_Int_7QNode_Int_10QNone_Int_1_argbuf_r) && (! lizzieLet17_5QNode_Int_7QNode_Int_10QNone_Int_bufchan_buf[0])))
        lizzieLet17_5QNode_Int_7QNode_Int_10QNone_Int_bufchan_buf <= lizzieLet17_5QNode_Int_7QNode_Int_10QNone_Int_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_QTree_Int) : (lizzieLet17_5QNode_Int_7QNode_Int_11,QTree_Int) (t1afa_destruct,Pointer_QTree_Int) > [(lizzieLet17_5QNode_Int_7QNode_Int_11QNone_Int,Pointer_QTree_Int),
                                                                                                                      (_202,Pointer_QTree_Int),
                                                                                                                      (lizzieLet17_5QNode_Int_7QNode_Int_11QNode_Int,Pointer_QTree_Int),
                                                                                                                      (_201,Pointer_QTree_Int)] */
  logic [3:0] t1afa_destruct_onehotd;
  always_comb
    if ((lizzieLet17_5QNode_Int_7QNode_Int_11_d[0] && t1afa_destruct_d[0]))
      unique case (lizzieLet17_5QNode_Int_7QNode_Int_11_d[2:1])
        2'd0: t1afa_destruct_onehotd = 4'd1;
        2'd1: t1afa_destruct_onehotd = 4'd2;
        2'd2: t1afa_destruct_onehotd = 4'd4;
        2'd3: t1afa_destruct_onehotd = 4'd8;
        default: t1afa_destruct_onehotd = 4'd0;
      endcase
    else t1afa_destruct_onehotd = 4'd0;
  assign lizzieLet17_5QNode_Int_7QNode_Int_11QNone_Int_d = {t1afa_destruct_d[16:1],
                                                            t1afa_destruct_onehotd[0]};
  assign _202_d = {t1afa_destruct_d[16:1],
                   t1afa_destruct_onehotd[1]};
  assign lizzieLet17_5QNode_Int_7QNode_Int_11QNode_Int_d = {t1afa_destruct_d[16:1],
                                                            t1afa_destruct_onehotd[2]};
  assign _201_d = {t1afa_destruct_d[16:1],
                   t1afa_destruct_onehotd[3]};
  assign t1afa_destruct_r = (| (t1afa_destruct_onehotd & {_201_r,
                                                          lizzieLet17_5QNode_Int_7QNode_Int_11QNode_Int_r,
                                                          _202_r,
                                                          lizzieLet17_5QNode_Int_7QNode_Int_11QNone_Int_r}));
  assign lizzieLet17_5QNode_Int_7QNode_Int_11_r = t1afa_destruct_r;
  
  /* buf (Ty Pointer_QTree_Int) : (lizzieLet17_5QNode_Int_7QNode_Int_11QNone_Int,Pointer_QTree_Int) > (lizzieLet17_5QNode_Int_7QNode_Int_11QNone_Int_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t lizzieLet17_5QNode_Int_7QNode_Int_11QNone_Int_bufchan_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_11QNone_Int_bufchan_r;
  assign lizzieLet17_5QNode_Int_7QNode_Int_11QNone_Int_r = ((! lizzieLet17_5QNode_Int_7QNode_Int_11QNone_Int_bufchan_d[0]) || lizzieLet17_5QNode_Int_7QNode_Int_11QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNode_Int_11QNone_Int_bufchan_d <= {16'd0,
                                                                  1'd0};
    else
      if (lizzieLet17_5QNode_Int_7QNode_Int_11QNone_Int_r)
        lizzieLet17_5QNode_Int_7QNode_Int_11QNone_Int_bufchan_d <= lizzieLet17_5QNode_Int_7QNode_Int_11QNone_Int_d;
  Pointer_QTree_Int_t lizzieLet17_5QNode_Int_7QNode_Int_11QNone_Int_bufchan_buf;
  assign lizzieLet17_5QNode_Int_7QNode_Int_11QNone_Int_bufchan_r = (! lizzieLet17_5QNode_Int_7QNode_Int_11QNone_Int_bufchan_buf[0]);
  assign lizzieLet17_5QNode_Int_7QNode_Int_11QNone_Int_1_argbuf_d = (lizzieLet17_5QNode_Int_7QNode_Int_11QNone_Int_bufchan_buf[0] ? lizzieLet17_5QNode_Int_7QNode_Int_11QNone_Int_bufchan_buf :
                                                                     lizzieLet17_5QNode_Int_7QNode_Int_11QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNode_Int_11QNone_Int_bufchan_buf <= {16'd0,
                                                                    1'd0};
    else
      if ((lizzieLet17_5QNode_Int_7QNode_Int_11QNone_Int_1_argbuf_r && lizzieLet17_5QNode_Int_7QNode_Int_11QNone_Int_bufchan_buf[0]))
        lizzieLet17_5QNode_Int_7QNode_Int_11QNone_Int_bufchan_buf <= {16'd0,
                                                                      1'd0};
      else if (((! lizzieLet17_5QNode_Int_7QNode_Int_11QNone_Int_1_argbuf_r) && (! lizzieLet17_5QNode_Int_7QNode_Int_11QNone_Int_bufchan_buf[0])))
        lizzieLet17_5QNode_Int_7QNode_Int_11QNone_Int_bufchan_buf <= lizzieLet17_5QNode_Int_7QNode_Int_11QNone_Int_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_QTree_Int) : (lizzieLet17_5QNode_Int_7QNode_Int_12,QTree_Int) (t2afb_destruct,Pointer_QTree_Int) > [(lizzieLet17_5QNode_Int_7QNode_Int_12QNone_Int,Pointer_QTree_Int),
                                                                                                                      (_200,Pointer_QTree_Int),
                                                                                                                      (lizzieLet17_5QNode_Int_7QNode_Int_12QNode_Int,Pointer_QTree_Int),
                                                                                                                      (_199,Pointer_QTree_Int)] */
  logic [3:0] t2afb_destruct_onehotd;
  always_comb
    if ((lizzieLet17_5QNode_Int_7QNode_Int_12_d[0] && t2afb_destruct_d[0]))
      unique case (lizzieLet17_5QNode_Int_7QNode_Int_12_d[2:1])
        2'd0: t2afb_destruct_onehotd = 4'd1;
        2'd1: t2afb_destruct_onehotd = 4'd2;
        2'd2: t2afb_destruct_onehotd = 4'd4;
        2'd3: t2afb_destruct_onehotd = 4'd8;
        default: t2afb_destruct_onehotd = 4'd0;
      endcase
    else t2afb_destruct_onehotd = 4'd0;
  assign lizzieLet17_5QNode_Int_7QNode_Int_12QNone_Int_d = {t2afb_destruct_d[16:1],
                                                            t2afb_destruct_onehotd[0]};
  assign _200_d = {t2afb_destruct_d[16:1],
                   t2afb_destruct_onehotd[1]};
  assign lizzieLet17_5QNode_Int_7QNode_Int_12QNode_Int_d = {t2afb_destruct_d[16:1],
                                                            t2afb_destruct_onehotd[2]};
  assign _199_d = {t2afb_destruct_d[16:1],
                   t2afb_destruct_onehotd[3]};
  assign t2afb_destruct_r = (| (t2afb_destruct_onehotd & {_199_r,
                                                          lizzieLet17_5QNode_Int_7QNode_Int_12QNode_Int_r,
                                                          _200_r,
                                                          lizzieLet17_5QNode_Int_7QNode_Int_12QNone_Int_r}));
  assign lizzieLet17_5QNode_Int_7QNode_Int_12_r = t2afb_destruct_r;
  
  /* buf (Ty Pointer_QTree_Int) : (lizzieLet17_5QNode_Int_7QNode_Int_12QNone_Int,Pointer_QTree_Int) > (lizzieLet17_5QNode_Int_7QNode_Int_12QNone_Int_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t lizzieLet17_5QNode_Int_7QNode_Int_12QNone_Int_bufchan_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_12QNone_Int_bufchan_r;
  assign lizzieLet17_5QNode_Int_7QNode_Int_12QNone_Int_r = ((! lizzieLet17_5QNode_Int_7QNode_Int_12QNone_Int_bufchan_d[0]) || lizzieLet17_5QNode_Int_7QNode_Int_12QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNode_Int_12QNone_Int_bufchan_d <= {16'd0,
                                                                  1'd0};
    else
      if (lizzieLet17_5QNode_Int_7QNode_Int_12QNone_Int_r)
        lizzieLet17_5QNode_Int_7QNode_Int_12QNone_Int_bufchan_d <= lizzieLet17_5QNode_Int_7QNode_Int_12QNone_Int_d;
  Pointer_QTree_Int_t lizzieLet17_5QNode_Int_7QNode_Int_12QNone_Int_bufchan_buf;
  assign lizzieLet17_5QNode_Int_7QNode_Int_12QNone_Int_bufchan_r = (! lizzieLet17_5QNode_Int_7QNode_Int_12QNone_Int_bufchan_buf[0]);
  assign lizzieLet17_5QNode_Int_7QNode_Int_12QNone_Int_1_argbuf_d = (lizzieLet17_5QNode_Int_7QNode_Int_12QNone_Int_bufchan_buf[0] ? lizzieLet17_5QNode_Int_7QNode_Int_12QNone_Int_bufchan_buf :
                                                                     lizzieLet17_5QNode_Int_7QNode_Int_12QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNode_Int_12QNone_Int_bufchan_buf <= {16'd0,
                                                                    1'd0};
    else
      if ((lizzieLet17_5QNode_Int_7QNode_Int_12QNone_Int_1_argbuf_r && lizzieLet17_5QNode_Int_7QNode_Int_12QNone_Int_bufchan_buf[0]))
        lizzieLet17_5QNode_Int_7QNode_Int_12QNone_Int_bufchan_buf <= {16'd0,
                                                                      1'd0};
      else if (((! lizzieLet17_5QNode_Int_7QNode_Int_12QNone_Int_1_argbuf_r) && (! lizzieLet17_5QNode_Int_7QNode_Int_12QNone_Int_bufchan_buf[0])))
        lizzieLet17_5QNode_Int_7QNode_Int_12QNone_Int_bufchan_buf <= lizzieLet17_5QNode_Int_7QNode_Int_12QNone_Int_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_QTree_Int) : (lizzieLet17_5QNode_Int_7QNode_Int_13,QTree_Int) (t3afc_destruct,Pointer_QTree_Int) > [(lizzieLet17_5QNode_Int_7QNode_Int_13QNone_Int,Pointer_QTree_Int),
                                                                                                                      (_198,Pointer_QTree_Int),
                                                                                                                      (lizzieLet17_5QNode_Int_7QNode_Int_13QNode_Int,Pointer_QTree_Int),
                                                                                                                      (_197,Pointer_QTree_Int)] */
  logic [3:0] t3afc_destruct_onehotd;
  always_comb
    if ((lizzieLet17_5QNode_Int_7QNode_Int_13_d[0] && t3afc_destruct_d[0]))
      unique case (lizzieLet17_5QNode_Int_7QNode_Int_13_d[2:1])
        2'd0: t3afc_destruct_onehotd = 4'd1;
        2'd1: t3afc_destruct_onehotd = 4'd2;
        2'd2: t3afc_destruct_onehotd = 4'd4;
        2'd3: t3afc_destruct_onehotd = 4'd8;
        default: t3afc_destruct_onehotd = 4'd0;
      endcase
    else t3afc_destruct_onehotd = 4'd0;
  assign lizzieLet17_5QNode_Int_7QNode_Int_13QNone_Int_d = {t3afc_destruct_d[16:1],
                                                            t3afc_destruct_onehotd[0]};
  assign _198_d = {t3afc_destruct_d[16:1],
                   t3afc_destruct_onehotd[1]};
  assign lizzieLet17_5QNode_Int_7QNode_Int_13QNode_Int_d = {t3afc_destruct_d[16:1],
                                                            t3afc_destruct_onehotd[2]};
  assign _197_d = {t3afc_destruct_d[16:1],
                   t3afc_destruct_onehotd[3]};
  assign t3afc_destruct_r = (| (t3afc_destruct_onehotd & {_197_r,
                                                          lizzieLet17_5QNode_Int_7QNode_Int_13QNode_Int_r,
                                                          _198_r,
                                                          lizzieLet17_5QNode_Int_7QNode_Int_13QNone_Int_r}));
  assign lizzieLet17_5QNode_Int_7QNode_Int_13_r = t3afc_destruct_r;
  
  /* buf (Ty Pointer_QTree_Int) : (lizzieLet17_5QNode_Int_7QNode_Int_13QNone_Int,Pointer_QTree_Int) > (lizzieLet17_5QNode_Int_7QNode_Int_13QNone_Int_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t lizzieLet17_5QNode_Int_7QNode_Int_13QNone_Int_bufchan_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_13QNone_Int_bufchan_r;
  assign lizzieLet17_5QNode_Int_7QNode_Int_13QNone_Int_r = ((! lizzieLet17_5QNode_Int_7QNode_Int_13QNone_Int_bufchan_d[0]) || lizzieLet17_5QNode_Int_7QNode_Int_13QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNode_Int_13QNone_Int_bufchan_d <= {16'd0,
                                                                  1'd0};
    else
      if (lizzieLet17_5QNode_Int_7QNode_Int_13QNone_Int_r)
        lizzieLet17_5QNode_Int_7QNode_Int_13QNone_Int_bufchan_d <= lizzieLet17_5QNode_Int_7QNode_Int_13QNone_Int_d;
  Pointer_QTree_Int_t lizzieLet17_5QNode_Int_7QNode_Int_13QNone_Int_bufchan_buf;
  assign lizzieLet17_5QNode_Int_7QNode_Int_13QNone_Int_bufchan_r = (! lizzieLet17_5QNode_Int_7QNode_Int_13QNone_Int_bufchan_buf[0]);
  assign lizzieLet17_5QNode_Int_7QNode_Int_13QNone_Int_1_argbuf_d = (lizzieLet17_5QNode_Int_7QNode_Int_13QNone_Int_bufchan_buf[0] ? lizzieLet17_5QNode_Int_7QNode_Int_13QNone_Int_bufchan_buf :
                                                                     lizzieLet17_5QNode_Int_7QNode_Int_13QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNode_Int_13QNone_Int_bufchan_buf <= {16'd0,
                                                                    1'd0};
    else
      if ((lizzieLet17_5QNode_Int_7QNode_Int_13QNone_Int_1_argbuf_r && lizzieLet17_5QNode_Int_7QNode_Int_13QNone_Int_bufchan_buf[0]))
        lizzieLet17_5QNode_Int_7QNode_Int_13QNone_Int_bufchan_buf <= {16'd0,
                                                                      1'd0};
      else if (((! lizzieLet17_5QNode_Int_7QNode_Int_13QNone_Int_1_argbuf_r) && (! lizzieLet17_5QNode_Int_7QNode_Int_13QNone_Int_bufchan_buf[0])))
        lizzieLet17_5QNode_Int_7QNode_Int_13QNone_Int_bufchan_buf <= lizzieLet17_5QNode_Int_7QNode_Int_13QNone_Int_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_QTree_Int) : (lizzieLet17_5QNode_Int_7QNode_Int_14,QTree_Int) (t4afd_destruct,Pointer_QTree_Int) > [(lizzieLet17_5QNode_Int_7QNode_Int_14QNone_Int,Pointer_QTree_Int),
                                                                                                                      (_196,Pointer_QTree_Int),
                                                                                                                      (lizzieLet17_5QNode_Int_7QNode_Int_14QNode_Int,Pointer_QTree_Int),
                                                                                                                      (_195,Pointer_QTree_Int)] */
  logic [3:0] t4afd_destruct_onehotd;
  always_comb
    if ((lizzieLet17_5QNode_Int_7QNode_Int_14_d[0] && t4afd_destruct_d[0]))
      unique case (lizzieLet17_5QNode_Int_7QNode_Int_14_d[2:1])
        2'd0: t4afd_destruct_onehotd = 4'd1;
        2'd1: t4afd_destruct_onehotd = 4'd2;
        2'd2: t4afd_destruct_onehotd = 4'd4;
        2'd3: t4afd_destruct_onehotd = 4'd8;
        default: t4afd_destruct_onehotd = 4'd0;
      endcase
    else t4afd_destruct_onehotd = 4'd0;
  assign lizzieLet17_5QNode_Int_7QNode_Int_14QNone_Int_d = {t4afd_destruct_d[16:1],
                                                            t4afd_destruct_onehotd[0]};
  assign _196_d = {t4afd_destruct_d[16:1],
                   t4afd_destruct_onehotd[1]};
  assign lizzieLet17_5QNode_Int_7QNode_Int_14QNode_Int_d = {t4afd_destruct_d[16:1],
                                                            t4afd_destruct_onehotd[2]};
  assign _195_d = {t4afd_destruct_d[16:1],
                   t4afd_destruct_onehotd[3]};
  assign t4afd_destruct_r = (| (t4afd_destruct_onehotd & {_195_r,
                                                          lizzieLet17_5QNode_Int_7QNode_Int_14QNode_Int_r,
                                                          _196_r,
                                                          lizzieLet17_5QNode_Int_7QNode_Int_14QNone_Int_r}));
  assign lizzieLet17_5QNode_Int_7QNode_Int_14_r = t4afd_destruct_r;
  
  /* buf (Ty Pointer_QTree_Int) : (lizzieLet17_5QNode_Int_7QNode_Int_14QNode_Int,Pointer_QTree_Int) > (lizzieLet17_5QNode_Int_7QNode_Int_14QNode_Int_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t lizzieLet17_5QNode_Int_7QNode_Int_14QNode_Int_bufchan_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_14QNode_Int_bufchan_r;
  assign lizzieLet17_5QNode_Int_7QNode_Int_14QNode_Int_r = ((! lizzieLet17_5QNode_Int_7QNode_Int_14QNode_Int_bufchan_d[0]) || lizzieLet17_5QNode_Int_7QNode_Int_14QNode_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNode_Int_14QNode_Int_bufchan_d <= {16'd0,
                                                                  1'd0};
    else
      if (lizzieLet17_5QNode_Int_7QNode_Int_14QNode_Int_r)
        lizzieLet17_5QNode_Int_7QNode_Int_14QNode_Int_bufchan_d <= lizzieLet17_5QNode_Int_7QNode_Int_14QNode_Int_d;
  Pointer_QTree_Int_t lizzieLet17_5QNode_Int_7QNode_Int_14QNode_Int_bufchan_buf;
  assign lizzieLet17_5QNode_Int_7QNode_Int_14QNode_Int_bufchan_r = (! lizzieLet17_5QNode_Int_7QNode_Int_14QNode_Int_bufchan_buf[0]);
  assign lizzieLet17_5QNode_Int_7QNode_Int_14QNode_Int_1_argbuf_d = (lizzieLet17_5QNode_Int_7QNode_Int_14QNode_Int_bufchan_buf[0] ? lizzieLet17_5QNode_Int_7QNode_Int_14QNode_Int_bufchan_buf :
                                                                     lizzieLet17_5QNode_Int_7QNode_Int_14QNode_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNode_Int_14QNode_Int_bufchan_buf <= {16'd0,
                                                                    1'd0};
    else
      if ((lizzieLet17_5QNode_Int_7QNode_Int_14QNode_Int_1_argbuf_r && lizzieLet17_5QNode_Int_7QNode_Int_14QNode_Int_bufchan_buf[0]))
        lizzieLet17_5QNode_Int_7QNode_Int_14QNode_Int_bufchan_buf <= {16'd0,
                                                                      1'd0};
      else if (((! lizzieLet17_5QNode_Int_7QNode_Int_14QNode_Int_1_argbuf_r) && (! lizzieLet17_5QNode_Int_7QNode_Int_14QNode_Int_bufchan_buf[0])))
        lizzieLet17_5QNode_Int_7QNode_Int_14QNode_Int_bufchan_buf <= lizzieLet17_5QNode_Int_7QNode_Int_14QNode_Int_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (lizzieLet17_5QNode_Int_7QNode_Int_14QNone_Int,Pointer_QTree_Int) > (lizzieLet17_5QNode_Int_7QNode_Int_14QNone_Int_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t lizzieLet17_5QNode_Int_7QNode_Int_14QNone_Int_bufchan_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_14QNone_Int_bufchan_r;
  assign lizzieLet17_5QNode_Int_7QNode_Int_14QNone_Int_r = ((! lizzieLet17_5QNode_Int_7QNode_Int_14QNone_Int_bufchan_d[0]) || lizzieLet17_5QNode_Int_7QNode_Int_14QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNode_Int_14QNone_Int_bufchan_d <= {16'd0,
                                                                  1'd0};
    else
      if (lizzieLet17_5QNode_Int_7QNode_Int_14QNone_Int_r)
        lizzieLet17_5QNode_Int_7QNode_Int_14QNone_Int_bufchan_d <= lizzieLet17_5QNode_Int_7QNode_Int_14QNone_Int_d;
  Pointer_QTree_Int_t lizzieLet17_5QNode_Int_7QNode_Int_14QNone_Int_bufchan_buf;
  assign lizzieLet17_5QNode_Int_7QNode_Int_14QNone_Int_bufchan_r = (! lizzieLet17_5QNode_Int_7QNode_Int_14QNone_Int_bufchan_buf[0]);
  assign lizzieLet17_5QNode_Int_7QNode_Int_14QNone_Int_1_argbuf_d = (lizzieLet17_5QNode_Int_7QNode_Int_14QNone_Int_bufchan_buf[0] ? lizzieLet17_5QNode_Int_7QNode_Int_14QNone_Int_bufchan_buf :
                                                                     lizzieLet17_5QNode_Int_7QNode_Int_14QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNode_Int_14QNone_Int_bufchan_buf <= {16'd0,
                                                                    1'd0};
    else
      if ((lizzieLet17_5QNode_Int_7QNode_Int_14QNone_Int_1_argbuf_r && lizzieLet17_5QNode_Int_7QNode_Int_14QNone_Int_bufchan_buf[0]))
        lizzieLet17_5QNode_Int_7QNode_Int_14QNone_Int_bufchan_buf <= {16'd0,
                                                                      1'd0};
      else if (((! lizzieLet17_5QNode_Int_7QNode_Int_14QNone_Int_1_argbuf_r) && (! lizzieLet17_5QNode_Int_7QNode_Int_14QNone_Int_bufchan_buf[0])))
        lizzieLet17_5QNode_Int_7QNode_Int_14QNone_Int_bufchan_buf <= lizzieLet17_5QNode_Int_7QNode_Int_14QNone_Int_bufchan_d;
  
  /* destruct (Ty QTree_Int,
          Dcon QNode_Int) : (lizzieLet17_5QNode_Int_7QNode_Int_1QNode_Int,QTree_Int) > [(t1'aff_destruct,Pointer_QTree_Int),
                                                                                        (t2'afg_destruct,Pointer_QTree_Int),
                                                                                        (t3'afh_destruct,Pointer_QTree_Int),
                                                                                        (t4'afi_destruct,Pointer_QTree_Int)] */
  logic [3:0] lizzieLet17_5QNode_Int_7QNode_Int_1QNode_Int_emitted;
  logic [3:0] lizzieLet17_5QNode_Int_7QNode_Int_1QNode_Int_done;
  assign \t1'aff_destruct_d  = {lizzieLet17_5QNode_Int_7QNode_Int_1QNode_Int_d[18:3],
                                (lizzieLet17_5QNode_Int_7QNode_Int_1QNode_Int_d[0] && (! lizzieLet17_5QNode_Int_7QNode_Int_1QNode_Int_emitted[0]))};
  assign \t2'afg_destruct_d  = {lizzieLet17_5QNode_Int_7QNode_Int_1QNode_Int_d[34:19],
                                (lizzieLet17_5QNode_Int_7QNode_Int_1QNode_Int_d[0] && (! lizzieLet17_5QNode_Int_7QNode_Int_1QNode_Int_emitted[1]))};
  assign \t3'afh_destruct_d  = {lizzieLet17_5QNode_Int_7QNode_Int_1QNode_Int_d[50:35],
                                (lizzieLet17_5QNode_Int_7QNode_Int_1QNode_Int_d[0] && (! lizzieLet17_5QNode_Int_7QNode_Int_1QNode_Int_emitted[2]))};
  assign \t4'afi_destruct_d  = {lizzieLet17_5QNode_Int_7QNode_Int_1QNode_Int_d[66:51],
                                (lizzieLet17_5QNode_Int_7QNode_Int_1QNode_Int_d[0] && (! lizzieLet17_5QNode_Int_7QNode_Int_1QNode_Int_emitted[3]))};
  assign lizzieLet17_5QNode_Int_7QNode_Int_1QNode_Int_done = (lizzieLet17_5QNode_Int_7QNode_Int_1QNode_Int_emitted | ({\t4'afi_destruct_d [0],
                                                                                                                       \t3'afh_destruct_d [0],
                                                                                                                       \t2'afg_destruct_d [0],
                                                                                                                       \t1'aff_destruct_d [0]} & {\t4'afi_destruct_r ,
                                                                                                                                                  \t3'afh_destruct_r ,
                                                                                                                                                  \t2'afg_destruct_r ,
                                                                                                                                                  \t1'aff_destruct_r }));
  assign lizzieLet17_5QNode_Int_7QNode_Int_1QNode_Int_r = (& lizzieLet17_5QNode_Int_7QNode_Int_1QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNode_Int_1QNode_Int_emitted <= 4'd0;
    else
      lizzieLet17_5QNode_Int_7QNode_Int_1QNode_Int_emitted <= (lizzieLet17_5QNode_Int_7QNode_Int_1QNode_Int_r ? 4'd0 :
                                                               lizzieLet17_5QNode_Int_7QNode_Int_1QNode_Int_done);
  
  /* demux (Ty QTree_Int,
       Ty QTree_Int) : (lizzieLet17_5QNode_Int_7QNode_Int_2,QTree_Int) (lizzieLet17_5QNode_Int_7QNode_Int_1,QTree_Int) > [(_194,QTree_Int),
                                                                                                                          (_193,QTree_Int),
                                                                                                                          (lizzieLet17_5QNode_Int_7QNode_Int_1QNode_Int,QTree_Int),
                                                                                                                          (_192,QTree_Int)] */
  logic [3:0] lizzieLet17_5QNode_Int_7QNode_Int_1_onehotd;
  always_comb
    if ((lizzieLet17_5QNode_Int_7QNode_Int_2_d[0] && lizzieLet17_5QNode_Int_7QNode_Int_1_d[0]))
      unique case (lizzieLet17_5QNode_Int_7QNode_Int_2_d[2:1])
        2'd0: lizzieLet17_5QNode_Int_7QNode_Int_1_onehotd = 4'd1;
        2'd1: lizzieLet17_5QNode_Int_7QNode_Int_1_onehotd = 4'd2;
        2'd2: lizzieLet17_5QNode_Int_7QNode_Int_1_onehotd = 4'd4;
        2'd3: lizzieLet17_5QNode_Int_7QNode_Int_1_onehotd = 4'd8;
        default: lizzieLet17_5QNode_Int_7QNode_Int_1_onehotd = 4'd0;
      endcase
    else lizzieLet17_5QNode_Int_7QNode_Int_1_onehotd = 4'd0;
  assign _194_d = {lizzieLet17_5QNode_Int_7QNode_Int_1_d[66:1],
                   lizzieLet17_5QNode_Int_7QNode_Int_1_onehotd[0]};
  assign _193_d = {lizzieLet17_5QNode_Int_7QNode_Int_1_d[66:1],
                   lizzieLet17_5QNode_Int_7QNode_Int_1_onehotd[1]};
  assign lizzieLet17_5QNode_Int_7QNode_Int_1QNode_Int_d = {lizzieLet17_5QNode_Int_7QNode_Int_1_d[66:1],
                                                           lizzieLet17_5QNode_Int_7QNode_Int_1_onehotd[2]};
  assign _192_d = {lizzieLet17_5QNode_Int_7QNode_Int_1_d[66:1],
                   lizzieLet17_5QNode_Int_7QNode_Int_1_onehotd[3]};
  assign lizzieLet17_5QNode_Int_7QNode_Int_1_r = (| (lizzieLet17_5QNode_Int_7QNode_Int_1_onehotd & {_192_r,
                                                                                                    lizzieLet17_5QNode_Int_7QNode_Int_1QNode_Int_r,
                                                                                                    _193_r,
                                                                                                    _194_r}));
  assign lizzieLet17_5QNode_Int_7QNode_Int_2_r = lizzieLet17_5QNode_Int_7QNode_Int_1_r;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_QTree_Int) : (lizzieLet17_5QNode_Int_7QNode_Int_3,QTree_Int) (lizzieLet17_5QNode_Int_10QNode_Int,Pointer_QTree_Int) > [(lizzieLet17_5QNode_Int_7QNode_Int_3QNone_Int,Pointer_QTree_Int),
                                                                                                                                         (_191,Pointer_QTree_Int),
                                                                                                                                         (lizzieLet17_5QNode_Int_7QNode_Int_3QNode_Int,Pointer_QTree_Int),
                                                                                                                                         (_190,Pointer_QTree_Int)] */
  logic [3:0] lizzieLet17_5QNode_Int_10QNode_Int_onehotd;
  always_comb
    if ((lizzieLet17_5QNode_Int_7QNode_Int_3_d[0] && lizzieLet17_5QNode_Int_10QNode_Int_d[0]))
      unique case (lizzieLet17_5QNode_Int_7QNode_Int_3_d[2:1])
        2'd0: lizzieLet17_5QNode_Int_10QNode_Int_onehotd = 4'd1;
        2'd1: lizzieLet17_5QNode_Int_10QNode_Int_onehotd = 4'd2;
        2'd2: lizzieLet17_5QNode_Int_10QNode_Int_onehotd = 4'd4;
        2'd3: lizzieLet17_5QNode_Int_10QNode_Int_onehotd = 4'd8;
        default: lizzieLet17_5QNode_Int_10QNode_Int_onehotd = 4'd0;
      endcase
    else lizzieLet17_5QNode_Int_10QNode_Int_onehotd = 4'd0;
  assign lizzieLet17_5QNode_Int_7QNode_Int_3QNone_Int_d = {lizzieLet17_5QNode_Int_10QNode_Int_d[16:1],
                                                           lizzieLet17_5QNode_Int_10QNode_Int_onehotd[0]};
  assign _191_d = {lizzieLet17_5QNode_Int_10QNode_Int_d[16:1],
                   lizzieLet17_5QNode_Int_10QNode_Int_onehotd[1]};
  assign lizzieLet17_5QNode_Int_7QNode_Int_3QNode_Int_d = {lizzieLet17_5QNode_Int_10QNode_Int_d[16:1],
                                                           lizzieLet17_5QNode_Int_10QNode_Int_onehotd[2]};
  assign _190_d = {lizzieLet17_5QNode_Int_10QNode_Int_d[16:1],
                   lizzieLet17_5QNode_Int_10QNode_Int_onehotd[3]};
  assign lizzieLet17_5QNode_Int_10QNode_Int_r = (| (lizzieLet17_5QNode_Int_10QNode_Int_onehotd & {_190_r,
                                                                                                  lizzieLet17_5QNode_Int_7QNode_Int_3QNode_Int_r,
                                                                                                  _191_r,
                                                                                                  lizzieLet17_5QNode_Int_7QNode_Int_3QNone_Int_r}));
  assign lizzieLet17_5QNode_Int_7QNode_Int_3_r = lizzieLet17_5QNode_Int_10QNode_Int_r;
  
  /* buf (Ty Pointer_QTree_Int) : (lizzieLet17_5QNode_Int_7QNode_Int_3QNone_Int,Pointer_QTree_Int) > (lizzieLet17_5QNode_Int_7QNode_Int_3QNone_Int_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t lizzieLet17_5QNode_Int_7QNode_Int_3QNone_Int_bufchan_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_3QNone_Int_bufchan_r;
  assign lizzieLet17_5QNode_Int_7QNode_Int_3QNone_Int_r = ((! lizzieLet17_5QNode_Int_7QNode_Int_3QNone_Int_bufchan_d[0]) || lizzieLet17_5QNode_Int_7QNode_Int_3QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNode_Int_3QNone_Int_bufchan_d <= {16'd0,
                                                                 1'd0};
    else
      if (lizzieLet17_5QNode_Int_7QNode_Int_3QNone_Int_r)
        lizzieLet17_5QNode_Int_7QNode_Int_3QNone_Int_bufchan_d <= lizzieLet17_5QNode_Int_7QNode_Int_3QNone_Int_d;
  Pointer_QTree_Int_t lizzieLet17_5QNode_Int_7QNode_Int_3QNone_Int_bufchan_buf;
  assign lizzieLet17_5QNode_Int_7QNode_Int_3QNone_Int_bufchan_r = (! lizzieLet17_5QNode_Int_7QNode_Int_3QNone_Int_bufchan_buf[0]);
  assign lizzieLet17_5QNode_Int_7QNode_Int_3QNone_Int_1_argbuf_d = (lizzieLet17_5QNode_Int_7QNode_Int_3QNone_Int_bufchan_buf[0] ? lizzieLet17_5QNode_Int_7QNode_Int_3QNone_Int_bufchan_buf :
                                                                    lizzieLet17_5QNode_Int_7QNode_Int_3QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNode_Int_3QNone_Int_bufchan_buf <= {16'd0,
                                                                   1'd0};
    else
      if ((lizzieLet17_5QNode_Int_7QNode_Int_3QNone_Int_1_argbuf_r && lizzieLet17_5QNode_Int_7QNode_Int_3QNone_Int_bufchan_buf[0]))
        lizzieLet17_5QNode_Int_7QNode_Int_3QNone_Int_bufchan_buf <= {16'd0,
                                                                     1'd0};
      else if (((! lizzieLet17_5QNode_Int_7QNode_Int_3QNone_Int_1_argbuf_r) && (! lizzieLet17_5QNode_Int_7QNode_Int_3QNone_Int_bufchan_buf[0])))
        lizzieLet17_5QNode_Int_7QNode_Int_3QNone_Int_bufchan_buf <= lizzieLet17_5QNode_Int_7QNode_Int_3QNone_Int_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_QTree_Int) : (lizzieLet17_5QNode_Int_7QNode_Int_4,QTree_Int) (lizzieLet17_5QNode_Int_11QNode_Int,Pointer_QTree_Int) > [(lizzieLet17_5QNode_Int_7QNode_Int_4QNone_Int,Pointer_QTree_Int),
                                                                                                                                         (_189,Pointer_QTree_Int),
                                                                                                                                         (lizzieLet17_5QNode_Int_7QNode_Int_4QNode_Int,Pointer_QTree_Int),
                                                                                                                                         (_188,Pointer_QTree_Int)] */
  logic [3:0] lizzieLet17_5QNode_Int_11QNode_Int_onehotd;
  always_comb
    if ((lizzieLet17_5QNode_Int_7QNode_Int_4_d[0] && lizzieLet17_5QNode_Int_11QNode_Int_d[0]))
      unique case (lizzieLet17_5QNode_Int_7QNode_Int_4_d[2:1])
        2'd0: lizzieLet17_5QNode_Int_11QNode_Int_onehotd = 4'd1;
        2'd1: lizzieLet17_5QNode_Int_11QNode_Int_onehotd = 4'd2;
        2'd2: lizzieLet17_5QNode_Int_11QNode_Int_onehotd = 4'd4;
        2'd3: lizzieLet17_5QNode_Int_11QNode_Int_onehotd = 4'd8;
        default: lizzieLet17_5QNode_Int_11QNode_Int_onehotd = 4'd0;
      endcase
    else lizzieLet17_5QNode_Int_11QNode_Int_onehotd = 4'd0;
  assign lizzieLet17_5QNode_Int_7QNode_Int_4QNone_Int_d = {lizzieLet17_5QNode_Int_11QNode_Int_d[16:1],
                                                           lizzieLet17_5QNode_Int_11QNode_Int_onehotd[0]};
  assign _189_d = {lizzieLet17_5QNode_Int_11QNode_Int_d[16:1],
                   lizzieLet17_5QNode_Int_11QNode_Int_onehotd[1]};
  assign lizzieLet17_5QNode_Int_7QNode_Int_4QNode_Int_d = {lizzieLet17_5QNode_Int_11QNode_Int_d[16:1],
                                                           lizzieLet17_5QNode_Int_11QNode_Int_onehotd[2]};
  assign _188_d = {lizzieLet17_5QNode_Int_11QNode_Int_d[16:1],
                   lizzieLet17_5QNode_Int_11QNode_Int_onehotd[3]};
  assign lizzieLet17_5QNode_Int_11QNode_Int_r = (| (lizzieLet17_5QNode_Int_11QNode_Int_onehotd & {_188_r,
                                                                                                  lizzieLet17_5QNode_Int_7QNode_Int_4QNode_Int_r,
                                                                                                  _189_r,
                                                                                                  lizzieLet17_5QNode_Int_7QNode_Int_4QNone_Int_r}));
  assign lizzieLet17_5QNode_Int_7QNode_Int_4_r = lizzieLet17_5QNode_Int_11QNode_Int_r;
  
  /* buf (Ty Pointer_QTree_Int) : (lizzieLet17_5QNode_Int_7QNode_Int_4QNone_Int,Pointer_QTree_Int) > (lizzieLet17_5QNode_Int_7QNode_Int_4QNone_Int_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t lizzieLet17_5QNode_Int_7QNode_Int_4QNone_Int_bufchan_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_4QNone_Int_bufchan_r;
  assign lizzieLet17_5QNode_Int_7QNode_Int_4QNone_Int_r = ((! lizzieLet17_5QNode_Int_7QNode_Int_4QNone_Int_bufchan_d[0]) || lizzieLet17_5QNode_Int_7QNode_Int_4QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNode_Int_4QNone_Int_bufchan_d <= {16'd0,
                                                                 1'd0};
    else
      if (lizzieLet17_5QNode_Int_7QNode_Int_4QNone_Int_r)
        lizzieLet17_5QNode_Int_7QNode_Int_4QNone_Int_bufchan_d <= lizzieLet17_5QNode_Int_7QNode_Int_4QNone_Int_d;
  Pointer_QTree_Int_t lizzieLet17_5QNode_Int_7QNode_Int_4QNone_Int_bufchan_buf;
  assign lizzieLet17_5QNode_Int_7QNode_Int_4QNone_Int_bufchan_r = (! lizzieLet17_5QNode_Int_7QNode_Int_4QNone_Int_bufchan_buf[0]);
  assign lizzieLet17_5QNode_Int_7QNode_Int_4QNone_Int_1_argbuf_d = (lizzieLet17_5QNode_Int_7QNode_Int_4QNone_Int_bufchan_buf[0] ? lizzieLet17_5QNode_Int_7QNode_Int_4QNone_Int_bufchan_buf :
                                                                    lizzieLet17_5QNode_Int_7QNode_Int_4QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNode_Int_4QNone_Int_bufchan_buf <= {16'd0,
                                                                   1'd0};
    else
      if ((lizzieLet17_5QNode_Int_7QNode_Int_4QNone_Int_1_argbuf_r && lizzieLet17_5QNode_Int_7QNode_Int_4QNone_Int_bufchan_buf[0]))
        lizzieLet17_5QNode_Int_7QNode_Int_4QNone_Int_bufchan_buf <= {16'd0,
                                                                     1'd0};
      else if (((! lizzieLet17_5QNode_Int_7QNode_Int_4QNone_Int_1_argbuf_r) && (! lizzieLet17_5QNode_Int_7QNode_Int_4QNone_Int_bufchan_buf[0])))
        lizzieLet17_5QNode_Int_7QNode_Int_4QNone_Int_bufchan_buf <= lizzieLet17_5QNode_Int_7QNode_Int_4QNone_Int_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_QTree_Int) : (lizzieLet17_5QNode_Int_7QNode_Int_5,QTree_Int) (lizzieLet17_5QNode_Int_12QNode_Int,Pointer_QTree_Int) > [(lizzieLet17_5QNode_Int_7QNode_Int_5QNone_Int,Pointer_QTree_Int),
                                                                                                                                         (_187,Pointer_QTree_Int),
                                                                                                                                         (lizzieLet17_5QNode_Int_7QNode_Int_5QNode_Int,Pointer_QTree_Int),
                                                                                                                                         (_186,Pointer_QTree_Int)] */
  logic [3:0] lizzieLet17_5QNode_Int_12QNode_Int_onehotd;
  always_comb
    if ((lizzieLet17_5QNode_Int_7QNode_Int_5_d[0] && lizzieLet17_5QNode_Int_12QNode_Int_d[0]))
      unique case (lizzieLet17_5QNode_Int_7QNode_Int_5_d[2:1])
        2'd0: lizzieLet17_5QNode_Int_12QNode_Int_onehotd = 4'd1;
        2'd1: lizzieLet17_5QNode_Int_12QNode_Int_onehotd = 4'd2;
        2'd2: lizzieLet17_5QNode_Int_12QNode_Int_onehotd = 4'd4;
        2'd3: lizzieLet17_5QNode_Int_12QNode_Int_onehotd = 4'd8;
        default: lizzieLet17_5QNode_Int_12QNode_Int_onehotd = 4'd0;
      endcase
    else lizzieLet17_5QNode_Int_12QNode_Int_onehotd = 4'd0;
  assign lizzieLet17_5QNode_Int_7QNode_Int_5QNone_Int_d = {lizzieLet17_5QNode_Int_12QNode_Int_d[16:1],
                                                           lizzieLet17_5QNode_Int_12QNode_Int_onehotd[0]};
  assign _187_d = {lizzieLet17_5QNode_Int_12QNode_Int_d[16:1],
                   lizzieLet17_5QNode_Int_12QNode_Int_onehotd[1]};
  assign lizzieLet17_5QNode_Int_7QNode_Int_5QNode_Int_d = {lizzieLet17_5QNode_Int_12QNode_Int_d[16:1],
                                                           lizzieLet17_5QNode_Int_12QNode_Int_onehotd[2]};
  assign _186_d = {lizzieLet17_5QNode_Int_12QNode_Int_d[16:1],
                   lizzieLet17_5QNode_Int_12QNode_Int_onehotd[3]};
  assign lizzieLet17_5QNode_Int_12QNode_Int_r = (| (lizzieLet17_5QNode_Int_12QNode_Int_onehotd & {_186_r,
                                                                                                  lizzieLet17_5QNode_Int_7QNode_Int_5QNode_Int_r,
                                                                                                  _187_r,
                                                                                                  lizzieLet17_5QNode_Int_7QNode_Int_5QNone_Int_r}));
  assign lizzieLet17_5QNode_Int_7QNode_Int_5_r = lizzieLet17_5QNode_Int_12QNode_Int_r;
  
  /* buf (Ty Pointer_QTree_Int) : (lizzieLet17_5QNode_Int_7QNode_Int_5QNode_Int,Pointer_QTree_Int) > (lizzieLet17_5QNode_Int_7QNode_Int_5QNode_Int_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t lizzieLet17_5QNode_Int_7QNode_Int_5QNode_Int_bufchan_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_5QNode_Int_bufchan_r;
  assign lizzieLet17_5QNode_Int_7QNode_Int_5QNode_Int_r = ((! lizzieLet17_5QNode_Int_7QNode_Int_5QNode_Int_bufchan_d[0]) || lizzieLet17_5QNode_Int_7QNode_Int_5QNode_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNode_Int_5QNode_Int_bufchan_d <= {16'd0,
                                                                 1'd0};
    else
      if (lizzieLet17_5QNode_Int_7QNode_Int_5QNode_Int_r)
        lizzieLet17_5QNode_Int_7QNode_Int_5QNode_Int_bufchan_d <= lizzieLet17_5QNode_Int_7QNode_Int_5QNode_Int_d;
  Pointer_QTree_Int_t lizzieLet17_5QNode_Int_7QNode_Int_5QNode_Int_bufchan_buf;
  assign lizzieLet17_5QNode_Int_7QNode_Int_5QNode_Int_bufchan_r = (! lizzieLet17_5QNode_Int_7QNode_Int_5QNode_Int_bufchan_buf[0]);
  assign lizzieLet17_5QNode_Int_7QNode_Int_5QNode_Int_1_argbuf_d = (lizzieLet17_5QNode_Int_7QNode_Int_5QNode_Int_bufchan_buf[0] ? lizzieLet17_5QNode_Int_7QNode_Int_5QNode_Int_bufchan_buf :
                                                                    lizzieLet17_5QNode_Int_7QNode_Int_5QNode_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNode_Int_5QNode_Int_bufchan_buf <= {16'd0,
                                                                   1'd0};
    else
      if ((lizzieLet17_5QNode_Int_7QNode_Int_5QNode_Int_1_argbuf_r && lizzieLet17_5QNode_Int_7QNode_Int_5QNode_Int_bufchan_buf[0]))
        lizzieLet17_5QNode_Int_7QNode_Int_5QNode_Int_bufchan_buf <= {16'd0,
                                                                     1'd0};
      else if (((! lizzieLet17_5QNode_Int_7QNode_Int_5QNode_Int_1_argbuf_r) && (! lizzieLet17_5QNode_Int_7QNode_Int_5QNode_Int_bufchan_buf[0])))
        lizzieLet17_5QNode_Int_7QNode_Int_5QNode_Int_bufchan_buf <= lizzieLet17_5QNode_Int_7QNode_Int_5QNode_Int_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (lizzieLet17_5QNode_Int_7QNode_Int_5QNone_Int,Pointer_QTree_Int) > (lizzieLet17_5QNode_Int_7QNode_Int_5QNone_Int_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t lizzieLet17_5QNode_Int_7QNode_Int_5QNone_Int_bufchan_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_5QNone_Int_bufchan_r;
  assign lizzieLet17_5QNode_Int_7QNode_Int_5QNone_Int_r = ((! lizzieLet17_5QNode_Int_7QNode_Int_5QNone_Int_bufchan_d[0]) || lizzieLet17_5QNode_Int_7QNode_Int_5QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNode_Int_5QNone_Int_bufchan_d <= {16'd0,
                                                                 1'd0};
    else
      if (lizzieLet17_5QNode_Int_7QNode_Int_5QNone_Int_r)
        lizzieLet17_5QNode_Int_7QNode_Int_5QNone_Int_bufchan_d <= lizzieLet17_5QNode_Int_7QNode_Int_5QNone_Int_d;
  Pointer_QTree_Int_t lizzieLet17_5QNode_Int_7QNode_Int_5QNone_Int_bufchan_buf;
  assign lizzieLet17_5QNode_Int_7QNode_Int_5QNone_Int_bufchan_r = (! lizzieLet17_5QNode_Int_7QNode_Int_5QNone_Int_bufchan_buf[0]);
  assign lizzieLet17_5QNode_Int_7QNode_Int_5QNone_Int_1_argbuf_d = (lizzieLet17_5QNode_Int_7QNode_Int_5QNone_Int_bufchan_buf[0] ? lizzieLet17_5QNode_Int_7QNode_Int_5QNone_Int_bufchan_buf :
                                                                    lizzieLet17_5QNode_Int_7QNode_Int_5QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNode_Int_5QNone_Int_bufchan_buf <= {16'd0,
                                                                   1'd0};
    else
      if ((lizzieLet17_5QNode_Int_7QNode_Int_5QNone_Int_1_argbuf_r && lizzieLet17_5QNode_Int_7QNode_Int_5QNone_Int_bufchan_buf[0]))
        lizzieLet17_5QNode_Int_7QNode_Int_5QNone_Int_bufchan_buf <= {16'd0,
                                                                     1'd0};
      else if (((! lizzieLet17_5QNode_Int_7QNode_Int_5QNone_Int_1_argbuf_r) && (! lizzieLet17_5QNode_Int_7QNode_Int_5QNone_Int_bufchan_buf[0])))
        lizzieLet17_5QNode_Int_7QNode_Int_5QNone_Int_bufchan_buf <= lizzieLet17_5QNode_Int_7QNode_Int_5QNone_Int_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty MyDTInt_Int_Int) : (lizzieLet17_5QNode_Int_7QNode_Int_6,QTree_Int) (lizzieLet17_5QNode_Int_3QNode_Int,MyDTInt_Int_Int) > [(lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int,MyDTInt_Int_Int),
                                                                                                                                    (_185,MyDTInt_Int_Int),
                                                                                                                                    (lizzieLet17_5QNode_Int_7QNode_Int_6QNode_Int,MyDTInt_Int_Int),
                                                                                                                                    (_184,MyDTInt_Int_Int)] */
  logic [3:0] lizzieLet17_5QNode_Int_3QNode_Int_onehotd;
  always_comb
    if ((lizzieLet17_5QNode_Int_7QNode_Int_6_d[0] && lizzieLet17_5QNode_Int_3QNode_Int_d[0]))
      unique case (lizzieLet17_5QNode_Int_7QNode_Int_6_d[2:1])
        2'd0: lizzieLet17_5QNode_Int_3QNode_Int_onehotd = 4'd1;
        2'd1: lizzieLet17_5QNode_Int_3QNode_Int_onehotd = 4'd2;
        2'd2: lizzieLet17_5QNode_Int_3QNode_Int_onehotd = 4'd4;
        2'd3: lizzieLet17_5QNode_Int_3QNode_Int_onehotd = 4'd8;
        default: lizzieLet17_5QNode_Int_3QNode_Int_onehotd = 4'd0;
      endcase
    else lizzieLet17_5QNode_Int_3QNode_Int_onehotd = 4'd0;
  assign lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_d = lizzieLet17_5QNode_Int_3QNode_Int_onehotd[0];
  assign _185_d = lizzieLet17_5QNode_Int_3QNode_Int_onehotd[1];
  assign lizzieLet17_5QNode_Int_7QNode_Int_6QNode_Int_d = lizzieLet17_5QNode_Int_3QNode_Int_onehotd[2];
  assign _184_d = lizzieLet17_5QNode_Int_3QNode_Int_onehotd[3];
  assign lizzieLet17_5QNode_Int_3QNode_Int_r = (| (lizzieLet17_5QNode_Int_3QNode_Int_onehotd & {_184_r,
                                                                                                lizzieLet17_5QNode_Int_7QNode_Int_6QNode_Int_r,
                                                                                                _185_r,
                                                                                                lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_r}));
  assign lizzieLet17_5QNode_Int_7QNode_Int_6_r = lizzieLet17_5QNode_Int_3QNode_Int_r;
  
  /* fork (Ty MyDTInt_Int_Int) : (lizzieLet17_5QNode_Int_7QNode_Int_6QNode_Int,MyDTInt_Int_Int) > [(lizzieLet17_5QNode_Int_7QNode_Int_6QNode_Int_1,MyDTInt_Int_Int),
                                                                                              (lizzieLet17_5QNode_Int_7QNode_Int_6QNode_Int_2,MyDTInt_Int_Int)] */
  logic [1:0] lizzieLet17_5QNode_Int_7QNode_Int_6QNode_Int_emitted;
  logic [1:0] lizzieLet17_5QNode_Int_7QNode_Int_6QNode_Int_done;
  assign lizzieLet17_5QNode_Int_7QNode_Int_6QNode_Int_1_d = (lizzieLet17_5QNode_Int_7QNode_Int_6QNode_Int_d[0] && (! lizzieLet17_5QNode_Int_7QNode_Int_6QNode_Int_emitted[0]));
  assign lizzieLet17_5QNode_Int_7QNode_Int_6QNode_Int_2_d = (lizzieLet17_5QNode_Int_7QNode_Int_6QNode_Int_d[0] && (! lizzieLet17_5QNode_Int_7QNode_Int_6QNode_Int_emitted[1]));
  assign lizzieLet17_5QNode_Int_7QNode_Int_6QNode_Int_done = (lizzieLet17_5QNode_Int_7QNode_Int_6QNode_Int_emitted | ({lizzieLet17_5QNode_Int_7QNode_Int_6QNode_Int_2_d[0],
                                                                                                                       lizzieLet17_5QNode_Int_7QNode_Int_6QNode_Int_1_d[0]} & {lizzieLet17_5QNode_Int_7QNode_Int_6QNode_Int_2_r,
                                                                                                                                                                               lizzieLet17_5QNode_Int_7QNode_Int_6QNode_Int_1_r}));
  assign lizzieLet17_5QNode_Int_7QNode_Int_6QNode_Int_r = (& lizzieLet17_5QNode_Int_7QNode_Int_6QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNode_Int_6QNode_Int_emitted <= 2'd0;
    else
      lizzieLet17_5QNode_Int_7QNode_Int_6QNode_Int_emitted <= (lizzieLet17_5QNode_Int_7QNode_Int_6QNode_Int_r ? 2'd0 :
                                                               lizzieLet17_5QNode_Int_7QNode_Int_6QNode_Int_done);
  
  /* buf (Ty MyDTInt_Int_Int) : (lizzieLet17_5QNode_Int_7QNode_Int_6QNode_Int_2,MyDTInt_Int_Int) > (lizzieLet17_5QNode_Int_7QNode_Int_6QNode_Int_2_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t lizzieLet17_5QNode_Int_7QNode_Int_6QNode_Int_2_bufchan_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_6QNode_Int_2_bufchan_r;
  assign lizzieLet17_5QNode_Int_7QNode_Int_6QNode_Int_2_r = ((! lizzieLet17_5QNode_Int_7QNode_Int_6QNode_Int_2_bufchan_d[0]) || lizzieLet17_5QNode_Int_7QNode_Int_6QNode_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNode_Int_6QNode_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet17_5QNode_Int_7QNode_Int_6QNode_Int_2_r)
        lizzieLet17_5QNode_Int_7QNode_Int_6QNode_Int_2_bufchan_d <= lizzieLet17_5QNode_Int_7QNode_Int_6QNode_Int_2_d;
  MyDTInt_Int_Int_t lizzieLet17_5QNode_Int_7QNode_Int_6QNode_Int_2_bufchan_buf;
  assign lizzieLet17_5QNode_Int_7QNode_Int_6QNode_Int_2_bufchan_r = (! lizzieLet17_5QNode_Int_7QNode_Int_6QNode_Int_2_bufchan_buf[0]);
  assign lizzieLet17_5QNode_Int_7QNode_Int_6QNode_Int_2_argbuf_d = (lizzieLet17_5QNode_Int_7QNode_Int_6QNode_Int_2_bufchan_buf[0] ? lizzieLet17_5QNode_Int_7QNode_Int_6QNode_Int_2_bufchan_buf :
                                                                    lizzieLet17_5QNode_Int_7QNode_Int_6QNode_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNode_Int_6QNode_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet17_5QNode_Int_7QNode_Int_6QNode_Int_2_argbuf_r && lizzieLet17_5QNode_Int_7QNode_Int_6QNode_Int_2_bufchan_buf[0]))
        lizzieLet17_5QNode_Int_7QNode_Int_6QNode_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet17_5QNode_Int_7QNode_Int_6QNode_Int_2_argbuf_r) && (! lizzieLet17_5QNode_Int_7QNode_Int_6QNode_Int_2_bufchan_buf[0])))
        lizzieLet17_5QNode_Int_7QNode_Int_6QNode_Int_2_bufchan_buf <= lizzieLet17_5QNode_Int_7QNode_Int_6QNode_Int_2_bufchan_d;
  
  /* fork (Ty MyDTInt_Int_Int) : (lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int,MyDTInt_Int_Int) > [(lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_1,MyDTInt_Int_Int),
                                                                                              (lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_2,MyDTInt_Int_Int),
                                                                                              (lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_3,MyDTInt_Int_Int),
                                                                                              (lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_4,MyDTInt_Int_Int)] */
  logic [3:0] lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_emitted;
  logic [3:0] lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_done;
  assign lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_1_d = (lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_d[0] && (! lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_emitted[0]));
  assign lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_2_d = (lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_d[0] && (! lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_emitted[1]));
  assign lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_3_d = (lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_d[0] && (! lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_emitted[2]));
  assign lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_4_d = (lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_d[0] && (! lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_emitted[3]));
  assign lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_done = (lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_emitted | ({lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_4_d[0],
                                                                                                                       lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_3_d[0],
                                                                                                                       lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_2_d[0],
                                                                                                                       lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_1_d[0]} & {lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_4_r,
                                                                                                                                                                               lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_3_r,
                                                                                                                                                                               lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_2_r,
                                                                                                                                                                               lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_1_r}));
  assign lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_r = (& lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_emitted <= 4'd0;
    else
      lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_emitted <= (lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_r ? 4'd0 :
                                                               lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_done);
  
  /* buf (Ty MyDTInt_Int_Int) : (lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_1,MyDTInt_Int_Int) > (lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_1_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_1_bufchan_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_1_bufchan_r;
  assign lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_1_r = ((! lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_1_bufchan_d[0]) || lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_1_bufchan_d <= 1'd0;
    else
      if (lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_1_r)
        lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_1_bufchan_d <= lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_1_d;
  MyDTInt_Int_Int_t lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_1_bufchan_buf;
  assign lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_1_bufchan_r = (! lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_1_bufchan_buf[0]);
  assign lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_1_argbuf_d = (lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_1_bufchan_buf[0] ? lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_1_bufchan_buf :
                                                                    lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_1_argbuf_r && lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_1_bufchan_buf[0]))
        lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_1_argbuf_r) && (! lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_1_bufchan_buf[0])))
        lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_1_bufchan_buf <= lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_1_bufchan_d;
  
  /* buf (Ty MyDTInt_Int_Int) : (lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_2,MyDTInt_Int_Int) > (lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_2_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_2_bufchan_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_2_bufchan_r;
  assign lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_2_r = ((! lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_2_bufchan_d[0]) || lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_2_r)
        lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_2_bufchan_d <= lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_2_d;
  MyDTInt_Int_Int_t lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_2_bufchan_buf;
  assign lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_2_bufchan_r = (! lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_2_bufchan_buf[0]);
  assign lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_2_argbuf_d = (lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_2_bufchan_buf[0] ? lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_2_bufchan_buf :
                                                                    lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_2_argbuf_r && lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_2_bufchan_buf[0]))
        lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_2_argbuf_r) && (! lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_2_bufchan_buf[0])))
        lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_2_bufchan_buf <= lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_2_bufchan_d;
  
  /* buf (Ty MyDTInt_Int_Int) : (lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_3,MyDTInt_Int_Int) > (lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_3_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_3_bufchan_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_3_bufchan_r;
  assign lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_3_r = ((! lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_3_bufchan_d[0]) || lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_3_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_3_bufchan_d <= 1'd0;
    else
      if (lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_3_r)
        lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_3_bufchan_d <= lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_3_d;
  MyDTInt_Int_Int_t lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_3_bufchan_buf;
  assign lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_3_bufchan_r = (! lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_3_bufchan_buf[0]);
  assign lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_3_argbuf_d = (lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_3_bufchan_buf[0] ? lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_3_bufchan_buf :
                                                                    lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_3_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_3_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_3_argbuf_r && lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_3_bufchan_buf[0]))
        lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_3_bufchan_buf <= 1'd0;
      else if (((! lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_3_argbuf_r) && (! lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_3_bufchan_buf[0])))
        lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_3_bufchan_buf <= lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_3_bufchan_d;
  
  /* buf (Ty MyDTInt_Int_Int) : (lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_4,MyDTInt_Int_Int) > (lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_4_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_4_bufchan_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_4_bufchan_r;
  assign lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_4_r = ((! lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_4_bufchan_d[0]) || lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_4_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_4_bufchan_d <= 1'd0;
    else
      if (lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_4_r)
        lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_4_bufchan_d <= lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_4_d;
  MyDTInt_Int_Int_t lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_4_bufchan_buf;
  assign lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_4_bufchan_r = (! lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_4_bufchan_buf[0]);
  assign lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_4_argbuf_d = (lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_4_bufchan_buf[0] ? lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_4_bufchan_buf :
                                                                    lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_4_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_4_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_4_argbuf_r && lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_4_bufchan_buf[0]))
        lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_4_bufchan_buf <= 1'd0;
      else if (((! lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_4_argbuf_r) && (! lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_4_bufchan_buf[0])))
        lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_4_bufchan_buf <= lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_4_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_CTf_f_Int) : (lizzieLet17_5QNode_Int_7QNode_Int_7,QTree_Int) (lizzieLet17_5QNode_Int_4QNode_Int,Pointer_CTf_f_Int) > [(lizzieLet17_5QNode_Int_7QNode_Int_7QNone_Int,Pointer_CTf_f_Int),
                                                                                                                                        (lizzieLet17_5QNode_Int_7QNode_Int_7QVal_Int,Pointer_CTf_f_Int),
                                                                                                                                        (lizzieLet17_5QNode_Int_7QNode_Int_7QNode_Int,Pointer_CTf_f_Int),
                                                                                                                                        (lizzieLet17_5QNode_Int_7QNode_Int_7QError_Int,Pointer_CTf_f_Int)] */
  logic [3:0] lizzieLet17_5QNode_Int_4QNode_Int_onehotd;
  always_comb
    if ((lizzieLet17_5QNode_Int_7QNode_Int_7_d[0] && lizzieLet17_5QNode_Int_4QNode_Int_d[0]))
      unique case (lizzieLet17_5QNode_Int_7QNode_Int_7_d[2:1])
        2'd0: lizzieLet17_5QNode_Int_4QNode_Int_onehotd = 4'd1;
        2'd1: lizzieLet17_5QNode_Int_4QNode_Int_onehotd = 4'd2;
        2'd2: lizzieLet17_5QNode_Int_4QNode_Int_onehotd = 4'd4;
        2'd3: lizzieLet17_5QNode_Int_4QNode_Int_onehotd = 4'd8;
        default: lizzieLet17_5QNode_Int_4QNode_Int_onehotd = 4'd0;
      endcase
    else lizzieLet17_5QNode_Int_4QNode_Int_onehotd = 4'd0;
  assign lizzieLet17_5QNode_Int_7QNode_Int_7QNone_Int_d = {lizzieLet17_5QNode_Int_4QNode_Int_d[16:1],
                                                           lizzieLet17_5QNode_Int_4QNode_Int_onehotd[0]};
  assign lizzieLet17_5QNode_Int_7QNode_Int_7QVal_Int_d = {lizzieLet17_5QNode_Int_4QNode_Int_d[16:1],
                                                          lizzieLet17_5QNode_Int_4QNode_Int_onehotd[1]};
  assign lizzieLet17_5QNode_Int_7QNode_Int_7QNode_Int_d = {lizzieLet17_5QNode_Int_4QNode_Int_d[16:1],
                                                           lizzieLet17_5QNode_Int_4QNode_Int_onehotd[2]};
  assign lizzieLet17_5QNode_Int_7QNode_Int_7QError_Int_d = {lizzieLet17_5QNode_Int_4QNode_Int_d[16:1],
                                                            lizzieLet17_5QNode_Int_4QNode_Int_onehotd[3]};
  assign lizzieLet17_5QNode_Int_4QNode_Int_r = (| (lizzieLet17_5QNode_Int_4QNode_Int_onehotd & {lizzieLet17_5QNode_Int_7QNode_Int_7QError_Int_r,
                                                                                                lizzieLet17_5QNode_Int_7QNode_Int_7QNode_Int_r,
                                                                                                lizzieLet17_5QNode_Int_7QNode_Int_7QVal_Int_r,
                                                                                                lizzieLet17_5QNode_Int_7QNode_Int_7QNone_Int_r}));
  assign lizzieLet17_5QNode_Int_7QNode_Int_7_r = lizzieLet17_5QNode_Int_4QNode_Int_r;
  
  /* buf (Ty Pointer_CTf_f_Int) : (lizzieLet17_5QNode_Int_7QNode_Int_7QError_Int,Pointer_CTf_f_Int) > (lizzieLet17_5QNode_Int_7QNode_Int_7QError_Int_1_argbuf,Pointer_CTf_f_Int) */
  Pointer_CTf_f_Int_t lizzieLet17_5QNode_Int_7QNode_Int_7QError_Int_bufchan_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_7QError_Int_bufchan_r;
  assign lizzieLet17_5QNode_Int_7QNode_Int_7QError_Int_r = ((! lizzieLet17_5QNode_Int_7QNode_Int_7QError_Int_bufchan_d[0]) || lizzieLet17_5QNode_Int_7QNode_Int_7QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNode_Int_7QError_Int_bufchan_d <= {16'd0,
                                                                  1'd0};
    else
      if (lizzieLet17_5QNode_Int_7QNode_Int_7QError_Int_r)
        lizzieLet17_5QNode_Int_7QNode_Int_7QError_Int_bufchan_d <= lizzieLet17_5QNode_Int_7QNode_Int_7QError_Int_d;
  Pointer_CTf_f_Int_t lizzieLet17_5QNode_Int_7QNode_Int_7QError_Int_bufchan_buf;
  assign lizzieLet17_5QNode_Int_7QNode_Int_7QError_Int_bufchan_r = (! lizzieLet17_5QNode_Int_7QNode_Int_7QError_Int_bufchan_buf[0]);
  assign lizzieLet17_5QNode_Int_7QNode_Int_7QError_Int_1_argbuf_d = (lizzieLet17_5QNode_Int_7QNode_Int_7QError_Int_bufchan_buf[0] ? lizzieLet17_5QNode_Int_7QNode_Int_7QError_Int_bufchan_buf :
                                                                     lizzieLet17_5QNode_Int_7QNode_Int_7QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNode_Int_7QError_Int_bufchan_buf <= {16'd0,
                                                                    1'd0};
    else
      if ((lizzieLet17_5QNode_Int_7QNode_Int_7QError_Int_1_argbuf_r && lizzieLet17_5QNode_Int_7QNode_Int_7QError_Int_bufchan_buf[0]))
        lizzieLet17_5QNode_Int_7QNode_Int_7QError_Int_bufchan_buf <= {16'd0,
                                                                      1'd0};
      else if (((! lizzieLet17_5QNode_Int_7QNode_Int_7QError_Int_1_argbuf_r) && (! lizzieLet17_5QNode_Int_7QNode_Int_7QError_Int_bufchan_buf[0])))
        lizzieLet17_5QNode_Int_7QNode_Int_7QError_Int_bufchan_buf <= lizzieLet17_5QNode_Int_7QNode_Int_7QError_Int_bufchan_d;
  
  /* dcon (Ty CTf_f_Int,
      Dcon Lcall_f_f_Int3) : [(lizzieLet17_5QNode_Int_7QNode_Int_7QNode_Int,Pointer_CTf_f_Int),
                              (lizzieLet17_5QNode_Int_7QNode_Int_10QNode_Int,Pointer_QTree_Int),
                              (lizzieLet17_5QNode_Int_7QNode_Int_11QNode_Int,Pointer_QTree_Int),
                              (t1'aff_destruct,Pointer_QTree_Int),
                              (lizzieLet17_5QNode_Int_7QNode_Int_9QNode_Int_1,MyDTInt_Bool),
                              (lizzieLet17_5QNode_Int_7QNode_Int_6QNode_Int_1,MyDTInt_Int_Int),
                              (lizzieLet17_5QNode_Int_7QNode_Int_3QNode_Int,Pointer_QTree_Int),
                              (lizzieLet17_5QNode_Int_7QNode_Int_12QNode_Int,Pointer_QTree_Int),
                              (t2'afg_destruct,Pointer_QTree_Int),
                              (lizzieLet17_5QNode_Int_7QNode_Int_4QNode_Int,Pointer_QTree_Int),
                              (lizzieLet17_5QNode_Int_7QNode_Int_13QNode_Int,Pointer_QTree_Int),
                              (t3'afh_destruct,Pointer_QTree_Int)] > (lizzieLet17_5QNode_Int_7QNode_Int_7QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_10QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_11QNode_Int_1t1'aff_1lizzieLet17_5QNode_Int_7QNode_Int_9QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_6QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_3QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_12QNode_Int_1t2'afg_1lizzieLet17_5QNode_Int_7QNode_Int_4QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_13QNode_Int_1t3'afh_1Lcall_f_f_Int3,CTf_f_Int) */
  assign \lizzieLet17_5QNode_Int_7QNode_Int_7QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_10QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_11QNode_Int_1t1'aff_1lizzieLet17_5QNode_Int_7QNode_Int_9QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_6QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_3QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_12QNode_Int_1t2'afg_1lizzieLet17_5QNode_Int_7QNode_Int_4QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_13QNode_Int_1t3'afh_1Lcall_f_f_Int3_d  = Lcall_f_f_Int3_dc((& {lizzieLet17_5QNode_Int_7QNode_Int_7QNode_Int_d[0],
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              lizzieLet17_5QNode_Int_7QNode_Int_10QNode_Int_d[0],
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              lizzieLet17_5QNode_Int_7QNode_Int_11QNode_Int_d[0],
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              \t1'aff_destruct_d [0],
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              lizzieLet17_5QNode_Int_7QNode_Int_9QNode_Int_1_d[0],
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              lizzieLet17_5QNode_Int_7QNode_Int_6QNode_Int_1_d[0],
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              lizzieLet17_5QNode_Int_7QNode_Int_3QNode_Int_d[0],
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              lizzieLet17_5QNode_Int_7QNode_Int_12QNode_Int_d[0],
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              \t2'afg_destruct_d [0],
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              lizzieLet17_5QNode_Int_7QNode_Int_4QNode_Int_d[0],
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              lizzieLet17_5QNode_Int_7QNode_Int_13QNode_Int_d[0],
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              \t3'afh_destruct_d [0]}), lizzieLet17_5QNode_Int_7QNode_Int_7QNode_Int_d, lizzieLet17_5QNode_Int_7QNode_Int_10QNode_Int_d, lizzieLet17_5QNode_Int_7QNode_Int_11QNode_Int_d, \t1'aff_destruct_d , lizzieLet17_5QNode_Int_7QNode_Int_9QNode_Int_1_d, lizzieLet17_5QNode_Int_7QNode_Int_6QNode_Int_1_d, lizzieLet17_5QNode_Int_7QNode_Int_3QNode_Int_d, lizzieLet17_5QNode_Int_7QNode_Int_12QNode_Int_d, \t2'afg_destruct_d , lizzieLet17_5QNode_Int_7QNode_Int_4QNode_Int_d, lizzieLet17_5QNode_Int_7QNode_Int_13QNode_Int_d, \t3'afh_destruct_d );
  assign {lizzieLet17_5QNode_Int_7QNode_Int_7QNode_Int_r,
          lizzieLet17_5QNode_Int_7QNode_Int_10QNode_Int_r,
          lizzieLet17_5QNode_Int_7QNode_Int_11QNode_Int_r,
          \t1'aff_destruct_r ,
          lizzieLet17_5QNode_Int_7QNode_Int_9QNode_Int_1_r,
          lizzieLet17_5QNode_Int_7QNode_Int_6QNode_Int_1_r,
          lizzieLet17_5QNode_Int_7QNode_Int_3QNode_Int_r,
          lizzieLet17_5QNode_Int_7QNode_Int_12QNode_Int_r,
          \t2'afg_destruct_r ,
          lizzieLet17_5QNode_Int_7QNode_Int_4QNode_Int_r,
          lizzieLet17_5QNode_Int_7QNode_Int_13QNode_Int_r,
          \t3'afh_destruct_r } = {12 {(\lizzieLet17_5QNode_Int_7QNode_Int_7QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_10QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_11QNode_Int_1t1'aff_1lizzieLet17_5QNode_Int_7QNode_Int_9QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_6QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_3QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_12QNode_Int_1t2'afg_1lizzieLet17_5QNode_Int_7QNode_Int_4QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_13QNode_Int_1t3'afh_1Lcall_f_f_Int3_r  && \lizzieLet17_5QNode_Int_7QNode_Int_7QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_10QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_11QNode_Int_1t1'aff_1lizzieLet17_5QNode_Int_7QNode_Int_9QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_6QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_3QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_12QNode_Int_1t2'afg_1lizzieLet17_5QNode_Int_7QNode_Int_4QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_13QNode_Int_1t3'afh_1Lcall_f_f_Int3_d [0])}};
  
  /* buf (Ty CTf_f_Int) : (lizzieLet17_5QNode_Int_7QNode_Int_7QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_10QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_11QNode_Int_1t1'aff_1lizzieLet17_5QNode_Int_7QNode_Int_9QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_6QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_3QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_12QNode_Int_1t2'afg_1lizzieLet17_5QNode_Int_7QNode_Int_4QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_13QNode_Int_1t3'afh_1Lcall_f_f_Int3,CTf_f_Int) > (lizzieLet52_1_argbuf,CTf_f_Int) */
  CTf_f_Int_t \lizzieLet17_5QNode_Int_7QNode_Int_7QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_10QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_11QNode_Int_1t1'aff_1lizzieLet17_5QNode_Int_7QNode_Int_9QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_6QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_3QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_12QNode_Int_1t2'afg_1lizzieLet17_5QNode_Int_7QNode_Int_4QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_13QNode_Int_1t3'afh_1Lcall_f_f_Int3_bufchan_d ;
  logic \lizzieLet17_5QNode_Int_7QNode_Int_7QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_10QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_11QNode_Int_1t1'aff_1lizzieLet17_5QNode_Int_7QNode_Int_9QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_6QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_3QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_12QNode_Int_1t2'afg_1lizzieLet17_5QNode_Int_7QNode_Int_4QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_13QNode_Int_1t3'afh_1Lcall_f_f_Int3_bufchan_r ;
  assign \lizzieLet17_5QNode_Int_7QNode_Int_7QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_10QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_11QNode_Int_1t1'aff_1lizzieLet17_5QNode_Int_7QNode_Int_9QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_6QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_3QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_12QNode_Int_1t2'afg_1lizzieLet17_5QNode_Int_7QNode_Int_4QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_13QNode_Int_1t3'afh_1Lcall_f_f_Int3_r  = ((! \lizzieLet17_5QNode_Int_7QNode_Int_7QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_10QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_11QNode_Int_1t1'aff_1lizzieLet17_5QNode_Int_7QNode_Int_9QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_6QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_3QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_12QNode_Int_1t2'afg_1lizzieLet17_5QNode_Int_7QNode_Int_4QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_13QNode_Int_1t3'afh_1Lcall_f_f_Int3_bufchan_d [0]) || \lizzieLet17_5QNode_Int_7QNode_Int_7QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_10QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_11QNode_Int_1t1'aff_1lizzieLet17_5QNode_Int_7QNode_Int_9QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_6QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_3QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_12QNode_Int_1t2'afg_1lizzieLet17_5QNode_Int_7QNode_Int_4QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_13QNode_Int_1t3'afh_1Lcall_f_f_Int3_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet17_5QNode_Int_7QNode_Int_7QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_10QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_11QNode_Int_1t1'aff_1lizzieLet17_5QNode_Int_7QNode_Int_9QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_6QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_3QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_12QNode_Int_1t2'afg_1lizzieLet17_5QNode_Int_7QNode_Int_4QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_13QNode_Int_1t3'afh_1Lcall_f_f_Int3_bufchan_d  <= {163'd0,
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               1'd0};
    else
      if (\lizzieLet17_5QNode_Int_7QNode_Int_7QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_10QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_11QNode_Int_1t1'aff_1lizzieLet17_5QNode_Int_7QNode_Int_9QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_6QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_3QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_12QNode_Int_1t2'afg_1lizzieLet17_5QNode_Int_7QNode_Int_4QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_13QNode_Int_1t3'afh_1Lcall_f_f_Int3_r )
        \lizzieLet17_5QNode_Int_7QNode_Int_7QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_10QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_11QNode_Int_1t1'aff_1lizzieLet17_5QNode_Int_7QNode_Int_9QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_6QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_3QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_12QNode_Int_1t2'afg_1lizzieLet17_5QNode_Int_7QNode_Int_4QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_13QNode_Int_1t3'afh_1Lcall_f_f_Int3_bufchan_d  <= \lizzieLet17_5QNode_Int_7QNode_Int_7QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_10QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_11QNode_Int_1t1'aff_1lizzieLet17_5QNode_Int_7QNode_Int_9QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_6QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_3QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_12QNode_Int_1t2'afg_1lizzieLet17_5QNode_Int_7QNode_Int_4QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_13QNode_Int_1t3'afh_1Lcall_f_f_Int3_d ;
  CTf_f_Int_t \lizzieLet17_5QNode_Int_7QNode_Int_7QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_10QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_11QNode_Int_1t1'aff_1lizzieLet17_5QNode_Int_7QNode_Int_9QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_6QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_3QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_12QNode_Int_1t2'afg_1lizzieLet17_5QNode_Int_7QNode_Int_4QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_13QNode_Int_1t3'afh_1Lcall_f_f_Int3_bufchan_buf ;
  assign \lizzieLet17_5QNode_Int_7QNode_Int_7QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_10QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_11QNode_Int_1t1'aff_1lizzieLet17_5QNode_Int_7QNode_Int_9QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_6QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_3QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_12QNode_Int_1t2'afg_1lizzieLet17_5QNode_Int_7QNode_Int_4QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_13QNode_Int_1t3'afh_1Lcall_f_f_Int3_bufchan_r  = (! \lizzieLet17_5QNode_Int_7QNode_Int_7QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_10QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_11QNode_Int_1t1'aff_1lizzieLet17_5QNode_Int_7QNode_Int_9QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_6QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_3QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_12QNode_Int_1t2'afg_1lizzieLet17_5QNode_Int_7QNode_Int_4QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_13QNode_Int_1t3'afh_1Lcall_f_f_Int3_bufchan_buf [0]);
  assign lizzieLet52_1_argbuf_d = (\lizzieLet17_5QNode_Int_7QNode_Int_7QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_10QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_11QNode_Int_1t1'aff_1lizzieLet17_5QNode_Int_7QNode_Int_9QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_6QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_3QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_12QNode_Int_1t2'afg_1lizzieLet17_5QNode_Int_7QNode_Int_4QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_13QNode_Int_1t3'afh_1Lcall_f_f_Int3_bufchan_buf [0] ? \lizzieLet17_5QNode_Int_7QNode_Int_7QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_10QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_11QNode_Int_1t1'aff_1lizzieLet17_5QNode_Int_7QNode_Int_9QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_6QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_3QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_12QNode_Int_1t2'afg_1lizzieLet17_5QNode_Int_7QNode_Int_4QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_13QNode_Int_1t3'afh_1Lcall_f_f_Int3_bufchan_buf  :
                                   \lizzieLet17_5QNode_Int_7QNode_Int_7QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_10QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_11QNode_Int_1t1'aff_1lizzieLet17_5QNode_Int_7QNode_Int_9QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_6QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_3QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_12QNode_Int_1t2'afg_1lizzieLet17_5QNode_Int_7QNode_Int_4QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_13QNode_Int_1t3'afh_1Lcall_f_f_Int3_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet17_5QNode_Int_7QNode_Int_7QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_10QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_11QNode_Int_1t1'aff_1lizzieLet17_5QNode_Int_7QNode_Int_9QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_6QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_3QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_12QNode_Int_1t2'afg_1lizzieLet17_5QNode_Int_7QNode_Int_4QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_13QNode_Int_1t3'afh_1Lcall_f_f_Int3_bufchan_buf  <= {163'd0,
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 1'd0};
    else
      if ((lizzieLet52_1_argbuf_r && \lizzieLet17_5QNode_Int_7QNode_Int_7QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_10QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_11QNode_Int_1t1'aff_1lizzieLet17_5QNode_Int_7QNode_Int_9QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_6QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_3QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_12QNode_Int_1t2'afg_1lizzieLet17_5QNode_Int_7QNode_Int_4QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_13QNode_Int_1t3'afh_1Lcall_f_f_Int3_bufchan_buf [0]))
        \lizzieLet17_5QNode_Int_7QNode_Int_7QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_10QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_11QNode_Int_1t1'aff_1lizzieLet17_5QNode_Int_7QNode_Int_9QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_6QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_3QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_12QNode_Int_1t2'afg_1lizzieLet17_5QNode_Int_7QNode_Int_4QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_13QNode_Int_1t3'afh_1Lcall_f_f_Int3_bufchan_buf  <= {163'd0,
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   1'd0};
      else if (((! lizzieLet52_1_argbuf_r) && (! \lizzieLet17_5QNode_Int_7QNode_Int_7QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_10QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_11QNode_Int_1t1'aff_1lizzieLet17_5QNode_Int_7QNode_Int_9QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_6QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_3QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_12QNode_Int_1t2'afg_1lizzieLet17_5QNode_Int_7QNode_Int_4QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_13QNode_Int_1t3'afh_1Lcall_f_f_Int3_bufchan_buf [0])))
        \lizzieLet17_5QNode_Int_7QNode_Int_7QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_10QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_11QNode_Int_1t1'aff_1lizzieLet17_5QNode_Int_7QNode_Int_9QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_6QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_3QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_12QNode_Int_1t2'afg_1lizzieLet17_5QNode_Int_7QNode_Int_4QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_13QNode_Int_1t3'afh_1Lcall_f_f_Int3_bufchan_buf  <= \lizzieLet17_5QNode_Int_7QNode_Int_7QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_10QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_11QNode_Int_1t1'aff_1lizzieLet17_5QNode_Int_7QNode_Int_9QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_6QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_3QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_12QNode_Int_1t2'afg_1lizzieLet17_5QNode_Int_7QNode_Int_4QNode_Int_1lizzieLet17_5QNode_Int_7QNode_Int_13QNode_Int_1t3'afh_1Lcall_f_f_Int3_bufchan_d ;
  
  /* buf (Ty Pointer_CTf_f_Int) : (lizzieLet17_5QNode_Int_7QNode_Int_7QNone_Int,Pointer_CTf_f_Int) > (lizzieLet17_5QNode_Int_7QNode_Int_7QNone_Int_1_argbuf,Pointer_CTf_f_Int) */
  Pointer_CTf_f_Int_t lizzieLet17_5QNode_Int_7QNode_Int_7QNone_Int_bufchan_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_7QNone_Int_bufchan_r;
  assign lizzieLet17_5QNode_Int_7QNode_Int_7QNone_Int_r = ((! lizzieLet17_5QNode_Int_7QNode_Int_7QNone_Int_bufchan_d[0]) || lizzieLet17_5QNode_Int_7QNode_Int_7QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNode_Int_7QNone_Int_bufchan_d <= {16'd0,
                                                                 1'd0};
    else
      if (lizzieLet17_5QNode_Int_7QNode_Int_7QNone_Int_r)
        lizzieLet17_5QNode_Int_7QNode_Int_7QNone_Int_bufchan_d <= lizzieLet17_5QNode_Int_7QNode_Int_7QNone_Int_d;
  Pointer_CTf_f_Int_t lizzieLet17_5QNode_Int_7QNode_Int_7QNone_Int_bufchan_buf;
  assign lizzieLet17_5QNode_Int_7QNode_Int_7QNone_Int_bufchan_r = (! lizzieLet17_5QNode_Int_7QNode_Int_7QNone_Int_bufchan_buf[0]);
  assign lizzieLet17_5QNode_Int_7QNode_Int_7QNone_Int_1_argbuf_d = (lizzieLet17_5QNode_Int_7QNode_Int_7QNone_Int_bufchan_buf[0] ? lizzieLet17_5QNode_Int_7QNode_Int_7QNone_Int_bufchan_buf :
                                                                    lizzieLet17_5QNode_Int_7QNode_Int_7QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNode_Int_7QNone_Int_bufchan_buf <= {16'd0,
                                                                   1'd0};
    else
      if ((lizzieLet17_5QNode_Int_7QNode_Int_7QNone_Int_1_argbuf_r && lizzieLet17_5QNode_Int_7QNode_Int_7QNone_Int_bufchan_buf[0]))
        lizzieLet17_5QNode_Int_7QNode_Int_7QNone_Int_bufchan_buf <= {16'd0,
                                                                     1'd0};
      else if (((! lizzieLet17_5QNode_Int_7QNode_Int_7QNone_Int_1_argbuf_r) && (! lizzieLet17_5QNode_Int_7QNode_Int_7QNone_Int_bufchan_buf[0])))
        lizzieLet17_5QNode_Int_7QNode_Int_7QNone_Int_bufchan_buf <= lizzieLet17_5QNode_Int_7QNode_Int_7QNone_Int_bufchan_d;
  
  /* buf (Ty Pointer_CTf_f_Int) : (lizzieLet17_5QNode_Int_7QNode_Int_7QVal_Int,Pointer_CTf_f_Int) > (lizzieLet17_5QNode_Int_7QNode_Int_7QVal_Int_1_argbuf,Pointer_CTf_f_Int) */
  Pointer_CTf_f_Int_t lizzieLet17_5QNode_Int_7QNode_Int_7QVal_Int_bufchan_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_7QVal_Int_bufchan_r;
  assign lizzieLet17_5QNode_Int_7QNode_Int_7QVal_Int_r = ((! lizzieLet17_5QNode_Int_7QNode_Int_7QVal_Int_bufchan_d[0]) || lizzieLet17_5QNode_Int_7QNode_Int_7QVal_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNode_Int_7QVal_Int_bufchan_d <= {16'd0,
                                                                1'd0};
    else
      if (lizzieLet17_5QNode_Int_7QNode_Int_7QVal_Int_r)
        lizzieLet17_5QNode_Int_7QNode_Int_7QVal_Int_bufchan_d <= lizzieLet17_5QNode_Int_7QNode_Int_7QVal_Int_d;
  Pointer_CTf_f_Int_t lizzieLet17_5QNode_Int_7QNode_Int_7QVal_Int_bufchan_buf;
  assign lizzieLet17_5QNode_Int_7QNode_Int_7QVal_Int_bufchan_r = (! lizzieLet17_5QNode_Int_7QNode_Int_7QVal_Int_bufchan_buf[0]);
  assign lizzieLet17_5QNode_Int_7QNode_Int_7QVal_Int_1_argbuf_d = (lizzieLet17_5QNode_Int_7QNode_Int_7QVal_Int_bufchan_buf[0] ? lizzieLet17_5QNode_Int_7QNode_Int_7QVal_Int_bufchan_buf :
                                                                   lizzieLet17_5QNode_Int_7QNode_Int_7QVal_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNode_Int_7QVal_Int_bufchan_buf <= {16'd0,
                                                                  1'd0};
    else
      if ((lizzieLet17_5QNode_Int_7QNode_Int_7QVal_Int_1_argbuf_r && lizzieLet17_5QNode_Int_7QNode_Int_7QVal_Int_bufchan_buf[0]))
        lizzieLet17_5QNode_Int_7QNode_Int_7QVal_Int_bufchan_buf <= {16'd0,
                                                                    1'd0};
      else if (((! lizzieLet17_5QNode_Int_7QNode_Int_7QVal_Int_1_argbuf_r) && (! lizzieLet17_5QNode_Int_7QNode_Int_7QVal_Int_bufchan_buf[0])))
        lizzieLet17_5QNode_Int_7QNode_Int_7QVal_Int_bufchan_buf <= lizzieLet17_5QNode_Int_7QNode_Int_7QVal_Int_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Go) : (lizzieLet17_5QNode_Int_7QNode_Int_8,QTree_Int) (lizzieLet17_5QNode_Int_5QNode_Int,Go) > [(lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int,Go),
                                                                                                          (lizzieLet17_5QNode_Int_7QNode_Int_8QVal_Int,Go),
                                                                                                          (lizzieLet17_5QNode_Int_7QNode_Int_8QNode_Int,Go),
                                                                                                          (lizzieLet17_5QNode_Int_7QNode_Int_8QError_Int,Go)] */
  logic [3:0] lizzieLet17_5QNode_Int_5QNode_Int_onehotd;
  always_comb
    if ((lizzieLet17_5QNode_Int_7QNode_Int_8_d[0] && lizzieLet17_5QNode_Int_5QNode_Int_d[0]))
      unique case (lizzieLet17_5QNode_Int_7QNode_Int_8_d[2:1])
        2'd0: lizzieLet17_5QNode_Int_5QNode_Int_onehotd = 4'd1;
        2'd1: lizzieLet17_5QNode_Int_5QNode_Int_onehotd = 4'd2;
        2'd2: lizzieLet17_5QNode_Int_5QNode_Int_onehotd = 4'd4;
        2'd3: lizzieLet17_5QNode_Int_5QNode_Int_onehotd = 4'd8;
        default: lizzieLet17_5QNode_Int_5QNode_Int_onehotd = 4'd0;
      endcase
    else lizzieLet17_5QNode_Int_5QNode_Int_onehotd = 4'd0;
  assign lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_d = lizzieLet17_5QNode_Int_5QNode_Int_onehotd[0];
  assign lizzieLet17_5QNode_Int_7QNode_Int_8QVal_Int_d = lizzieLet17_5QNode_Int_5QNode_Int_onehotd[1];
  assign lizzieLet17_5QNode_Int_7QNode_Int_8QNode_Int_d = lizzieLet17_5QNode_Int_5QNode_Int_onehotd[2];
  assign lizzieLet17_5QNode_Int_7QNode_Int_8QError_Int_d = lizzieLet17_5QNode_Int_5QNode_Int_onehotd[3];
  assign lizzieLet17_5QNode_Int_5QNode_Int_r = (| (lizzieLet17_5QNode_Int_5QNode_Int_onehotd & {lizzieLet17_5QNode_Int_7QNode_Int_8QError_Int_r,
                                                                                                lizzieLet17_5QNode_Int_7QNode_Int_8QNode_Int_r,
                                                                                                lizzieLet17_5QNode_Int_7QNode_Int_8QVal_Int_r,
                                                                                                lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_r}));
  assign lizzieLet17_5QNode_Int_7QNode_Int_8_r = lizzieLet17_5QNode_Int_5QNode_Int_r;
  
  /* fork (Ty Go) : (lizzieLet17_5QNode_Int_7QNode_Int_8QError_Int,Go) > [(lizzieLet17_5QNode_Int_7QNode_Int_8QError_Int_1,Go),
                                                                     (lizzieLet17_5QNode_Int_7QNode_Int_8QError_Int_2,Go)] */
  logic [1:0] lizzieLet17_5QNode_Int_7QNode_Int_8QError_Int_emitted;
  logic [1:0] lizzieLet17_5QNode_Int_7QNode_Int_8QError_Int_done;
  assign lizzieLet17_5QNode_Int_7QNode_Int_8QError_Int_1_d = (lizzieLet17_5QNode_Int_7QNode_Int_8QError_Int_d[0] && (! lizzieLet17_5QNode_Int_7QNode_Int_8QError_Int_emitted[0]));
  assign lizzieLet17_5QNode_Int_7QNode_Int_8QError_Int_2_d = (lizzieLet17_5QNode_Int_7QNode_Int_8QError_Int_d[0] && (! lizzieLet17_5QNode_Int_7QNode_Int_8QError_Int_emitted[1]));
  assign lizzieLet17_5QNode_Int_7QNode_Int_8QError_Int_done = (lizzieLet17_5QNode_Int_7QNode_Int_8QError_Int_emitted | ({lizzieLet17_5QNode_Int_7QNode_Int_8QError_Int_2_d[0],
                                                                                                                         lizzieLet17_5QNode_Int_7QNode_Int_8QError_Int_1_d[0]} & {lizzieLet17_5QNode_Int_7QNode_Int_8QError_Int_2_r,
                                                                                                                                                                                  lizzieLet17_5QNode_Int_7QNode_Int_8QError_Int_1_r}));
  assign lizzieLet17_5QNode_Int_7QNode_Int_8QError_Int_r = (& lizzieLet17_5QNode_Int_7QNode_Int_8QError_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNode_Int_8QError_Int_emitted <= 2'd0;
    else
      lizzieLet17_5QNode_Int_7QNode_Int_8QError_Int_emitted <= (lizzieLet17_5QNode_Int_7QNode_Int_8QError_Int_r ? 2'd0 :
                                                                lizzieLet17_5QNode_Int_7QNode_Int_8QError_Int_done);
  
  /* dcon (Ty QTree_Int,
      Dcon QError_Int) : [(lizzieLet17_5QNode_Int_7QNode_Int_8QError_Int_1,Go)] > (lizzieLet17_5QNode_Int_7QNode_Int_8QError_Int_1QError_Int,QTree_Int) */
  assign lizzieLet17_5QNode_Int_7QNode_Int_8QError_Int_1QError_Int_d = QError_Int_dc((& {lizzieLet17_5QNode_Int_7QNode_Int_8QError_Int_1_d[0]}), lizzieLet17_5QNode_Int_7QNode_Int_8QError_Int_1_d);
  assign {lizzieLet17_5QNode_Int_7QNode_Int_8QError_Int_1_r} = {1 {(lizzieLet17_5QNode_Int_7QNode_Int_8QError_Int_1QError_Int_r && lizzieLet17_5QNode_Int_7QNode_Int_8QError_Int_1QError_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (lizzieLet17_5QNode_Int_7QNode_Int_8QError_Int_1QError_Int,QTree_Int) > (lizzieLet53_1_argbuf,QTree_Int) */
  QTree_Int_t lizzieLet17_5QNode_Int_7QNode_Int_8QError_Int_1QError_Int_bufchan_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_8QError_Int_1QError_Int_bufchan_r;
  assign lizzieLet17_5QNode_Int_7QNode_Int_8QError_Int_1QError_Int_r = ((! lizzieLet17_5QNode_Int_7QNode_Int_8QError_Int_1QError_Int_bufchan_d[0]) || lizzieLet17_5QNode_Int_7QNode_Int_8QError_Int_1QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNode_Int_8QError_Int_1QError_Int_bufchan_d <= {66'd0,
                                                                              1'd0};
    else
      if (lizzieLet17_5QNode_Int_7QNode_Int_8QError_Int_1QError_Int_r)
        lizzieLet17_5QNode_Int_7QNode_Int_8QError_Int_1QError_Int_bufchan_d <= lizzieLet17_5QNode_Int_7QNode_Int_8QError_Int_1QError_Int_d;
  QTree_Int_t lizzieLet17_5QNode_Int_7QNode_Int_8QError_Int_1QError_Int_bufchan_buf;
  assign lizzieLet17_5QNode_Int_7QNode_Int_8QError_Int_1QError_Int_bufchan_r = (! lizzieLet17_5QNode_Int_7QNode_Int_8QError_Int_1QError_Int_bufchan_buf[0]);
  assign lizzieLet53_1_argbuf_d = (lizzieLet17_5QNode_Int_7QNode_Int_8QError_Int_1QError_Int_bufchan_buf[0] ? lizzieLet17_5QNode_Int_7QNode_Int_8QError_Int_1QError_Int_bufchan_buf :
                                   lizzieLet17_5QNode_Int_7QNode_Int_8QError_Int_1QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNode_Int_8QError_Int_1QError_Int_bufchan_buf <= {66'd0,
                                                                                1'd0};
    else
      if ((lizzieLet53_1_argbuf_r && lizzieLet17_5QNode_Int_7QNode_Int_8QError_Int_1QError_Int_bufchan_buf[0]))
        lizzieLet17_5QNode_Int_7QNode_Int_8QError_Int_1QError_Int_bufchan_buf <= {66'd0,
                                                                                  1'd0};
      else if (((! lizzieLet53_1_argbuf_r) && (! lizzieLet17_5QNode_Int_7QNode_Int_8QError_Int_1QError_Int_bufchan_buf[0])))
        lizzieLet17_5QNode_Int_7QNode_Int_8QError_Int_1QError_Int_bufchan_buf <= lizzieLet17_5QNode_Int_7QNode_Int_8QError_Int_1QError_Int_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet17_5QNode_Int_7QNode_Int_8QError_Int_2,Go) > (lizzieLet17_5QNode_Int_7QNode_Int_8QError_Int_2_argbuf,Go) */
  Go_t lizzieLet17_5QNode_Int_7QNode_Int_8QError_Int_2_bufchan_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_8QError_Int_2_bufchan_r;
  assign lizzieLet17_5QNode_Int_7QNode_Int_8QError_Int_2_r = ((! lizzieLet17_5QNode_Int_7QNode_Int_8QError_Int_2_bufchan_d[0]) || lizzieLet17_5QNode_Int_7QNode_Int_8QError_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNode_Int_8QError_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet17_5QNode_Int_7QNode_Int_8QError_Int_2_r)
        lizzieLet17_5QNode_Int_7QNode_Int_8QError_Int_2_bufchan_d <= lizzieLet17_5QNode_Int_7QNode_Int_8QError_Int_2_d;
  Go_t lizzieLet17_5QNode_Int_7QNode_Int_8QError_Int_2_bufchan_buf;
  assign lizzieLet17_5QNode_Int_7QNode_Int_8QError_Int_2_bufchan_r = (! lizzieLet17_5QNode_Int_7QNode_Int_8QError_Int_2_bufchan_buf[0]);
  assign lizzieLet17_5QNode_Int_7QNode_Int_8QError_Int_2_argbuf_d = (lizzieLet17_5QNode_Int_7QNode_Int_8QError_Int_2_bufchan_buf[0] ? lizzieLet17_5QNode_Int_7QNode_Int_8QError_Int_2_bufchan_buf :
                                                                     lizzieLet17_5QNode_Int_7QNode_Int_8QError_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNode_Int_8QError_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet17_5QNode_Int_7QNode_Int_8QError_Int_2_argbuf_r && lizzieLet17_5QNode_Int_7QNode_Int_8QError_Int_2_bufchan_buf[0]))
        lizzieLet17_5QNode_Int_7QNode_Int_8QError_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet17_5QNode_Int_7QNode_Int_8QError_Int_2_argbuf_r) && (! lizzieLet17_5QNode_Int_7QNode_Int_8QError_Int_2_bufchan_buf[0])))
        lizzieLet17_5QNode_Int_7QNode_Int_8QError_Int_2_bufchan_buf <= lizzieLet17_5QNode_Int_7QNode_Int_8QError_Int_2_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet17_5QNode_Int_7QNode_Int_8QNode_Int,Go) > (lizzieLet17_5QNode_Int_7QNode_Int_8QNode_Int_1_argbuf,Go) */
  Go_t lizzieLet17_5QNode_Int_7QNode_Int_8QNode_Int_bufchan_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_8QNode_Int_bufchan_r;
  assign lizzieLet17_5QNode_Int_7QNode_Int_8QNode_Int_r = ((! lizzieLet17_5QNode_Int_7QNode_Int_8QNode_Int_bufchan_d[0]) || lizzieLet17_5QNode_Int_7QNode_Int_8QNode_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNode_Int_8QNode_Int_bufchan_d <= 1'd0;
    else
      if (lizzieLet17_5QNode_Int_7QNode_Int_8QNode_Int_r)
        lizzieLet17_5QNode_Int_7QNode_Int_8QNode_Int_bufchan_d <= lizzieLet17_5QNode_Int_7QNode_Int_8QNode_Int_d;
  Go_t lizzieLet17_5QNode_Int_7QNode_Int_8QNode_Int_bufchan_buf;
  assign lizzieLet17_5QNode_Int_7QNode_Int_8QNode_Int_bufchan_r = (! lizzieLet17_5QNode_Int_7QNode_Int_8QNode_Int_bufchan_buf[0]);
  assign lizzieLet17_5QNode_Int_7QNode_Int_8QNode_Int_1_argbuf_d = (lizzieLet17_5QNode_Int_7QNode_Int_8QNode_Int_bufchan_buf[0] ? lizzieLet17_5QNode_Int_7QNode_Int_8QNode_Int_bufchan_buf :
                                                                    lizzieLet17_5QNode_Int_7QNode_Int_8QNode_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNode_Int_8QNode_Int_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet17_5QNode_Int_7QNode_Int_8QNode_Int_1_argbuf_r && lizzieLet17_5QNode_Int_7QNode_Int_8QNode_Int_bufchan_buf[0]))
        lizzieLet17_5QNode_Int_7QNode_Int_8QNode_Int_bufchan_buf <= 1'd0;
      else if (((! lizzieLet17_5QNode_Int_7QNode_Int_8QNode_Int_1_argbuf_r) && (! lizzieLet17_5QNode_Int_7QNode_Int_8QNode_Int_bufchan_buf[0])))
        lizzieLet17_5QNode_Int_7QNode_Int_8QNode_Int_bufchan_buf <= lizzieLet17_5QNode_Int_7QNode_Int_8QNode_Int_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int,Go) > [(lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_1,Go),
                                                                    (lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_2,Go),
                                                                    (lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_3,Go),
                                                                    (lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_4,Go),
                                                                    (lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_5,Go)] */
  logic [4:0] lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_emitted;
  logic [4:0] lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_done;
  assign lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_1_d = (lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_d[0] && (! lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_emitted[0]));
  assign lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_2_d = (lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_d[0] && (! lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_emitted[1]));
  assign lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_3_d = (lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_d[0] && (! lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_emitted[2]));
  assign lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_4_d = (lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_d[0] && (! lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_emitted[3]));
  assign lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_5_d = (lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_d[0] && (! lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_emitted[4]));
  assign lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_done = (lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_emitted | ({lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_5_d[0],
                                                                                                                       lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_4_d[0],
                                                                                                                       lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_3_d[0],
                                                                                                                       lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_2_d[0],
                                                                                                                       lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_1_d[0]} & {lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_5_r,
                                                                                                                                                                               lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_4_r,
                                                                                                                                                                               lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_3_r,
                                                                                                                                                                               lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_2_r,
                                                                                                                                                                               lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_1_r}));
  assign lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_r = (& lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_emitted <= 5'd0;
    else
      lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_emitted <= (lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_r ? 5'd0 :
                                                               lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_done);
  
  /* buf (Ty Go) : (lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_1,Go) > (lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_1_argbuf,Go) */
  Go_t lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_1_bufchan_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_1_bufchan_r;
  assign lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_1_r = ((! lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_1_bufchan_d[0]) || lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_1_bufchan_d <= 1'd0;
    else
      if (lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_1_r)
        lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_1_bufchan_d <= lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_1_d;
  Go_t lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_1_bufchan_buf;
  assign lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_1_bufchan_r = (! lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_1_bufchan_buf[0]);
  assign lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_1_argbuf_d = (lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_1_bufchan_buf[0] ? lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_1_bufchan_buf :
                                                                    lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_1_argbuf_r && lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_1_bufchan_buf[0]))
        lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_1_argbuf_r) && (! lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_1_bufchan_buf[0])))
        lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_1_bufchan_buf <= lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_1_bufchan_d;
  
  /* dcon (Ty TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int,
      Dcon TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int) : [(lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_1_argbuf,Go),
                                                                                              (lizzieLet17_5QNode_Int_7QNode_Int_5QNone_Int_1_argbuf,Pointer_QTree_Int),
                                                                                              (lizzieLet17_5QNode_Int_7QNode_Int_14QNone_Int_1_argbuf,Pointer_QTree_Int),
                                                                                              (lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_1_argbuf,MyDTInt_Bool),
                                                                                              (lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_1_argbuf,MyDTInt_Int_Int)] > (f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int9,TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int) */
  assign \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int9_d  = TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_dc((& {lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_1_argbuf_d[0],
                                                                                                                                                                                                                    lizzieLet17_5QNode_Int_7QNode_Int_5QNone_Int_1_argbuf_d[0],
                                                                                                                                                                                                                    lizzieLet17_5QNode_Int_7QNode_Int_14QNone_Int_1_argbuf_d[0],
                                                                                                                                                                                                                    lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_1_argbuf_d[0],
                                                                                                                                                                                                                    lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_1_argbuf_d[0]}), lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_1_argbuf_d, lizzieLet17_5QNode_Int_7QNode_Int_5QNone_Int_1_argbuf_d, lizzieLet17_5QNode_Int_7QNode_Int_14QNone_Int_1_argbuf_d, lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_1_argbuf_d, lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_1_argbuf_d);
  assign {lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_1_argbuf_r,
          lizzieLet17_5QNode_Int_7QNode_Int_5QNone_Int_1_argbuf_r,
          lizzieLet17_5QNode_Int_7QNode_Int_14QNone_Int_1_argbuf_r,
          lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_1_argbuf_r,
          lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_1_argbuf_r} = {5 {(\f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int9_r  && \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int9_d [0])}};
  
  /* buf (Ty Go) : (lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_2,Go) > (lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_2_argbuf,Go) */
  Go_t lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_2_bufchan_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_2_bufchan_r;
  assign lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_2_r = ((! lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_2_bufchan_d[0]) || lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_2_r)
        lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_2_bufchan_d <= lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_2_d;
  Go_t lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_2_bufchan_buf;
  assign lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_2_bufchan_r = (! lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_2_bufchan_buf[0]);
  assign lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_2_argbuf_d = (lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_2_bufchan_buf[0] ? lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_2_bufchan_buf :
                                                                    lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_2_argbuf_r && lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_2_bufchan_buf[0]))
        lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_2_argbuf_r) && (! lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_2_bufchan_buf[0])))
        lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_2_bufchan_buf <= lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_2_bufchan_d;
  
  /* dcon (Ty TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int,
      Dcon TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int) : [(lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_2_argbuf,Go),
                                                                                              (lizzieLet17_5QNode_Int_7QNode_Int_4QNone_Int_1_argbuf,Pointer_QTree_Int),
                                                                                              (lizzieLet17_5QNode_Int_7QNode_Int_13QNone_Int_1_argbuf,Pointer_QTree_Int),
                                                                                              (lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_2_argbuf,MyDTInt_Bool),
                                                                                              (lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_2_argbuf,MyDTInt_Int_Int)] > (f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int10,TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int) */
  assign \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int10_d  = TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_dc((& {lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_2_argbuf_d[0],
                                                                                                                                                                                                                     lizzieLet17_5QNode_Int_7QNode_Int_4QNone_Int_1_argbuf_d[0],
                                                                                                                                                                                                                     lizzieLet17_5QNode_Int_7QNode_Int_13QNone_Int_1_argbuf_d[0],
                                                                                                                                                                                                                     lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_2_argbuf_d[0],
                                                                                                                                                                                                                     lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_2_argbuf_d[0]}), lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_2_argbuf_d, lizzieLet17_5QNode_Int_7QNode_Int_4QNone_Int_1_argbuf_d, lizzieLet17_5QNode_Int_7QNode_Int_13QNone_Int_1_argbuf_d, lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_2_argbuf_d, lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_2_argbuf_d);
  assign {lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_2_argbuf_r,
          lizzieLet17_5QNode_Int_7QNode_Int_4QNone_Int_1_argbuf_r,
          lizzieLet17_5QNode_Int_7QNode_Int_13QNone_Int_1_argbuf_r,
          lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_2_argbuf_r,
          lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_2_argbuf_r} = {5 {(\f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int10_r  && \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int10_d [0])}};
  
  /* buf (Ty Go) : (lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_3,Go) > (lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_3_argbuf,Go) */
  Go_t lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_3_bufchan_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_3_bufchan_r;
  assign lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_3_r = ((! lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_3_bufchan_d[0]) || lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_3_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_3_bufchan_d <= 1'd0;
    else
      if (lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_3_r)
        lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_3_bufchan_d <= lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_3_d;
  Go_t lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_3_bufchan_buf;
  assign lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_3_bufchan_r = (! lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_3_bufchan_buf[0]);
  assign lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_3_argbuf_d = (lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_3_bufchan_buf[0] ? lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_3_bufchan_buf :
                                                                    lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_3_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_3_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_3_argbuf_r && lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_3_bufchan_buf[0]))
        lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_3_bufchan_buf <= 1'd0;
      else if (((! lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_3_argbuf_r) && (! lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_3_bufchan_buf[0])))
        lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_3_bufchan_buf <= lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_3_bufchan_d;
  
  /* dcon (Ty TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int,
      Dcon TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int) : [(lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_3_argbuf,Go),
                                                                                              (lizzieLet17_5QNode_Int_7QNode_Int_3QNone_Int_1_argbuf,Pointer_QTree_Int),
                                                                                              (lizzieLet17_5QNode_Int_7QNode_Int_12QNone_Int_1_argbuf,Pointer_QTree_Int),
                                                                                              (lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_3_argbuf,MyDTInt_Bool),
                                                                                              (lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_3_argbuf,MyDTInt_Int_Int)] > (f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int11,TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int) */
  assign \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int11_d  = TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_dc((& {lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_3_argbuf_d[0],
                                                                                                                                                                                                                     lizzieLet17_5QNode_Int_7QNode_Int_3QNone_Int_1_argbuf_d[0],
                                                                                                                                                                                                                     lizzieLet17_5QNode_Int_7QNode_Int_12QNone_Int_1_argbuf_d[0],
                                                                                                                                                                                                                     lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_3_argbuf_d[0],
                                                                                                                                                                                                                     lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_3_argbuf_d[0]}), lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_3_argbuf_d, lizzieLet17_5QNode_Int_7QNode_Int_3QNone_Int_1_argbuf_d, lizzieLet17_5QNode_Int_7QNode_Int_12QNone_Int_1_argbuf_d, lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_3_argbuf_d, lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_3_argbuf_d);
  assign {lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_3_argbuf_r,
          lizzieLet17_5QNode_Int_7QNode_Int_3QNone_Int_1_argbuf_r,
          lizzieLet17_5QNode_Int_7QNode_Int_12QNone_Int_1_argbuf_r,
          lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_3_argbuf_r,
          lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_3_argbuf_r} = {5 {(\f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int11_r  && \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int11_d [0])}};
  
  /* buf (Ty Go) : (lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_4,Go) > (lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_4_argbuf,Go) */
  Go_t lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_4_bufchan_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_4_bufchan_r;
  assign lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_4_r = ((! lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_4_bufchan_d[0]) || lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_4_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_4_bufchan_d <= 1'd0;
    else
      if (lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_4_r)
        lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_4_bufchan_d <= lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_4_d;
  Go_t lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_4_bufchan_buf;
  assign lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_4_bufchan_r = (! lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_4_bufchan_buf[0]);
  assign lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_4_argbuf_d = (lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_4_bufchan_buf[0] ? lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_4_bufchan_buf :
                                                                    lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_4_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_4_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_4_argbuf_r && lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_4_bufchan_buf[0]))
        lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_4_bufchan_buf <= 1'd0;
      else if (((! lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_4_argbuf_r) && (! lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_4_bufchan_buf[0])))
        lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_4_bufchan_buf <= lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_4_bufchan_d;
  
  /* dcon (Ty TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int,
      Dcon TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int) : [(lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_4_argbuf,Go),
                                                                                              (lizzieLet17_5QNode_Int_7QNode_Int_10QNone_Int_1_argbuf,Pointer_QTree_Int),
                                                                                              (lizzieLet17_5QNode_Int_7QNode_Int_11QNone_Int_1_argbuf,Pointer_QTree_Int),
                                                                                              (lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_4_argbuf,MyDTInt_Bool),
                                                                                              (lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_4_argbuf,MyDTInt_Int_Int)] > (f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int12,TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int) */
  assign \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int12_d  = TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_dc((& {lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_4_argbuf_d[0],
                                                                                                                                                                                                                     lizzieLet17_5QNode_Int_7QNode_Int_10QNone_Int_1_argbuf_d[0],
                                                                                                                                                                                                                     lizzieLet17_5QNode_Int_7QNode_Int_11QNone_Int_1_argbuf_d[0],
                                                                                                                                                                                                                     lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_4_argbuf_d[0],
                                                                                                                                                                                                                     lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_4_argbuf_d[0]}), lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_4_argbuf_d, lizzieLet17_5QNode_Int_7QNode_Int_10QNone_Int_1_argbuf_d, lizzieLet17_5QNode_Int_7QNode_Int_11QNone_Int_1_argbuf_d, lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_4_argbuf_d, lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_4_argbuf_d);
  assign {lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_4_argbuf_r,
          lizzieLet17_5QNode_Int_7QNode_Int_10QNone_Int_1_argbuf_r,
          lizzieLet17_5QNode_Int_7QNode_Int_11QNone_Int_1_argbuf_r,
          lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_4_argbuf_r,
          lizzieLet17_5QNode_Int_7QNode_Int_6QNone_Int_4_argbuf_r} = {5 {(\f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int12_r  && \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int12_d [0])}};
  
  /* buf (Ty Go) : (lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_5,Go) > (lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_5_argbuf,Go) */
  Go_t lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_5_bufchan_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_5_bufchan_r;
  assign lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_5_r = ((! lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_5_bufchan_d[0]) || lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_5_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_5_bufchan_d <= 1'd0;
    else
      if (lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_5_r)
        lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_5_bufchan_d <= lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_5_d;
  Go_t lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_5_bufchan_buf;
  assign lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_5_bufchan_r = (! lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_5_bufchan_buf[0]);
  assign lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_5_argbuf_d = (lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_5_bufchan_buf[0] ? lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_5_bufchan_buf :
                                                                    lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_5_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_5_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_5_argbuf_r && lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_5_bufchan_buf[0]))
        lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_5_bufchan_buf <= 1'd0;
      else if (((! lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_5_argbuf_r) && (! lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_5_bufchan_buf[0])))
        lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_5_bufchan_buf <= lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_5_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet17_5QNode_Int_7QNode_Int_8QVal_Int,Go) > [(lizzieLet17_5QNode_Int_7QNode_Int_8QVal_Int_1,Go),
                                                                   (lizzieLet17_5QNode_Int_7QNode_Int_8QVal_Int_2,Go)] */
  logic [1:0] lizzieLet17_5QNode_Int_7QNode_Int_8QVal_Int_emitted;
  logic [1:0] lizzieLet17_5QNode_Int_7QNode_Int_8QVal_Int_done;
  assign lizzieLet17_5QNode_Int_7QNode_Int_8QVal_Int_1_d = (lizzieLet17_5QNode_Int_7QNode_Int_8QVal_Int_d[0] && (! lizzieLet17_5QNode_Int_7QNode_Int_8QVal_Int_emitted[0]));
  assign lizzieLet17_5QNode_Int_7QNode_Int_8QVal_Int_2_d = (lizzieLet17_5QNode_Int_7QNode_Int_8QVal_Int_d[0] && (! lizzieLet17_5QNode_Int_7QNode_Int_8QVal_Int_emitted[1]));
  assign lizzieLet17_5QNode_Int_7QNode_Int_8QVal_Int_done = (lizzieLet17_5QNode_Int_7QNode_Int_8QVal_Int_emitted | ({lizzieLet17_5QNode_Int_7QNode_Int_8QVal_Int_2_d[0],
                                                                                                                     lizzieLet17_5QNode_Int_7QNode_Int_8QVal_Int_1_d[0]} & {lizzieLet17_5QNode_Int_7QNode_Int_8QVal_Int_2_r,
                                                                                                                                                                            lizzieLet17_5QNode_Int_7QNode_Int_8QVal_Int_1_r}));
  assign lizzieLet17_5QNode_Int_7QNode_Int_8QVal_Int_r = (& lizzieLet17_5QNode_Int_7QNode_Int_8QVal_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNode_Int_8QVal_Int_emitted <= 2'd0;
    else
      lizzieLet17_5QNode_Int_7QNode_Int_8QVal_Int_emitted <= (lizzieLet17_5QNode_Int_7QNode_Int_8QVal_Int_r ? 2'd0 :
                                                              lizzieLet17_5QNode_Int_7QNode_Int_8QVal_Int_done);
  
  /* dcon (Ty QTree_Int,
      Dcon QError_Int) : [(lizzieLet17_5QNode_Int_7QNode_Int_8QVal_Int_1,Go)] > (lizzieLet17_5QNode_Int_7QNode_Int_8QVal_Int_1QError_Int,QTree_Int) */
  assign lizzieLet17_5QNode_Int_7QNode_Int_8QVal_Int_1QError_Int_d = QError_Int_dc((& {lizzieLet17_5QNode_Int_7QNode_Int_8QVal_Int_1_d[0]}), lizzieLet17_5QNode_Int_7QNode_Int_8QVal_Int_1_d);
  assign {lizzieLet17_5QNode_Int_7QNode_Int_8QVal_Int_1_r} = {1 {(lizzieLet17_5QNode_Int_7QNode_Int_8QVal_Int_1QError_Int_r && lizzieLet17_5QNode_Int_7QNode_Int_8QVal_Int_1QError_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (lizzieLet17_5QNode_Int_7QNode_Int_8QVal_Int_1QError_Int,QTree_Int) > (lizzieLet51_1_argbuf,QTree_Int) */
  QTree_Int_t lizzieLet17_5QNode_Int_7QNode_Int_8QVal_Int_1QError_Int_bufchan_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_8QVal_Int_1QError_Int_bufchan_r;
  assign lizzieLet17_5QNode_Int_7QNode_Int_8QVal_Int_1QError_Int_r = ((! lizzieLet17_5QNode_Int_7QNode_Int_8QVal_Int_1QError_Int_bufchan_d[0]) || lizzieLet17_5QNode_Int_7QNode_Int_8QVal_Int_1QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNode_Int_8QVal_Int_1QError_Int_bufchan_d <= {66'd0,
                                                                            1'd0};
    else
      if (lizzieLet17_5QNode_Int_7QNode_Int_8QVal_Int_1QError_Int_r)
        lizzieLet17_5QNode_Int_7QNode_Int_8QVal_Int_1QError_Int_bufchan_d <= lizzieLet17_5QNode_Int_7QNode_Int_8QVal_Int_1QError_Int_d;
  QTree_Int_t lizzieLet17_5QNode_Int_7QNode_Int_8QVal_Int_1QError_Int_bufchan_buf;
  assign lizzieLet17_5QNode_Int_7QNode_Int_8QVal_Int_1QError_Int_bufchan_r = (! lizzieLet17_5QNode_Int_7QNode_Int_8QVal_Int_1QError_Int_bufchan_buf[0]);
  assign lizzieLet51_1_argbuf_d = (lizzieLet17_5QNode_Int_7QNode_Int_8QVal_Int_1QError_Int_bufchan_buf[0] ? lizzieLet17_5QNode_Int_7QNode_Int_8QVal_Int_1QError_Int_bufchan_buf :
                                   lizzieLet17_5QNode_Int_7QNode_Int_8QVal_Int_1QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNode_Int_8QVal_Int_1QError_Int_bufchan_buf <= {66'd0,
                                                                              1'd0};
    else
      if ((lizzieLet51_1_argbuf_r && lizzieLet17_5QNode_Int_7QNode_Int_8QVal_Int_1QError_Int_bufchan_buf[0]))
        lizzieLet17_5QNode_Int_7QNode_Int_8QVal_Int_1QError_Int_bufchan_buf <= {66'd0,
                                                                                1'd0};
      else if (((! lizzieLet51_1_argbuf_r) && (! lizzieLet17_5QNode_Int_7QNode_Int_8QVal_Int_1QError_Int_bufchan_buf[0])))
        lizzieLet17_5QNode_Int_7QNode_Int_8QVal_Int_1QError_Int_bufchan_buf <= lizzieLet17_5QNode_Int_7QNode_Int_8QVal_Int_1QError_Int_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet17_5QNode_Int_7QNode_Int_8QVal_Int_2,Go) > (lizzieLet17_5QNode_Int_7QNode_Int_8QVal_Int_2_argbuf,Go) */
  Go_t lizzieLet17_5QNode_Int_7QNode_Int_8QVal_Int_2_bufchan_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_8QVal_Int_2_bufchan_r;
  assign lizzieLet17_5QNode_Int_7QNode_Int_8QVal_Int_2_r = ((! lizzieLet17_5QNode_Int_7QNode_Int_8QVal_Int_2_bufchan_d[0]) || lizzieLet17_5QNode_Int_7QNode_Int_8QVal_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNode_Int_8QVal_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet17_5QNode_Int_7QNode_Int_8QVal_Int_2_r)
        lizzieLet17_5QNode_Int_7QNode_Int_8QVal_Int_2_bufchan_d <= lizzieLet17_5QNode_Int_7QNode_Int_8QVal_Int_2_d;
  Go_t lizzieLet17_5QNode_Int_7QNode_Int_8QVal_Int_2_bufchan_buf;
  assign lizzieLet17_5QNode_Int_7QNode_Int_8QVal_Int_2_bufchan_r = (! lizzieLet17_5QNode_Int_7QNode_Int_8QVal_Int_2_bufchan_buf[0]);
  assign lizzieLet17_5QNode_Int_7QNode_Int_8QVal_Int_2_argbuf_d = (lizzieLet17_5QNode_Int_7QNode_Int_8QVal_Int_2_bufchan_buf[0] ? lizzieLet17_5QNode_Int_7QNode_Int_8QVal_Int_2_bufchan_buf :
                                                                   lizzieLet17_5QNode_Int_7QNode_Int_8QVal_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNode_Int_8QVal_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet17_5QNode_Int_7QNode_Int_8QVal_Int_2_argbuf_r && lizzieLet17_5QNode_Int_7QNode_Int_8QVal_Int_2_bufchan_buf[0]))
        lizzieLet17_5QNode_Int_7QNode_Int_8QVal_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet17_5QNode_Int_7QNode_Int_8QVal_Int_2_argbuf_r) && (! lizzieLet17_5QNode_Int_7QNode_Int_8QVal_Int_2_bufchan_buf[0])))
        lizzieLet17_5QNode_Int_7QNode_Int_8QVal_Int_2_bufchan_buf <= lizzieLet17_5QNode_Int_7QNode_Int_8QVal_Int_2_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty MyDTInt_Bool) : (lizzieLet17_5QNode_Int_7QNode_Int_9,QTree_Int) (lizzieLet17_5QNode_Int_6QNode_Int,MyDTInt_Bool) > [(lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int,MyDTInt_Bool),
                                                                                                                              (_183,MyDTInt_Bool),
                                                                                                                              (lizzieLet17_5QNode_Int_7QNode_Int_9QNode_Int,MyDTInt_Bool),
                                                                                                                              (_182,MyDTInt_Bool)] */
  logic [3:0] lizzieLet17_5QNode_Int_6QNode_Int_onehotd;
  always_comb
    if ((lizzieLet17_5QNode_Int_7QNode_Int_9_d[0] && lizzieLet17_5QNode_Int_6QNode_Int_d[0]))
      unique case (lizzieLet17_5QNode_Int_7QNode_Int_9_d[2:1])
        2'd0: lizzieLet17_5QNode_Int_6QNode_Int_onehotd = 4'd1;
        2'd1: lizzieLet17_5QNode_Int_6QNode_Int_onehotd = 4'd2;
        2'd2: lizzieLet17_5QNode_Int_6QNode_Int_onehotd = 4'd4;
        2'd3: lizzieLet17_5QNode_Int_6QNode_Int_onehotd = 4'd8;
        default: lizzieLet17_5QNode_Int_6QNode_Int_onehotd = 4'd0;
      endcase
    else lizzieLet17_5QNode_Int_6QNode_Int_onehotd = 4'd0;
  assign lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_d = lizzieLet17_5QNode_Int_6QNode_Int_onehotd[0];
  assign _183_d = lizzieLet17_5QNode_Int_6QNode_Int_onehotd[1];
  assign lizzieLet17_5QNode_Int_7QNode_Int_9QNode_Int_d = lizzieLet17_5QNode_Int_6QNode_Int_onehotd[2];
  assign _182_d = lizzieLet17_5QNode_Int_6QNode_Int_onehotd[3];
  assign lizzieLet17_5QNode_Int_6QNode_Int_r = (| (lizzieLet17_5QNode_Int_6QNode_Int_onehotd & {_182_r,
                                                                                                lizzieLet17_5QNode_Int_7QNode_Int_9QNode_Int_r,
                                                                                                _183_r,
                                                                                                lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_r}));
  assign lizzieLet17_5QNode_Int_7QNode_Int_9_r = lizzieLet17_5QNode_Int_6QNode_Int_r;
  
  /* fork (Ty MyDTInt_Bool) : (lizzieLet17_5QNode_Int_7QNode_Int_9QNode_Int,MyDTInt_Bool) > [(lizzieLet17_5QNode_Int_7QNode_Int_9QNode_Int_1,MyDTInt_Bool),
                                                                                        (lizzieLet17_5QNode_Int_7QNode_Int_9QNode_Int_2,MyDTInt_Bool)] */
  logic [1:0] lizzieLet17_5QNode_Int_7QNode_Int_9QNode_Int_emitted;
  logic [1:0] lizzieLet17_5QNode_Int_7QNode_Int_9QNode_Int_done;
  assign lizzieLet17_5QNode_Int_7QNode_Int_9QNode_Int_1_d = (lizzieLet17_5QNode_Int_7QNode_Int_9QNode_Int_d[0] && (! lizzieLet17_5QNode_Int_7QNode_Int_9QNode_Int_emitted[0]));
  assign lizzieLet17_5QNode_Int_7QNode_Int_9QNode_Int_2_d = (lizzieLet17_5QNode_Int_7QNode_Int_9QNode_Int_d[0] && (! lizzieLet17_5QNode_Int_7QNode_Int_9QNode_Int_emitted[1]));
  assign lizzieLet17_5QNode_Int_7QNode_Int_9QNode_Int_done = (lizzieLet17_5QNode_Int_7QNode_Int_9QNode_Int_emitted | ({lizzieLet17_5QNode_Int_7QNode_Int_9QNode_Int_2_d[0],
                                                                                                                       lizzieLet17_5QNode_Int_7QNode_Int_9QNode_Int_1_d[0]} & {lizzieLet17_5QNode_Int_7QNode_Int_9QNode_Int_2_r,
                                                                                                                                                                               lizzieLet17_5QNode_Int_7QNode_Int_9QNode_Int_1_r}));
  assign lizzieLet17_5QNode_Int_7QNode_Int_9QNode_Int_r = (& lizzieLet17_5QNode_Int_7QNode_Int_9QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNode_Int_9QNode_Int_emitted <= 2'd0;
    else
      lizzieLet17_5QNode_Int_7QNode_Int_9QNode_Int_emitted <= (lizzieLet17_5QNode_Int_7QNode_Int_9QNode_Int_r ? 2'd0 :
                                                               lizzieLet17_5QNode_Int_7QNode_Int_9QNode_Int_done);
  
  /* buf (Ty MyDTInt_Bool) : (lizzieLet17_5QNode_Int_7QNode_Int_9QNode_Int_2,MyDTInt_Bool) > (lizzieLet17_5QNode_Int_7QNode_Int_9QNode_Int_2_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t lizzieLet17_5QNode_Int_7QNode_Int_9QNode_Int_2_bufchan_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_9QNode_Int_2_bufchan_r;
  assign lizzieLet17_5QNode_Int_7QNode_Int_9QNode_Int_2_r = ((! lizzieLet17_5QNode_Int_7QNode_Int_9QNode_Int_2_bufchan_d[0]) || lizzieLet17_5QNode_Int_7QNode_Int_9QNode_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNode_Int_9QNode_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet17_5QNode_Int_7QNode_Int_9QNode_Int_2_r)
        lizzieLet17_5QNode_Int_7QNode_Int_9QNode_Int_2_bufchan_d <= lizzieLet17_5QNode_Int_7QNode_Int_9QNode_Int_2_d;
  MyDTInt_Bool_t lizzieLet17_5QNode_Int_7QNode_Int_9QNode_Int_2_bufchan_buf;
  assign lizzieLet17_5QNode_Int_7QNode_Int_9QNode_Int_2_bufchan_r = (! lizzieLet17_5QNode_Int_7QNode_Int_9QNode_Int_2_bufchan_buf[0]);
  assign lizzieLet17_5QNode_Int_7QNode_Int_9QNode_Int_2_argbuf_d = (lizzieLet17_5QNode_Int_7QNode_Int_9QNode_Int_2_bufchan_buf[0] ? lizzieLet17_5QNode_Int_7QNode_Int_9QNode_Int_2_bufchan_buf :
                                                                    lizzieLet17_5QNode_Int_7QNode_Int_9QNode_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNode_Int_9QNode_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet17_5QNode_Int_7QNode_Int_9QNode_Int_2_argbuf_r && lizzieLet17_5QNode_Int_7QNode_Int_9QNode_Int_2_bufchan_buf[0]))
        lizzieLet17_5QNode_Int_7QNode_Int_9QNode_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet17_5QNode_Int_7QNode_Int_9QNode_Int_2_argbuf_r) && (! lizzieLet17_5QNode_Int_7QNode_Int_9QNode_Int_2_bufchan_buf[0])))
        lizzieLet17_5QNode_Int_7QNode_Int_9QNode_Int_2_bufchan_buf <= lizzieLet17_5QNode_Int_7QNode_Int_9QNode_Int_2_bufchan_d;
  
  /* fork (Ty MyDTInt_Bool) : (lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int,MyDTInt_Bool) > [(lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_1,MyDTInt_Bool),
                                                                                        (lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_2,MyDTInt_Bool),
                                                                                        (lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_3,MyDTInt_Bool),
                                                                                        (lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_4,MyDTInt_Bool)] */
  logic [3:0] lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_emitted;
  logic [3:0] lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_done;
  assign lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_1_d = (lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_d[0] && (! lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_emitted[0]));
  assign lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_2_d = (lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_d[0] && (! lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_emitted[1]));
  assign lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_3_d = (lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_d[0] && (! lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_emitted[2]));
  assign lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_4_d = (lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_d[0] && (! lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_emitted[3]));
  assign lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_done = (lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_emitted | ({lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_4_d[0],
                                                                                                                       lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_3_d[0],
                                                                                                                       lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_2_d[0],
                                                                                                                       lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_1_d[0]} & {lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_4_r,
                                                                                                                                                                               lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_3_r,
                                                                                                                                                                               lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_2_r,
                                                                                                                                                                               lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_1_r}));
  assign lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_r = (& lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_emitted <= 4'd0;
    else
      lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_emitted <= (lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_r ? 4'd0 :
                                                               lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_done);
  
  /* buf (Ty MyDTInt_Bool) : (lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_1,MyDTInt_Bool) > (lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_1_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_1_bufchan_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_1_bufchan_r;
  assign lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_1_r = ((! lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_1_bufchan_d[0]) || lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_1_bufchan_d <= 1'd0;
    else
      if (lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_1_r)
        lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_1_bufchan_d <= lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_1_d;
  MyDTInt_Bool_t lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_1_bufchan_buf;
  assign lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_1_bufchan_r = (! lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_1_bufchan_buf[0]);
  assign lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_1_argbuf_d = (lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_1_bufchan_buf[0] ? lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_1_bufchan_buf :
                                                                    lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_1_argbuf_r && lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_1_bufchan_buf[0]))
        lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_1_argbuf_r) && (! lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_1_bufchan_buf[0])))
        lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_1_bufchan_buf <= lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_1_bufchan_d;
  
  /* buf (Ty MyDTInt_Bool) : (lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_2,MyDTInt_Bool) > (lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_2_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_2_bufchan_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_2_bufchan_r;
  assign lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_2_r = ((! lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_2_bufchan_d[0]) || lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_2_r)
        lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_2_bufchan_d <= lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_2_d;
  MyDTInt_Bool_t lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_2_bufchan_buf;
  assign lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_2_bufchan_r = (! lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_2_bufchan_buf[0]);
  assign lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_2_argbuf_d = (lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_2_bufchan_buf[0] ? lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_2_bufchan_buf :
                                                                    lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_2_argbuf_r && lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_2_bufchan_buf[0]))
        lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_2_argbuf_r) && (! lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_2_bufchan_buf[0])))
        lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_2_bufchan_buf <= lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_2_bufchan_d;
  
  /* buf (Ty MyDTInt_Bool) : (lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_3,MyDTInt_Bool) > (lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_3_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_3_bufchan_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_3_bufchan_r;
  assign lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_3_r = ((! lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_3_bufchan_d[0]) || lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_3_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_3_bufchan_d <= 1'd0;
    else
      if (lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_3_r)
        lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_3_bufchan_d <= lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_3_d;
  MyDTInt_Bool_t lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_3_bufchan_buf;
  assign lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_3_bufchan_r = (! lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_3_bufchan_buf[0]);
  assign lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_3_argbuf_d = (lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_3_bufchan_buf[0] ? lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_3_bufchan_buf :
                                                                    lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_3_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_3_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_3_argbuf_r && lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_3_bufchan_buf[0]))
        lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_3_bufchan_buf <= 1'd0;
      else if (((! lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_3_argbuf_r) && (! lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_3_bufchan_buf[0])))
        lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_3_bufchan_buf <= lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_3_bufchan_d;
  
  /* buf (Ty MyDTInt_Bool) : (lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_4,MyDTInt_Bool) > (lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_4_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_4_bufchan_d;
  logic lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_4_bufchan_r;
  assign lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_4_r = ((! lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_4_bufchan_d[0]) || lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_4_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_4_bufchan_d <= 1'd0;
    else
      if (lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_4_r)
        lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_4_bufchan_d <= lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_4_d;
  MyDTInt_Bool_t lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_4_bufchan_buf;
  assign lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_4_bufchan_r = (! lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_4_bufchan_buf[0]);
  assign lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_4_argbuf_d = (lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_4_bufchan_buf[0] ? lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_4_bufchan_buf :
                                                                    lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_4_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_4_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_4_argbuf_r && lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_4_bufchan_buf[0]))
        lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_4_bufchan_buf <= 1'd0;
      else if (((! lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_4_argbuf_r) && (! lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_4_bufchan_buf[0])))
        lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_4_bufchan_buf <= lizzieLet17_5QNode_Int_7QNode_Int_9QNone_Int_4_bufchan_d;
  
  /* fork (Ty QTree_Int) : (lizzieLet17_5QNode_Int_7QNone_Int,QTree_Int) > [(lizzieLet17_5QNode_Int_7QNone_Int_1,QTree_Int),
                                                                       (lizzieLet17_5QNode_Int_7QNone_Int_2,QTree_Int),
                                                                       (lizzieLet17_5QNode_Int_7QNone_Int_3,QTree_Int),
                                                                       (lizzieLet17_5QNode_Int_7QNone_Int_4,QTree_Int),
                                                                       (lizzieLet17_5QNode_Int_7QNone_Int_5,QTree_Int),
                                                                       (lizzieLet17_5QNode_Int_7QNone_Int_6,QTree_Int),
                                                                       (lizzieLet17_5QNode_Int_7QNone_Int_7,QTree_Int),
                                                                       (lizzieLet17_5QNode_Int_7QNone_Int_8,QTree_Int),
                                                                       (lizzieLet17_5QNode_Int_7QNone_Int_9,QTree_Int),
                                                                       (lizzieLet17_5QNode_Int_7QNone_Int_10,QTree_Int),
                                                                       (lizzieLet17_5QNode_Int_7QNone_Int_11,QTree_Int)] */
  logic [10:0] lizzieLet17_5QNode_Int_7QNone_Int_emitted;
  logic [10:0] lizzieLet17_5QNode_Int_7QNone_Int_done;
  assign lizzieLet17_5QNode_Int_7QNone_Int_1_d = {lizzieLet17_5QNode_Int_7QNone_Int_d[66:1],
                                                  (lizzieLet17_5QNode_Int_7QNone_Int_d[0] && (! lizzieLet17_5QNode_Int_7QNone_Int_emitted[0]))};
  assign lizzieLet17_5QNode_Int_7QNone_Int_2_d = {lizzieLet17_5QNode_Int_7QNone_Int_d[66:1],
                                                  (lizzieLet17_5QNode_Int_7QNone_Int_d[0] && (! lizzieLet17_5QNode_Int_7QNone_Int_emitted[1]))};
  assign lizzieLet17_5QNode_Int_7QNone_Int_3_d = {lizzieLet17_5QNode_Int_7QNone_Int_d[66:1],
                                                  (lizzieLet17_5QNode_Int_7QNone_Int_d[0] && (! lizzieLet17_5QNode_Int_7QNone_Int_emitted[2]))};
  assign lizzieLet17_5QNode_Int_7QNone_Int_4_d = {lizzieLet17_5QNode_Int_7QNone_Int_d[66:1],
                                                  (lizzieLet17_5QNode_Int_7QNone_Int_d[0] && (! lizzieLet17_5QNode_Int_7QNone_Int_emitted[3]))};
  assign lizzieLet17_5QNode_Int_7QNone_Int_5_d = {lizzieLet17_5QNode_Int_7QNone_Int_d[66:1],
                                                  (lizzieLet17_5QNode_Int_7QNone_Int_d[0] && (! lizzieLet17_5QNode_Int_7QNone_Int_emitted[4]))};
  assign lizzieLet17_5QNode_Int_7QNone_Int_6_d = {lizzieLet17_5QNode_Int_7QNone_Int_d[66:1],
                                                  (lizzieLet17_5QNode_Int_7QNone_Int_d[0] && (! lizzieLet17_5QNode_Int_7QNone_Int_emitted[5]))};
  assign lizzieLet17_5QNode_Int_7QNone_Int_7_d = {lizzieLet17_5QNode_Int_7QNone_Int_d[66:1],
                                                  (lizzieLet17_5QNode_Int_7QNone_Int_d[0] && (! lizzieLet17_5QNode_Int_7QNone_Int_emitted[6]))};
  assign lizzieLet17_5QNode_Int_7QNone_Int_8_d = {lizzieLet17_5QNode_Int_7QNone_Int_d[66:1],
                                                  (lizzieLet17_5QNode_Int_7QNone_Int_d[0] && (! lizzieLet17_5QNode_Int_7QNone_Int_emitted[7]))};
  assign lizzieLet17_5QNode_Int_7QNone_Int_9_d = {lizzieLet17_5QNode_Int_7QNone_Int_d[66:1],
                                                  (lizzieLet17_5QNode_Int_7QNone_Int_d[0] && (! lizzieLet17_5QNode_Int_7QNone_Int_emitted[8]))};
  assign lizzieLet17_5QNode_Int_7QNone_Int_10_d = {lizzieLet17_5QNode_Int_7QNone_Int_d[66:1],
                                                   (lizzieLet17_5QNode_Int_7QNone_Int_d[0] && (! lizzieLet17_5QNode_Int_7QNone_Int_emitted[9]))};
  assign lizzieLet17_5QNode_Int_7QNone_Int_11_d = {lizzieLet17_5QNode_Int_7QNone_Int_d[66:1],
                                                   (lizzieLet17_5QNode_Int_7QNone_Int_d[0] && (! lizzieLet17_5QNode_Int_7QNone_Int_emitted[10]))};
  assign lizzieLet17_5QNode_Int_7QNone_Int_done = (lizzieLet17_5QNode_Int_7QNone_Int_emitted | ({lizzieLet17_5QNode_Int_7QNone_Int_11_d[0],
                                                                                                 lizzieLet17_5QNode_Int_7QNone_Int_10_d[0],
                                                                                                 lizzieLet17_5QNode_Int_7QNone_Int_9_d[0],
                                                                                                 lizzieLet17_5QNode_Int_7QNone_Int_8_d[0],
                                                                                                 lizzieLet17_5QNode_Int_7QNone_Int_7_d[0],
                                                                                                 lizzieLet17_5QNode_Int_7QNone_Int_6_d[0],
                                                                                                 lizzieLet17_5QNode_Int_7QNone_Int_5_d[0],
                                                                                                 lizzieLet17_5QNode_Int_7QNone_Int_4_d[0],
                                                                                                 lizzieLet17_5QNode_Int_7QNone_Int_3_d[0],
                                                                                                 lizzieLet17_5QNode_Int_7QNone_Int_2_d[0],
                                                                                                 lizzieLet17_5QNode_Int_7QNone_Int_1_d[0]} & {lizzieLet17_5QNode_Int_7QNone_Int_11_r,
                                                                                                                                              lizzieLet17_5QNode_Int_7QNone_Int_10_r,
                                                                                                                                              lizzieLet17_5QNode_Int_7QNone_Int_9_r,
                                                                                                                                              lizzieLet17_5QNode_Int_7QNone_Int_8_r,
                                                                                                                                              lizzieLet17_5QNode_Int_7QNone_Int_7_r,
                                                                                                                                              lizzieLet17_5QNode_Int_7QNone_Int_6_r,
                                                                                                                                              lizzieLet17_5QNode_Int_7QNone_Int_5_r,
                                                                                                                                              lizzieLet17_5QNode_Int_7QNone_Int_4_r,
                                                                                                                                              lizzieLet17_5QNode_Int_7QNone_Int_3_r,
                                                                                                                                              lizzieLet17_5QNode_Int_7QNone_Int_2_r,
                                                                                                                                              lizzieLet17_5QNode_Int_7QNone_Int_1_r}));
  assign lizzieLet17_5QNode_Int_7QNone_Int_r = (& lizzieLet17_5QNode_Int_7QNone_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNone_Int_emitted <= 11'd0;
    else
      lizzieLet17_5QNode_Int_7QNone_Int_emitted <= (lizzieLet17_5QNode_Int_7QNone_Int_r ? 11'd0 :
                                                    lizzieLet17_5QNode_Int_7QNone_Int_done);
  
  /* demux (Ty QTree_Int,
       Ty Pointer_QTree_Int) : (lizzieLet17_5QNode_Int_7QNone_Int_10,QTree_Int) (lizzieLet17_5QNode_Int_8QNone_Int,Pointer_QTree_Int) > [(lizzieLet17_5QNode_Int_7QNone_Int_10QNone_Int,Pointer_QTree_Int),
                                                                                                                                         (_181,Pointer_QTree_Int),
                                                                                                                                         (_180,Pointer_QTree_Int),
                                                                                                                                         (_179,Pointer_QTree_Int)] */
  logic [3:0] lizzieLet17_5QNode_Int_8QNone_Int_onehotd;
  always_comb
    if ((lizzieLet17_5QNode_Int_7QNone_Int_10_d[0] && lizzieLet17_5QNode_Int_8QNone_Int_d[0]))
      unique case (lizzieLet17_5QNode_Int_7QNone_Int_10_d[2:1])
        2'd0: lizzieLet17_5QNode_Int_8QNone_Int_onehotd = 4'd1;
        2'd1: lizzieLet17_5QNode_Int_8QNone_Int_onehotd = 4'd2;
        2'd2: lizzieLet17_5QNode_Int_8QNone_Int_onehotd = 4'd4;
        2'd3: lizzieLet17_5QNode_Int_8QNone_Int_onehotd = 4'd8;
        default: lizzieLet17_5QNode_Int_8QNone_Int_onehotd = 4'd0;
      endcase
    else lizzieLet17_5QNode_Int_8QNone_Int_onehotd = 4'd0;
  assign lizzieLet17_5QNode_Int_7QNone_Int_10QNone_Int_d = {lizzieLet17_5QNode_Int_8QNone_Int_d[16:1],
                                                            lizzieLet17_5QNode_Int_8QNone_Int_onehotd[0]};
  assign _181_d = {lizzieLet17_5QNode_Int_8QNone_Int_d[16:1],
                   lizzieLet17_5QNode_Int_8QNone_Int_onehotd[1]};
  assign _180_d = {lizzieLet17_5QNode_Int_8QNone_Int_d[16:1],
                   lizzieLet17_5QNode_Int_8QNone_Int_onehotd[2]};
  assign _179_d = {lizzieLet17_5QNode_Int_8QNone_Int_d[16:1],
                   lizzieLet17_5QNode_Int_8QNone_Int_onehotd[3]};
  assign lizzieLet17_5QNode_Int_8QNone_Int_r = (| (lizzieLet17_5QNode_Int_8QNone_Int_onehotd & {_179_r,
                                                                                                _180_r,
                                                                                                _181_r,
                                                                                                lizzieLet17_5QNode_Int_7QNone_Int_10QNone_Int_r}));
  assign lizzieLet17_5QNode_Int_7QNone_Int_10_r = lizzieLet17_5QNode_Int_8QNone_Int_r;
  
  /* buf (Ty Pointer_QTree_Int) : (lizzieLet17_5QNode_Int_7QNone_Int_10QNone_Int,Pointer_QTree_Int) > (lizzieLet17_5QNode_Int_7QNone_Int_10QNone_Int_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t lizzieLet17_5QNode_Int_7QNone_Int_10QNone_Int_bufchan_d;
  logic lizzieLet17_5QNode_Int_7QNone_Int_10QNone_Int_bufchan_r;
  assign lizzieLet17_5QNode_Int_7QNone_Int_10QNone_Int_r = ((! lizzieLet17_5QNode_Int_7QNone_Int_10QNone_Int_bufchan_d[0]) || lizzieLet17_5QNode_Int_7QNone_Int_10QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNone_Int_10QNone_Int_bufchan_d <= {16'd0,
                                                                  1'd0};
    else
      if (lizzieLet17_5QNode_Int_7QNone_Int_10QNone_Int_r)
        lizzieLet17_5QNode_Int_7QNone_Int_10QNone_Int_bufchan_d <= lizzieLet17_5QNode_Int_7QNone_Int_10QNone_Int_d;
  Pointer_QTree_Int_t lizzieLet17_5QNode_Int_7QNone_Int_10QNone_Int_bufchan_buf;
  assign lizzieLet17_5QNode_Int_7QNone_Int_10QNone_Int_bufchan_r = (! lizzieLet17_5QNode_Int_7QNone_Int_10QNone_Int_bufchan_buf[0]);
  assign lizzieLet17_5QNode_Int_7QNone_Int_10QNone_Int_1_argbuf_d = (lizzieLet17_5QNode_Int_7QNone_Int_10QNone_Int_bufchan_buf[0] ? lizzieLet17_5QNode_Int_7QNone_Int_10QNone_Int_bufchan_buf :
                                                                     lizzieLet17_5QNode_Int_7QNone_Int_10QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNone_Int_10QNone_Int_bufchan_buf <= {16'd0,
                                                                    1'd0};
    else
      if ((lizzieLet17_5QNode_Int_7QNone_Int_10QNone_Int_1_argbuf_r && lizzieLet17_5QNode_Int_7QNone_Int_10QNone_Int_bufchan_buf[0]))
        lizzieLet17_5QNode_Int_7QNone_Int_10QNone_Int_bufchan_buf <= {16'd0,
                                                                      1'd0};
      else if (((! lizzieLet17_5QNode_Int_7QNone_Int_10QNone_Int_1_argbuf_r) && (! lizzieLet17_5QNode_Int_7QNone_Int_10QNone_Int_bufchan_buf[0])))
        lizzieLet17_5QNode_Int_7QNone_Int_10QNone_Int_bufchan_buf <= lizzieLet17_5QNode_Int_7QNone_Int_10QNone_Int_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_QTree_Int) : (lizzieLet17_5QNode_Int_7QNone_Int_11,QTree_Int) (lizzieLet17_5QNode_Int_9QNone_Int,Pointer_QTree_Int) > [(_178,Pointer_QTree_Int),
                                                                                                                                         (_177,Pointer_QTree_Int),
                                                                                                                                         (lizzieLet17_5QNode_Int_7QNone_Int_11QNode_Int,Pointer_QTree_Int),
                                                                                                                                         (_176,Pointer_QTree_Int)] */
  logic [3:0] lizzieLet17_5QNode_Int_9QNone_Int_onehotd;
  always_comb
    if ((lizzieLet17_5QNode_Int_7QNone_Int_11_d[0] && lizzieLet17_5QNode_Int_9QNone_Int_d[0]))
      unique case (lizzieLet17_5QNode_Int_7QNone_Int_11_d[2:1])
        2'd0: lizzieLet17_5QNode_Int_9QNone_Int_onehotd = 4'd1;
        2'd1: lizzieLet17_5QNode_Int_9QNone_Int_onehotd = 4'd2;
        2'd2: lizzieLet17_5QNode_Int_9QNone_Int_onehotd = 4'd4;
        2'd3: lizzieLet17_5QNode_Int_9QNone_Int_onehotd = 4'd8;
        default: lizzieLet17_5QNode_Int_9QNone_Int_onehotd = 4'd0;
      endcase
    else lizzieLet17_5QNode_Int_9QNone_Int_onehotd = 4'd0;
  assign _178_d = {lizzieLet17_5QNode_Int_9QNone_Int_d[16:1],
                   lizzieLet17_5QNode_Int_9QNone_Int_onehotd[0]};
  assign _177_d = {lizzieLet17_5QNode_Int_9QNone_Int_d[16:1],
                   lizzieLet17_5QNode_Int_9QNone_Int_onehotd[1]};
  assign lizzieLet17_5QNode_Int_7QNone_Int_11QNode_Int_d = {lizzieLet17_5QNode_Int_9QNone_Int_d[16:1],
                                                            lizzieLet17_5QNode_Int_9QNone_Int_onehotd[2]};
  assign _176_d = {lizzieLet17_5QNode_Int_9QNone_Int_d[16:1],
                   lizzieLet17_5QNode_Int_9QNone_Int_onehotd[3]};
  assign lizzieLet17_5QNode_Int_9QNone_Int_r = (| (lizzieLet17_5QNode_Int_9QNone_Int_onehotd & {_176_r,
                                                                                                lizzieLet17_5QNode_Int_7QNone_Int_11QNode_Int_r,
                                                                                                _177_r,
                                                                                                _178_r}));
  assign lizzieLet17_5QNode_Int_7QNone_Int_11_r = lizzieLet17_5QNode_Int_9QNone_Int_r;
  
  /* buf (Ty Pointer_QTree_Int) : (lizzieLet17_5QNode_Int_7QNone_Int_11QNode_Int,Pointer_QTree_Int) > (lizzieLet17_5QNode_Int_7QNone_Int_11QNode_Int_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t lizzieLet17_5QNode_Int_7QNone_Int_11QNode_Int_bufchan_d;
  logic lizzieLet17_5QNode_Int_7QNone_Int_11QNode_Int_bufchan_r;
  assign lizzieLet17_5QNode_Int_7QNone_Int_11QNode_Int_r = ((! lizzieLet17_5QNode_Int_7QNone_Int_11QNode_Int_bufchan_d[0]) || lizzieLet17_5QNode_Int_7QNone_Int_11QNode_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNone_Int_11QNode_Int_bufchan_d <= {16'd0,
                                                                  1'd0};
    else
      if (lizzieLet17_5QNode_Int_7QNone_Int_11QNode_Int_r)
        lizzieLet17_5QNode_Int_7QNone_Int_11QNode_Int_bufchan_d <= lizzieLet17_5QNode_Int_7QNone_Int_11QNode_Int_d;
  Pointer_QTree_Int_t lizzieLet17_5QNode_Int_7QNone_Int_11QNode_Int_bufchan_buf;
  assign lizzieLet17_5QNode_Int_7QNone_Int_11QNode_Int_bufchan_r = (! lizzieLet17_5QNode_Int_7QNone_Int_11QNode_Int_bufchan_buf[0]);
  assign lizzieLet17_5QNode_Int_7QNone_Int_11QNode_Int_1_argbuf_d = (lizzieLet17_5QNode_Int_7QNone_Int_11QNode_Int_bufchan_buf[0] ? lizzieLet17_5QNode_Int_7QNone_Int_11QNode_Int_bufchan_buf :
                                                                     lizzieLet17_5QNode_Int_7QNone_Int_11QNode_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNone_Int_11QNode_Int_bufchan_buf <= {16'd0,
                                                                    1'd0};
    else
      if ((lizzieLet17_5QNode_Int_7QNone_Int_11QNode_Int_1_argbuf_r && lizzieLet17_5QNode_Int_7QNone_Int_11QNode_Int_bufchan_buf[0]))
        lizzieLet17_5QNode_Int_7QNone_Int_11QNode_Int_bufchan_buf <= {16'd0,
                                                                      1'd0};
      else if (((! lizzieLet17_5QNode_Int_7QNone_Int_11QNode_Int_1_argbuf_r) && (! lizzieLet17_5QNode_Int_7QNone_Int_11QNode_Int_bufchan_buf[0])))
        lizzieLet17_5QNode_Int_7QNone_Int_11QNode_Int_bufchan_buf <= lizzieLet17_5QNode_Int_7QNone_Int_11QNode_Int_bufchan_d;
  
  /* destruct (Ty QTree_Int,
          Dcon QNode_Int) : (lizzieLet17_5QNode_Int_7QNone_Int_1QNode_Int,QTree_Int) > [(t1af5_destruct,Pointer_QTree_Int),
                                                                                        (t2af6_destruct,Pointer_QTree_Int),
                                                                                        (t3af7_destruct,Pointer_QTree_Int),
                                                                                        (t4af8_destruct,Pointer_QTree_Int)] */
  logic [3:0] lizzieLet17_5QNode_Int_7QNone_Int_1QNode_Int_emitted;
  logic [3:0] lizzieLet17_5QNode_Int_7QNone_Int_1QNode_Int_done;
  assign t1af5_destruct_d = {lizzieLet17_5QNode_Int_7QNone_Int_1QNode_Int_d[18:3],
                             (lizzieLet17_5QNode_Int_7QNone_Int_1QNode_Int_d[0] && (! lizzieLet17_5QNode_Int_7QNone_Int_1QNode_Int_emitted[0]))};
  assign t2af6_destruct_d = {lizzieLet17_5QNode_Int_7QNone_Int_1QNode_Int_d[34:19],
                             (lizzieLet17_5QNode_Int_7QNone_Int_1QNode_Int_d[0] && (! lizzieLet17_5QNode_Int_7QNone_Int_1QNode_Int_emitted[1]))};
  assign t3af7_destruct_d = {lizzieLet17_5QNode_Int_7QNone_Int_1QNode_Int_d[50:35],
                             (lizzieLet17_5QNode_Int_7QNone_Int_1QNode_Int_d[0] && (! lizzieLet17_5QNode_Int_7QNone_Int_1QNode_Int_emitted[2]))};
  assign t4af8_destruct_d = {lizzieLet17_5QNode_Int_7QNone_Int_1QNode_Int_d[66:51],
                             (lizzieLet17_5QNode_Int_7QNone_Int_1QNode_Int_d[0] && (! lizzieLet17_5QNode_Int_7QNone_Int_1QNode_Int_emitted[3]))};
  assign lizzieLet17_5QNode_Int_7QNone_Int_1QNode_Int_done = (lizzieLet17_5QNode_Int_7QNone_Int_1QNode_Int_emitted | ({t4af8_destruct_d[0],
                                                                                                                       t3af7_destruct_d[0],
                                                                                                                       t2af6_destruct_d[0],
                                                                                                                       t1af5_destruct_d[0]} & {t4af8_destruct_r,
                                                                                                                                               t3af7_destruct_r,
                                                                                                                                               t2af6_destruct_r,
                                                                                                                                               t1af5_destruct_r}));
  assign lizzieLet17_5QNode_Int_7QNone_Int_1QNode_Int_r = (& lizzieLet17_5QNode_Int_7QNone_Int_1QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNone_Int_1QNode_Int_emitted <= 4'd0;
    else
      lizzieLet17_5QNode_Int_7QNone_Int_1QNode_Int_emitted <= (lizzieLet17_5QNode_Int_7QNone_Int_1QNode_Int_r ? 4'd0 :
                                                               lizzieLet17_5QNode_Int_7QNone_Int_1QNode_Int_done);
  
  /* demux (Ty QTree_Int,
       Ty QTree_Int) : (lizzieLet17_5QNode_Int_7QNone_Int_2,QTree_Int) (lizzieLet17_5QNode_Int_7QNone_Int_1,QTree_Int) > [(_175,QTree_Int),
                                                                                                                          (_174,QTree_Int),
                                                                                                                          (lizzieLet17_5QNode_Int_7QNone_Int_1QNode_Int,QTree_Int),
                                                                                                                          (_173,QTree_Int)] */
  logic [3:0] lizzieLet17_5QNode_Int_7QNone_Int_1_onehotd;
  always_comb
    if ((lizzieLet17_5QNode_Int_7QNone_Int_2_d[0] && lizzieLet17_5QNode_Int_7QNone_Int_1_d[0]))
      unique case (lizzieLet17_5QNode_Int_7QNone_Int_2_d[2:1])
        2'd0: lizzieLet17_5QNode_Int_7QNone_Int_1_onehotd = 4'd1;
        2'd1: lizzieLet17_5QNode_Int_7QNone_Int_1_onehotd = 4'd2;
        2'd2: lizzieLet17_5QNode_Int_7QNone_Int_1_onehotd = 4'd4;
        2'd3: lizzieLet17_5QNode_Int_7QNone_Int_1_onehotd = 4'd8;
        default: lizzieLet17_5QNode_Int_7QNone_Int_1_onehotd = 4'd0;
      endcase
    else lizzieLet17_5QNode_Int_7QNone_Int_1_onehotd = 4'd0;
  assign _175_d = {lizzieLet17_5QNode_Int_7QNone_Int_1_d[66:1],
                   lizzieLet17_5QNode_Int_7QNone_Int_1_onehotd[0]};
  assign _174_d = {lizzieLet17_5QNode_Int_7QNone_Int_1_d[66:1],
                   lizzieLet17_5QNode_Int_7QNone_Int_1_onehotd[1]};
  assign lizzieLet17_5QNode_Int_7QNone_Int_1QNode_Int_d = {lizzieLet17_5QNode_Int_7QNone_Int_1_d[66:1],
                                                           lizzieLet17_5QNode_Int_7QNone_Int_1_onehotd[2]};
  assign _173_d = {lizzieLet17_5QNode_Int_7QNone_Int_1_d[66:1],
                   lizzieLet17_5QNode_Int_7QNone_Int_1_onehotd[3]};
  assign lizzieLet17_5QNode_Int_7QNone_Int_1_r = (| (lizzieLet17_5QNode_Int_7QNone_Int_1_onehotd & {_173_r,
                                                                                                    lizzieLet17_5QNode_Int_7QNone_Int_1QNode_Int_r,
                                                                                                    _174_r,
                                                                                                    _175_r}));
  assign lizzieLet17_5QNode_Int_7QNone_Int_2_r = lizzieLet17_5QNode_Int_7QNone_Int_1_r;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_QTree_Int) : (lizzieLet17_5QNode_Int_7QNone_Int_3,QTree_Int) (lizzieLet17_5QNode_Int_10QNone_Int,Pointer_QTree_Int) > [(_172,Pointer_QTree_Int),
                                                                                                                                         (_171,Pointer_QTree_Int),
                                                                                                                                         (lizzieLet17_5QNode_Int_7QNone_Int_3QNode_Int,Pointer_QTree_Int),
                                                                                                                                         (_170,Pointer_QTree_Int)] */
  logic [3:0] lizzieLet17_5QNode_Int_10QNone_Int_onehotd;
  always_comb
    if ((lizzieLet17_5QNode_Int_7QNone_Int_3_d[0] && lizzieLet17_5QNode_Int_10QNone_Int_d[0]))
      unique case (lizzieLet17_5QNode_Int_7QNone_Int_3_d[2:1])
        2'd0: lizzieLet17_5QNode_Int_10QNone_Int_onehotd = 4'd1;
        2'd1: lizzieLet17_5QNode_Int_10QNone_Int_onehotd = 4'd2;
        2'd2: lizzieLet17_5QNode_Int_10QNone_Int_onehotd = 4'd4;
        2'd3: lizzieLet17_5QNode_Int_10QNone_Int_onehotd = 4'd8;
        default: lizzieLet17_5QNode_Int_10QNone_Int_onehotd = 4'd0;
      endcase
    else lizzieLet17_5QNode_Int_10QNone_Int_onehotd = 4'd0;
  assign _172_d = {lizzieLet17_5QNode_Int_10QNone_Int_d[16:1],
                   lizzieLet17_5QNode_Int_10QNone_Int_onehotd[0]};
  assign _171_d = {lizzieLet17_5QNode_Int_10QNone_Int_d[16:1],
                   lizzieLet17_5QNode_Int_10QNone_Int_onehotd[1]};
  assign lizzieLet17_5QNode_Int_7QNone_Int_3QNode_Int_d = {lizzieLet17_5QNode_Int_10QNone_Int_d[16:1],
                                                           lizzieLet17_5QNode_Int_10QNone_Int_onehotd[2]};
  assign _170_d = {lizzieLet17_5QNode_Int_10QNone_Int_d[16:1],
                   lizzieLet17_5QNode_Int_10QNone_Int_onehotd[3]};
  assign lizzieLet17_5QNode_Int_10QNone_Int_r = (| (lizzieLet17_5QNode_Int_10QNone_Int_onehotd & {_170_r,
                                                                                                  lizzieLet17_5QNode_Int_7QNone_Int_3QNode_Int_r,
                                                                                                  _171_r,
                                                                                                  _172_r}));
  assign lizzieLet17_5QNode_Int_7QNone_Int_3_r = lizzieLet17_5QNode_Int_10QNone_Int_r;
  
  /* buf (Ty Pointer_QTree_Int) : (lizzieLet17_5QNode_Int_7QNone_Int_3QNode_Int,Pointer_QTree_Int) > (lizzieLet17_5QNode_Int_7QNone_Int_3QNode_Int_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t lizzieLet17_5QNode_Int_7QNone_Int_3QNode_Int_bufchan_d;
  logic lizzieLet17_5QNode_Int_7QNone_Int_3QNode_Int_bufchan_r;
  assign lizzieLet17_5QNode_Int_7QNone_Int_3QNode_Int_r = ((! lizzieLet17_5QNode_Int_7QNone_Int_3QNode_Int_bufchan_d[0]) || lizzieLet17_5QNode_Int_7QNone_Int_3QNode_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNone_Int_3QNode_Int_bufchan_d <= {16'd0,
                                                                 1'd0};
    else
      if (lizzieLet17_5QNode_Int_7QNone_Int_3QNode_Int_r)
        lizzieLet17_5QNode_Int_7QNone_Int_3QNode_Int_bufchan_d <= lizzieLet17_5QNode_Int_7QNone_Int_3QNode_Int_d;
  Pointer_QTree_Int_t lizzieLet17_5QNode_Int_7QNone_Int_3QNode_Int_bufchan_buf;
  assign lizzieLet17_5QNode_Int_7QNone_Int_3QNode_Int_bufchan_r = (! lizzieLet17_5QNode_Int_7QNone_Int_3QNode_Int_bufchan_buf[0]);
  assign lizzieLet17_5QNode_Int_7QNone_Int_3QNode_Int_1_argbuf_d = (lizzieLet17_5QNode_Int_7QNone_Int_3QNode_Int_bufchan_buf[0] ? lizzieLet17_5QNode_Int_7QNone_Int_3QNode_Int_bufchan_buf :
                                                                    lizzieLet17_5QNode_Int_7QNone_Int_3QNode_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNone_Int_3QNode_Int_bufchan_buf <= {16'd0,
                                                                   1'd0};
    else
      if ((lizzieLet17_5QNode_Int_7QNone_Int_3QNode_Int_1_argbuf_r && lizzieLet17_5QNode_Int_7QNone_Int_3QNode_Int_bufchan_buf[0]))
        lizzieLet17_5QNode_Int_7QNone_Int_3QNode_Int_bufchan_buf <= {16'd0,
                                                                     1'd0};
      else if (((! lizzieLet17_5QNode_Int_7QNone_Int_3QNode_Int_1_argbuf_r) && (! lizzieLet17_5QNode_Int_7QNone_Int_3QNode_Int_bufchan_buf[0])))
        lizzieLet17_5QNode_Int_7QNone_Int_3QNode_Int_bufchan_buf <= lizzieLet17_5QNode_Int_7QNone_Int_3QNode_Int_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_QTree_Int) : (lizzieLet17_5QNode_Int_7QNone_Int_4,QTree_Int) (lizzieLet17_5QNode_Int_11QNone_Int,Pointer_QTree_Int) > [(_169,Pointer_QTree_Int),
                                                                                                                                         (_168,Pointer_QTree_Int),
                                                                                                                                         (lizzieLet17_5QNode_Int_7QNone_Int_4QNode_Int,Pointer_QTree_Int),
                                                                                                                                         (_167,Pointer_QTree_Int)] */
  logic [3:0] lizzieLet17_5QNode_Int_11QNone_Int_onehotd;
  always_comb
    if ((lizzieLet17_5QNode_Int_7QNone_Int_4_d[0] && lizzieLet17_5QNode_Int_11QNone_Int_d[0]))
      unique case (lizzieLet17_5QNode_Int_7QNone_Int_4_d[2:1])
        2'd0: lizzieLet17_5QNode_Int_11QNone_Int_onehotd = 4'd1;
        2'd1: lizzieLet17_5QNode_Int_11QNone_Int_onehotd = 4'd2;
        2'd2: lizzieLet17_5QNode_Int_11QNone_Int_onehotd = 4'd4;
        2'd3: lizzieLet17_5QNode_Int_11QNone_Int_onehotd = 4'd8;
        default: lizzieLet17_5QNode_Int_11QNone_Int_onehotd = 4'd0;
      endcase
    else lizzieLet17_5QNode_Int_11QNone_Int_onehotd = 4'd0;
  assign _169_d = {lizzieLet17_5QNode_Int_11QNone_Int_d[16:1],
                   lizzieLet17_5QNode_Int_11QNone_Int_onehotd[0]};
  assign _168_d = {lizzieLet17_5QNode_Int_11QNone_Int_d[16:1],
                   lizzieLet17_5QNode_Int_11QNone_Int_onehotd[1]};
  assign lizzieLet17_5QNode_Int_7QNone_Int_4QNode_Int_d = {lizzieLet17_5QNode_Int_11QNone_Int_d[16:1],
                                                           lizzieLet17_5QNode_Int_11QNone_Int_onehotd[2]};
  assign _167_d = {lizzieLet17_5QNode_Int_11QNone_Int_d[16:1],
                   lizzieLet17_5QNode_Int_11QNone_Int_onehotd[3]};
  assign lizzieLet17_5QNode_Int_11QNone_Int_r = (| (lizzieLet17_5QNode_Int_11QNone_Int_onehotd & {_167_r,
                                                                                                  lizzieLet17_5QNode_Int_7QNone_Int_4QNode_Int_r,
                                                                                                  _168_r,
                                                                                                  _169_r}));
  assign lizzieLet17_5QNode_Int_7QNone_Int_4_r = lizzieLet17_5QNode_Int_11QNone_Int_r;
  
  /* buf (Ty Pointer_QTree_Int) : (lizzieLet17_5QNode_Int_7QNone_Int_4QNode_Int,Pointer_QTree_Int) > (lizzieLet17_5QNode_Int_7QNone_Int_4QNode_Int_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t lizzieLet17_5QNode_Int_7QNone_Int_4QNode_Int_bufchan_d;
  logic lizzieLet17_5QNode_Int_7QNone_Int_4QNode_Int_bufchan_r;
  assign lizzieLet17_5QNode_Int_7QNone_Int_4QNode_Int_r = ((! lizzieLet17_5QNode_Int_7QNone_Int_4QNode_Int_bufchan_d[0]) || lizzieLet17_5QNode_Int_7QNone_Int_4QNode_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNone_Int_4QNode_Int_bufchan_d <= {16'd0,
                                                                 1'd0};
    else
      if (lizzieLet17_5QNode_Int_7QNone_Int_4QNode_Int_r)
        lizzieLet17_5QNode_Int_7QNone_Int_4QNode_Int_bufchan_d <= lizzieLet17_5QNode_Int_7QNone_Int_4QNode_Int_d;
  Pointer_QTree_Int_t lizzieLet17_5QNode_Int_7QNone_Int_4QNode_Int_bufchan_buf;
  assign lizzieLet17_5QNode_Int_7QNone_Int_4QNode_Int_bufchan_r = (! lizzieLet17_5QNode_Int_7QNone_Int_4QNode_Int_bufchan_buf[0]);
  assign lizzieLet17_5QNode_Int_7QNone_Int_4QNode_Int_1_argbuf_d = (lizzieLet17_5QNode_Int_7QNone_Int_4QNode_Int_bufchan_buf[0] ? lizzieLet17_5QNode_Int_7QNone_Int_4QNode_Int_bufchan_buf :
                                                                    lizzieLet17_5QNode_Int_7QNone_Int_4QNode_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNone_Int_4QNode_Int_bufchan_buf <= {16'd0,
                                                                   1'd0};
    else
      if ((lizzieLet17_5QNode_Int_7QNone_Int_4QNode_Int_1_argbuf_r && lizzieLet17_5QNode_Int_7QNone_Int_4QNode_Int_bufchan_buf[0]))
        lizzieLet17_5QNode_Int_7QNone_Int_4QNode_Int_bufchan_buf <= {16'd0,
                                                                     1'd0};
      else if (((! lizzieLet17_5QNode_Int_7QNone_Int_4QNode_Int_1_argbuf_r) && (! lizzieLet17_5QNode_Int_7QNone_Int_4QNode_Int_bufchan_buf[0])))
        lizzieLet17_5QNode_Int_7QNone_Int_4QNode_Int_bufchan_buf <= lizzieLet17_5QNode_Int_7QNone_Int_4QNode_Int_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_QTree_Int) : (lizzieLet17_5QNode_Int_7QNone_Int_5,QTree_Int) (lizzieLet17_5QNode_Int_12QNone_Int,Pointer_QTree_Int) > [(_166,Pointer_QTree_Int),
                                                                                                                                         (_165,Pointer_QTree_Int),
                                                                                                                                         (lizzieLet17_5QNode_Int_7QNone_Int_5QNode_Int,Pointer_QTree_Int),
                                                                                                                                         (_164,Pointer_QTree_Int)] */
  logic [3:0] lizzieLet17_5QNode_Int_12QNone_Int_onehotd;
  always_comb
    if ((lizzieLet17_5QNode_Int_7QNone_Int_5_d[0] && lizzieLet17_5QNode_Int_12QNone_Int_d[0]))
      unique case (lizzieLet17_5QNode_Int_7QNone_Int_5_d[2:1])
        2'd0: lizzieLet17_5QNode_Int_12QNone_Int_onehotd = 4'd1;
        2'd1: lizzieLet17_5QNode_Int_12QNone_Int_onehotd = 4'd2;
        2'd2: lizzieLet17_5QNode_Int_12QNone_Int_onehotd = 4'd4;
        2'd3: lizzieLet17_5QNode_Int_12QNone_Int_onehotd = 4'd8;
        default: lizzieLet17_5QNode_Int_12QNone_Int_onehotd = 4'd0;
      endcase
    else lizzieLet17_5QNode_Int_12QNone_Int_onehotd = 4'd0;
  assign _166_d = {lizzieLet17_5QNode_Int_12QNone_Int_d[16:1],
                   lizzieLet17_5QNode_Int_12QNone_Int_onehotd[0]};
  assign _165_d = {lizzieLet17_5QNode_Int_12QNone_Int_d[16:1],
                   lizzieLet17_5QNode_Int_12QNone_Int_onehotd[1]};
  assign lizzieLet17_5QNode_Int_7QNone_Int_5QNode_Int_d = {lizzieLet17_5QNode_Int_12QNone_Int_d[16:1],
                                                           lizzieLet17_5QNode_Int_12QNone_Int_onehotd[2]};
  assign _164_d = {lizzieLet17_5QNode_Int_12QNone_Int_d[16:1],
                   lizzieLet17_5QNode_Int_12QNone_Int_onehotd[3]};
  assign lizzieLet17_5QNode_Int_12QNone_Int_r = (| (lizzieLet17_5QNode_Int_12QNone_Int_onehotd & {_164_r,
                                                                                                  lizzieLet17_5QNode_Int_7QNone_Int_5QNode_Int_r,
                                                                                                  _165_r,
                                                                                                  _166_r}));
  assign lizzieLet17_5QNode_Int_7QNone_Int_5_r = lizzieLet17_5QNode_Int_12QNone_Int_r;
  
  /* buf (Ty Pointer_QTree_Int) : (lizzieLet17_5QNode_Int_7QNone_Int_5QNode_Int,Pointer_QTree_Int) > (lizzieLet17_5QNode_Int_7QNone_Int_5QNode_Int_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t lizzieLet17_5QNode_Int_7QNone_Int_5QNode_Int_bufchan_d;
  logic lizzieLet17_5QNode_Int_7QNone_Int_5QNode_Int_bufchan_r;
  assign lizzieLet17_5QNode_Int_7QNone_Int_5QNode_Int_r = ((! lizzieLet17_5QNode_Int_7QNone_Int_5QNode_Int_bufchan_d[0]) || lizzieLet17_5QNode_Int_7QNone_Int_5QNode_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNone_Int_5QNode_Int_bufchan_d <= {16'd0,
                                                                 1'd0};
    else
      if (lizzieLet17_5QNode_Int_7QNone_Int_5QNode_Int_r)
        lizzieLet17_5QNode_Int_7QNone_Int_5QNode_Int_bufchan_d <= lizzieLet17_5QNode_Int_7QNone_Int_5QNode_Int_d;
  Pointer_QTree_Int_t lizzieLet17_5QNode_Int_7QNone_Int_5QNode_Int_bufchan_buf;
  assign lizzieLet17_5QNode_Int_7QNone_Int_5QNode_Int_bufchan_r = (! lizzieLet17_5QNode_Int_7QNone_Int_5QNode_Int_bufchan_buf[0]);
  assign lizzieLet17_5QNode_Int_7QNone_Int_5QNode_Int_1_argbuf_d = (lizzieLet17_5QNode_Int_7QNone_Int_5QNode_Int_bufchan_buf[0] ? lizzieLet17_5QNode_Int_7QNone_Int_5QNode_Int_bufchan_buf :
                                                                    lizzieLet17_5QNode_Int_7QNone_Int_5QNode_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNone_Int_5QNode_Int_bufchan_buf <= {16'd0,
                                                                   1'd0};
    else
      if ((lizzieLet17_5QNode_Int_7QNone_Int_5QNode_Int_1_argbuf_r && lizzieLet17_5QNode_Int_7QNone_Int_5QNode_Int_bufchan_buf[0]))
        lizzieLet17_5QNode_Int_7QNone_Int_5QNode_Int_bufchan_buf <= {16'd0,
                                                                     1'd0};
      else if (((! lizzieLet17_5QNode_Int_7QNone_Int_5QNode_Int_1_argbuf_r) && (! lizzieLet17_5QNode_Int_7QNone_Int_5QNode_Int_bufchan_buf[0])))
        lizzieLet17_5QNode_Int_7QNone_Int_5QNode_Int_bufchan_buf <= lizzieLet17_5QNode_Int_7QNone_Int_5QNode_Int_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty MyDTInt_Int_Int) : (lizzieLet17_5QNode_Int_7QNone_Int_6,QTree_Int) (lizzieLet17_5QNode_Int_3QNone_Int,MyDTInt_Int_Int) > [(_163,MyDTInt_Int_Int),
                                                                                                                                    (_162,MyDTInt_Int_Int),
                                                                                                                                    (lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int,MyDTInt_Int_Int),
                                                                                                                                    (_161,MyDTInt_Int_Int)] */
  logic [3:0] lizzieLet17_5QNode_Int_3QNone_Int_onehotd;
  always_comb
    if ((lizzieLet17_5QNode_Int_7QNone_Int_6_d[0] && lizzieLet17_5QNode_Int_3QNone_Int_d[0]))
      unique case (lizzieLet17_5QNode_Int_7QNone_Int_6_d[2:1])
        2'd0: lizzieLet17_5QNode_Int_3QNone_Int_onehotd = 4'd1;
        2'd1: lizzieLet17_5QNode_Int_3QNone_Int_onehotd = 4'd2;
        2'd2: lizzieLet17_5QNode_Int_3QNone_Int_onehotd = 4'd4;
        2'd3: lizzieLet17_5QNode_Int_3QNone_Int_onehotd = 4'd8;
        default: lizzieLet17_5QNode_Int_3QNone_Int_onehotd = 4'd0;
      endcase
    else lizzieLet17_5QNode_Int_3QNone_Int_onehotd = 4'd0;
  assign _163_d = lizzieLet17_5QNode_Int_3QNone_Int_onehotd[0];
  assign _162_d = lizzieLet17_5QNode_Int_3QNone_Int_onehotd[1];
  assign lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_d = lizzieLet17_5QNode_Int_3QNone_Int_onehotd[2];
  assign _161_d = lizzieLet17_5QNode_Int_3QNone_Int_onehotd[3];
  assign lizzieLet17_5QNode_Int_3QNone_Int_r = (| (lizzieLet17_5QNode_Int_3QNone_Int_onehotd & {_161_r,
                                                                                                lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_r,
                                                                                                _162_r,
                                                                                                _163_r}));
  assign lizzieLet17_5QNode_Int_7QNone_Int_6_r = lizzieLet17_5QNode_Int_3QNone_Int_r;
  
  /* fork (Ty MyDTInt_Int_Int) : (lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int,MyDTInt_Int_Int) > [(lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_1,MyDTInt_Int_Int),
                                                                                              (lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_2,MyDTInt_Int_Int),
                                                                                              (lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_3,MyDTInt_Int_Int),
                                                                                              (lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_4,MyDTInt_Int_Int)] */
  logic [3:0] lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_emitted;
  logic [3:0] lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_done;
  assign lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_1_d = (lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_d[0] && (! lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_emitted[0]));
  assign lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_2_d = (lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_d[0] && (! lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_emitted[1]));
  assign lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_3_d = (lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_d[0] && (! lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_emitted[2]));
  assign lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_4_d = (lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_d[0] && (! lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_emitted[3]));
  assign lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_done = (lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_emitted | ({lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_4_d[0],
                                                                                                                       lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_3_d[0],
                                                                                                                       lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_2_d[0],
                                                                                                                       lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_1_d[0]} & {lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_4_r,
                                                                                                                                                                               lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_3_r,
                                                                                                                                                                               lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_2_r,
                                                                                                                                                                               lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_1_r}));
  assign lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_r = (& lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_emitted <= 4'd0;
    else
      lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_emitted <= (lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_r ? 4'd0 :
                                                               lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_done);
  
  /* buf (Ty MyDTInt_Int_Int) : (lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_1,MyDTInt_Int_Int) > (lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_1_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_1_bufchan_d;
  logic lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_1_bufchan_r;
  assign lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_1_r = ((! lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_1_bufchan_d[0]) || lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_1_bufchan_d <= 1'd0;
    else
      if (lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_1_r)
        lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_1_bufchan_d <= lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_1_d;
  MyDTInt_Int_Int_t lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_1_bufchan_buf;
  assign lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_1_bufchan_r = (! lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_1_bufchan_buf[0]);
  assign lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_1_argbuf_d = (lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_1_bufchan_buf[0] ? lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_1_bufchan_buf :
                                                                    lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_1_argbuf_r && lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_1_bufchan_buf[0]))
        lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_1_argbuf_r) && (! lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_1_bufchan_buf[0])))
        lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_1_bufchan_buf <= lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_1_bufchan_d;
  
  /* buf (Ty MyDTInt_Int_Int) : (lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_2,MyDTInt_Int_Int) > (lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_2_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_2_bufchan_d;
  logic lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_2_bufchan_r;
  assign lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_2_r = ((! lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_2_bufchan_d[0]) || lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_2_r)
        lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_2_bufchan_d <= lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_2_d;
  MyDTInt_Int_Int_t lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_2_bufchan_buf;
  assign lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_2_bufchan_r = (! lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_2_bufchan_buf[0]);
  assign lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_2_argbuf_d = (lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_2_bufchan_buf[0] ? lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_2_bufchan_buf :
                                                                    lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_2_argbuf_r && lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_2_bufchan_buf[0]))
        lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_2_argbuf_r) && (! lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_2_bufchan_buf[0])))
        lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_2_bufchan_buf <= lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_2_bufchan_d;
  
  /* buf (Ty MyDTInt_Int_Int) : (lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_3,MyDTInt_Int_Int) > (lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_3_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_3_bufchan_d;
  logic lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_3_bufchan_r;
  assign lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_3_r = ((! lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_3_bufchan_d[0]) || lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_3_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_3_bufchan_d <= 1'd0;
    else
      if (lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_3_r)
        lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_3_bufchan_d <= lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_3_d;
  MyDTInt_Int_Int_t lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_3_bufchan_buf;
  assign lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_3_bufchan_r = (! lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_3_bufchan_buf[0]);
  assign lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_3_argbuf_d = (lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_3_bufchan_buf[0] ? lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_3_bufchan_buf :
                                                                    lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_3_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_3_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_3_argbuf_r && lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_3_bufchan_buf[0]))
        lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_3_bufchan_buf <= 1'd0;
      else if (((! lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_3_argbuf_r) && (! lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_3_bufchan_buf[0])))
        lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_3_bufchan_buf <= lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_3_bufchan_d;
  
  /* buf (Ty MyDTInt_Int_Int) : (lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_4,MyDTInt_Int_Int) > (lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_4_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_4_bufchan_d;
  logic lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_4_bufchan_r;
  assign lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_4_r = ((! lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_4_bufchan_d[0]) || lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_4_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_4_bufchan_d <= 1'd0;
    else
      if (lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_4_r)
        lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_4_bufchan_d <= lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_4_d;
  MyDTInt_Int_Int_t lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_4_bufchan_buf;
  assign lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_4_bufchan_r = (! lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_4_bufchan_buf[0]);
  assign lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_4_argbuf_d = (lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_4_bufchan_buf[0] ? lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_4_bufchan_buf :
                                                                    lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_4_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_4_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_4_argbuf_r && lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_4_bufchan_buf[0]))
        lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_4_bufchan_buf <= 1'd0;
      else if (((! lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_4_argbuf_r) && (! lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_4_bufchan_buf[0])))
        lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_4_bufchan_buf <= lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_4_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_CTf_f_Int) : (lizzieLet17_5QNode_Int_7QNone_Int_7,QTree_Int) (lizzieLet17_5QNode_Int_4QNone_Int,Pointer_CTf_f_Int) > [(lizzieLet17_5QNode_Int_7QNone_Int_7QNone_Int,Pointer_CTf_f_Int),
                                                                                                                                        (lizzieLet17_5QNode_Int_7QNone_Int_7QVal_Int,Pointer_CTf_f_Int),
                                                                                                                                        (lizzieLet17_5QNode_Int_7QNone_Int_7QNode_Int,Pointer_CTf_f_Int),
                                                                                                                                        (lizzieLet17_5QNode_Int_7QNone_Int_7QError_Int,Pointer_CTf_f_Int)] */
  logic [3:0] lizzieLet17_5QNode_Int_4QNone_Int_onehotd;
  always_comb
    if ((lizzieLet17_5QNode_Int_7QNone_Int_7_d[0] && lizzieLet17_5QNode_Int_4QNone_Int_d[0]))
      unique case (lizzieLet17_5QNode_Int_7QNone_Int_7_d[2:1])
        2'd0: lizzieLet17_5QNode_Int_4QNone_Int_onehotd = 4'd1;
        2'd1: lizzieLet17_5QNode_Int_4QNone_Int_onehotd = 4'd2;
        2'd2: lizzieLet17_5QNode_Int_4QNone_Int_onehotd = 4'd4;
        2'd3: lizzieLet17_5QNode_Int_4QNone_Int_onehotd = 4'd8;
        default: lizzieLet17_5QNode_Int_4QNone_Int_onehotd = 4'd0;
      endcase
    else lizzieLet17_5QNode_Int_4QNone_Int_onehotd = 4'd0;
  assign lizzieLet17_5QNode_Int_7QNone_Int_7QNone_Int_d = {lizzieLet17_5QNode_Int_4QNone_Int_d[16:1],
                                                           lizzieLet17_5QNode_Int_4QNone_Int_onehotd[0]};
  assign lizzieLet17_5QNode_Int_7QNone_Int_7QVal_Int_d = {lizzieLet17_5QNode_Int_4QNone_Int_d[16:1],
                                                          lizzieLet17_5QNode_Int_4QNone_Int_onehotd[1]};
  assign lizzieLet17_5QNode_Int_7QNone_Int_7QNode_Int_d = {lizzieLet17_5QNode_Int_4QNone_Int_d[16:1],
                                                           lizzieLet17_5QNode_Int_4QNone_Int_onehotd[2]};
  assign lizzieLet17_5QNode_Int_7QNone_Int_7QError_Int_d = {lizzieLet17_5QNode_Int_4QNone_Int_d[16:1],
                                                            lizzieLet17_5QNode_Int_4QNone_Int_onehotd[3]};
  assign lizzieLet17_5QNode_Int_4QNone_Int_r = (| (lizzieLet17_5QNode_Int_4QNone_Int_onehotd & {lizzieLet17_5QNode_Int_7QNone_Int_7QError_Int_r,
                                                                                                lizzieLet17_5QNode_Int_7QNone_Int_7QNode_Int_r,
                                                                                                lizzieLet17_5QNode_Int_7QNone_Int_7QVal_Int_r,
                                                                                                lizzieLet17_5QNode_Int_7QNone_Int_7QNone_Int_r}));
  assign lizzieLet17_5QNode_Int_7QNone_Int_7_r = lizzieLet17_5QNode_Int_4QNone_Int_r;
  
  /* buf (Ty Pointer_CTf_f_Int) : (lizzieLet17_5QNode_Int_7QNone_Int_7QError_Int,Pointer_CTf_f_Int) > (lizzieLet17_5QNode_Int_7QNone_Int_7QError_Int_1_argbuf,Pointer_CTf_f_Int) */
  Pointer_CTf_f_Int_t lizzieLet17_5QNode_Int_7QNone_Int_7QError_Int_bufchan_d;
  logic lizzieLet17_5QNode_Int_7QNone_Int_7QError_Int_bufchan_r;
  assign lizzieLet17_5QNode_Int_7QNone_Int_7QError_Int_r = ((! lizzieLet17_5QNode_Int_7QNone_Int_7QError_Int_bufchan_d[0]) || lizzieLet17_5QNode_Int_7QNone_Int_7QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNone_Int_7QError_Int_bufchan_d <= {16'd0,
                                                                  1'd0};
    else
      if (lizzieLet17_5QNode_Int_7QNone_Int_7QError_Int_r)
        lizzieLet17_5QNode_Int_7QNone_Int_7QError_Int_bufchan_d <= lizzieLet17_5QNode_Int_7QNone_Int_7QError_Int_d;
  Pointer_CTf_f_Int_t lizzieLet17_5QNode_Int_7QNone_Int_7QError_Int_bufchan_buf;
  assign lizzieLet17_5QNode_Int_7QNone_Int_7QError_Int_bufchan_r = (! lizzieLet17_5QNode_Int_7QNone_Int_7QError_Int_bufchan_buf[0]);
  assign lizzieLet17_5QNode_Int_7QNone_Int_7QError_Int_1_argbuf_d = (lizzieLet17_5QNode_Int_7QNone_Int_7QError_Int_bufchan_buf[0] ? lizzieLet17_5QNode_Int_7QNone_Int_7QError_Int_bufchan_buf :
                                                                     lizzieLet17_5QNode_Int_7QNone_Int_7QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNone_Int_7QError_Int_bufchan_buf <= {16'd0,
                                                                    1'd0};
    else
      if ((lizzieLet17_5QNode_Int_7QNone_Int_7QError_Int_1_argbuf_r && lizzieLet17_5QNode_Int_7QNone_Int_7QError_Int_bufchan_buf[0]))
        lizzieLet17_5QNode_Int_7QNone_Int_7QError_Int_bufchan_buf <= {16'd0,
                                                                      1'd0};
      else if (((! lizzieLet17_5QNode_Int_7QNone_Int_7QError_Int_1_argbuf_r) && (! lizzieLet17_5QNode_Int_7QNone_Int_7QError_Int_bufchan_buf[0])))
        lizzieLet17_5QNode_Int_7QNone_Int_7QError_Int_bufchan_buf <= lizzieLet17_5QNode_Int_7QNone_Int_7QError_Int_bufchan_d;
  
  /* buf (Ty Pointer_CTf_f_Int) : (lizzieLet17_5QNode_Int_7QNone_Int_7QNode_Int,Pointer_CTf_f_Int) > (lizzieLet17_5QNode_Int_7QNone_Int_7QNode_Int_1_argbuf,Pointer_CTf_f_Int) */
  Pointer_CTf_f_Int_t lizzieLet17_5QNode_Int_7QNone_Int_7QNode_Int_bufchan_d;
  logic lizzieLet17_5QNode_Int_7QNone_Int_7QNode_Int_bufchan_r;
  assign lizzieLet17_5QNode_Int_7QNone_Int_7QNode_Int_r = ((! lizzieLet17_5QNode_Int_7QNone_Int_7QNode_Int_bufchan_d[0]) || lizzieLet17_5QNode_Int_7QNone_Int_7QNode_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNone_Int_7QNode_Int_bufchan_d <= {16'd0,
                                                                 1'd0};
    else
      if (lizzieLet17_5QNode_Int_7QNone_Int_7QNode_Int_r)
        lizzieLet17_5QNode_Int_7QNone_Int_7QNode_Int_bufchan_d <= lizzieLet17_5QNode_Int_7QNone_Int_7QNode_Int_d;
  Pointer_CTf_f_Int_t lizzieLet17_5QNode_Int_7QNone_Int_7QNode_Int_bufchan_buf;
  assign lizzieLet17_5QNode_Int_7QNone_Int_7QNode_Int_bufchan_r = (! lizzieLet17_5QNode_Int_7QNone_Int_7QNode_Int_bufchan_buf[0]);
  assign lizzieLet17_5QNode_Int_7QNone_Int_7QNode_Int_1_argbuf_d = (lizzieLet17_5QNode_Int_7QNone_Int_7QNode_Int_bufchan_buf[0] ? lizzieLet17_5QNode_Int_7QNone_Int_7QNode_Int_bufchan_buf :
                                                                    lizzieLet17_5QNode_Int_7QNone_Int_7QNode_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNone_Int_7QNode_Int_bufchan_buf <= {16'd0,
                                                                   1'd0};
    else
      if ((lizzieLet17_5QNode_Int_7QNone_Int_7QNode_Int_1_argbuf_r && lizzieLet17_5QNode_Int_7QNone_Int_7QNode_Int_bufchan_buf[0]))
        lizzieLet17_5QNode_Int_7QNone_Int_7QNode_Int_bufchan_buf <= {16'd0,
                                                                     1'd0};
      else if (((! lizzieLet17_5QNode_Int_7QNone_Int_7QNode_Int_1_argbuf_r) && (! lizzieLet17_5QNode_Int_7QNone_Int_7QNode_Int_bufchan_buf[0])))
        lizzieLet17_5QNode_Int_7QNone_Int_7QNode_Int_bufchan_buf <= lizzieLet17_5QNode_Int_7QNone_Int_7QNode_Int_bufchan_d;
  
  /* buf (Ty Pointer_CTf_f_Int) : (lizzieLet17_5QNode_Int_7QNone_Int_7QNone_Int,Pointer_CTf_f_Int) > (lizzieLet17_5QNode_Int_7QNone_Int_7QNone_Int_1_argbuf,Pointer_CTf_f_Int) */
  Pointer_CTf_f_Int_t lizzieLet17_5QNode_Int_7QNone_Int_7QNone_Int_bufchan_d;
  logic lizzieLet17_5QNode_Int_7QNone_Int_7QNone_Int_bufchan_r;
  assign lizzieLet17_5QNode_Int_7QNone_Int_7QNone_Int_r = ((! lizzieLet17_5QNode_Int_7QNone_Int_7QNone_Int_bufchan_d[0]) || lizzieLet17_5QNode_Int_7QNone_Int_7QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNone_Int_7QNone_Int_bufchan_d <= {16'd0,
                                                                 1'd0};
    else
      if (lizzieLet17_5QNode_Int_7QNone_Int_7QNone_Int_r)
        lizzieLet17_5QNode_Int_7QNone_Int_7QNone_Int_bufchan_d <= lizzieLet17_5QNode_Int_7QNone_Int_7QNone_Int_d;
  Pointer_CTf_f_Int_t lizzieLet17_5QNode_Int_7QNone_Int_7QNone_Int_bufchan_buf;
  assign lizzieLet17_5QNode_Int_7QNone_Int_7QNone_Int_bufchan_r = (! lizzieLet17_5QNode_Int_7QNone_Int_7QNone_Int_bufchan_buf[0]);
  assign lizzieLet17_5QNode_Int_7QNone_Int_7QNone_Int_1_argbuf_d = (lizzieLet17_5QNode_Int_7QNone_Int_7QNone_Int_bufchan_buf[0] ? lizzieLet17_5QNode_Int_7QNone_Int_7QNone_Int_bufchan_buf :
                                                                    lizzieLet17_5QNode_Int_7QNone_Int_7QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNone_Int_7QNone_Int_bufchan_buf <= {16'd0,
                                                                   1'd0};
    else
      if ((lizzieLet17_5QNode_Int_7QNone_Int_7QNone_Int_1_argbuf_r && lizzieLet17_5QNode_Int_7QNone_Int_7QNone_Int_bufchan_buf[0]))
        lizzieLet17_5QNode_Int_7QNone_Int_7QNone_Int_bufchan_buf <= {16'd0,
                                                                     1'd0};
      else if (((! lizzieLet17_5QNode_Int_7QNone_Int_7QNone_Int_1_argbuf_r) && (! lizzieLet17_5QNode_Int_7QNone_Int_7QNone_Int_bufchan_buf[0])))
        lizzieLet17_5QNode_Int_7QNone_Int_7QNone_Int_bufchan_buf <= lizzieLet17_5QNode_Int_7QNone_Int_7QNone_Int_bufchan_d;
  
  /* buf (Ty Pointer_CTf_f_Int) : (lizzieLet17_5QNode_Int_7QNone_Int_7QVal_Int,Pointer_CTf_f_Int) > (lizzieLet17_5QNode_Int_7QNone_Int_7QVal_Int_1_argbuf,Pointer_CTf_f_Int) */
  Pointer_CTf_f_Int_t lizzieLet17_5QNode_Int_7QNone_Int_7QVal_Int_bufchan_d;
  logic lizzieLet17_5QNode_Int_7QNone_Int_7QVal_Int_bufchan_r;
  assign lizzieLet17_5QNode_Int_7QNone_Int_7QVal_Int_r = ((! lizzieLet17_5QNode_Int_7QNone_Int_7QVal_Int_bufchan_d[0]) || lizzieLet17_5QNode_Int_7QNone_Int_7QVal_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNone_Int_7QVal_Int_bufchan_d <= {16'd0,
                                                                1'd0};
    else
      if (lizzieLet17_5QNode_Int_7QNone_Int_7QVal_Int_r)
        lizzieLet17_5QNode_Int_7QNone_Int_7QVal_Int_bufchan_d <= lizzieLet17_5QNode_Int_7QNone_Int_7QVal_Int_d;
  Pointer_CTf_f_Int_t lizzieLet17_5QNode_Int_7QNone_Int_7QVal_Int_bufchan_buf;
  assign lizzieLet17_5QNode_Int_7QNone_Int_7QVal_Int_bufchan_r = (! lizzieLet17_5QNode_Int_7QNone_Int_7QVal_Int_bufchan_buf[0]);
  assign lizzieLet17_5QNode_Int_7QNone_Int_7QVal_Int_1_argbuf_d = (lizzieLet17_5QNode_Int_7QNone_Int_7QVal_Int_bufchan_buf[0] ? lizzieLet17_5QNode_Int_7QNone_Int_7QVal_Int_bufchan_buf :
                                                                   lizzieLet17_5QNode_Int_7QNone_Int_7QVal_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNone_Int_7QVal_Int_bufchan_buf <= {16'd0,
                                                                  1'd0};
    else
      if ((lizzieLet17_5QNode_Int_7QNone_Int_7QVal_Int_1_argbuf_r && lizzieLet17_5QNode_Int_7QNone_Int_7QVal_Int_bufchan_buf[0]))
        lizzieLet17_5QNode_Int_7QNone_Int_7QVal_Int_bufchan_buf <= {16'd0,
                                                                    1'd0};
      else if (((! lizzieLet17_5QNode_Int_7QNone_Int_7QVal_Int_1_argbuf_r) && (! lizzieLet17_5QNode_Int_7QNone_Int_7QVal_Int_bufchan_buf[0])))
        lizzieLet17_5QNode_Int_7QNone_Int_7QVal_Int_bufchan_buf <= lizzieLet17_5QNode_Int_7QNone_Int_7QVal_Int_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Go) : (lizzieLet17_5QNode_Int_7QNone_Int_8,QTree_Int) (lizzieLet17_5QNode_Int_5QNone_Int,Go) > [(lizzieLet17_5QNode_Int_7QNone_Int_8QNone_Int,Go),
                                                                                                          (lizzieLet17_5QNode_Int_7QNone_Int_8QVal_Int,Go),
                                                                                                          (lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int,Go),
                                                                                                          (lizzieLet17_5QNode_Int_7QNone_Int_8QError_Int,Go)] */
  logic [3:0] lizzieLet17_5QNode_Int_5QNone_Int_onehotd;
  always_comb
    if ((lizzieLet17_5QNode_Int_7QNone_Int_8_d[0] && lizzieLet17_5QNode_Int_5QNone_Int_d[0]))
      unique case (lizzieLet17_5QNode_Int_7QNone_Int_8_d[2:1])
        2'd0: lizzieLet17_5QNode_Int_5QNone_Int_onehotd = 4'd1;
        2'd1: lizzieLet17_5QNode_Int_5QNone_Int_onehotd = 4'd2;
        2'd2: lizzieLet17_5QNode_Int_5QNone_Int_onehotd = 4'd4;
        2'd3: lizzieLet17_5QNode_Int_5QNone_Int_onehotd = 4'd8;
        default: lizzieLet17_5QNode_Int_5QNone_Int_onehotd = 4'd0;
      endcase
    else lizzieLet17_5QNode_Int_5QNone_Int_onehotd = 4'd0;
  assign lizzieLet17_5QNode_Int_7QNone_Int_8QNone_Int_d = lizzieLet17_5QNode_Int_5QNone_Int_onehotd[0];
  assign lizzieLet17_5QNode_Int_7QNone_Int_8QVal_Int_d = lizzieLet17_5QNode_Int_5QNone_Int_onehotd[1];
  assign lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_d = lizzieLet17_5QNode_Int_5QNone_Int_onehotd[2];
  assign lizzieLet17_5QNode_Int_7QNone_Int_8QError_Int_d = lizzieLet17_5QNode_Int_5QNone_Int_onehotd[3];
  assign lizzieLet17_5QNode_Int_5QNone_Int_r = (| (lizzieLet17_5QNode_Int_5QNone_Int_onehotd & {lizzieLet17_5QNode_Int_7QNone_Int_8QError_Int_r,
                                                                                                lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_r,
                                                                                                lizzieLet17_5QNode_Int_7QNone_Int_8QVal_Int_r,
                                                                                                lizzieLet17_5QNode_Int_7QNone_Int_8QNone_Int_r}));
  assign lizzieLet17_5QNode_Int_7QNone_Int_8_r = lizzieLet17_5QNode_Int_5QNone_Int_r;
  
  /* fork (Ty Go) : (lizzieLet17_5QNode_Int_7QNone_Int_8QError_Int,Go) > [(lizzieLet17_5QNode_Int_7QNone_Int_8QError_Int_1,Go),
                                                                     (lizzieLet17_5QNode_Int_7QNone_Int_8QError_Int_2,Go)] */
  logic [1:0] lizzieLet17_5QNode_Int_7QNone_Int_8QError_Int_emitted;
  logic [1:0] lizzieLet17_5QNode_Int_7QNone_Int_8QError_Int_done;
  assign lizzieLet17_5QNode_Int_7QNone_Int_8QError_Int_1_d = (lizzieLet17_5QNode_Int_7QNone_Int_8QError_Int_d[0] && (! lizzieLet17_5QNode_Int_7QNone_Int_8QError_Int_emitted[0]));
  assign lizzieLet17_5QNode_Int_7QNone_Int_8QError_Int_2_d = (lizzieLet17_5QNode_Int_7QNone_Int_8QError_Int_d[0] && (! lizzieLet17_5QNode_Int_7QNone_Int_8QError_Int_emitted[1]));
  assign lizzieLet17_5QNode_Int_7QNone_Int_8QError_Int_done = (lizzieLet17_5QNode_Int_7QNone_Int_8QError_Int_emitted | ({lizzieLet17_5QNode_Int_7QNone_Int_8QError_Int_2_d[0],
                                                                                                                         lizzieLet17_5QNode_Int_7QNone_Int_8QError_Int_1_d[0]} & {lizzieLet17_5QNode_Int_7QNone_Int_8QError_Int_2_r,
                                                                                                                                                                                  lizzieLet17_5QNode_Int_7QNone_Int_8QError_Int_1_r}));
  assign lizzieLet17_5QNode_Int_7QNone_Int_8QError_Int_r = (& lizzieLet17_5QNode_Int_7QNone_Int_8QError_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNone_Int_8QError_Int_emitted <= 2'd0;
    else
      lizzieLet17_5QNode_Int_7QNone_Int_8QError_Int_emitted <= (lizzieLet17_5QNode_Int_7QNone_Int_8QError_Int_r ? 2'd0 :
                                                                lizzieLet17_5QNode_Int_7QNone_Int_8QError_Int_done);
  
  /* dcon (Ty QTree_Int,
      Dcon QError_Int) : [(lizzieLet17_5QNode_Int_7QNone_Int_8QError_Int_1,Go)] > (lizzieLet17_5QNode_Int_7QNone_Int_8QError_Int_1QError_Int,QTree_Int) */
  assign lizzieLet17_5QNode_Int_7QNone_Int_8QError_Int_1QError_Int_d = QError_Int_dc((& {lizzieLet17_5QNode_Int_7QNone_Int_8QError_Int_1_d[0]}), lizzieLet17_5QNode_Int_7QNone_Int_8QError_Int_1_d);
  assign {lizzieLet17_5QNode_Int_7QNone_Int_8QError_Int_1_r} = {1 {(lizzieLet17_5QNode_Int_7QNone_Int_8QError_Int_1QError_Int_r && lizzieLet17_5QNode_Int_7QNone_Int_8QError_Int_1QError_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (lizzieLet17_5QNode_Int_7QNone_Int_8QError_Int_1QError_Int,QTree_Int) > (lizzieLet47_1_argbuf,QTree_Int) */
  QTree_Int_t lizzieLet17_5QNode_Int_7QNone_Int_8QError_Int_1QError_Int_bufchan_d;
  logic lizzieLet17_5QNode_Int_7QNone_Int_8QError_Int_1QError_Int_bufchan_r;
  assign lizzieLet17_5QNode_Int_7QNone_Int_8QError_Int_1QError_Int_r = ((! lizzieLet17_5QNode_Int_7QNone_Int_8QError_Int_1QError_Int_bufchan_d[0]) || lizzieLet17_5QNode_Int_7QNone_Int_8QError_Int_1QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNone_Int_8QError_Int_1QError_Int_bufchan_d <= {66'd0,
                                                                              1'd0};
    else
      if (lizzieLet17_5QNode_Int_7QNone_Int_8QError_Int_1QError_Int_r)
        lizzieLet17_5QNode_Int_7QNone_Int_8QError_Int_1QError_Int_bufchan_d <= lizzieLet17_5QNode_Int_7QNone_Int_8QError_Int_1QError_Int_d;
  QTree_Int_t lizzieLet17_5QNode_Int_7QNone_Int_8QError_Int_1QError_Int_bufchan_buf;
  assign lizzieLet17_5QNode_Int_7QNone_Int_8QError_Int_1QError_Int_bufchan_r = (! lizzieLet17_5QNode_Int_7QNone_Int_8QError_Int_1QError_Int_bufchan_buf[0]);
  assign lizzieLet47_1_argbuf_d = (lizzieLet17_5QNode_Int_7QNone_Int_8QError_Int_1QError_Int_bufchan_buf[0] ? lizzieLet17_5QNode_Int_7QNone_Int_8QError_Int_1QError_Int_bufchan_buf :
                                   lizzieLet17_5QNode_Int_7QNone_Int_8QError_Int_1QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNone_Int_8QError_Int_1QError_Int_bufchan_buf <= {66'd0,
                                                                                1'd0};
    else
      if ((lizzieLet47_1_argbuf_r && lizzieLet17_5QNode_Int_7QNone_Int_8QError_Int_1QError_Int_bufchan_buf[0]))
        lizzieLet17_5QNode_Int_7QNone_Int_8QError_Int_1QError_Int_bufchan_buf <= {66'd0,
                                                                                  1'd0};
      else if (((! lizzieLet47_1_argbuf_r) && (! lizzieLet17_5QNode_Int_7QNone_Int_8QError_Int_1QError_Int_bufchan_buf[0])))
        lizzieLet17_5QNode_Int_7QNone_Int_8QError_Int_1QError_Int_bufchan_buf <= lizzieLet17_5QNode_Int_7QNone_Int_8QError_Int_1QError_Int_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet17_5QNode_Int_7QNone_Int_8QError_Int_2,Go) > (lizzieLet17_5QNode_Int_7QNone_Int_8QError_Int_2_argbuf,Go) */
  Go_t lizzieLet17_5QNode_Int_7QNone_Int_8QError_Int_2_bufchan_d;
  logic lizzieLet17_5QNode_Int_7QNone_Int_8QError_Int_2_bufchan_r;
  assign lizzieLet17_5QNode_Int_7QNone_Int_8QError_Int_2_r = ((! lizzieLet17_5QNode_Int_7QNone_Int_8QError_Int_2_bufchan_d[0]) || lizzieLet17_5QNode_Int_7QNone_Int_8QError_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNone_Int_8QError_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet17_5QNode_Int_7QNone_Int_8QError_Int_2_r)
        lizzieLet17_5QNode_Int_7QNone_Int_8QError_Int_2_bufchan_d <= lizzieLet17_5QNode_Int_7QNone_Int_8QError_Int_2_d;
  Go_t lizzieLet17_5QNode_Int_7QNone_Int_8QError_Int_2_bufchan_buf;
  assign lizzieLet17_5QNode_Int_7QNone_Int_8QError_Int_2_bufchan_r = (! lizzieLet17_5QNode_Int_7QNone_Int_8QError_Int_2_bufchan_buf[0]);
  assign lizzieLet17_5QNode_Int_7QNone_Int_8QError_Int_2_argbuf_d = (lizzieLet17_5QNode_Int_7QNone_Int_8QError_Int_2_bufchan_buf[0] ? lizzieLet17_5QNode_Int_7QNone_Int_8QError_Int_2_bufchan_buf :
                                                                     lizzieLet17_5QNode_Int_7QNone_Int_8QError_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNone_Int_8QError_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet17_5QNode_Int_7QNone_Int_8QError_Int_2_argbuf_r && lizzieLet17_5QNode_Int_7QNone_Int_8QError_Int_2_bufchan_buf[0]))
        lizzieLet17_5QNode_Int_7QNone_Int_8QError_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet17_5QNode_Int_7QNone_Int_8QError_Int_2_argbuf_r) && (! lizzieLet17_5QNode_Int_7QNone_Int_8QError_Int_2_bufchan_buf[0])))
        lizzieLet17_5QNode_Int_7QNone_Int_8QError_Int_2_bufchan_buf <= lizzieLet17_5QNode_Int_7QNone_Int_8QError_Int_2_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int,Go) > [(lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_1,Go),
                                                                    (lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_2,Go),
                                                                    (lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_3,Go),
                                                                    (lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_4,Go),
                                                                    (lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_5,Go)] */
  logic [4:0] lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_emitted;
  logic [4:0] lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_done;
  assign lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_1_d = (lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_d[0] && (! lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_emitted[0]));
  assign lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_2_d = (lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_d[0] && (! lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_emitted[1]));
  assign lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_3_d = (lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_d[0] && (! lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_emitted[2]));
  assign lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_4_d = (lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_d[0] && (! lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_emitted[3]));
  assign lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_5_d = (lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_d[0] && (! lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_emitted[4]));
  assign lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_done = (lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_emitted | ({lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_5_d[0],
                                                                                                                       lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_4_d[0],
                                                                                                                       lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_3_d[0],
                                                                                                                       lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_2_d[0],
                                                                                                                       lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_1_d[0]} & {lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_5_r,
                                                                                                                                                                               lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_4_r,
                                                                                                                                                                               lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_3_r,
                                                                                                                                                                               lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_2_r,
                                                                                                                                                                               lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_1_r}));
  assign lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_r = (& lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_emitted <= 5'd0;
    else
      lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_emitted <= (lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_r ? 5'd0 :
                                                               lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_done);
  
  /* buf (Ty Go) : (lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_1,Go) > (lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_1_argbuf,Go) */
  Go_t lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_1_bufchan_d;
  logic lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_1_bufchan_r;
  assign lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_1_r = ((! lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_1_bufchan_d[0]) || lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_1_bufchan_d <= 1'd0;
    else
      if (lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_1_r)
        lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_1_bufchan_d <= lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_1_d;
  Go_t lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_1_bufchan_buf;
  assign lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_1_bufchan_r = (! lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_1_bufchan_buf[0]);
  assign lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_1_argbuf_d = (lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_1_bufchan_buf[0] ? lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_1_bufchan_buf :
                                                                    lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_1_argbuf_r && lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_1_bufchan_buf[0]))
        lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_1_argbuf_r) && (! lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_1_bufchan_buf[0])))
        lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_1_bufchan_buf <= lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_1_bufchan_d;
  
  /* dcon (Ty TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int,
      Dcon TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int) : [(lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_1_argbuf,Go),
                                                                                              (lizzieLet17_5QNode_Int_7QNone_Int_5QNode_Int_1_argbuf,Pointer_QTree_Int),
                                                                                              (t4af8_1_argbuf,Pointer_QTree_Int),
                                                                                              (lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_1_argbuf,MyDTInt_Bool),
                                                                                              (lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_1_argbuf,MyDTInt_Int_Int)] > (f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int5,TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int) */
  assign \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int5_d  = TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_dc((& {lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_1_argbuf_d[0],
                                                                                                                                                                                                                    lizzieLet17_5QNode_Int_7QNone_Int_5QNode_Int_1_argbuf_d[0],
                                                                                                                                                                                                                    t4af8_1_argbuf_d[0],
                                                                                                                                                                                                                    lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_1_argbuf_d[0],
                                                                                                                                                                                                                    lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_1_argbuf_d[0]}), lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_1_argbuf_d, lizzieLet17_5QNode_Int_7QNone_Int_5QNode_Int_1_argbuf_d, t4af8_1_argbuf_d, lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_1_argbuf_d, lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_1_argbuf_d);
  assign {lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_1_argbuf_r,
          lizzieLet17_5QNode_Int_7QNone_Int_5QNode_Int_1_argbuf_r,
          t4af8_1_argbuf_r,
          lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_1_argbuf_r,
          lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_1_argbuf_r} = {5 {(\f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int5_r  && \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int5_d [0])}};
  
  /* buf (Ty Go) : (lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_2,Go) > (lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_2_argbuf,Go) */
  Go_t lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_2_bufchan_d;
  logic lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_2_bufchan_r;
  assign lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_2_r = ((! lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_2_bufchan_d[0]) || lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_2_r)
        lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_2_bufchan_d <= lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_2_d;
  Go_t lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_2_bufchan_buf;
  assign lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_2_bufchan_r = (! lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_2_bufchan_buf[0]);
  assign lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_2_argbuf_d = (lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_2_bufchan_buf[0] ? lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_2_bufchan_buf :
                                                                    lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_2_argbuf_r && lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_2_bufchan_buf[0]))
        lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_2_argbuf_r) && (! lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_2_bufchan_buf[0])))
        lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_2_bufchan_buf <= lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_2_bufchan_d;
  
  /* dcon (Ty TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int,
      Dcon TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int) : [(lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_2_argbuf,Go),
                                                                                              (lizzieLet17_5QNode_Int_7QNone_Int_4QNode_Int_1_argbuf,Pointer_QTree_Int),
                                                                                              (t3af7_1_argbuf,Pointer_QTree_Int),
                                                                                              (lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_2_argbuf,MyDTInt_Bool),
                                                                                              (lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_2_argbuf,MyDTInt_Int_Int)] > (f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int6,TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int) */
  assign \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int6_d  = TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_dc((& {lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_2_argbuf_d[0],
                                                                                                                                                                                                                    lizzieLet17_5QNode_Int_7QNone_Int_4QNode_Int_1_argbuf_d[0],
                                                                                                                                                                                                                    t3af7_1_argbuf_d[0],
                                                                                                                                                                                                                    lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_2_argbuf_d[0],
                                                                                                                                                                                                                    lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_2_argbuf_d[0]}), lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_2_argbuf_d, lizzieLet17_5QNode_Int_7QNone_Int_4QNode_Int_1_argbuf_d, t3af7_1_argbuf_d, lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_2_argbuf_d, lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_2_argbuf_d);
  assign {lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_2_argbuf_r,
          lizzieLet17_5QNode_Int_7QNone_Int_4QNode_Int_1_argbuf_r,
          t3af7_1_argbuf_r,
          lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_2_argbuf_r,
          lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_2_argbuf_r} = {5 {(\f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int6_r  && \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int6_d [0])}};
  
  /* buf (Ty Go) : (lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_3,Go) > (lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_3_argbuf,Go) */
  Go_t lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_3_bufchan_d;
  logic lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_3_bufchan_r;
  assign lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_3_r = ((! lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_3_bufchan_d[0]) || lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_3_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_3_bufchan_d <= 1'd0;
    else
      if (lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_3_r)
        lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_3_bufchan_d <= lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_3_d;
  Go_t lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_3_bufchan_buf;
  assign lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_3_bufchan_r = (! lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_3_bufchan_buf[0]);
  assign lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_3_argbuf_d = (lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_3_bufchan_buf[0] ? lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_3_bufchan_buf :
                                                                    lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_3_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_3_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_3_argbuf_r && lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_3_bufchan_buf[0]))
        lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_3_bufchan_buf <= 1'd0;
      else if (((! lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_3_argbuf_r) && (! lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_3_bufchan_buf[0])))
        lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_3_bufchan_buf <= lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_3_bufchan_d;
  
  /* dcon (Ty TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int,
      Dcon TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int) : [(lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_3_argbuf,Go),
                                                                                              (lizzieLet17_5QNode_Int_7QNone_Int_3QNode_Int_1_argbuf,Pointer_QTree_Int),
                                                                                              (t2af6_1_argbuf,Pointer_QTree_Int),
                                                                                              (lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_3_argbuf,MyDTInt_Bool),
                                                                                              (lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_3_argbuf,MyDTInt_Int_Int)] > (f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int7,TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int) */
  assign \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int7_d  = TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_dc((& {lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_3_argbuf_d[0],
                                                                                                                                                                                                                    lizzieLet17_5QNode_Int_7QNone_Int_3QNode_Int_1_argbuf_d[0],
                                                                                                                                                                                                                    t2af6_1_argbuf_d[0],
                                                                                                                                                                                                                    lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_3_argbuf_d[0],
                                                                                                                                                                                                                    lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_3_argbuf_d[0]}), lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_3_argbuf_d, lizzieLet17_5QNode_Int_7QNone_Int_3QNode_Int_1_argbuf_d, t2af6_1_argbuf_d, lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_3_argbuf_d, lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_3_argbuf_d);
  assign {lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_3_argbuf_r,
          lizzieLet17_5QNode_Int_7QNone_Int_3QNode_Int_1_argbuf_r,
          t2af6_1_argbuf_r,
          lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_3_argbuf_r,
          lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_3_argbuf_r} = {5 {(\f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int7_r  && \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int7_d [0])}};
  
  /* buf (Ty Go) : (lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_4,Go) > (lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_4_argbuf,Go) */
  Go_t lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_4_bufchan_d;
  logic lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_4_bufchan_r;
  assign lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_4_r = ((! lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_4_bufchan_d[0]) || lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_4_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_4_bufchan_d <= 1'd0;
    else
      if (lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_4_r)
        lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_4_bufchan_d <= lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_4_d;
  Go_t lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_4_bufchan_buf;
  assign lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_4_bufchan_r = (! lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_4_bufchan_buf[0]);
  assign lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_4_argbuf_d = (lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_4_bufchan_buf[0] ? lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_4_bufchan_buf :
                                                                    lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_4_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_4_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_4_argbuf_r && lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_4_bufchan_buf[0]))
        lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_4_bufchan_buf <= 1'd0;
      else if (((! lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_4_argbuf_r) && (! lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_4_bufchan_buf[0])))
        lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_4_bufchan_buf <= lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_4_bufchan_d;
  
  /* dcon (Ty TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int,
      Dcon TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int) : [(lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_4_argbuf,Go),
                                                                                              (lizzieLet17_5QNode_Int_7QNone_Int_11QNode_Int_1_argbuf,Pointer_QTree_Int),
                                                                                              (t1af5_1_argbuf,Pointer_QTree_Int),
                                                                                              (lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_4_argbuf,MyDTInt_Bool),
                                                                                              (lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_4_argbuf,MyDTInt_Int_Int)] > (f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int8,TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int) */
  assign \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int8_d  = TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_dc((& {lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_4_argbuf_d[0],
                                                                                                                                                                                                                    lizzieLet17_5QNode_Int_7QNone_Int_11QNode_Int_1_argbuf_d[0],
                                                                                                                                                                                                                    t1af5_1_argbuf_d[0],
                                                                                                                                                                                                                    lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_4_argbuf_d[0],
                                                                                                                                                                                                                    lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_4_argbuf_d[0]}), lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_4_argbuf_d, lizzieLet17_5QNode_Int_7QNone_Int_11QNode_Int_1_argbuf_d, t1af5_1_argbuf_d, lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_4_argbuf_d, lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_4_argbuf_d);
  assign {lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_4_argbuf_r,
          lizzieLet17_5QNode_Int_7QNone_Int_11QNode_Int_1_argbuf_r,
          t1af5_1_argbuf_r,
          lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_4_argbuf_r,
          lizzieLet17_5QNode_Int_7QNone_Int_6QNode_Int_4_argbuf_r} = {5 {(\f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int8_r  && \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int8_d [0])}};
  
  /* buf (Ty Go) : (lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_5,Go) > (lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_5_argbuf,Go) */
  Go_t lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_5_bufchan_d;
  logic lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_5_bufchan_r;
  assign lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_5_r = ((! lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_5_bufchan_d[0]) || lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_5_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_5_bufchan_d <= 1'd0;
    else
      if (lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_5_r)
        lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_5_bufchan_d <= lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_5_d;
  Go_t lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_5_bufchan_buf;
  assign lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_5_bufchan_r = (! lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_5_bufchan_buf[0]);
  assign lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_5_argbuf_d = (lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_5_bufchan_buf[0] ? lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_5_bufchan_buf :
                                                                    lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_5_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_5_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_5_argbuf_r && lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_5_bufchan_buf[0]))
        lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_5_bufchan_buf <= 1'd0;
      else if (((! lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_5_argbuf_r) && (! lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_5_bufchan_buf[0])))
        lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_5_bufchan_buf <= lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_5_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet17_5QNode_Int_7QNone_Int_8QNone_Int,Go) > (lizzieLet17_5QNode_Int_7QNone_Int_8QNone_Int_1_argbuf,Go) */
  Go_t lizzieLet17_5QNode_Int_7QNone_Int_8QNone_Int_bufchan_d;
  logic lizzieLet17_5QNode_Int_7QNone_Int_8QNone_Int_bufchan_r;
  assign lizzieLet17_5QNode_Int_7QNone_Int_8QNone_Int_r = ((! lizzieLet17_5QNode_Int_7QNone_Int_8QNone_Int_bufchan_d[0]) || lizzieLet17_5QNode_Int_7QNone_Int_8QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNone_Int_8QNone_Int_bufchan_d <= 1'd0;
    else
      if (lizzieLet17_5QNode_Int_7QNone_Int_8QNone_Int_r)
        lizzieLet17_5QNode_Int_7QNone_Int_8QNone_Int_bufchan_d <= lizzieLet17_5QNode_Int_7QNone_Int_8QNone_Int_d;
  Go_t lizzieLet17_5QNode_Int_7QNone_Int_8QNone_Int_bufchan_buf;
  assign lizzieLet17_5QNode_Int_7QNone_Int_8QNone_Int_bufchan_r = (! lizzieLet17_5QNode_Int_7QNone_Int_8QNone_Int_bufchan_buf[0]);
  assign lizzieLet17_5QNode_Int_7QNone_Int_8QNone_Int_1_argbuf_d = (lizzieLet17_5QNode_Int_7QNone_Int_8QNone_Int_bufchan_buf[0] ? lizzieLet17_5QNode_Int_7QNone_Int_8QNone_Int_bufchan_buf :
                                                                    lizzieLet17_5QNode_Int_7QNone_Int_8QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNone_Int_8QNone_Int_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet17_5QNode_Int_7QNone_Int_8QNone_Int_1_argbuf_r && lizzieLet17_5QNode_Int_7QNone_Int_8QNone_Int_bufchan_buf[0]))
        lizzieLet17_5QNode_Int_7QNone_Int_8QNone_Int_bufchan_buf <= 1'd0;
      else if (((! lizzieLet17_5QNode_Int_7QNone_Int_8QNone_Int_1_argbuf_r) && (! lizzieLet17_5QNode_Int_7QNone_Int_8QNone_Int_bufchan_buf[0])))
        lizzieLet17_5QNode_Int_7QNone_Int_8QNone_Int_bufchan_buf <= lizzieLet17_5QNode_Int_7QNone_Int_8QNone_Int_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet17_5QNode_Int_7QNone_Int_8QVal_Int,Go) > [(lizzieLet17_5QNode_Int_7QNone_Int_8QVal_Int_1,Go),
                                                                   (lizzieLet17_5QNode_Int_7QNone_Int_8QVal_Int_2,Go)] */
  logic [1:0] lizzieLet17_5QNode_Int_7QNone_Int_8QVal_Int_emitted;
  logic [1:0] lizzieLet17_5QNode_Int_7QNone_Int_8QVal_Int_done;
  assign lizzieLet17_5QNode_Int_7QNone_Int_8QVal_Int_1_d = (lizzieLet17_5QNode_Int_7QNone_Int_8QVal_Int_d[0] && (! lizzieLet17_5QNode_Int_7QNone_Int_8QVal_Int_emitted[0]));
  assign lizzieLet17_5QNode_Int_7QNone_Int_8QVal_Int_2_d = (lizzieLet17_5QNode_Int_7QNone_Int_8QVal_Int_d[0] && (! lizzieLet17_5QNode_Int_7QNone_Int_8QVal_Int_emitted[1]));
  assign lizzieLet17_5QNode_Int_7QNone_Int_8QVal_Int_done = (lizzieLet17_5QNode_Int_7QNone_Int_8QVal_Int_emitted | ({lizzieLet17_5QNode_Int_7QNone_Int_8QVal_Int_2_d[0],
                                                                                                                     lizzieLet17_5QNode_Int_7QNone_Int_8QVal_Int_1_d[0]} & {lizzieLet17_5QNode_Int_7QNone_Int_8QVal_Int_2_r,
                                                                                                                                                                            lizzieLet17_5QNode_Int_7QNone_Int_8QVal_Int_1_r}));
  assign lizzieLet17_5QNode_Int_7QNone_Int_8QVal_Int_r = (& lizzieLet17_5QNode_Int_7QNone_Int_8QVal_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNone_Int_8QVal_Int_emitted <= 2'd0;
    else
      lizzieLet17_5QNode_Int_7QNone_Int_8QVal_Int_emitted <= (lizzieLet17_5QNode_Int_7QNone_Int_8QVal_Int_r ? 2'd0 :
                                                              lizzieLet17_5QNode_Int_7QNone_Int_8QVal_Int_done);
  
  /* dcon (Ty QTree_Int,
      Dcon QError_Int) : [(lizzieLet17_5QNode_Int_7QNone_Int_8QVal_Int_1,Go)] > (lizzieLet17_5QNode_Int_7QNone_Int_8QVal_Int_1QError_Int,QTree_Int) */
  assign lizzieLet17_5QNode_Int_7QNone_Int_8QVal_Int_1QError_Int_d = QError_Int_dc((& {lizzieLet17_5QNode_Int_7QNone_Int_8QVal_Int_1_d[0]}), lizzieLet17_5QNode_Int_7QNone_Int_8QVal_Int_1_d);
  assign {lizzieLet17_5QNode_Int_7QNone_Int_8QVal_Int_1_r} = {1 {(lizzieLet17_5QNode_Int_7QNone_Int_8QVal_Int_1QError_Int_r && lizzieLet17_5QNode_Int_7QNone_Int_8QVal_Int_1QError_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (lizzieLet17_5QNode_Int_7QNone_Int_8QVal_Int_1QError_Int,QTree_Int) > (lizzieLet45_1_argbuf,QTree_Int) */
  QTree_Int_t lizzieLet17_5QNode_Int_7QNone_Int_8QVal_Int_1QError_Int_bufchan_d;
  logic lizzieLet17_5QNode_Int_7QNone_Int_8QVal_Int_1QError_Int_bufchan_r;
  assign lizzieLet17_5QNode_Int_7QNone_Int_8QVal_Int_1QError_Int_r = ((! lizzieLet17_5QNode_Int_7QNone_Int_8QVal_Int_1QError_Int_bufchan_d[0]) || lizzieLet17_5QNode_Int_7QNone_Int_8QVal_Int_1QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNone_Int_8QVal_Int_1QError_Int_bufchan_d <= {66'd0,
                                                                            1'd0};
    else
      if (lizzieLet17_5QNode_Int_7QNone_Int_8QVal_Int_1QError_Int_r)
        lizzieLet17_5QNode_Int_7QNone_Int_8QVal_Int_1QError_Int_bufchan_d <= lizzieLet17_5QNode_Int_7QNone_Int_8QVal_Int_1QError_Int_d;
  QTree_Int_t lizzieLet17_5QNode_Int_7QNone_Int_8QVal_Int_1QError_Int_bufchan_buf;
  assign lizzieLet17_5QNode_Int_7QNone_Int_8QVal_Int_1QError_Int_bufchan_r = (! lizzieLet17_5QNode_Int_7QNone_Int_8QVal_Int_1QError_Int_bufchan_buf[0]);
  assign lizzieLet45_1_argbuf_d = (lizzieLet17_5QNode_Int_7QNone_Int_8QVal_Int_1QError_Int_bufchan_buf[0] ? lizzieLet17_5QNode_Int_7QNone_Int_8QVal_Int_1QError_Int_bufchan_buf :
                                   lizzieLet17_5QNode_Int_7QNone_Int_8QVal_Int_1QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNone_Int_8QVal_Int_1QError_Int_bufchan_buf <= {66'd0,
                                                                              1'd0};
    else
      if ((lizzieLet45_1_argbuf_r && lizzieLet17_5QNode_Int_7QNone_Int_8QVal_Int_1QError_Int_bufchan_buf[0]))
        lizzieLet17_5QNode_Int_7QNone_Int_8QVal_Int_1QError_Int_bufchan_buf <= {66'd0,
                                                                                1'd0};
      else if (((! lizzieLet45_1_argbuf_r) && (! lizzieLet17_5QNode_Int_7QNone_Int_8QVal_Int_1QError_Int_bufchan_buf[0])))
        lizzieLet17_5QNode_Int_7QNone_Int_8QVal_Int_1QError_Int_bufchan_buf <= lizzieLet17_5QNode_Int_7QNone_Int_8QVal_Int_1QError_Int_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet17_5QNode_Int_7QNone_Int_8QVal_Int_2,Go) > (lizzieLet17_5QNode_Int_7QNone_Int_8QVal_Int_2_argbuf,Go) */
  Go_t lizzieLet17_5QNode_Int_7QNone_Int_8QVal_Int_2_bufchan_d;
  logic lizzieLet17_5QNode_Int_7QNone_Int_8QVal_Int_2_bufchan_r;
  assign lizzieLet17_5QNode_Int_7QNone_Int_8QVal_Int_2_r = ((! lizzieLet17_5QNode_Int_7QNone_Int_8QVal_Int_2_bufchan_d[0]) || lizzieLet17_5QNode_Int_7QNone_Int_8QVal_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNone_Int_8QVal_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet17_5QNode_Int_7QNone_Int_8QVal_Int_2_r)
        lizzieLet17_5QNode_Int_7QNone_Int_8QVal_Int_2_bufchan_d <= lizzieLet17_5QNode_Int_7QNone_Int_8QVal_Int_2_d;
  Go_t lizzieLet17_5QNode_Int_7QNone_Int_8QVal_Int_2_bufchan_buf;
  assign lizzieLet17_5QNode_Int_7QNone_Int_8QVal_Int_2_bufchan_r = (! lizzieLet17_5QNode_Int_7QNone_Int_8QVal_Int_2_bufchan_buf[0]);
  assign lizzieLet17_5QNode_Int_7QNone_Int_8QVal_Int_2_argbuf_d = (lizzieLet17_5QNode_Int_7QNone_Int_8QVal_Int_2_bufchan_buf[0] ? lizzieLet17_5QNode_Int_7QNone_Int_8QVal_Int_2_bufchan_buf :
                                                                   lizzieLet17_5QNode_Int_7QNone_Int_8QVal_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNone_Int_8QVal_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet17_5QNode_Int_7QNone_Int_8QVal_Int_2_argbuf_r && lizzieLet17_5QNode_Int_7QNone_Int_8QVal_Int_2_bufchan_buf[0]))
        lizzieLet17_5QNode_Int_7QNone_Int_8QVal_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet17_5QNode_Int_7QNone_Int_8QVal_Int_2_argbuf_r) && (! lizzieLet17_5QNode_Int_7QNone_Int_8QVal_Int_2_bufchan_buf[0])))
        lizzieLet17_5QNode_Int_7QNone_Int_8QVal_Int_2_bufchan_buf <= lizzieLet17_5QNode_Int_7QNone_Int_8QVal_Int_2_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty MyDTInt_Bool) : (lizzieLet17_5QNode_Int_7QNone_Int_9,QTree_Int) (lizzieLet17_5QNode_Int_6QNone_Int,MyDTInt_Bool) > [(_160,MyDTInt_Bool),
                                                                                                                              (_159,MyDTInt_Bool),
                                                                                                                              (lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int,MyDTInt_Bool),
                                                                                                                              (_158,MyDTInt_Bool)] */
  logic [3:0] lizzieLet17_5QNode_Int_6QNone_Int_onehotd;
  always_comb
    if ((lizzieLet17_5QNode_Int_7QNone_Int_9_d[0] && lizzieLet17_5QNode_Int_6QNone_Int_d[0]))
      unique case (lizzieLet17_5QNode_Int_7QNone_Int_9_d[2:1])
        2'd0: lizzieLet17_5QNode_Int_6QNone_Int_onehotd = 4'd1;
        2'd1: lizzieLet17_5QNode_Int_6QNone_Int_onehotd = 4'd2;
        2'd2: lizzieLet17_5QNode_Int_6QNone_Int_onehotd = 4'd4;
        2'd3: lizzieLet17_5QNode_Int_6QNone_Int_onehotd = 4'd8;
        default: lizzieLet17_5QNode_Int_6QNone_Int_onehotd = 4'd0;
      endcase
    else lizzieLet17_5QNode_Int_6QNone_Int_onehotd = 4'd0;
  assign _160_d = lizzieLet17_5QNode_Int_6QNone_Int_onehotd[0];
  assign _159_d = lizzieLet17_5QNode_Int_6QNone_Int_onehotd[1];
  assign lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_d = lizzieLet17_5QNode_Int_6QNone_Int_onehotd[2];
  assign _158_d = lizzieLet17_5QNode_Int_6QNone_Int_onehotd[3];
  assign lizzieLet17_5QNode_Int_6QNone_Int_r = (| (lizzieLet17_5QNode_Int_6QNone_Int_onehotd & {_158_r,
                                                                                                lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_r,
                                                                                                _159_r,
                                                                                                _160_r}));
  assign lizzieLet17_5QNode_Int_7QNone_Int_9_r = lizzieLet17_5QNode_Int_6QNone_Int_r;
  
  /* fork (Ty MyDTInt_Bool) : (lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int,MyDTInt_Bool) > [(lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_1,MyDTInt_Bool),
                                                                                        (lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_2,MyDTInt_Bool),
                                                                                        (lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_3,MyDTInt_Bool),
                                                                                        (lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_4,MyDTInt_Bool)] */
  logic [3:0] lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_emitted;
  logic [3:0] lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_done;
  assign lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_1_d = (lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_d[0] && (! lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_emitted[0]));
  assign lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_2_d = (lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_d[0] && (! lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_emitted[1]));
  assign lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_3_d = (lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_d[0] && (! lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_emitted[2]));
  assign lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_4_d = (lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_d[0] && (! lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_emitted[3]));
  assign lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_done = (lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_emitted | ({lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_4_d[0],
                                                                                                                       lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_3_d[0],
                                                                                                                       lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_2_d[0],
                                                                                                                       lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_1_d[0]} & {lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_4_r,
                                                                                                                                                                               lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_3_r,
                                                                                                                                                                               lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_2_r,
                                                                                                                                                                               lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_1_r}));
  assign lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_r = (& lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_emitted <= 4'd0;
    else
      lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_emitted <= (lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_r ? 4'd0 :
                                                               lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_done);
  
  /* buf (Ty MyDTInt_Bool) : (lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_1,MyDTInt_Bool) > (lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_1_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_1_bufchan_d;
  logic lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_1_bufchan_r;
  assign lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_1_r = ((! lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_1_bufchan_d[0]) || lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_1_bufchan_d <= 1'd0;
    else
      if (lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_1_r)
        lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_1_bufchan_d <= lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_1_d;
  MyDTInt_Bool_t lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_1_bufchan_buf;
  assign lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_1_bufchan_r = (! lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_1_bufchan_buf[0]);
  assign lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_1_argbuf_d = (lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_1_bufchan_buf[0] ? lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_1_bufchan_buf :
                                                                    lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_1_argbuf_r && lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_1_bufchan_buf[0]))
        lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_1_argbuf_r) && (! lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_1_bufchan_buf[0])))
        lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_1_bufchan_buf <= lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_1_bufchan_d;
  
  /* buf (Ty MyDTInt_Bool) : (lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_2,MyDTInt_Bool) > (lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_2_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_2_bufchan_d;
  logic lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_2_bufchan_r;
  assign lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_2_r = ((! lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_2_bufchan_d[0]) || lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_2_r)
        lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_2_bufchan_d <= lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_2_d;
  MyDTInt_Bool_t lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_2_bufchan_buf;
  assign lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_2_bufchan_r = (! lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_2_bufchan_buf[0]);
  assign lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_2_argbuf_d = (lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_2_bufchan_buf[0] ? lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_2_bufchan_buf :
                                                                    lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_2_argbuf_r && lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_2_bufchan_buf[0]))
        lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_2_argbuf_r) && (! lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_2_bufchan_buf[0])))
        lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_2_bufchan_buf <= lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_2_bufchan_d;
  
  /* buf (Ty MyDTInt_Bool) : (lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_3,MyDTInt_Bool) > (lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_3_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_3_bufchan_d;
  logic lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_3_bufchan_r;
  assign lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_3_r = ((! lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_3_bufchan_d[0]) || lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_3_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_3_bufchan_d <= 1'd0;
    else
      if (lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_3_r)
        lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_3_bufchan_d <= lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_3_d;
  MyDTInt_Bool_t lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_3_bufchan_buf;
  assign lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_3_bufchan_r = (! lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_3_bufchan_buf[0]);
  assign lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_3_argbuf_d = (lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_3_bufchan_buf[0] ? lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_3_bufchan_buf :
                                                                    lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_3_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_3_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_3_argbuf_r && lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_3_bufchan_buf[0]))
        lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_3_bufchan_buf <= 1'd0;
      else if (((! lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_3_argbuf_r) && (! lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_3_bufchan_buf[0])))
        lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_3_bufchan_buf <= lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_3_bufchan_d;
  
  /* buf (Ty MyDTInt_Bool) : (lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_4,MyDTInt_Bool) > (lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_4_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_4_bufchan_d;
  logic lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_4_bufchan_r;
  assign lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_4_r = ((! lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_4_bufchan_d[0]) || lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_4_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_4_bufchan_d <= 1'd0;
    else
      if (lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_4_r)
        lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_4_bufchan_d <= lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_4_d;
  MyDTInt_Bool_t lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_4_bufchan_buf;
  assign lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_4_bufchan_r = (! lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_4_bufchan_buf[0]);
  assign lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_4_argbuf_d = (lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_4_bufchan_buf[0] ? lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_4_bufchan_buf :
                                                                    lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_4_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_4_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_4_argbuf_r && lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_4_bufchan_buf[0]))
        lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_4_bufchan_buf <= 1'd0;
      else if (((! lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_4_argbuf_r) && (! lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_4_bufchan_buf[0])))
        lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_4_bufchan_buf <= lizzieLet17_5QNode_Int_7QNone_Int_9QNode_Int_4_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_QTree_Int) : (lizzieLet17_5QNode_Int_8,QTree_Int) (lizzieLet17_7QNode_Int,Pointer_QTree_Int) > [(lizzieLet17_5QNode_Int_8QNone_Int,Pointer_QTree_Int),
                                                                                                                  (_157,Pointer_QTree_Int),
                                                                                                                  (_156,Pointer_QTree_Int),
                                                                                                                  (_155,Pointer_QTree_Int)] */
  logic [3:0] lizzieLet17_7QNode_Int_onehotd;
  always_comb
    if ((lizzieLet17_5QNode_Int_8_d[0] && lizzieLet17_7QNode_Int_d[0]))
      unique case (lizzieLet17_5QNode_Int_8_d[2:1])
        2'd0: lizzieLet17_7QNode_Int_onehotd = 4'd1;
        2'd1: lizzieLet17_7QNode_Int_onehotd = 4'd2;
        2'd2: lizzieLet17_7QNode_Int_onehotd = 4'd4;
        2'd3: lizzieLet17_7QNode_Int_onehotd = 4'd8;
        default: lizzieLet17_7QNode_Int_onehotd = 4'd0;
      endcase
    else lizzieLet17_7QNode_Int_onehotd = 4'd0;
  assign lizzieLet17_5QNode_Int_8QNone_Int_d = {lizzieLet17_7QNode_Int_d[16:1],
                                                lizzieLet17_7QNode_Int_onehotd[0]};
  assign _157_d = {lizzieLet17_7QNode_Int_d[16:1],
                   lizzieLet17_7QNode_Int_onehotd[1]};
  assign _156_d = {lizzieLet17_7QNode_Int_d[16:1],
                   lizzieLet17_7QNode_Int_onehotd[2]};
  assign _155_d = {lizzieLet17_7QNode_Int_d[16:1],
                   lizzieLet17_7QNode_Int_onehotd[3]};
  assign lizzieLet17_7QNode_Int_r = (| (lizzieLet17_7QNode_Int_onehotd & {_155_r,
                                                                          _156_r,
                                                                          _157_r,
                                                                          lizzieLet17_5QNode_Int_8QNone_Int_r}));
  assign lizzieLet17_5QNode_Int_8_r = lizzieLet17_7QNode_Int_r;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_QTree_Int) : (lizzieLet17_5QNode_Int_9,QTree_Int) (q1af0_destruct,Pointer_QTree_Int) > [(lizzieLet17_5QNode_Int_9QNone_Int,Pointer_QTree_Int),
                                                                                                          (_154,Pointer_QTree_Int),
                                                                                                          (lizzieLet17_5QNode_Int_9QNode_Int,Pointer_QTree_Int),
                                                                                                          (_153,Pointer_QTree_Int)] */
  logic [3:0] q1af0_destruct_onehotd;
  always_comb
    if ((lizzieLet17_5QNode_Int_9_d[0] && q1af0_destruct_d[0]))
      unique case (lizzieLet17_5QNode_Int_9_d[2:1])
        2'd0: q1af0_destruct_onehotd = 4'd1;
        2'd1: q1af0_destruct_onehotd = 4'd2;
        2'd2: q1af0_destruct_onehotd = 4'd4;
        2'd3: q1af0_destruct_onehotd = 4'd8;
        default: q1af0_destruct_onehotd = 4'd0;
      endcase
    else q1af0_destruct_onehotd = 4'd0;
  assign lizzieLet17_5QNode_Int_9QNone_Int_d = {q1af0_destruct_d[16:1],
                                                q1af0_destruct_onehotd[0]};
  assign _154_d = {q1af0_destruct_d[16:1],
                   q1af0_destruct_onehotd[1]};
  assign lizzieLet17_5QNode_Int_9QNode_Int_d = {q1af0_destruct_d[16:1],
                                                q1af0_destruct_onehotd[2]};
  assign _153_d = {q1af0_destruct_d[16:1],
                   q1af0_destruct_onehotd[3]};
  assign q1af0_destruct_r = (| (q1af0_destruct_onehotd & {_153_r,
                                                          lizzieLet17_5QNode_Int_9QNode_Int_r,
                                                          _154_r,
                                                          lizzieLet17_5QNode_Int_9QNone_Int_r}));
  assign lizzieLet17_5QNode_Int_9_r = q1af0_destruct_r;
  
  /* fork (Ty QTree_Int) : (lizzieLet17_5QNone_Int,QTree_Int) > [(lizzieLet17_5QNone_Int_1,QTree_Int),
                                                            (lizzieLet17_5QNone_Int_2,QTree_Int),
                                                            (lizzieLet17_5QNone_Int_3,QTree_Int),
                                                            (lizzieLet17_5QNone_Int_4,QTree_Int),
                                                            (lizzieLet17_5QNone_Int_5,QTree_Int),
                                                            (lizzieLet17_5QNone_Int_6,QTree_Int),
                                                            (lizzieLet17_5QNone_Int_7,QTree_Int),
                                                            (lizzieLet17_5QNone_Int_8,QTree_Int),
                                                            (lizzieLet17_5QNone_Int_9,QTree_Int)] */
  logic [8:0] lizzieLet17_5QNone_Int_emitted;
  logic [8:0] lizzieLet17_5QNone_Int_done;
  assign lizzieLet17_5QNone_Int_1_d = {lizzieLet17_5QNone_Int_d[66:1],
                                       (lizzieLet17_5QNone_Int_d[0] && (! lizzieLet17_5QNone_Int_emitted[0]))};
  assign lizzieLet17_5QNone_Int_2_d = {lizzieLet17_5QNone_Int_d[66:1],
                                       (lizzieLet17_5QNone_Int_d[0] && (! lizzieLet17_5QNone_Int_emitted[1]))};
  assign lizzieLet17_5QNone_Int_3_d = {lizzieLet17_5QNone_Int_d[66:1],
                                       (lizzieLet17_5QNone_Int_d[0] && (! lizzieLet17_5QNone_Int_emitted[2]))};
  assign lizzieLet17_5QNone_Int_4_d = {lizzieLet17_5QNone_Int_d[66:1],
                                       (lizzieLet17_5QNone_Int_d[0] && (! lizzieLet17_5QNone_Int_emitted[3]))};
  assign lizzieLet17_5QNone_Int_5_d = {lizzieLet17_5QNone_Int_d[66:1],
                                       (lizzieLet17_5QNone_Int_d[0] && (! lizzieLet17_5QNone_Int_emitted[4]))};
  assign lizzieLet17_5QNone_Int_6_d = {lizzieLet17_5QNone_Int_d[66:1],
                                       (lizzieLet17_5QNone_Int_d[0] && (! lizzieLet17_5QNone_Int_emitted[5]))};
  assign lizzieLet17_5QNone_Int_7_d = {lizzieLet17_5QNone_Int_d[66:1],
                                       (lizzieLet17_5QNone_Int_d[0] && (! lizzieLet17_5QNone_Int_emitted[6]))};
  assign lizzieLet17_5QNone_Int_8_d = {lizzieLet17_5QNone_Int_d[66:1],
                                       (lizzieLet17_5QNone_Int_d[0] && (! lizzieLet17_5QNone_Int_emitted[7]))};
  assign lizzieLet17_5QNone_Int_9_d = {lizzieLet17_5QNone_Int_d[66:1],
                                       (lizzieLet17_5QNone_Int_d[0] && (! lizzieLet17_5QNone_Int_emitted[8]))};
  assign lizzieLet17_5QNone_Int_done = (lizzieLet17_5QNone_Int_emitted | ({lizzieLet17_5QNone_Int_9_d[0],
                                                                           lizzieLet17_5QNone_Int_8_d[0],
                                                                           lizzieLet17_5QNone_Int_7_d[0],
                                                                           lizzieLet17_5QNone_Int_6_d[0],
                                                                           lizzieLet17_5QNone_Int_5_d[0],
                                                                           lizzieLet17_5QNone_Int_4_d[0],
                                                                           lizzieLet17_5QNone_Int_3_d[0],
                                                                           lizzieLet17_5QNone_Int_2_d[0],
                                                                           lizzieLet17_5QNone_Int_1_d[0]} & {lizzieLet17_5QNone_Int_9_r,
                                                                                                             lizzieLet17_5QNone_Int_8_r,
                                                                                                             lizzieLet17_5QNone_Int_7_r,
                                                                                                             lizzieLet17_5QNone_Int_6_r,
                                                                                                             lizzieLet17_5QNone_Int_5_r,
                                                                                                             lizzieLet17_5QNone_Int_4_r,
                                                                                                             lizzieLet17_5QNone_Int_3_r,
                                                                                                             lizzieLet17_5QNone_Int_2_r,
                                                                                                             lizzieLet17_5QNone_Int_1_r}));
  assign lizzieLet17_5QNone_Int_r = (& lizzieLet17_5QNone_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet17_5QNone_Int_emitted <= 9'd0;
    else
      lizzieLet17_5QNone_Int_emitted <= (lizzieLet17_5QNone_Int_r ? 9'd0 :
                                         lizzieLet17_5QNone_Int_done);
  
  /* destruct (Ty QTree_Int,
          Dcon QNode_Int) : (lizzieLet17_5QNone_Int_1QNode_Int,QTree_Int) > [(q1aeB_destruct,Pointer_QTree_Int),
                                                                             (q2aeC_destruct,Pointer_QTree_Int),
                                                                             (q3aeD_destruct,Pointer_QTree_Int),
                                                                             (q4aeE_destruct,Pointer_QTree_Int)] */
  logic [3:0] lizzieLet17_5QNone_Int_1QNode_Int_emitted;
  logic [3:0] lizzieLet17_5QNone_Int_1QNode_Int_done;
  assign q1aeB_destruct_d = {lizzieLet17_5QNone_Int_1QNode_Int_d[18:3],
                             (lizzieLet17_5QNone_Int_1QNode_Int_d[0] && (! lizzieLet17_5QNone_Int_1QNode_Int_emitted[0]))};
  assign q2aeC_destruct_d = {lizzieLet17_5QNone_Int_1QNode_Int_d[34:19],
                             (lizzieLet17_5QNone_Int_1QNode_Int_d[0] && (! lizzieLet17_5QNone_Int_1QNode_Int_emitted[1]))};
  assign q3aeD_destruct_d = {lizzieLet17_5QNone_Int_1QNode_Int_d[50:35],
                             (lizzieLet17_5QNone_Int_1QNode_Int_d[0] && (! lizzieLet17_5QNone_Int_1QNode_Int_emitted[2]))};
  assign q4aeE_destruct_d = {lizzieLet17_5QNone_Int_1QNode_Int_d[66:51],
                             (lizzieLet17_5QNone_Int_1QNode_Int_d[0] && (! lizzieLet17_5QNone_Int_1QNode_Int_emitted[3]))};
  assign lizzieLet17_5QNone_Int_1QNode_Int_done = (lizzieLet17_5QNone_Int_1QNode_Int_emitted | ({q4aeE_destruct_d[0],
                                                                                                 q3aeD_destruct_d[0],
                                                                                                 q2aeC_destruct_d[0],
                                                                                                 q1aeB_destruct_d[0]} & {q4aeE_destruct_r,
                                                                                                                         q3aeD_destruct_r,
                                                                                                                         q2aeC_destruct_r,
                                                                                                                         q1aeB_destruct_r}));
  assign lizzieLet17_5QNone_Int_1QNode_Int_r = (& lizzieLet17_5QNone_Int_1QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNone_Int_1QNode_Int_emitted <= 4'd0;
    else
      lizzieLet17_5QNone_Int_1QNode_Int_emitted <= (lizzieLet17_5QNone_Int_1QNode_Int_r ? 4'd0 :
                                                    lizzieLet17_5QNone_Int_1QNode_Int_done);
  
  /* destruct (Ty QTree_Int,
          Dcon QVal_Int) : (lizzieLet17_5QNone_Int_1QVal_Int,QTree_Int) > [(v1aev_destruct,Int)] */
  assign v1aev_destruct_d = {lizzieLet17_5QNone_Int_1QVal_Int_d[34:3],
                             lizzieLet17_5QNone_Int_1QVal_Int_d[0]};
  assign lizzieLet17_5QNone_Int_1QVal_Int_r = v1aev_destruct_r;
  
  /* demux (Ty QTree_Int,
       Ty QTree_Int) : (lizzieLet17_5QNone_Int_2,QTree_Int) (lizzieLet17_5QNone_Int_1,QTree_Int) > [(_152,QTree_Int),
                                                                                                    (lizzieLet17_5QNone_Int_1QVal_Int,QTree_Int),
                                                                                                    (lizzieLet17_5QNone_Int_1QNode_Int,QTree_Int),
                                                                                                    (_151,QTree_Int)] */
  logic [3:0] lizzieLet17_5QNone_Int_1_onehotd;
  always_comb
    if ((lizzieLet17_5QNone_Int_2_d[0] && lizzieLet17_5QNone_Int_1_d[0]))
      unique case (lizzieLet17_5QNone_Int_2_d[2:1])
        2'd0: lizzieLet17_5QNone_Int_1_onehotd = 4'd1;
        2'd1: lizzieLet17_5QNone_Int_1_onehotd = 4'd2;
        2'd2: lizzieLet17_5QNone_Int_1_onehotd = 4'd4;
        2'd3: lizzieLet17_5QNone_Int_1_onehotd = 4'd8;
        default: lizzieLet17_5QNone_Int_1_onehotd = 4'd0;
      endcase
    else lizzieLet17_5QNone_Int_1_onehotd = 4'd0;
  assign _152_d = {lizzieLet17_5QNone_Int_1_d[66:1],
                   lizzieLet17_5QNone_Int_1_onehotd[0]};
  assign lizzieLet17_5QNone_Int_1QVal_Int_d = {lizzieLet17_5QNone_Int_1_d[66:1],
                                               lizzieLet17_5QNone_Int_1_onehotd[1]};
  assign lizzieLet17_5QNone_Int_1QNode_Int_d = {lizzieLet17_5QNone_Int_1_d[66:1],
                                                lizzieLet17_5QNone_Int_1_onehotd[2]};
  assign _151_d = {lizzieLet17_5QNone_Int_1_d[66:1],
                   lizzieLet17_5QNone_Int_1_onehotd[3]};
  assign lizzieLet17_5QNone_Int_1_r = (| (lizzieLet17_5QNone_Int_1_onehotd & {_151_r,
                                                                              lizzieLet17_5QNone_Int_1QNode_Int_r,
                                                                              lizzieLet17_5QNone_Int_1QVal_Int_r,
                                                                              _152_r}));
  assign lizzieLet17_5QNone_Int_2_r = lizzieLet17_5QNone_Int_1_r;
  
  /* demux (Ty QTree_Int,
       Ty MyDTInt_Int_Int) : (lizzieLet17_5QNone_Int_3,QTree_Int) (lizzieLet17_10QNone_Int,MyDTInt_Int_Int) > [(_150,MyDTInt_Int_Int),
                                                                                                               (lizzieLet17_5QNone_Int_3QVal_Int,MyDTInt_Int_Int),
                                                                                                               (lizzieLet17_5QNone_Int_3QNode_Int,MyDTInt_Int_Int),
                                                                                                               (_149,MyDTInt_Int_Int)] */
  logic [3:0] lizzieLet17_10QNone_Int_onehotd;
  always_comb
    if ((lizzieLet17_5QNone_Int_3_d[0] && lizzieLet17_10QNone_Int_d[0]))
      unique case (lizzieLet17_5QNone_Int_3_d[2:1])
        2'd0: lizzieLet17_10QNone_Int_onehotd = 4'd1;
        2'd1: lizzieLet17_10QNone_Int_onehotd = 4'd2;
        2'd2: lizzieLet17_10QNone_Int_onehotd = 4'd4;
        2'd3: lizzieLet17_10QNone_Int_onehotd = 4'd8;
        default: lizzieLet17_10QNone_Int_onehotd = 4'd0;
      endcase
    else lizzieLet17_10QNone_Int_onehotd = 4'd0;
  assign _150_d = lizzieLet17_10QNone_Int_onehotd[0];
  assign lizzieLet17_5QNone_Int_3QVal_Int_d = lizzieLet17_10QNone_Int_onehotd[1];
  assign lizzieLet17_5QNone_Int_3QNode_Int_d = lizzieLet17_10QNone_Int_onehotd[2];
  assign _149_d = lizzieLet17_10QNone_Int_onehotd[3];
  assign lizzieLet17_10QNone_Int_r = (| (lizzieLet17_10QNone_Int_onehotd & {_149_r,
                                                                            lizzieLet17_5QNone_Int_3QNode_Int_r,
                                                                            lizzieLet17_5QNone_Int_3QVal_Int_r,
                                                                            _150_r}));
  assign lizzieLet17_5QNone_Int_3_r = lizzieLet17_10QNone_Int_r;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_CTf_f_Int) : (lizzieLet17_5QNone_Int_4,QTree_Int) (lizzieLet17_11QNone_Int,Pointer_CTf_f_Int) > [(lizzieLet17_5QNone_Int_4QNone_Int,Pointer_CTf_f_Int),
                                                                                                                   (lizzieLet17_5QNone_Int_4QVal_Int,Pointer_CTf_f_Int),
                                                                                                                   (lizzieLet17_5QNone_Int_4QNode_Int,Pointer_CTf_f_Int),
                                                                                                                   (lizzieLet17_5QNone_Int_4QError_Int,Pointer_CTf_f_Int)] */
  logic [3:0] lizzieLet17_11QNone_Int_onehotd;
  always_comb
    if ((lizzieLet17_5QNone_Int_4_d[0] && lizzieLet17_11QNone_Int_d[0]))
      unique case (lizzieLet17_5QNone_Int_4_d[2:1])
        2'd0: lizzieLet17_11QNone_Int_onehotd = 4'd1;
        2'd1: lizzieLet17_11QNone_Int_onehotd = 4'd2;
        2'd2: lizzieLet17_11QNone_Int_onehotd = 4'd4;
        2'd3: lizzieLet17_11QNone_Int_onehotd = 4'd8;
        default: lizzieLet17_11QNone_Int_onehotd = 4'd0;
      endcase
    else lizzieLet17_11QNone_Int_onehotd = 4'd0;
  assign lizzieLet17_5QNone_Int_4QNone_Int_d = {lizzieLet17_11QNone_Int_d[16:1],
                                                lizzieLet17_11QNone_Int_onehotd[0]};
  assign lizzieLet17_5QNone_Int_4QVal_Int_d = {lizzieLet17_11QNone_Int_d[16:1],
                                               lizzieLet17_11QNone_Int_onehotd[1]};
  assign lizzieLet17_5QNone_Int_4QNode_Int_d = {lizzieLet17_11QNone_Int_d[16:1],
                                                lizzieLet17_11QNone_Int_onehotd[2]};
  assign lizzieLet17_5QNone_Int_4QError_Int_d = {lizzieLet17_11QNone_Int_d[16:1],
                                                 lizzieLet17_11QNone_Int_onehotd[3]};
  assign lizzieLet17_11QNone_Int_r = (| (lizzieLet17_11QNone_Int_onehotd & {lizzieLet17_5QNone_Int_4QError_Int_r,
                                                                            lizzieLet17_5QNone_Int_4QNode_Int_r,
                                                                            lizzieLet17_5QNone_Int_4QVal_Int_r,
                                                                            lizzieLet17_5QNone_Int_4QNone_Int_r}));
  assign lizzieLet17_5QNone_Int_4_r = lizzieLet17_11QNone_Int_r;
  
  /* buf (Ty Pointer_CTf_f_Int) : (lizzieLet17_5QNone_Int_4QError_Int,Pointer_CTf_f_Int) > (lizzieLet17_5QNone_Int_4QError_Int_1_argbuf,Pointer_CTf_f_Int) */
  Pointer_CTf_f_Int_t lizzieLet17_5QNone_Int_4QError_Int_bufchan_d;
  logic lizzieLet17_5QNone_Int_4QError_Int_bufchan_r;
  assign lizzieLet17_5QNone_Int_4QError_Int_r = ((! lizzieLet17_5QNone_Int_4QError_Int_bufchan_d[0]) || lizzieLet17_5QNone_Int_4QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNone_Int_4QError_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet17_5QNone_Int_4QError_Int_r)
        lizzieLet17_5QNone_Int_4QError_Int_bufchan_d <= lizzieLet17_5QNone_Int_4QError_Int_d;
  Pointer_CTf_f_Int_t lizzieLet17_5QNone_Int_4QError_Int_bufchan_buf;
  assign lizzieLet17_5QNone_Int_4QError_Int_bufchan_r = (! lizzieLet17_5QNone_Int_4QError_Int_bufchan_buf[0]);
  assign lizzieLet17_5QNone_Int_4QError_Int_1_argbuf_d = (lizzieLet17_5QNone_Int_4QError_Int_bufchan_buf[0] ? lizzieLet17_5QNone_Int_4QError_Int_bufchan_buf :
                                                          lizzieLet17_5QNone_Int_4QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNone_Int_4QError_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet17_5QNone_Int_4QError_Int_1_argbuf_r && lizzieLet17_5QNone_Int_4QError_Int_bufchan_buf[0]))
        lizzieLet17_5QNone_Int_4QError_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet17_5QNone_Int_4QError_Int_1_argbuf_r) && (! lizzieLet17_5QNone_Int_4QError_Int_bufchan_buf[0])))
        lizzieLet17_5QNone_Int_4QError_Int_bufchan_buf <= lizzieLet17_5QNone_Int_4QError_Int_bufchan_d;
  
  /* buf (Ty Pointer_CTf_f_Int) : (lizzieLet17_5QNone_Int_4QNone_Int,Pointer_CTf_f_Int) > (lizzieLet17_5QNone_Int_4QNone_Int_1_argbuf,Pointer_CTf_f_Int) */
  Pointer_CTf_f_Int_t lizzieLet17_5QNone_Int_4QNone_Int_bufchan_d;
  logic lizzieLet17_5QNone_Int_4QNone_Int_bufchan_r;
  assign lizzieLet17_5QNone_Int_4QNone_Int_r = ((! lizzieLet17_5QNone_Int_4QNone_Int_bufchan_d[0]) || lizzieLet17_5QNone_Int_4QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNone_Int_4QNone_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet17_5QNone_Int_4QNone_Int_r)
        lizzieLet17_5QNone_Int_4QNone_Int_bufchan_d <= lizzieLet17_5QNone_Int_4QNone_Int_d;
  Pointer_CTf_f_Int_t lizzieLet17_5QNone_Int_4QNone_Int_bufchan_buf;
  assign lizzieLet17_5QNone_Int_4QNone_Int_bufchan_r = (! lizzieLet17_5QNone_Int_4QNone_Int_bufchan_buf[0]);
  assign lizzieLet17_5QNone_Int_4QNone_Int_1_argbuf_d = (lizzieLet17_5QNone_Int_4QNone_Int_bufchan_buf[0] ? lizzieLet17_5QNone_Int_4QNone_Int_bufchan_buf :
                                                         lizzieLet17_5QNone_Int_4QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNone_Int_4QNone_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet17_5QNone_Int_4QNone_Int_1_argbuf_r && lizzieLet17_5QNone_Int_4QNone_Int_bufchan_buf[0]))
        lizzieLet17_5QNone_Int_4QNone_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet17_5QNone_Int_4QNone_Int_1_argbuf_r) && (! lizzieLet17_5QNone_Int_4QNone_Int_bufchan_buf[0])))
        lizzieLet17_5QNone_Int_4QNone_Int_bufchan_buf <= lizzieLet17_5QNone_Int_4QNone_Int_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Go) : (lizzieLet17_5QNone_Int_5,QTree_Int) (lizzieLet17_3QNone_Int,Go) > [(lizzieLet17_5QNone_Int_5QNone_Int,Go),
                                                                                    (lizzieLet17_5QNone_Int_5QVal_Int,Go),
                                                                                    (lizzieLet17_5QNone_Int_5QNode_Int,Go),
                                                                                    (lizzieLet17_5QNone_Int_5QError_Int,Go)] */
  logic [3:0] lizzieLet17_3QNone_Int_onehotd;
  always_comb
    if ((lizzieLet17_5QNone_Int_5_d[0] && lizzieLet17_3QNone_Int_d[0]))
      unique case (lizzieLet17_5QNone_Int_5_d[2:1])
        2'd0: lizzieLet17_3QNone_Int_onehotd = 4'd1;
        2'd1: lizzieLet17_3QNone_Int_onehotd = 4'd2;
        2'd2: lizzieLet17_3QNone_Int_onehotd = 4'd4;
        2'd3: lizzieLet17_3QNone_Int_onehotd = 4'd8;
        default: lizzieLet17_3QNone_Int_onehotd = 4'd0;
      endcase
    else lizzieLet17_3QNone_Int_onehotd = 4'd0;
  assign lizzieLet17_5QNone_Int_5QNone_Int_d = lizzieLet17_3QNone_Int_onehotd[0];
  assign lizzieLet17_5QNone_Int_5QVal_Int_d = lizzieLet17_3QNone_Int_onehotd[1];
  assign lizzieLet17_5QNone_Int_5QNode_Int_d = lizzieLet17_3QNone_Int_onehotd[2];
  assign lizzieLet17_5QNone_Int_5QError_Int_d = lizzieLet17_3QNone_Int_onehotd[3];
  assign lizzieLet17_3QNone_Int_r = (| (lizzieLet17_3QNone_Int_onehotd & {lizzieLet17_5QNone_Int_5QError_Int_r,
                                                                          lizzieLet17_5QNone_Int_5QNode_Int_r,
                                                                          lizzieLet17_5QNone_Int_5QVal_Int_r,
                                                                          lizzieLet17_5QNone_Int_5QNone_Int_r}));
  assign lizzieLet17_5QNone_Int_5_r = lizzieLet17_3QNone_Int_r;
  
  /* fork (Ty Go) : (lizzieLet17_5QNone_Int_5QError_Int,Go) > [(lizzieLet17_5QNone_Int_5QError_Int_1,Go),
                                                          (lizzieLet17_5QNone_Int_5QError_Int_2,Go)] */
  logic [1:0] lizzieLet17_5QNone_Int_5QError_Int_emitted;
  logic [1:0] lizzieLet17_5QNone_Int_5QError_Int_done;
  assign lizzieLet17_5QNone_Int_5QError_Int_1_d = (lizzieLet17_5QNone_Int_5QError_Int_d[0] && (! lizzieLet17_5QNone_Int_5QError_Int_emitted[0]));
  assign lizzieLet17_5QNone_Int_5QError_Int_2_d = (lizzieLet17_5QNone_Int_5QError_Int_d[0] && (! lizzieLet17_5QNone_Int_5QError_Int_emitted[1]));
  assign lizzieLet17_5QNone_Int_5QError_Int_done = (lizzieLet17_5QNone_Int_5QError_Int_emitted | ({lizzieLet17_5QNone_Int_5QError_Int_2_d[0],
                                                                                                   lizzieLet17_5QNone_Int_5QError_Int_1_d[0]} & {lizzieLet17_5QNone_Int_5QError_Int_2_r,
                                                                                                                                                 lizzieLet17_5QNone_Int_5QError_Int_1_r}));
  assign lizzieLet17_5QNone_Int_5QError_Int_r = (& lizzieLet17_5QNone_Int_5QError_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNone_Int_5QError_Int_emitted <= 2'd0;
    else
      lizzieLet17_5QNone_Int_5QError_Int_emitted <= (lizzieLet17_5QNone_Int_5QError_Int_r ? 2'd0 :
                                                     lizzieLet17_5QNone_Int_5QError_Int_done);
  
  /* dcon (Ty QTree_Int,
      Dcon QError_Int) : [(lizzieLet17_5QNone_Int_5QError_Int_1,Go)] > (lizzieLet17_5QNone_Int_5QError_Int_1QError_Int,QTree_Int) */
  assign lizzieLet17_5QNone_Int_5QError_Int_1QError_Int_d = QError_Int_dc((& {lizzieLet17_5QNone_Int_5QError_Int_1_d[0]}), lizzieLet17_5QNone_Int_5QError_Int_1_d);
  assign {lizzieLet17_5QNone_Int_5QError_Int_1_r} = {1 {(lizzieLet17_5QNone_Int_5QError_Int_1QError_Int_r && lizzieLet17_5QNone_Int_5QError_Int_1QError_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (lizzieLet17_5QNone_Int_5QError_Int_1QError_Int,QTree_Int) > (lizzieLet28_1_argbuf,QTree_Int) */
  QTree_Int_t lizzieLet17_5QNone_Int_5QError_Int_1QError_Int_bufchan_d;
  logic lizzieLet17_5QNone_Int_5QError_Int_1QError_Int_bufchan_r;
  assign lizzieLet17_5QNone_Int_5QError_Int_1QError_Int_r = ((! lizzieLet17_5QNone_Int_5QError_Int_1QError_Int_bufchan_d[0]) || lizzieLet17_5QNone_Int_5QError_Int_1QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNone_Int_5QError_Int_1QError_Int_bufchan_d <= {66'd0,
                                                                   1'd0};
    else
      if (lizzieLet17_5QNone_Int_5QError_Int_1QError_Int_r)
        lizzieLet17_5QNone_Int_5QError_Int_1QError_Int_bufchan_d <= lizzieLet17_5QNone_Int_5QError_Int_1QError_Int_d;
  QTree_Int_t lizzieLet17_5QNone_Int_5QError_Int_1QError_Int_bufchan_buf;
  assign lizzieLet17_5QNone_Int_5QError_Int_1QError_Int_bufchan_r = (! lizzieLet17_5QNone_Int_5QError_Int_1QError_Int_bufchan_buf[0]);
  assign lizzieLet28_1_argbuf_d = (lizzieLet17_5QNone_Int_5QError_Int_1QError_Int_bufchan_buf[0] ? lizzieLet17_5QNone_Int_5QError_Int_1QError_Int_bufchan_buf :
                                   lizzieLet17_5QNone_Int_5QError_Int_1QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNone_Int_5QError_Int_1QError_Int_bufchan_buf <= {66'd0,
                                                                     1'd0};
    else
      if ((lizzieLet28_1_argbuf_r && lizzieLet17_5QNone_Int_5QError_Int_1QError_Int_bufchan_buf[0]))
        lizzieLet17_5QNone_Int_5QError_Int_1QError_Int_bufchan_buf <= {66'd0,
                                                                       1'd0};
      else if (((! lizzieLet28_1_argbuf_r) && (! lizzieLet17_5QNone_Int_5QError_Int_1QError_Int_bufchan_buf[0])))
        lizzieLet17_5QNone_Int_5QError_Int_1QError_Int_bufchan_buf <= lizzieLet17_5QNone_Int_5QError_Int_1QError_Int_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet17_5QNone_Int_5QError_Int_2,Go) > (lizzieLet17_5QNone_Int_5QError_Int_2_argbuf,Go) */
  Go_t lizzieLet17_5QNone_Int_5QError_Int_2_bufchan_d;
  logic lizzieLet17_5QNone_Int_5QError_Int_2_bufchan_r;
  assign lizzieLet17_5QNone_Int_5QError_Int_2_r = ((! lizzieLet17_5QNone_Int_5QError_Int_2_bufchan_d[0]) || lizzieLet17_5QNone_Int_5QError_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNone_Int_5QError_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet17_5QNone_Int_5QError_Int_2_r)
        lizzieLet17_5QNone_Int_5QError_Int_2_bufchan_d <= lizzieLet17_5QNone_Int_5QError_Int_2_d;
  Go_t lizzieLet17_5QNone_Int_5QError_Int_2_bufchan_buf;
  assign lizzieLet17_5QNone_Int_5QError_Int_2_bufchan_r = (! lizzieLet17_5QNone_Int_5QError_Int_2_bufchan_buf[0]);
  assign lizzieLet17_5QNone_Int_5QError_Int_2_argbuf_d = (lizzieLet17_5QNone_Int_5QError_Int_2_bufchan_buf[0] ? lizzieLet17_5QNone_Int_5QError_Int_2_bufchan_buf :
                                                          lizzieLet17_5QNone_Int_5QError_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNone_Int_5QError_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet17_5QNone_Int_5QError_Int_2_argbuf_r && lizzieLet17_5QNone_Int_5QError_Int_2_bufchan_buf[0]))
        lizzieLet17_5QNone_Int_5QError_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet17_5QNone_Int_5QError_Int_2_argbuf_r) && (! lizzieLet17_5QNone_Int_5QError_Int_2_bufchan_buf[0])))
        lizzieLet17_5QNone_Int_5QError_Int_2_bufchan_buf <= lizzieLet17_5QNone_Int_5QError_Int_2_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet17_5QNone_Int_5QNone_Int,Go) > (lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf,Go) */
  Go_t lizzieLet17_5QNone_Int_5QNone_Int_bufchan_d;
  logic lizzieLet17_5QNone_Int_5QNone_Int_bufchan_r;
  assign lizzieLet17_5QNone_Int_5QNone_Int_r = ((! lizzieLet17_5QNone_Int_5QNone_Int_bufchan_d[0]) || lizzieLet17_5QNone_Int_5QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNone_Int_5QNone_Int_bufchan_d <= 1'd0;
    else
      if (lizzieLet17_5QNone_Int_5QNone_Int_r)
        lizzieLet17_5QNone_Int_5QNone_Int_bufchan_d <= lizzieLet17_5QNone_Int_5QNone_Int_d;
  Go_t lizzieLet17_5QNone_Int_5QNone_Int_bufchan_buf;
  assign lizzieLet17_5QNone_Int_5QNone_Int_bufchan_r = (! lizzieLet17_5QNone_Int_5QNone_Int_bufchan_buf[0]);
  assign lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_d = (lizzieLet17_5QNone_Int_5QNone_Int_bufchan_buf[0] ? lizzieLet17_5QNone_Int_5QNone_Int_bufchan_buf :
                                                         lizzieLet17_5QNone_Int_5QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNone_Int_5QNone_Int_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_r && lizzieLet17_5QNone_Int_5QNone_Int_bufchan_buf[0]))
        lizzieLet17_5QNone_Int_5QNone_Int_bufchan_buf <= 1'd0;
      else if (((! lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_r) && (! lizzieLet17_5QNone_Int_5QNone_Int_bufchan_buf[0])))
        lizzieLet17_5QNone_Int_5QNone_Int_bufchan_buf <= lizzieLet17_5QNone_Int_5QNone_Int_bufchan_d;
  
  /* mergectrl (Ty C35,
           Ty Go) : [(lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf,Go),
                     (lizzieLet67_3Lcall_f_f_Int0_1_argbuf,Go),
                     (lizzieLet17_5QNone_Int_7QVal_Int_5QNone_Int_1_argbuf,Go),
                     (es_2_1_3MyFalse_1_argbuf,Go),
                     (es_2_1_3MyTrue_2_argbuf,Go),
                     (lizzieLet17_5QNone_Int_7QVal_Int_5QNode_Int_2_argbuf,Go),
                     (lizzieLet17_5QNone_Int_7QVal_Int_5QError_Int_2_argbuf,Go),
                     (lizzieLet17_5QNone_Int_7QNode_Int_5QNone_Int_1_argbuf,Go),
                     (lizzieLet17_5QNone_Int_7QNode_Int_5QVal_Int_2_argbuf,Go),
                     (lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_5_argbuf,Go),
                     (lizzieLet17_5QNone_Int_7QNode_Int_5QError_Int_2_argbuf,Go),
                     (lizzieLet17_5QNone_Int_5QError_Int_2_argbuf,Go),
                     (lizzieLet17_5QVal_Int_7QNone_Int_6QNone_Int_1_argbuf,Go),
                     (es_10_4MyFalse_1_argbuf,Go),
                     (es_10_4MyTrue_2_argbuf,Go),
                     (lizzieLet17_5QVal_Int_7QNone_Int_6QNode_Int_2_argbuf,Go),
                     (lizzieLet17_5QVal_Int_7QNone_Int_6QError_Int_2_argbuf,Go),
                     (es_14_6MyFalse_6QNone_Int_1_argbuf,Go),
                     (es_21_4MyFalse_1_argbuf,Go),
                     (es_21_4MyTrue_2_argbuf,Go),
                     (es_14_6MyFalse_6QNode_Int_2_argbuf,Go),
                     (es_14_6MyFalse_6QError_Int_2_argbuf,Go),
                     (es_14_4MyTrue_1_argbuf,Go),
                     (lizzieLet17_5QVal_Int_5QNode_Int_2_argbuf,Go),
                     (lizzieLet17_5QVal_Int_5QError_Int_2_argbuf,Go),
                     (lizzieLet17_5QNode_Int_7QNone_Int_8QNone_Int_1_argbuf,Go),
                     (lizzieLet17_5QNode_Int_7QNone_Int_8QVal_Int_2_argbuf,Go),
                     (lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_5_argbuf,Go),
                     (lizzieLet17_5QNode_Int_7QNone_Int_8QError_Int_2_argbuf,Go),
                     (lizzieLet17_5QNode_Int_5QVal_Int_2_argbuf,Go),
                     (lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_5_argbuf,Go),
                     (lizzieLet17_5QNode_Int_7QNode_Int_8QVal_Int_2_argbuf,Go),
                     (lizzieLet17_5QNode_Int_7QNode_Int_8QError_Int_2_argbuf,Go),
                     (lizzieLet17_5QNode_Int_5QError_Int_2_argbuf,Go),
                     (lizzieLet17_3QError_Int_2_argbuf,Go)] > (go_15_goMux_choice,C35) (go_15_goMux_data,Go) */
  logic [34:0] lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_select_d;
  assign lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_select_d = ((| lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_select_q) ? lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_select_q :
                                                                (lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_d[0] ? 35'd1 :
                                                                 (lizzieLet67_3Lcall_f_f_Int0_1_argbuf_d[0] ? 35'd2 :
                                                                  (lizzieLet17_5QNone_Int_7QVal_Int_5QNone_Int_1_argbuf_d[0] ? 35'd4 :
                                                                   (es_2_1_3MyFalse_1_argbuf_d[0] ? 35'd8 :
                                                                    (es_2_1_3MyTrue_2_argbuf_d[0] ? 35'd16 :
                                                                     (lizzieLet17_5QNone_Int_7QVal_Int_5QNode_Int_2_argbuf_d[0] ? 35'd32 :
                                                                      (lizzieLet17_5QNone_Int_7QVal_Int_5QError_Int_2_argbuf_d[0] ? 35'd64 :
                                                                       (lizzieLet17_5QNone_Int_7QNode_Int_5QNone_Int_1_argbuf_d[0] ? 35'd128 :
                                                                        (lizzieLet17_5QNone_Int_7QNode_Int_5QVal_Int_2_argbuf_d[0] ? 35'd256 :
                                                                         (lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_5_argbuf_d[0] ? 35'd512 :
                                                                          (lizzieLet17_5QNone_Int_7QNode_Int_5QError_Int_2_argbuf_d[0] ? 35'd1024 :
                                                                           (lizzieLet17_5QNone_Int_5QError_Int_2_argbuf_d[0] ? 35'd2048 :
                                                                            (lizzieLet17_5QVal_Int_7QNone_Int_6QNone_Int_1_argbuf_d[0] ? 35'd4096 :
                                                                             (es_10_4MyFalse_1_argbuf_d[0] ? 35'd8192 :
                                                                              (es_10_4MyTrue_2_argbuf_d[0] ? 35'd16384 :
                                                                               (lizzieLet17_5QVal_Int_7QNone_Int_6QNode_Int_2_argbuf_d[0] ? 35'd32768 :
                                                                                (lizzieLet17_5QVal_Int_7QNone_Int_6QError_Int_2_argbuf_d[0] ? 35'd65536 :
                                                                                 (es_14_6MyFalse_6QNone_Int_1_argbuf_d[0] ? 35'd131072 :
                                                                                  (es_21_4MyFalse_1_argbuf_d[0] ? 35'd262144 :
                                                                                   (es_21_4MyTrue_2_argbuf_d[0] ? 35'd524288 :
                                                                                    (es_14_6MyFalse_6QNode_Int_2_argbuf_d[0] ? 35'd1048576 :
                                                                                     (es_14_6MyFalse_6QError_Int_2_argbuf_d[0] ? 35'd2097152 :
                                                                                      (es_14_4MyTrue_1_argbuf_d[0] ? 35'd4194304 :
                                                                                       (lizzieLet17_5QVal_Int_5QNode_Int_2_argbuf_d[0] ? 35'd8388608 :
                                                                                        (lizzieLet17_5QVal_Int_5QError_Int_2_argbuf_d[0] ? 35'd16777216 :
                                                                                         (lizzieLet17_5QNode_Int_7QNone_Int_8QNone_Int_1_argbuf_d[0] ? 35'd33554432 :
                                                                                          (lizzieLet17_5QNode_Int_7QNone_Int_8QVal_Int_2_argbuf_d[0] ? 35'd67108864 :
                                                                                           (lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_5_argbuf_d[0] ? 35'd134217728 :
                                                                                            (lizzieLet17_5QNode_Int_7QNone_Int_8QError_Int_2_argbuf_d[0] ? 35'd268435456 :
                                                                                             (lizzieLet17_5QNode_Int_5QVal_Int_2_argbuf_d[0] ? 35'd536870912 :
                                                                                              (lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_5_argbuf_d[0] ? 35'd1073741824 :
                                                                                               (lizzieLet17_5QNode_Int_7QNode_Int_8QVal_Int_2_argbuf_d[0] ? 35'd2147483648 :
                                                                                                (lizzieLet17_5QNode_Int_7QNode_Int_8QError_Int_2_argbuf_d[0] ? 35'd4294967296 :
                                                                                                 (lizzieLet17_5QNode_Int_5QError_Int_2_argbuf_d[0] ? 35'd8589934592 :
                                                                                                  (lizzieLet17_3QError_Int_2_argbuf_d[0] ? 35'd17179869184 :
                                                                                                   35'd0))))))))))))))))))))))))))))))))))));
  logic [34:0] lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_select_q <= 35'd0;
    else
      lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_select_q <= (lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_done ? 35'd0 :
                                                              lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_select_d);
  logic [1:0] lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_emit_q <= 2'd0;
    else
      lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_emit_q <= (lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_done ? 2'd0 :
                                                            lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_emit_d);
  logic [1:0] lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_emit_d;
  assign lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_emit_d = (lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_emit_q | ({go_15_goMux_choice_d[0],
                                                                                                                    go_15_goMux_data_d[0]} & {go_15_goMux_choice_r,
                                                                                                                                              go_15_goMux_data_r}));
  logic lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_done;
  assign lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_done = (& lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_emit_d);
  assign {lizzieLet17_3QError_Int_2_argbuf_r,
          lizzieLet17_5QNode_Int_5QError_Int_2_argbuf_r,
          lizzieLet17_5QNode_Int_7QNode_Int_8QError_Int_2_argbuf_r,
          lizzieLet17_5QNode_Int_7QNode_Int_8QVal_Int_2_argbuf_r,
          lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_5_argbuf_r,
          lizzieLet17_5QNode_Int_5QVal_Int_2_argbuf_r,
          lizzieLet17_5QNode_Int_7QNone_Int_8QError_Int_2_argbuf_r,
          lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_5_argbuf_r,
          lizzieLet17_5QNode_Int_7QNone_Int_8QVal_Int_2_argbuf_r,
          lizzieLet17_5QNode_Int_7QNone_Int_8QNone_Int_1_argbuf_r,
          lizzieLet17_5QVal_Int_5QError_Int_2_argbuf_r,
          lizzieLet17_5QVal_Int_5QNode_Int_2_argbuf_r,
          es_14_4MyTrue_1_argbuf_r,
          es_14_6MyFalse_6QError_Int_2_argbuf_r,
          es_14_6MyFalse_6QNode_Int_2_argbuf_r,
          es_21_4MyTrue_2_argbuf_r,
          es_21_4MyFalse_1_argbuf_r,
          es_14_6MyFalse_6QNone_Int_1_argbuf_r,
          lizzieLet17_5QVal_Int_7QNone_Int_6QError_Int_2_argbuf_r,
          lizzieLet17_5QVal_Int_7QNone_Int_6QNode_Int_2_argbuf_r,
          es_10_4MyTrue_2_argbuf_r,
          es_10_4MyFalse_1_argbuf_r,
          lizzieLet17_5QVal_Int_7QNone_Int_6QNone_Int_1_argbuf_r,
          lizzieLet17_5QNone_Int_5QError_Int_2_argbuf_r,
          lizzieLet17_5QNone_Int_7QNode_Int_5QError_Int_2_argbuf_r,
          lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_5_argbuf_r,
          lizzieLet17_5QNone_Int_7QNode_Int_5QVal_Int_2_argbuf_r,
          lizzieLet17_5QNone_Int_7QNode_Int_5QNone_Int_1_argbuf_r,
          lizzieLet17_5QNone_Int_7QVal_Int_5QError_Int_2_argbuf_r,
          lizzieLet17_5QNone_Int_7QVal_Int_5QNode_Int_2_argbuf_r,
          es_2_1_3MyTrue_2_argbuf_r,
          es_2_1_3MyFalse_1_argbuf_r,
          lizzieLet17_5QNone_Int_7QVal_Int_5QNone_Int_1_argbuf_r,
          lizzieLet67_3Lcall_f_f_Int0_1_argbuf_r,
          lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_r} = (lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_done ? lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_select_d :
                                                           35'd0);
  assign go_15_goMux_data_d = ((lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_select_d[0] && (! lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_emit_q[0])) ? lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_d :
                               ((lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_select_d[1] && (! lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_emit_q[0])) ? lizzieLet67_3Lcall_f_f_Int0_1_argbuf_d :
                                ((lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_select_d[2] && (! lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_emit_q[0])) ? lizzieLet17_5QNone_Int_7QVal_Int_5QNone_Int_1_argbuf_d :
                                 ((lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_select_d[3] && (! lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_emit_q[0])) ? es_2_1_3MyFalse_1_argbuf_d :
                                  ((lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_select_d[4] && (! lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_emit_q[0])) ? es_2_1_3MyTrue_2_argbuf_d :
                                   ((lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_select_d[5] && (! lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_emit_q[0])) ? lizzieLet17_5QNone_Int_7QVal_Int_5QNode_Int_2_argbuf_d :
                                    ((lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_select_d[6] && (! lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_emit_q[0])) ? lizzieLet17_5QNone_Int_7QVal_Int_5QError_Int_2_argbuf_d :
                                     ((lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_select_d[7] && (! lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_emit_q[0])) ? lizzieLet17_5QNone_Int_7QNode_Int_5QNone_Int_1_argbuf_d :
                                      ((lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_select_d[8] && (! lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_emit_q[0])) ? lizzieLet17_5QNone_Int_7QNode_Int_5QVal_Int_2_argbuf_d :
                                       ((lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_select_d[9] && (! lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_emit_q[0])) ? lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_5_argbuf_d :
                                        ((lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_select_d[10] && (! lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_emit_q[0])) ? lizzieLet17_5QNone_Int_7QNode_Int_5QError_Int_2_argbuf_d :
                                         ((lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_select_d[11] && (! lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_emit_q[0])) ? lizzieLet17_5QNone_Int_5QError_Int_2_argbuf_d :
                                          ((lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_select_d[12] && (! lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_emit_q[0])) ? lizzieLet17_5QVal_Int_7QNone_Int_6QNone_Int_1_argbuf_d :
                                           ((lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_select_d[13] && (! lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_emit_q[0])) ? es_10_4MyFalse_1_argbuf_d :
                                            ((lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_select_d[14] && (! lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_emit_q[0])) ? es_10_4MyTrue_2_argbuf_d :
                                             ((lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_select_d[15] && (! lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_emit_q[0])) ? lizzieLet17_5QVal_Int_7QNone_Int_6QNode_Int_2_argbuf_d :
                                              ((lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_select_d[16] && (! lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_emit_q[0])) ? lizzieLet17_5QVal_Int_7QNone_Int_6QError_Int_2_argbuf_d :
                                               ((lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_select_d[17] && (! lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_emit_q[0])) ? es_14_6MyFalse_6QNone_Int_1_argbuf_d :
                                                ((lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_select_d[18] && (! lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_emit_q[0])) ? es_21_4MyFalse_1_argbuf_d :
                                                 ((lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_select_d[19] && (! lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_emit_q[0])) ? es_21_4MyTrue_2_argbuf_d :
                                                  ((lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_select_d[20] && (! lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_emit_q[0])) ? es_14_6MyFalse_6QNode_Int_2_argbuf_d :
                                                   ((lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_select_d[21] && (! lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_emit_q[0])) ? es_14_6MyFalse_6QError_Int_2_argbuf_d :
                                                    ((lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_select_d[22] && (! lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_emit_q[0])) ? es_14_4MyTrue_1_argbuf_d :
                                                     ((lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_select_d[23] && (! lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_emit_q[0])) ? lizzieLet17_5QVal_Int_5QNode_Int_2_argbuf_d :
                                                      ((lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_select_d[24] && (! lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_emit_q[0])) ? lizzieLet17_5QVal_Int_5QError_Int_2_argbuf_d :
                                                       ((lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_select_d[25] && (! lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_emit_q[0])) ? lizzieLet17_5QNode_Int_7QNone_Int_8QNone_Int_1_argbuf_d :
                                                        ((lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_select_d[26] && (! lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_emit_q[0])) ? lizzieLet17_5QNode_Int_7QNone_Int_8QVal_Int_2_argbuf_d :
                                                         ((lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_select_d[27] && (! lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_emit_q[0])) ? lizzieLet17_5QNode_Int_7QNone_Int_8QNode_Int_5_argbuf_d :
                                                          ((lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_select_d[28] && (! lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_emit_q[0])) ? lizzieLet17_5QNode_Int_7QNone_Int_8QError_Int_2_argbuf_d :
                                                           ((lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_select_d[29] && (! lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_emit_q[0])) ? lizzieLet17_5QNode_Int_5QVal_Int_2_argbuf_d :
                                                            ((lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_select_d[30] && (! lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_emit_q[0])) ? lizzieLet17_5QNode_Int_7QNode_Int_8QNone_Int_5_argbuf_d :
                                                             ((lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_select_d[31] && (! lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_emit_q[0])) ? lizzieLet17_5QNode_Int_7QNode_Int_8QVal_Int_2_argbuf_d :
                                                              ((lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_select_d[32] && (! lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_emit_q[0])) ? lizzieLet17_5QNode_Int_7QNode_Int_8QError_Int_2_argbuf_d :
                                                               ((lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_select_d[33] && (! lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_emit_q[0])) ? lizzieLet17_5QNode_Int_5QError_Int_2_argbuf_d :
                                                                ((lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_select_d[34] && (! lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_emit_q[0])) ? lizzieLet17_3QError_Int_2_argbuf_d :
                                                                 1'd0)))))))))))))))))))))))))))))))))));
  assign go_15_goMux_choice_d = ((lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_select_d[0] && (! lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_emit_q[1])) ? C1_35_dc(1'd1) :
                                 ((lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_select_d[1] && (! lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_emit_q[1])) ? C2_35_dc(1'd1) :
                                  ((lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_select_d[2] && (! lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_emit_q[1])) ? C3_35_dc(1'd1) :
                                   ((lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_select_d[3] && (! lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_emit_q[1])) ? C4_35_dc(1'd1) :
                                    ((lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_select_d[4] && (! lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_emit_q[1])) ? C5_35_dc(1'd1) :
                                     ((lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_select_d[5] && (! lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_emit_q[1])) ? C6_35_dc(1'd1) :
                                      ((lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_select_d[6] && (! lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_emit_q[1])) ? C7_35_dc(1'd1) :
                                       ((lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_select_d[7] && (! lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_emit_q[1])) ? C8_35_dc(1'd1) :
                                        ((lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_select_d[8] && (! lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_emit_q[1])) ? C9_35_dc(1'd1) :
                                         ((lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_select_d[9] && (! lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_emit_q[1])) ? C10_35_dc(1'd1) :
                                          ((lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_select_d[10] && (! lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_emit_q[1])) ? C11_35_dc(1'd1) :
                                           ((lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_select_d[11] && (! lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_emit_q[1])) ? C12_35_dc(1'd1) :
                                            ((lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_select_d[12] && (! lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_emit_q[1])) ? C13_35_dc(1'd1) :
                                             ((lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_select_d[13] && (! lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_emit_q[1])) ? C14_35_dc(1'd1) :
                                              ((lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_select_d[14] && (! lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_emit_q[1])) ? C15_35_dc(1'd1) :
                                               ((lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_select_d[15] && (! lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_emit_q[1])) ? C16_35_dc(1'd1) :
                                                ((lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_select_d[16] && (! lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_emit_q[1])) ? C17_35_dc(1'd1) :
                                                 ((lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_select_d[17] && (! lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_emit_q[1])) ? C18_35_dc(1'd1) :
                                                  ((lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_select_d[18] && (! lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_emit_q[1])) ? C19_35_dc(1'd1) :
                                                   ((lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_select_d[19] && (! lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_emit_q[1])) ? C20_35_dc(1'd1) :
                                                    ((lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_select_d[20] && (! lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_emit_q[1])) ? C21_35_dc(1'd1) :
                                                     ((lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_select_d[21] && (! lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_emit_q[1])) ? C22_35_dc(1'd1) :
                                                      ((lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_select_d[22] && (! lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_emit_q[1])) ? C23_35_dc(1'd1) :
                                                       ((lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_select_d[23] && (! lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_emit_q[1])) ? C24_35_dc(1'd1) :
                                                        ((lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_select_d[24] && (! lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_emit_q[1])) ? C25_35_dc(1'd1) :
                                                         ((lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_select_d[25] && (! lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_emit_q[1])) ? C26_35_dc(1'd1) :
                                                          ((lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_select_d[26] && (! lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_emit_q[1])) ? C27_35_dc(1'd1) :
                                                           ((lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_select_d[27] && (! lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_emit_q[1])) ? C28_35_dc(1'd1) :
                                                            ((lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_select_d[28] && (! lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_emit_q[1])) ? C29_35_dc(1'd1) :
                                                             ((lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_select_d[29] && (! lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_emit_q[1])) ? C30_35_dc(1'd1) :
                                                              ((lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_select_d[30] && (! lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_emit_q[1])) ? C31_35_dc(1'd1) :
                                                               ((lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_select_d[31] && (! lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_emit_q[1])) ? C32_35_dc(1'd1) :
                                                                ((lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_select_d[32] && (! lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_emit_q[1])) ? C33_35_dc(1'd1) :
                                                                 ((lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_select_d[33] && (! lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_emit_q[1])) ? C34_35_dc(1'd1) :
                                                                  ((lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_select_d[34] && (! lizzieLet17_5QNone_Int_5QNone_Int_1_argbuf_emit_q[1])) ? C35_35_dc(1'd1) :
                                                                   {6'd0,
                                                                    1'd0})))))))))))))))))))))))))))))))))));
  
  /* demux (Ty QTree_Int,
       Ty MyDTInt_Bool) : (lizzieLet17_5QNone_Int_6,QTree_Int) (lizzieLet17_4QNone_Int,MyDTInt_Bool) > [(_148,MyDTInt_Bool),
                                                                                                        (lizzieLet17_5QNone_Int_6QVal_Int,MyDTInt_Bool),
                                                                                                        (lizzieLet17_5QNone_Int_6QNode_Int,MyDTInt_Bool),
                                                                                                        (_147,MyDTInt_Bool)] */
  logic [3:0] lizzieLet17_4QNone_Int_onehotd;
  always_comb
    if ((lizzieLet17_5QNone_Int_6_d[0] && lizzieLet17_4QNone_Int_d[0]))
      unique case (lizzieLet17_5QNone_Int_6_d[2:1])
        2'd0: lizzieLet17_4QNone_Int_onehotd = 4'd1;
        2'd1: lizzieLet17_4QNone_Int_onehotd = 4'd2;
        2'd2: lizzieLet17_4QNone_Int_onehotd = 4'd4;
        2'd3: lizzieLet17_4QNone_Int_onehotd = 4'd8;
        default: lizzieLet17_4QNone_Int_onehotd = 4'd0;
      endcase
    else lizzieLet17_4QNone_Int_onehotd = 4'd0;
  assign _148_d = lizzieLet17_4QNone_Int_onehotd[0];
  assign lizzieLet17_5QNone_Int_6QVal_Int_d = lizzieLet17_4QNone_Int_onehotd[1];
  assign lizzieLet17_5QNone_Int_6QNode_Int_d = lizzieLet17_4QNone_Int_onehotd[2];
  assign _147_d = lizzieLet17_4QNone_Int_onehotd[3];
  assign lizzieLet17_4QNone_Int_r = (| (lizzieLet17_4QNone_Int_onehotd & {_147_r,
                                                                          lizzieLet17_5QNone_Int_6QNode_Int_r,
                                                                          lizzieLet17_5QNone_Int_6QVal_Int_r,
                                                                          _148_r}));
  assign lizzieLet17_5QNone_Int_6_r = lizzieLet17_4QNone_Int_r;
  
  /* demux (Ty QTree_Int,
       Ty QTree_Int) : (lizzieLet17_5QNone_Int_7,QTree_Int) (lizzieLet17_6QNone_Int,QTree_Int) > [(_146,QTree_Int),
                                                                                                  (lizzieLet17_5QNone_Int_7QVal_Int,QTree_Int),
                                                                                                  (lizzieLet17_5QNone_Int_7QNode_Int,QTree_Int),
                                                                                                  (_145,QTree_Int)] */
  logic [3:0] lizzieLet17_6QNone_Int_onehotd;
  always_comb
    if ((lizzieLet17_5QNone_Int_7_d[0] && lizzieLet17_6QNone_Int_d[0]))
      unique case (lizzieLet17_5QNone_Int_7_d[2:1])
        2'd0: lizzieLet17_6QNone_Int_onehotd = 4'd1;
        2'd1: lizzieLet17_6QNone_Int_onehotd = 4'd2;
        2'd2: lizzieLet17_6QNone_Int_onehotd = 4'd4;
        2'd3: lizzieLet17_6QNone_Int_onehotd = 4'd8;
        default: lizzieLet17_6QNone_Int_onehotd = 4'd0;
      endcase
    else lizzieLet17_6QNone_Int_onehotd = 4'd0;
  assign _146_d = {lizzieLet17_6QNone_Int_d[66:1],
                   lizzieLet17_6QNone_Int_onehotd[0]};
  assign lizzieLet17_5QNone_Int_7QVal_Int_d = {lizzieLet17_6QNone_Int_d[66:1],
                                               lizzieLet17_6QNone_Int_onehotd[1]};
  assign lizzieLet17_5QNone_Int_7QNode_Int_d = {lizzieLet17_6QNone_Int_d[66:1],
                                                lizzieLet17_6QNone_Int_onehotd[2]};
  assign _145_d = {lizzieLet17_6QNone_Int_d[66:1],
                   lizzieLet17_6QNone_Int_onehotd[3]};
  assign lizzieLet17_6QNone_Int_r = (| (lizzieLet17_6QNone_Int_onehotd & {_145_r,
                                                                          lizzieLet17_5QNone_Int_7QNode_Int_r,
                                                                          lizzieLet17_5QNone_Int_7QVal_Int_r,
                                                                          _146_r}));
  assign lizzieLet17_5QNone_Int_7_r = lizzieLet17_6QNone_Int_r;
  
  /* fork (Ty QTree_Int) : (lizzieLet17_5QNone_Int_7QNode_Int,QTree_Int) > [(lizzieLet17_5QNone_Int_7QNode_Int_1,QTree_Int),
                                                                       (lizzieLet17_5QNone_Int_7QNode_Int_2,QTree_Int),
                                                                       (lizzieLet17_5QNone_Int_7QNode_Int_3,QTree_Int),
                                                                       (lizzieLet17_5QNone_Int_7QNode_Int_4,QTree_Int),
                                                                       (lizzieLet17_5QNone_Int_7QNode_Int_5,QTree_Int),
                                                                       (lizzieLet17_5QNone_Int_7QNode_Int_6,QTree_Int),
                                                                       (lizzieLet17_5QNone_Int_7QNode_Int_7,QTree_Int),
                                                                       (lizzieLet17_5QNone_Int_7QNode_Int_8,QTree_Int),
                                                                       (lizzieLet17_5QNone_Int_7QNode_Int_9,QTree_Int),
                                                                       (lizzieLet17_5QNone_Int_7QNode_Int_10,QTree_Int),
                                                                       (lizzieLet17_5QNone_Int_7QNode_Int_11,QTree_Int)] */
  logic [10:0] lizzieLet17_5QNone_Int_7QNode_Int_emitted;
  logic [10:0] lizzieLet17_5QNone_Int_7QNode_Int_done;
  assign lizzieLet17_5QNone_Int_7QNode_Int_1_d = {lizzieLet17_5QNone_Int_7QNode_Int_d[66:1],
                                                  (lizzieLet17_5QNone_Int_7QNode_Int_d[0] && (! lizzieLet17_5QNone_Int_7QNode_Int_emitted[0]))};
  assign lizzieLet17_5QNone_Int_7QNode_Int_2_d = {lizzieLet17_5QNone_Int_7QNode_Int_d[66:1],
                                                  (lizzieLet17_5QNone_Int_7QNode_Int_d[0] && (! lizzieLet17_5QNone_Int_7QNode_Int_emitted[1]))};
  assign lizzieLet17_5QNone_Int_7QNode_Int_3_d = {lizzieLet17_5QNone_Int_7QNode_Int_d[66:1],
                                                  (lizzieLet17_5QNone_Int_7QNode_Int_d[0] && (! lizzieLet17_5QNone_Int_7QNode_Int_emitted[2]))};
  assign lizzieLet17_5QNone_Int_7QNode_Int_4_d = {lizzieLet17_5QNone_Int_7QNode_Int_d[66:1],
                                                  (lizzieLet17_5QNone_Int_7QNode_Int_d[0] && (! lizzieLet17_5QNone_Int_7QNode_Int_emitted[3]))};
  assign lizzieLet17_5QNone_Int_7QNode_Int_5_d = {lizzieLet17_5QNone_Int_7QNode_Int_d[66:1],
                                                  (lizzieLet17_5QNone_Int_7QNode_Int_d[0] && (! lizzieLet17_5QNone_Int_7QNode_Int_emitted[4]))};
  assign lizzieLet17_5QNone_Int_7QNode_Int_6_d = {lizzieLet17_5QNone_Int_7QNode_Int_d[66:1],
                                                  (lizzieLet17_5QNone_Int_7QNode_Int_d[0] && (! lizzieLet17_5QNone_Int_7QNode_Int_emitted[5]))};
  assign lizzieLet17_5QNone_Int_7QNode_Int_7_d = {lizzieLet17_5QNone_Int_7QNode_Int_d[66:1],
                                                  (lizzieLet17_5QNone_Int_7QNode_Int_d[0] && (! lizzieLet17_5QNone_Int_7QNode_Int_emitted[6]))};
  assign lizzieLet17_5QNone_Int_7QNode_Int_8_d = {lizzieLet17_5QNone_Int_7QNode_Int_d[66:1],
                                                  (lizzieLet17_5QNone_Int_7QNode_Int_d[0] && (! lizzieLet17_5QNone_Int_7QNode_Int_emitted[7]))};
  assign lizzieLet17_5QNone_Int_7QNode_Int_9_d = {lizzieLet17_5QNone_Int_7QNode_Int_d[66:1],
                                                  (lizzieLet17_5QNone_Int_7QNode_Int_d[0] && (! lizzieLet17_5QNone_Int_7QNode_Int_emitted[8]))};
  assign lizzieLet17_5QNone_Int_7QNode_Int_10_d = {lizzieLet17_5QNone_Int_7QNode_Int_d[66:1],
                                                   (lizzieLet17_5QNone_Int_7QNode_Int_d[0] && (! lizzieLet17_5QNone_Int_7QNode_Int_emitted[9]))};
  assign lizzieLet17_5QNone_Int_7QNode_Int_11_d = {lizzieLet17_5QNone_Int_7QNode_Int_d[66:1],
                                                   (lizzieLet17_5QNone_Int_7QNode_Int_d[0] && (! lizzieLet17_5QNone_Int_7QNode_Int_emitted[10]))};
  assign lizzieLet17_5QNone_Int_7QNode_Int_done = (lizzieLet17_5QNone_Int_7QNode_Int_emitted | ({lizzieLet17_5QNone_Int_7QNode_Int_11_d[0],
                                                                                                 lizzieLet17_5QNone_Int_7QNode_Int_10_d[0],
                                                                                                 lizzieLet17_5QNone_Int_7QNode_Int_9_d[0],
                                                                                                 lizzieLet17_5QNone_Int_7QNode_Int_8_d[0],
                                                                                                 lizzieLet17_5QNone_Int_7QNode_Int_7_d[0],
                                                                                                 lizzieLet17_5QNone_Int_7QNode_Int_6_d[0],
                                                                                                 lizzieLet17_5QNone_Int_7QNode_Int_5_d[0],
                                                                                                 lizzieLet17_5QNone_Int_7QNode_Int_4_d[0],
                                                                                                 lizzieLet17_5QNone_Int_7QNode_Int_3_d[0],
                                                                                                 lizzieLet17_5QNone_Int_7QNode_Int_2_d[0],
                                                                                                 lizzieLet17_5QNone_Int_7QNode_Int_1_d[0]} & {lizzieLet17_5QNone_Int_7QNode_Int_11_r,
                                                                                                                                              lizzieLet17_5QNone_Int_7QNode_Int_10_r,
                                                                                                                                              lizzieLet17_5QNone_Int_7QNode_Int_9_r,
                                                                                                                                              lizzieLet17_5QNone_Int_7QNode_Int_8_r,
                                                                                                                                              lizzieLet17_5QNone_Int_7QNode_Int_7_r,
                                                                                                                                              lizzieLet17_5QNone_Int_7QNode_Int_6_r,
                                                                                                                                              lizzieLet17_5QNone_Int_7QNode_Int_5_r,
                                                                                                                                              lizzieLet17_5QNone_Int_7QNode_Int_4_r,
                                                                                                                                              lizzieLet17_5QNone_Int_7QNode_Int_3_r,
                                                                                                                                              lizzieLet17_5QNone_Int_7QNode_Int_2_r,
                                                                                                                                              lizzieLet17_5QNone_Int_7QNode_Int_1_r}));
  assign lizzieLet17_5QNone_Int_7QNode_Int_r = (& lizzieLet17_5QNone_Int_7QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNone_Int_7QNode_Int_emitted <= 11'd0;
    else
      lizzieLet17_5QNone_Int_7QNode_Int_emitted <= (lizzieLet17_5QNone_Int_7QNode_Int_r ? 11'd0 :
                                                    lizzieLet17_5QNone_Int_7QNode_Int_done);
  
  /* demux (Ty QTree_Int,
       Ty Pointer_QTree_Int) : (lizzieLet17_5QNone_Int_7QNode_Int_10,QTree_Int) (q3aeD_destruct,Pointer_QTree_Int) > [(_144,Pointer_QTree_Int),
                                                                                                                      (_143,Pointer_QTree_Int),
                                                                                                                      (lizzieLet17_5QNone_Int_7QNode_Int_10QNode_Int,Pointer_QTree_Int),
                                                                                                                      (_142,Pointer_QTree_Int)] */
  logic [3:0] q3aeD_destruct_onehotd;
  always_comb
    if ((lizzieLet17_5QNone_Int_7QNode_Int_10_d[0] && q3aeD_destruct_d[0]))
      unique case (lizzieLet17_5QNone_Int_7QNode_Int_10_d[2:1])
        2'd0: q3aeD_destruct_onehotd = 4'd1;
        2'd1: q3aeD_destruct_onehotd = 4'd2;
        2'd2: q3aeD_destruct_onehotd = 4'd4;
        2'd3: q3aeD_destruct_onehotd = 4'd8;
        default: q3aeD_destruct_onehotd = 4'd0;
      endcase
    else q3aeD_destruct_onehotd = 4'd0;
  assign _144_d = {q3aeD_destruct_d[16:1],
                   q3aeD_destruct_onehotd[0]};
  assign _143_d = {q3aeD_destruct_d[16:1],
                   q3aeD_destruct_onehotd[1]};
  assign lizzieLet17_5QNone_Int_7QNode_Int_10QNode_Int_d = {q3aeD_destruct_d[16:1],
                                                            q3aeD_destruct_onehotd[2]};
  assign _142_d = {q3aeD_destruct_d[16:1],
                   q3aeD_destruct_onehotd[3]};
  assign q3aeD_destruct_r = (| (q3aeD_destruct_onehotd & {_142_r,
                                                          lizzieLet17_5QNone_Int_7QNode_Int_10QNode_Int_r,
                                                          _143_r,
                                                          _144_r}));
  assign lizzieLet17_5QNone_Int_7QNode_Int_10_r = q3aeD_destruct_r;
  
  /* buf (Ty Pointer_QTree_Int) : (lizzieLet17_5QNone_Int_7QNode_Int_10QNode_Int,Pointer_QTree_Int) > (lizzieLet17_5QNone_Int_7QNode_Int_10QNode_Int_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t lizzieLet17_5QNone_Int_7QNode_Int_10QNode_Int_bufchan_d;
  logic lizzieLet17_5QNone_Int_7QNode_Int_10QNode_Int_bufchan_r;
  assign lizzieLet17_5QNone_Int_7QNode_Int_10QNode_Int_r = ((! lizzieLet17_5QNone_Int_7QNode_Int_10QNode_Int_bufchan_d[0]) || lizzieLet17_5QNone_Int_7QNode_Int_10QNode_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNone_Int_7QNode_Int_10QNode_Int_bufchan_d <= {16'd0,
                                                                  1'd0};
    else
      if (lizzieLet17_5QNone_Int_7QNode_Int_10QNode_Int_r)
        lizzieLet17_5QNone_Int_7QNode_Int_10QNode_Int_bufchan_d <= lizzieLet17_5QNone_Int_7QNode_Int_10QNode_Int_d;
  Pointer_QTree_Int_t lizzieLet17_5QNone_Int_7QNode_Int_10QNode_Int_bufchan_buf;
  assign lizzieLet17_5QNone_Int_7QNode_Int_10QNode_Int_bufchan_r = (! lizzieLet17_5QNone_Int_7QNode_Int_10QNode_Int_bufchan_buf[0]);
  assign lizzieLet17_5QNone_Int_7QNode_Int_10QNode_Int_1_argbuf_d = (lizzieLet17_5QNone_Int_7QNode_Int_10QNode_Int_bufchan_buf[0] ? lizzieLet17_5QNone_Int_7QNode_Int_10QNode_Int_bufchan_buf :
                                                                     lizzieLet17_5QNone_Int_7QNode_Int_10QNode_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNone_Int_7QNode_Int_10QNode_Int_bufchan_buf <= {16'd0,
                                                                    1'd0};
    else
      if ((lizzieLet17_5QNone_Int_7QNode_Int_10QNode_Int_1_argbuf_r && lizzieLet17_5QNone_Int_7QNode_Int_10QNode_Int_bufchan_buf[0]))
        lizzieLet17_5QNone_Int_7QNode_Int_10QNode_Int_bufchan_buf <= {16'd0,
                                                                      1'd0};
      else if (((! lizzieLet17_5QNone_Int_7QNode_Int_10QNode_Int_1_argbuf_r) && (! lizzieLet17_5QNone_Int_7QNode_Int_10QNode_Int_bufchan_buf[0])))
        lizzieLet17_5QNone_Int_7QNode_Int_10QNode_Int_bufchan_buf <= lizzieLet17_5QNone_Int_7QNode_Int_10QNode_Int_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_QTree_Int) : (lizzieLet17_5QNone_Int_7QNode_Int_11,QTree_Int) (q4aeE_destruct,Pointer_QTree_Int) > [(_141,Pointer_QTree_Int),
                                                                                                                      (_140,Pointer_QTree_Int),
                                                                                                                      (lizzieLet17_5QNone_Int_7QNode_Int_11QNode_Int,Pointer_QTree_Int),
                                                                                                                      (_139,Pointer_QTree_Int)] */
  logic [3:0] q4aeE_destruct_onehotd;
  always_comb
    if ((lizzieLet17_5QNone_Int_7QNode_Int_11_d[0] && q4aeE_destruct_d[0]))
      unique case (lizzieLet17_5QNone_Int_7QNode_Int_11_d[2:1])
        2'd0: q4aeE_destruct_onehotd = 4'd1;
        2'd1: q4aeE_destruct_onehotd = 4'd2;
        2'd2: q4aeE_destruct_onehotd = 4'd4;
        2'd3: q4aeE_destruct_onehotd = 4'd8;
        default: q4aeE_destruct_onehotd = 4'd0;
      endcase
    else q4aeE_destruct_onehotd = 4'd0;
  assign _141_d = {q4aeE_destruct_d[16:1],
                   q4aeE_destruct_onehotd[0]};
  assign _140_d = {q4aeE_destruct_d[16:1],
                   q4aeE_destruct_onehotd[1]};
  assign lizzieLet17_5QNone_Int_7QNode_Int_11QNode_Int_d = {q4aeE_destruct_d[16:1],
                                                            q4aeE_destruct_onehotd[2]};
  assign _139_d = {q4aeE_destruct_d[16:1],
                   q4aeE_destruct_onehotd[3]};
  assign q4aeE_destruct_r = (| (q4aeE_destruct_onehotd & {_139_r,
                                                          lizzieLet17_5QNone_Int_7QNode_Int_11QNode_Int_r,
                                                          _140_r,
                                                          _141_r}));
  assign lizzieLet17_5QNone_Int_7QNode_Int_11_r = q4aeE_destruct_r;
  
  /* buf (Ty Pointer_QTree_Int) : (lizzieLet17_5QNone_Int_7QNode_Int_11QNode_Int,Pointer_QTree_Int) > (lizzieLet17_5QNone_Int_7QNode_Int_11QNode_Int_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t lizzieLet17_5QNone_Int_7QNode_Int_11QNode_Int_bufchan_d;
  logic lizzieLet17_5QNone_Int_7QNode_Int_11QNode_Int_bufchan_r;
  assign lizzieLet17_5QNone_Int_7QNode_Int_11QNode_Int_r = ((! lizzieLet17_5QNone_Int_7QNode_Int_11QNode_Int_bufchan_d[0]) || lizzieLet17_5QNone_Int_7QNode_Int_11QNode_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNone_Int_7QNode_Int_11QNode_Int_bufchan_d <= {16'd0,
                                                                  1'd0};
    else
      if (lizzieLet17_5QNone_Int_7QNode_Int_11QNode_Int_r)
        lizzieLet17_5QNone_Int_7QNode_Int_11QNode_Int_bufchan_d <= lizzieLet17_5QNone_Int_7QNode_Int_11QNode_Int_d;
  Pointer_QTree_Int_t lizzieLet17_5QNone_Int_7QNode_Int_11QNode_Int_bufchan_buf;
  assign lizzieLet17_5QNone_Int_7QNode_Int_11QNode_Int_bufchan_r = (! lizzieLet17_5QNone_Int_7QNode_Int_11QNode_Int_bufchan_buf[0]);
  assign lizzieLet17_5QNone_Int_7QNode_Int_11QNode_Int_1_argbuf_d = (lizzieLet17_5QNone_Int_7QNode_Int_11QNode_Int_bufchan_buf[0] ? lizzieLet17_5QNone_Int_7QNode_Int_11QNode_Int_bufchan_buf :
                                                                     lizzieLet17_5QNone_Int_7QNode_Int_11QNode_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNone_Int_7QNode_Int_11QNode_Int_bufchan_buf <= {16'd0,
                                                                    1'd0};
    else
      if ((lizzieLet17_5QNone_Int_7QNode_Int_11QNode_Int_1_argbuf_r && lizzieLet17_5QNone_Int_7QNode_Int_11QNode_Int_bufchan_buf[0]))
        lizzieLet17_5QNone_Int_7QNode_Int_11QNode_Int_bufchan_buf <= {16'd0,
                                                                      1'd0};
      else if (((! lizzieLet17_5QNone_Int_7QNode_Int_11QNode_Int_1_argbuf_r) && (! lizzieLet17_5QNone_Int_7QNode_Int_11QNode_Int_bufchan_buf[0])))
        lizzieLet17_5QNone_Int_7QNode_Int_11QNode_Int_bufchan_buf <= lizzieLet17_5QNone_Int_7QNode_Int_11QNode_Int_bufchan_d;
  
  /* destruct (Ty QTree_Int,
          Dcon QNode_Int) : (lizzieLet17_5QNone_Int_7QNode_Int_1QNode_Int,QTree_Int) > [(t1aeG_destruct,Pointer_QTree_Int),
                                                                                        (t2aeH_destruct,Pointer_QTree_Int),
                                                                                        (t3aeI_destruct,Pointer_QTree_Int),
                                                                                        (t4aeJ_destruct,Pointer_QTree_Int)] */
  logic [3:0] lizzieLet17_5QNone_Int_7QNode_Int_1QNode_Int_emitted;
  logic [3:0] lizzieLet17_5QNone_Int_7QNode_Int_1QNode_Int_done;
  assign t1aeG_destruct_d = {lizzieLet17_5QNone_Int_7QNode_Int_1QNode_Int_d[18:3],
                             (lizzieLet17_5QNone_Int_7QNode_Int_1QNode_Int_d[0] && (! lizzieLet17_5QNone_Int_7QNode_Int_1QNode_Int_emitted[0]))};
  assign t2aeH_destruct_d = {lizzieLet17_5QNone_Int_7QNode_Int_1QNode_Int_d[34:19],
                             (lizzieLet17_5QNone_Int_7QNode_Int_1QNode_Int_d[0] && (! lizzieLet17_5QNone_Int_7QNode_Int_1QNode_Int_emitted[1]))};
  assign t3aeI_destruct_d = {lizzieLet17_5QNone_Int_7QNode_Int_1QNode_Int_d[50:35],
                             (lizzieLet17_5QNone_Int_7QNode_Int_1QNode_Int_d[0] && (! lizzieLet17_5QNone_Int_7QNode_Int_1QNode_Int_emitted[2]))};
  assign t4aeJ_destruct_d = {lizzieLet17_5QNone_Int_7QNode_Int_1QNode_Int_d[66:51],
                             (lizzieLet17_5QNone_Int_7QNode_Int_1QNode_Int_d[0] && (! lizzieLet17_5QNone_Int_7QNode_Int_1QNode_Int_emitted[3]))};
  assign lizzieLet17_5QNone_Int_7QNode_Int_1QNode_Int_done = (lizzieLet17_5QNone_Int_7QNode_Int_1QNode_Int_emitted | ({t4aeJ_destruct_d[0],
                                                                                                                       t3aeI_destruct_d[0],
                                                                                                                       t2aeH_destruct_d[0],
                                                                                                                       t1aeG_destruct_d[0]} & {t4aeJ_destruct_r,
                                                                                                                                               t3aeI_destruct_r,
                                                                                                                                               t2aeH_destruct_r,
                                                                                                                                               t1aeG_destruct_r}));
  assign lizzieLet17_5QNone_Int_7QNode_Int_1QNode_Int_r = (& lizzieLet17_5QNone_Int_7QNode_Int_1QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNone_Int_7QNode_Int_1QNode_Int_emitted <= 4'd0;
    else
      lizzieLet17_5QNone_Int_7QNode_Int_1QNode_Int_emitted <= (lizzieLet17_5QNone_Int_7QNode_Int_1QNode_Int_r ? 4'd0 :
                                                               lizzieLet17_5QNone_Int_7QNode_Int_1QNode_Int_done);
  
  /* demux (Ty QTree_Int,
       Ty QTree_Int) : (lizzieLet17_5QNone_Int_7QNode_Int_2,QTree_Int) (lizzieLet17_5QNone_Int_7QNode_Int_1,QTree_Int) > [(_138,QTree_Int),
                                                                                                                          (_137,QTree_Int),
                                                                                                                          (lizzieLet17_5QNone_Int_7QNode_Int_1QNode_Int,QTree_Int),
                                                                                                                          (_136,QTree_Int)] */
  logic [3:0] lizzieLet17_5QNone_Int_7QNode_Int_1_onehotd;
  always_comb
    if ((lizzieLet17_5QNone_Int_7QNode_Int_2_d[0] && lizzieLet17_5QNone_Int_7QNode_Int_1_d[0]))
      unique case (lizzieLet17_5QNone_Int_7QNode_Int_2_d[2:1])
        2'd0: lizzieLet17_5QNone_Int_7QNode_Int_1_onehotd = 4'd1;
        2'd1: lizzieLet17_5QNone_Int_7QNode_Int_1_onehotd = 4'd2;
        2'd2: lizzieLet17_5QNone_Int_7QNode_Int_1_onehotd = 4'd4;
        2'd3: lizzieLet17_5QNone_Int_7QNode_Int_1_onehotd = 4'd8;
        default: lizzieLet17_5QNone_Int_7QNode_Int_1_onehotd = 4'd0;
      endcase
    else lizzieLet17_5QNone_Int_7QNode_Int_1_onehotd = 4'd0;
  assign _138_d = {lizzieLet17_5QNone_Int_7QNode_Int_1_d[66:1],
                   lizzieLet17_5QNone_Int_7QNode_Int_1_onehotd[0]};
  assign _137_d = {lizzieLet17_5QNone_Int_7QNode_Int_1_d[66:1],
                   lizzieLet17_5QNone_Int_7QNode_Int_1_onehotd[1]};
  assign lizzieLet17_5QNone_Int_7QNode_Int_1QNode_Int_d = {lizzieLet17_5QNone_Int_7QNode_Int_1_d[66:1],
                                                           lizzieLet17_5QNone_Int_7QNode_Int_1_onehotd[2]};
  assign _136_d = {lizzieLet17_5QNone_Int_7QNode_Int_1_d[66:1],
                   lizzieLet17_5QNone_Int_7QNode_Int_1_onehotd[3]};
  assign lizzieLet17_5QNone_Int_7QNode_Int_1_r = (| (lizzieLet17_5QNone_Int_7QNode_Int_1_onehotd & {_136_r,
                                                                                                    lizzieLet17_5QNone_Int_7QNode_Int_1QNode_Int_r,
                                                                                                    _137_r,
                                                                                                    _138_r}));
  assign lizzieLet17_5QNone_Int_7QNode_Int_2_r = lizzieLet17_5QNone_Int_7QNode_Int_1_r;
  
  /* demux (Ty QTree_Int,
       Ty MyDTInt_Int_Int) : (lizzieLet17_5QNone_Int_7QNode_Int_3,QTree_Int) (lizzieLet17_5QNone_Int_3QNode_Int,MyDTInt_Int_Int) > [(_135,MyDTInt_Int_Int),
                                                                                                                                    (_134,MyDTInt_Int_Int),
                                                                                                                                    (lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int,MyDTInt_Int_Int),
                                                                                                                                    (_133,MyDTInt_Int_Int)] */
  logic [3:0] lizzieLet17_5QNone_Int_3QNode_Int_onehotd;
  always_comb
    if ((lizzieLet17_5QNone_Int_7QNode_Int_3_d[0] && lizzieLet17_5QNone_Int_3QNode_Int_d[0]))
      unique case (lizzieLet17_5QNone_Int_7QNode_Int_3_d[2:1])
        2'd0: lizzieLet17_5QNone_Int_3QNode_Int_onehotd = 4'd1;
        2'd1: lizzieLet17_5QNone_Int_3QNode_Int_onehotd = 4'd2;
        2'd2: lizzieLet17_5QNone_Int_3QNode_Int_onehotd = 4'd4;
        2'd3: lizzieLet17_5QNone_Int_3QNode_Int_onehotd = 4'd8;
        default: lizzieLet17_5QNone_Int_3QNode_Int_onehotd = 4'd0;
      endcase
    else lizzieLet17_5QNone_Int_3QNode_Int_onehotd = 4'd0;
  assign _135_d = lizzieLet17_5QNone_Int_3QNode_Int_onehotd[0];
  assign _134_d = lizzieLet17_5QNone_Int_3QNode_Int_onehotd[1];
  assign lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_d = lizzieLet17_5QNone_Int_3QNode_Int_onehotd[2];
  assign _133_d = lizzieLet17_5QNone_Int_3QNode_Int_onehotd[3];
  assign lizzieLet17_5QNone_Int_3QNode_Int_r = (| (lizzieLet17_5QNone_Int_3QNode_Int_onehotd & {_133_r,
                                                                                                lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_r,
                                                                                                _134_r,
                                                                                                _135_r}));
  assign lizzieLet17_5QNone_Int_7QNode_Int_3_r = lizzieLet17_5QNone_Int_3QNode_Int_r;
  
  /* fork (Ty MyDTInt_Int_Int) : (lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int,MyDTInt_Int_Int) > [(lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_1,MyDTInt_Int_Int),
                                                                                              (lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_2,MyDTInt_Int_Int),
                                                                                              (lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_3,MyDTInt_Int_Int),
                                                                                              (lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_4,MyDTInt_Int_Int)] */
  logic [3:0] lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_emitted;
  logic [3:0] lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_done;
  assign lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_1_d = (lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_d[0] && (! lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_emitted[0]));
  assign lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_2_d = (lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_d[0] && (! lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_emitted[1]));
  assign lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_3_d = (lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_d[0] && (! lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_emitted[2]));
  assign lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_4_d = (lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_d[0] && (! lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_emitted[3]));
  assign lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_done = (lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_emitted | ({lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_4_d[0],
                                                                                                                       lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_3_d[0],
                                                                                                                       lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_2_d[0],
                                                                                                                       lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_1_d[0]} & {lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_4_r,
                                                                                                                                                                               lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_3_r,
                                                                                                                                                                               lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_2_r,
                                                                                                                                                                               lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_1_r}));
  assign lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_r = (& lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_emitted <= 4'd0;
    else
      lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_emitted <= (lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_r ? 4'd0 :
                                                               lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_done);
  
  /* buf (Ty MyDTInt_Int_Int) : (lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_1,MyDTInt_Int_Int) > (lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_1_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_1_bufchan_d;
  logic lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_1_bufchan_r;
  assign lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_1_r = ((! lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_1_bufchan_d[0]) || lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_1_bufchan_d <= 1'd0;
    else
      if (lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_1_r)
        lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_1_bufchan_d <= lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_1_d;
  MyDTInt_Int_Int_t lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_1_bufchan_buf;
  assign lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_1_bufchan_r = (! lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_1_bufchan_buf[0]);
  assign lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_1_argbuf_d = (lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_1_bufchan_buf[0] ? lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_1_bufchan_buf :
                                                                    lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_1_argbuf_r && lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_1_bufchan_buf[0]))
        lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_1_argbuf_r) && (! lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_1_bufchan_buf[0])))
        lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_1_bufchan_buf <= lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_1_bufchan_d;
  
  /* buf (Ty MyDTInt_Int_Int) : (lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_2,MyDTInt_Int_Int) > (lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_2_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_2_bufchan_d;
  logic lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_2_bufchan_r;
  assign lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_2_r = ((! lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_2_bufchan_d[0]) || lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_2_r)
        lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_2_bufchan_d <= lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_2_d;
  MyDTInt_Int_Int_t lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_2_bufchan_buf;
  assign lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_2_bufchan_r = (! lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_2_bufchan_buf[0]);
  assign lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_2_argbuf_d = (lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_2_bufchan_buf[0] ? lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_2_bufchan_buf :
                                                                    lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_2_argbuf_r && lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_2_bufchan_buf[0]))
        lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_2_argbuf_r) && (! lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_2_bufchan_buf[0])))
        lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_2_bufchan_buf <= lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_2_bufchan_d;
  
  /* buf (Ty MyDTInt_Int_Int) : (lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_3,MyDTInt_Int_Int) > (lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_3_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_3_bufchan_d;
  logic lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_3_bufchan_r;
  assign lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_3_r = ((! lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_3_bufchan_d[0]) || lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_3_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_3_bufchan_d <= 1'd0;
    else
      if (lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_3_r)
        lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_3_bufchan_d <= lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_3_d;
  MyDTInt_Int_Int_t lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_3_bufchan_buf;
  assign lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_3_bufchan_r = (! lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_3_bufchan_buf[0]);
  assign lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_3_argbuf_d = (lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_3_bufchan_buf[0] ? lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_3_bufchan_buf :
                                                                    lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_3_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_3_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_3_argbuf_r && lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_3_bufchan_buf[0]))
        lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_3_bufchan_buf <= 1'd0;
      else if (((! lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_3_argbuf_r) && (! lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_3_bufchan_buf[0])))
        lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_3_bufchan_buf <= lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_3_bufchan_d;
  
  /* buf (Ty MyDTInt_Int_Int) : (lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_4,MyDTInt_Int_Int) > (lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_4_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_4_bufchan_d;
  logic lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_4_bufchan_r;
  assign lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_4_r = ((! lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_4_bufchan_d[0]) || lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_4_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_4_bufchan_d <= 1'd0;
    else
      if (lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_4_r)
        lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_4_bufchan_d <= lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_4_d;
  MyDTInt_Int_Int_t lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_4_bufchan_buf;
  assign lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_4_bufchan_r = (! lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_4_bufchan_buf[0]);
  assign lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_4_argbuf_d = (lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_4_bufchan_buf[0] ? lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_4_bufchan_buf :
                                                                    lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_4_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_4_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_4_argbuf_r && lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_4_bufchan_buf[0]))
        lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_4_bufchan_buf <= 1'd0;
      else if (((! lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_4_argbuf_r) && (! lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_4_bufchan_buf[0])))
        lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_4_bufchan_buf <= lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_4_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_CTf_f_Int) : (lizzieLet17_5QNone_Int_7QNode_Int_4,QTree_Int) (lizzieLet17_5QNone_Int_4QNode_Int,Pointer_CTf_f_Int) > [(lizzieLet17_5QNone_Int_7QNode_Int_4QNone_Int,Pointer_CTf_f_Int),
                                                                                                                                        (lizzieLet17_5QNone_Int_7QNode_Int_4QVal_Int,Pointer_CTf_f_Int),
                                                                                                                                        (lizzieLet17_5QNone_Int_7QNode_Int_4QNode_Int,Pointer_CTf_f_Int),
                                                                                                                                        (lizzieLet17_5QNone_Int_7QNode_Int_4QError_Int,Pointer_CTf_f_Int)] */
  logic [3:0] lizzieLet17_5QNone_Int_4QNode_Int_onehotd;
  always_comb
    if ((lizzieLet17_5QNone_Int_7QNode_Int_4_d[0] && lizzieLet17_5QNone_Int_4QNode_Int_d[0]))
      unique case (lizzieLet17_5QNone_Int_7QNode_Int_4_d[2:1])
        2'd0: lizzieLet17_5QNone_Int_4QNode_Int_onehotd = 4'd1;
        2'd1: lizzieLet17_5QNone_Int_4QNode_Int_onehotd = 4'd2;
        2'd2: lizzieLet17_5QNone_Int_4QNode_Int_onehotd = 4'd4;
        2'd3: lizzieLet17_5QNone_Int_4QNode_Int_onehotd = 4'd8;
        default: lizzieLet17_5QNone_Int_4QNode_Int_onehotd = 4'd0;
      endcase
    else lizzieLet17_5QNone_Int_4QNode_Int_onehotd = 4'd0;
  assign lizzieLet17_5QNone_Int_7QNode_Int_4QNone_Int_d = {lizzieLet17_5QNone_Int_4QNode_Int_d[16:1],
                                                           lizzieLet17_5QNone_Int_4QNode_Int_onehotd[0]};
  assign lizzieLet17_5QNone_Int_7QNode_Int_4QVal_Int_d = {lizzieLet17_5QNone_Int_4QNode_Int_d[16:1],
                                                          lizzieLet17_5QNone_Int_4QNode_Int_onehotd[1]};
  assign lizzieLet17_5QNone_Int_7QNode_Int_4QNode_Int_d = {lizzieLet17_5QNone_Int_4QNode_Int_d[16:1],
                                                           lizzieLet17_5QNone_Int_4QNode_Int_onehotd[2]};
  assign lizzieLet17_5QNone_Int_7QNode_Int_4QError_Int_d = {lizzieLet17_5QNone_Int_4QNode_Int_d[16:1],
                                                            lizzieLet17_5QNone_Int_4QNode_Int_onehotd[3]};
  assign lizzieLet17_5QNone_Int_4QNode_Int_r = (| (lizzieLet17_5QNone_Int_4QNode_Int_onehotd & {lizzieLet17_5QNone_Int_7QNode_Int_4QError_Int_r,
                                                                                                lizzieLet17_5QNone_Int_7QNode_Int_4QNode_Int_r,
                                                                                                lizzieLet17_5QNone_Int_7QNode_Int_4QVal_Int_r,
                                                                                                lizzieLet17_5QNone_Int_7QNode_Int_4QNone_Int_r}));
  assign lizzieLet17_5QNone_Int_7QNode_Int_4_r = lizzieLet17_5QNone_Int_4QNode_Int_r;
  
  /* buf (Ty Pointer_CTf_f_Int) : (lizzieLet17_5QNone_Int_7QNode_Int_4QError_Int,Pointer_CTf_f_Int) > (lizzieLet17_5QNone_Int_7QNode_Int_4QError_Int_1_argbuf,Pointer_CTf_f_Int) */
  Pointer_CTf_f_Int_t lizzieLet17_5QNone_Int_7QNode_Int_4QError_Int_bufchan_d;
  logic lizzieLet17_5QNone_Int_7QNode_Int_4QError_Int_bufchan_r;
  assign lizzieLet17_5QNone_Int_7QNode_Int_4QError_Int_r = ((! lizzieLet17_5QNone_Int_7QNode_Int_4QError_Int_bufchan_d[0]) || lizzieLet17_5QNone_Int_7QNode_Int_4QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNone_Int_7QNode_Int_4QError_Int_bufchan_d <= {16'd0,
                                                                  1'd0};
    else
      if (lizzieLet17_5QNone_Int_7QNode_Int_4QError_Int_r)
        lizzieLet17_5QNone_Int_7QNode_Int_4QError_Int_bufchan_d <= lizzieLet17_5QNone_Int_7QNode_Int_4QError_Int_d;
  Pointer_CTf_f_Int_t lizzieLet17_5QNone_Int_7QNode_Int_4QError_Int_bufchan_buf;
  assign lizzieLet17_5QNone_Int_7QNode_Int_4QError_Int_bufchan_r = (! lizzieLet17_5QNone_Int_7QNode_Int_4QError_Int_bufchan_buf[0]);
  assign lizzieLet17_5QNone_Int_7QNode_Int_4QError_Int_1_argbuf_d = (lizzieLet17_5QNone_Int_7QNode_Int_4QError_Int_bufchan_buf[0] ? lizzieLet17_5QNone_Int_7QNode_Int_4QError_Int_bufchan_buf :
                                                                     lizzieLet17_5QNone_Int_7QNode_Int_4QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNone_Int_7QNode_Int_4QError_Int_bufchan_buf <= {16'd0,
                                                                    1'd0};
    else
      if ((lizzieLet17_5QNone_Int_7QNode_Int_4QError_Int_1_argbuf_r && lizzieLet17_5QNone_Int_7QNode_Int_4QError_Int_bufchan_buf[0]))
        lizzieLet17_5QNone_Int_7QNode_Int_4QError_Int_bufchan_buf <= {16'd0,
                                                                      1'd0};
      else if (((! lizzieLet17_5QNone_Int_7QNode_Int_4QError_Int_1_argbuf_r) && (! lizzieLet17_5QNone_Int_7QNode_Int_4QError_Int_bufchan_buf[0])))
        lizzieLet17_5QNone_Int_7QNode_Int_4QError_Int_bufchan_buf <= lizzieLet17_5QNone_Int_7QNode_Int_4QError_Int_bufchan_d;
  
  /* buf (Ty Pointer_CTf_f_Int) : (lizzieLet17_5QNone_Int_7QNode_Int_4QNode_Int,Pointer_CTf_f_Int) > (lizzieLet17_5QNone_Int_7QNode_Int_4QNode_Int_1_argbuf,Pointer_CTf_f_Int) */
  Pointer_CTf_f_Int_t lizzieLet17_5QNone_Int_7QNode_Int_4QNode_Int_bufchan_d;
  logic lizzieLet17_5QNone_Int_7QNode_Int_4QNode_Int_bufchan_r;
  assign lizzieLet17_5QNone_Int_7QNode_Int_4QNode_Int_r = ((! lizzieLet17_5QNone_Int_7QNode_Int_4QNode_Int_bufchan_d[0]) || lizzieLet17_5QNone_Int_7QNode_Int_4QNode_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNone_Int_7QNode_Int_4QNode_Int_bufchan_d <= {16'd0,
                                                                 1'd0};
    else
      if (lizzieLet17_5QNone_Int_7QNode_Int_4QNode_Int_r)
        lizzieLet17_5QNone_Int_7QNode_Int_4QNode_Int_bufchan_d <= lizzieLet17_5QNone_Int_7QNode_Int_4QNode_Int_d;
  Pointer_CTf_f_Int_t lizzieLet17_5QNone_Int_7QNode_Int_4QNode_Int_bufchan_buf;
  assign lizzieLet17_5QNone_Int_7QNode_Int_4QNode_Int_bufchan_r = (! lizzieLet17_5QNone_Int_7QNode_Int_4QNode_Int_bufchan_buf[0]);
  assign lizzieLet17_5QNone_Int_7QNode_Int_4QNode_Int_1_argbuf_d = (lizzieLet17_5QNone_Int_7QNode_Int_4QNode_Int_bufchan_buf[0] ? lizzieLet17_5QNone_Int_7QNode_Int_4QNode_Int_bufchan_buf :
                                                                    lizzieLet17_5QNone_Int_7QNode_Int_4QNode_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNone_Int_7QNode_Int_4QNode_Int_bufchan_buf <= {16'd0,
                                                                   1'd0};
    else
      if ((lizzieLet17_5QNone_Int_7QNode_Int_4QNode_Int_1_argbuf_r && lizzieLet17_5QNone_Int_7QNode_Int_4QNode_Int_bufchan_buf[0]))
        lizzieLet17_5QNone_Int_7QNode_Int_4QNode_Int_bufchan_buf <= {16'd0,
                                                                     1'd0};
      else if (((! lizzieLet17_5QNone_Int_7QNode_Int_4QNode_Int_1_argbuf_r) && (! lizzieLet17_5QNone_Int_7QNode_Int_4QNode_Int_bufchan_buf[0])))
        lizzieLet17_5QNone_Int_7QNode_Int_4QNode_Int_bufchan_buf <= lizzieLet17_5QNone_Int_7QNode_Int_4QNode_Int_bufchan_d;
  
  /* buf (Ty Pointer_CTf_f_Int) : (lizzieLet17_5QNone_Int_7QNode_Int_4QNone_Int,Pointer_CTf_f_Int) > (lizzieLet17_5QNone_Int_7QNode_Int_4QNone_Int_1_argbuf,Pointer_CTf_f_Int) */
  Pointer_CTf_f_Int_t lizzieLet17_5QNone_Int_7QNode_Int_4QNone_Int_bufchan_d;
  logic lizzieLet17_5QNone_Int_7QNode_Int_4QNone_Int_bufchan_r;
  assign lizzieLet17_5QNone_Int_7QNode_Int_4QNone_Int_r = ((! lizzieLet17_5QNone_Int_7QNode_Int_4QNone_Int_bufchan_d[0]) || lizzieLet17_5QNone_Int_7QNode_Int_4QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNone_Int_7QNode_Int_4QNone_Int_bufchan_d <= {16'd0,
                                                                 1'd0};
    else
      if (lizzieLet17_5QNone_Int_7QNode_Int_4QNone_Int_r)
        lizzieLet17_5QNone_Int_7QNode_Int_4QNone_Int_bufchan_d <= lizzieLet17_5QNone_Int_7QNode_Int_4QNone_Int_d;
  Pointer_CTf_f_Int_t lizzieLet17_5QNone_Int_7QNode_Int_4QNone_Int_bufchan_buf;
  assign lizzieLet17_5QNone_Int_7QNode_Int_4QNone_Int_bufchan_r = (! lizzieLet17_5QNone_Int_7QNode_Int_4QNone_Int_bufchan_buf[0]);
  assign lizzieLet17_5QNone_Int_7QNode_Int_4QNone_Int_1_argbuf_d = (lizzieLet17_5QNone_Int_7QNode_Int_4QNone_Int_bufchan_buf[0] ? lizzieLet17_5QNone_Int_7QNode_Int_4QNone_Int_bufchan_buf :
                                                                    lizzieLet17_5QNone_Int_7QNode_Int_4QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNone_Int_7QNode_Int_4QNone_Int_bufchan_buf <= {16'd0,
                                                                   1'd0};
    else
      if ((lizzieLet17_5QNone_Int_7QNode_Int_4QNone_Int_1_argbuf_r && lizzieLet17_5QNone_Int_7QNode_Int_4QNone_Int_bufchan_buf[0]))
        lizzieLet17_5QNone_Int_7QNode_Int_4QNone_Int_bufchan_buf <= {16'd0,
                                                                     1'd0};
      else if (((! lizzieLet17_5QNone_Int_7QNode_Int_4QNone_Int_1_argbuf_r) && (! lizzieLet17_5QNone_Int_7QNode_Int_4QNone_Int_bufchan_buf[0])))
        lizzieLet17_5QNone_Int_7QNode_Int_4QNone_Int_bufchan_buf <= lizzieLet17_5QNone_Int_7QNode_Int_4QNone_Int_bufchan_d;
  
  /* buf (Ty Pointer_CTf_f_Int) : (lizzieLet17_5QNone_Int_7QNode_Int_4QVal_Int,Pointer_CTf_f_Int) > (lizzieLet17_5QNone_Int_7QNode_Int_4QVal_Int_1_argbuf,Pointer_CTf_f_Int) */
  Pointer_CTf_f_Int_t lizzieLet17_5QNone_Int_7QNode_Int_4QVal_Int_bufchan_d;
  logic lizzieLet17_5QNone_Int_7QNode_Int_4QVal_Int_bufchan_r;
  assign lizzieLet17_5QNone_Int_7QNode_Int_4QVal_Int_r = ((! lizzieLet17_5QNone_Int_7QNode_Int_4QVal_Int_bufchan_d[0]) || lizzieLet17_5QNone_Int_7QNode_Int_4QVal_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNone_Int_7QNode_Int_4QVal_Int_bufchan_d <= {16'd0,
                                                                1'd0};
    else
      if (lizzieLet17_5QNone_Int_7QNode_Int_4QVal_Int_r)
        lizzieLet17_5QNone_Int_7QNode_Int_4QVal_Int_bufchan_d <= lizzieLet17_5QNone_Int_7QNode_Int_4QVal_Int_d;
  Pointer_CTf_f_Int_t lizzieLet17_5QNone_Int_7QNode_Int_4QVal_Int_bufchan_buf;
  assign lizzieLet17_5QNone_Int_7QNode_Int_4QVal_Int_bufchan_r = (! lizzieLet17_5QNone_Int_7QNode_Int_4QVal_Int_bufchan_buf[0]);
  assign lizzieLet17_5QNone_Int_7QNode_Int_4QVal_Int_1_argbuf_d = (lizzieLet17_5QNone_Int_7QNode_Int_4QVal_Int_bufchan_buf[0] ? lizzieLet17_5QNone_Int_7QNode_Int_4QVal_Int_bufchan_buf :
                                                                   lizzieLet17_5QNone_Int_7QNode_Int_4QVal_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNone_Int_7QNode_Int_4QVal_Int_bufchan_buf <= {16'd0,
                                                                  1'd0};
    else
      if ((lizzieLet17_5QNone_Int_7QNode_Int_4QVal_Int_1_argbuf_r && lizzieLet17_5QNone_Int_7QNode_Int_4QVal_Int_bufchan_buf[0]))
        lizzieLet17_5QNone_Int_7QNode_Int_4QVal_Int_bufchan_buf <= {16'd0,
                                                                    1'd0};
      else if (((! lizzieLet17_5QNone_Int_7QNode_Int_4QVal_Int_1_argbuf_r) && (! lizzieLet17_5QNone_Int_7QNode_Int_4QVal_Int_bufchan_buf[0])))
        lizzieLet17_5QNone_Int_7QNode_Int_4QVal_Int_bufchan_buf <= lizzieLet17_5QNone_Int_7QNode_Int_4QVal_Int_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Go) : (lizzieLet17_5QNone_Int_7QNode_Int_5,QTree_Int) (lizzieLet17_5QNone_Int_5QNode_Int,Go) > [(lizzieLet17_5QNone_Int_7QNode_Int_5QNone_Int,Go),
                                                                                                          (lizzieLet17_5QNone_Int_7QNode_Int_5QVal_Int,Go),
                                                                                                          (lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int,Go),
                                                                                                          (lizzieLet17_5QNone_Int_7QNode_Int_5QError_Int,Go)] */
  logic [3:0] lizzieLet17_5QNone_Int_5QNode_Int_onehotd;
  always_comb
    if ((lizzieLet17_5QNone_Int_7QNode_Int_5_d[0] && lizzieLet17_5QNone_Int_5QNode_Int_d[0]))
      unique case (lizzieLet17_5QNone_Int_7QNode_Int_5_d[2:1])
        2'd0: lizzieLet17_5QNone_Int_5QNode_Int_onehotd = 4'd1;
        2'd1: lizzieLet17_5QNone_Int_5QNode_Int_onehotd = 4'd2;
        2'd2: lizzieLet17_5QNone_Int_5QNode_Int_onehotd = 4'd4;
        2'd3: lizzieLet17_5QNone_Int_5QNode_Int_onehotd = 4'd8;
        default: lizzieLet17_5QNone_Int_5QNode_Int_onehotd = 4'd0;
      endcase
    else lizzieLet17_5QNone_Int_5QNode_Int_onehotd = 4'd0;
  assign lizzieLet17_5QNone_Int_7QNode_Int_5QNone_Int_d = lizzieLet17_5QNone_Int_5QNode_Int_onehotd[0];
  assign lizzieLet17_5QNone_Int_7QNode_Int_5QVal_Int_d = lizzieLet17_5QNone_Int_5QNode_Int_onehotd[1];
  assign lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_d = lizzieLet17_5QNone_Int_5QNode_Int_onehotd[2];
  assign lizzieLet17_5QNone_Int_7QNode_Int_5QError_Int_d = lizzieLet17_5QNone_Int_5QNode_Int_onehotd[3];
  assign lizzieLet17_5QNone_Int_5QNode_Int_r = (| (lizzieLet17_5QNone_Int_5QNode_Int_onehotd & {lizzieLet17_5QNone_Int_7QNode_Int_5QError_Int_r,
                                                                                                lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_r,
                                                                                                lizzieLet17_5QNone_Int_7QNode_Int_5QVal_Int_r,
                                                                                                lizzieLet17_5QNone_Int_7QNode_Int_5QNone_Int_r}));
  assign lizzieLet17_5QNone_Int_7QNode_Int_5_r = lizzieLet17_5QNone_Int_5QNode_Int_r;
  
  /* fork (Ty Go) : (lizzieLet17_5QNone_Int_7QNode_Int_5QError_Int,Go) > [(lizzieLet17_5QNone_Int_7QNode_Int_5QError_Int_1,Go),
                                                                     (lizzieLet17_5QNone_Int_7QNode_Int_5QError_Int_2,Go)] */
  logic [1:0] lizzieLet17_5QNone_Int_7QNode_Int_5QError_Int_emitted;
  logic [1:0] lizzieLet17_5QNone_Int_7QNode_Int_5QError_Int_done;
  assign lizzieLet17_5QNone_Int_7QNode_Int_5QError_Int_1_d = (lizzieLet17_5QNone_Int_7QNode_Int_5QError_Int_d[0] && (! lizzieLet17_5QNone_Int_7QNode_Int_5QError_Int_emitted[0]));
  assign lizzieLet17_5QNone_Int_7QNode_Int_5QError_Int_2_d = (lizzieLet17_5QNone_Int_7QNode_Int_5QError_Int_d[0] && (! lizzieLet17_5QNone_Int_7QNode_Int_5QError_Int_emitted[1]));
  assign lizzieLet17_5QNone_Int_7QNode_Int_5QError_Int_done = (lizzieLet17_5QNone_Int_7QNode_Int_5QError_Int_emitted | ({lizzieLet17_5QNone_Int_7QNode_Int_5QError_Int_2_d[0],
                                                                                                                         lizzieLet17_5QNone_Int_7QNode_Int_5QError_Int_1_d[0]} & {lizzieLet17_5QNone_Int_7QNode_Int_5QError_Int_2_r,
                                                                                                                                                                                  lizzieLet17_5QNone_Int_7QNode_Int_5QError_Int_1_r}));
  assign lizzieLet17_5QNone_Int_7QNode_Int_5QError_Int_r = (& lizzieLet17_5QNone_Int_7QNode_Int_5QError_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNone_Int_7QNode_Int_5QError_Int_emitted <= 2'd0;
    else
      lizzieLet17_5QNone_Int_7QNode_Int_5QError_Int_emitted <= (lizzieLet17_5QNone_Int_7QNode_Int_5QError_Int_r ? 2'd0 :
                                                                lizzieLet17_5QNone_Int_7QNode_Int_5QError_Int_done);
  
  /* dcon (Ty QTree_Int,
      Dcon QError_Int) : [(lizzieLet17_5QNone_Int_7QNode_Int_5QError_Int_1,Go)] > (lizzieLet17_5QNone_Int_7QNode_Int_5QError_Int_1QError_Int,QTree_Int) */
  assign lizzieLet17_5QNone_Int_7QNode_Int_5QError_Int_1QError_Int_d = QError_Int_dc((& {lizzieLet17_5QNone_Int_7QNode_Int_5QError_Int_1_d[0]}), lizzieLet17_5QNone_Int_7QNode_Int_5QError_Int_1_d);
  assign {lizzieLet17_5QNone_Int_7QNode_Int_5QError_Int_1_r} = {1 {(lizzieLet17_5QNone_Int_7QNode_Int_5QError_Int_1QError_Int_r && lizzieLet17_5QNone_Int_7QNode_Int_5QError_Int_1QError_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (lizzieLet17_5QNone_Int_7QNode_Int_5QError_Int_1QError_Int,QTree_Int) > (lizzieLet27_1_argbuf,QTree_Int) */
  QTree_Int_t lizzieLet17_5QNone_Int_7QNode_Int_5QError_Int_1QError_Int_bufchan_d;
  logic lizzieLet17_5QNone_Int_7QNode_Int_5QError_Int_1QError_Int_bufchan_r;
  assign lizzieLet17_5QNone_Int_7QNode_Int_5QError_Int_1QError_Int_r = ((! lizzieLet17_5QNone_Int_7QNode_Int_5QError_Int_1QError_Int_bufchan_d[0]) || lizzieLet17_5QNone_Int_7QNode_Int_5QError_Int_1QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNone_Int_7QNode_Int_5QError_Int_1QError_Int_bufchan_d <= {66'd0,
                                                                              1'd0};
    else
      if (lizzieLet17_5QNone_Int_7QNode_Int_5QError_Int_1QError_Int_r)
        lizzieLet17_5QNone_Int_7QNode_Int_5QError_Int_1QError_Int_bufchan_d <= lizzieLet17_5QNone_Int_7QNode_Int_5QError_Int_1QError_Int_d;
  QTree_Int_t lizzieLet17_5QNone_Int_7QNode_Int_5QError_Int_1QError_Int_bufchan_buf;
  assign lizzieLet17_5QNone_Int_7QNode_Int_5QError_Int_1QError_Int_bufchan_r = (! lizzieLet17_5QNone_Int_7QNode_Int_5QError_Int_1QError_Int_bufchan_buf[0]);
  assign lizzieLet27_1_argbuf_d = (lizzieLet17_5QNone_Int_7QNode_Int_5QError_Int_1QError_Int_bufchan_buf[0] ? lizzieLet17_5QNone_Int_7QNode_Int_5QError_Int_1QError_Int_bufchan_buf :
                                   lizzieLet17_5QNone_Int_7QNode_Int_5QError_Int_1QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNone_Int_7QNode_Int_5QError_Int_1QError_Int_bufchan_buf <= {66'd0,
                                                                                1'd0};
    else
      if ((lizzieLet27_1_argbuf_r && lizzieLet17_5QNone_Int_7QNode_Int_5QError_Int_1QError_Int_bufchan_buf[0]))
        lizzieLet17_5QNone_Int_7QNode_Int_5QError_Int_1QError_Int_bufchan_buf <= {66'd0,
                                                                                  1'd0};
      else if (((! lizzieLet27_1_argbuf_r) && (! lizzieLet17_5QNone_Int_7QNode_Int_5QError_Int_1QError_Int_bufchan_buf[0])))
        lizzieLet17_5QNone_Int_7QNode_Int_5QError_Int_1QError_Int_bufchan_buf <= lizzieLet17_5QNone_Int_7QNode_Int_5QError_Int_1QError_Int_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet17_5QNone_Int_7QNode_Int_5QError_Int_2,Go) > (lizzieLet17_5QNone_Int_7QNode_Int_5QError_Int_2_argbuf,Go) */
  Go_t lizzieLet17_5QNone_Int_7QNode_Int_5QError_Int_2_bufchan_d;
  logic lizzieLet17_5QNone_Int_7QNode_Int_5QError_Int_2_bufchan_r;
  assign lizzieLet17_5QNone_Int_7QNode_Int_5QError_Int_2_r = ((! lizzieLet17_5QNone_Int_7QNode_Int_5QError_Int_2_bufchan_d[0]) || lizzieLet17_5QNone_Int_7QNode_Int_5QError_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNone_Int_7QNode_Int_5QError_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet17_5QNone_Int_7QNode_Int_5QError_Int_2_r)
        lizzieLet17_5QNone_Int_7QNode_Int_5QError_Int_2_bufchan_d <= lizzieLet17_5QNone_Int_7QNode_Int_5QError_Int_2_d;
  Go_t lizzieLet17_5QNone_Int_7QNode_Int_5QError_Int_2_bufchan_buf;
  assign lizzieLet17_5QNone_Int_7QNode_Int_5QError_Int_2_bufchan_r = (! lizzieLet17_5QNone_Int_7QNode_Int_5QError_Int_2_bufchan_buf[0]);
  assign lizzieLet17_5QNone_Int_7QNode_Int_5QError_Int_2_argbuf_d = (lizzieLet17_5QNone_Int_7QNode_Int_5QError_Int_2_bufchan_buf[0] ? lizzieLet17_5QNone_Int_7QNode_Int_5QError_Int_2_bufchan_buf :
                                                                     lizzieLet17_5QNone_Int_7QNode_Int_5QError_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNone_Int_7QNode_Int_5QError_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet17_5QNone_Int_7QNode_Int_5QError_Int_2_argbuf_r && lizzieLet17_5QNone_Int_7QNode_Int_5QError_Int_2_bufchan_buf[0]))
        lizzieLet17_5QNone_Int_7QNode_Int_5QError_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet17_5QNone_Int_7QNode_Int_5QError_Int_2_argbuf_r) && (! lizzieLet17_5QNone_Int_7QNode_Int_5QError_Int_2_bufchan_buf[0])))
        lizzieLet17_5QNone_Int_7QNode_Int_5QError_Int_2_bufchan_buf <= lizzieLet17_5QNone_Int_7QNode_Int_5QError_Int_2_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int,Go) > [(lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_1,Go),
                                                                    (lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_2,Go),
                                                                    (lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_3,Go),
                                                                    (lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_4,Go),
                                                                    (lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_5,Go)] */
  logic [4:0] lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_emitted;
  logic [4:0] lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_done;
  assign lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_1_d = (lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_d[0] && (! lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_emitted[0]));
  assign lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_2_d = (lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_d[0] && (! lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_emitted[1]));
  assign lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_3_d = (lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_d[0] && (! lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_emitted[2]));
  assign lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_4_d = (lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_d[0] && (! lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_emitted[3]));
  assign lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_5_d = (lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_d[0] && (! lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_emitted[4]));
  assign lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_done = (lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_emitted | ({lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_5_d[0],
                                                                                                                       lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_4_d[0],
                                                                                                                       lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_3_d[0],
                                                                                                                       lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_2_d[0],
                                                                                                                       lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_1_d[0]} & {lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_5_r,
                                                                                                                                                                               lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_4_r,
                                                                                                                                                                               lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_3_r,
                                                                                                                                                                               lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_2_r,
                                                                                                                                                                               lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_1_r}));
  assign lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_r = (& lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_emitted <= 5'd0;
    else
      lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_emitted <= (lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_r ? 5'd0 :
                                                               lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_done);
  
  /* buf (Ty Go) : (lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_1,Go) > (lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_1_argbuf,Go) */
  Go_t lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_1_bufchan_d;
  logic lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_1_bufchan_r;
  assign lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_1_r = ((! lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_1_bufchan_d[0]) || lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_1_bufchan_d <= 1'd0;
    else
      if (lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_1_r)
        lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_1_bufchan_d <= lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_1_d;
  Go_t lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_1_bufchan_buf;
  assign lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_1_bufchan_r = (! lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_1_bufchan_buf[0]);
  assign lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_1_argbuf_d = (lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_1_bufchan_buf[0] ? lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_1_bufchan_buf :
                                                                    lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_1_argbuf_r && lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_1_bufchan_buf[0]))
        lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_1_argbuf_r) && (! lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_1_bufchan_buf[0])))
        lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_1_bufchan_buf <= lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_1_bufchan_d;
  
  /* dcon (Ty TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int,
      Dcon TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int) : [(lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_1_argbuf,Go),
                                                                                              (lizzieLet17_5QNone_Int_7QNode_Int_11QNode_Int_1_argbuf,Pointer_QTree_Int),
                                                                                              (t4aeJ_1_argbuf,Pointer_QTree_Int),
                                                                                              (lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_1_argbuf,MyDTInt_Bool),
                                                                                              (lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_1_argbuf,MyDTInt_Int_Int)] > (f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1,TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int) */
  assign \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_d  = TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_dc((& {lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_1_argbuf_d[0],
                                                                                                                                                                                                                     lizzieLet17_5QNone_Int_7QNode_Int_11QNode_Int_1_argbuf_d[0],
                                                                                                                                                                                                                     t4aeJ_1_argbuf_d[0],
                                                                                                                                                                                                                     lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_1_argbuf_d[0],
                                                                                                                                                                                                                     lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_1_argbuf_d[0]}), lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_1_argbuf_d, lizzieLet17_5QNone_Int_7QNode_Int_11QNode_Int_1_argbuf_d, t4aeJ_1_argbuf_d, lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_1_argbuf_d, lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_1_argbuf_d);
  assign {lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_1_argbuf_r,
          lizzieLet17_5QNone_Int_7QNode_Int_11QNode_Int_1_argbuf_r,
          t4aeJ_1_argbuf_r,
          lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_1_argbuf_r,
          lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_1_argbuf_r} = {5 {(\f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_r  && \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_d [0])}};
  
  /* buf (Ty Go) : (lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_2,Go) > (lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_2_argbuf,Go) */
  Go_t lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_2_bufchan_d;
  logic lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_2_bufchan_r;
  assign lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_2_r = ((! lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_2_bufchan_d[0]) || lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_2_r)
        lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_2_bufchan_d <= lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_2_d;
  Go_t lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_2_bufchan_buf;
  assign lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_2_bufchan_r = (! lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_2_bufchan_buf[0]);
  assign lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_2_argbuf_d = (lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_2_bufchan_buf[0] ? lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_2_bufchan_buf :
                                                                    lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_2_argbuf_r && lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_2_bufchan_buf[0]))
        lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_2_argbuf_r) && (! lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_2_bufchan_buf[0])))
        lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_2_bufchan_buf <= lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_2_bufchan_d;
  
  /* dcon (Ty TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int,
      Dcon TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int) : [(lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_2_argbuf,Go),
                                                                                              (lizzieLet17_5QNone_Int_7QNode_Int_10QNode_Int_1_argbuf,Pointer_QTree_Int),
                                                                                              (t3aeI_1_argbuf,Pointer_QTree_Int),
                                                                                              (lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_2_argbuf,MyDTInt_Bool),
                                                                                              (lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_2_argbuf,MyDTInt_Int_Int)] > (f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int2,TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int) */
  assign \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int2_d  = TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_dc((& {lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_2_argbuf_d[0],
                                                                                                                                                                                                                    lizzieLet17_5QNone_Int_7QNode_Int_10QNode_Int_1_argbuf_d[0],
                                                                                                                                                                                                                    t3aeI_1_argbuf_d[0],
                                                                                                                                                                                                                    lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_2_argbuf_d[0],
                                                                                                                                                                                                                    lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_2_argbuf_d[0]}), lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_2_argbuf_d, lizzieLet17_5QNone_Int_7QNode_Int_10QNode_Int_1_argbuf_d, t3aeI_1_argbuf_d, lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_2_argbuf_d, lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_2_argbuf_d);
  assign {lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_2_argbuf_r,
          lizzieLet17_5QNone_Int_7QNode_Int_10QNode_Int_1_argbuf_r,
          t3aeI_1_argbuf_r,
          lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_2_argbuf_r,
          lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_2_argbuf_r} = {5 {(\f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int2_r  && \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int2_d [0])}};
  
  /* buf (Ty Go) : (lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_3,Go) > (lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_3_argbuf,Go) */
  Go_t lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_3_bufchan_d;
  logic lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_3_bufchan_r;
  assign lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_3_r = ((! lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_3_bufchan_d[0]) || lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_3_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_3_bufchan_d <= 1'd0;
    else
      if (lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_3_r)
        lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_3_bufchan_d <= lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_3_d;
  Go_t lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_3_bufchan_buf;
  assign lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_3_bufchan_r = (! lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_3_bufchan_buf[0]);
  assign lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_3_argbuf_d = (lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_3_bufchan_buf[0] ? lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_3_bufchan_buf :
                                                                    lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_3_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_3_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_3_argbuf_r && lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_3_bufchan_buf[0]))
        lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_3_bufchan_buf <= 1'd0;
      else if (((! lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_3_argbuf_r) && (! lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_3_bufchan_buf[0])))
        lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_3_bufchan_buf <= lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_3_bufchan_d;
  
  /* dcon (Ty TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int,
      Dcon TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int) : [(lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_3_argbuf,Go),
                                                                                              (lizzieLet17_5QNone_Int_7QNode_Int_9QNode_Int_1_argbuf,Pointer_QTree_Int),
                                                                                              (t2aeH_1_argbuf,Pointer_QTree_Int),
                                                                                              (lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_3_argbuf,MyDTInt_Bool),
                                                                                              (lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_3_argbuf,MyDTInt_Int_Int)] > (f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int3,TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int) */
  assign \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int3_d  = TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_dc((& {lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_3_argbuf_d[0],
                                                                                                                                                                                                                    lizzieLet17_5QNone_Int_7QNode_Int_9QNode_Int_1_argbuf_d[0],
                                                                                                                                                                                                                    t2aeH_1_argbuf_d[0],
                                                                                                                                                                                                                    lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_3_argbuf_d[0],
                                                                                                                                                                                                                    lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_3_argbuf_d[0]}), lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_3_argbuf_d, lizzieLet17_5QNone_Int_7QNode_Int_9QNode_Int_1_argbuf_d, t2aeH_1_argbuf_d, lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_3_argbuf_d, lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_3_argbuf_d);
  assign {lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_3_argbuf_r,
          lizzieLet17_5QNone_Int_7QNode_Int_9QNode_Int_1_argbuf_r,
          t2aeH_1_argbuf_r,
          lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_3_argbuf_r,
          lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_3_argbuf_r} = {5 {(\f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int3_r  && \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int3_d [0])}};
  
  /* buf (Ty Go) : (lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_4,Go) > (lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_4_argbuf,Go) */
  Go_t lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_4_bufchan_d;
  logic lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_4_bufchan_r;
  assign lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_4_r = ((! lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_4_bufchan_d[0]) || lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_4_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_4_bufchan_d <= 1'd0;
    else
      if (lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_4_r)
        lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_4_bufchan_d <= lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_4_d;
  Go_t lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_4_bufchan_buf;
  assign lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_4_bufchan_r = (! lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_4_bufchan_buf[0]);
  assign lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_4_argbuf_d = (lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_4_bufchan_buf[0] ? lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_4_bufchan_buf :
                                                                    lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_4_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_4_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_4_argbuf_r && lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_4_bufchan_buf[0]))
        lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_4_bufchan_buf <= 1'd0;
      else if (((! lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_4_argbuf_r) && (! lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_4_bufchan_buf[0])))
        lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_4_bufchan_buf <= lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_4_bufchan_d;
  
  /* dcon (Ty TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int,
      Dcon TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int) : [(lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_4_argbuf,Go),
                                                                                              (lizzieLet17_5QNone_Int_7QNode_Int_8QNode_Int_1_argbuf,Pointer_QTree_Int),
                                                                                              (t1aeG_1_argbuf,Pointer_QTree_Int),
                                                                                              (lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_4_argbuf,MyDTInt_Bool),
                                                                                              (lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_4_argbuf,MyDTInt_Int_Int)] > (f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int4,TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int) */
  assign \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int4_d  = TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_dc((& {lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_4_argbuf_d[0],
                                                                                                                                                                                                                    lizzieLet17_5QNone_Int_7QNode_Int_8QNode_Int_1_argbuf_d[0],
                                                                                                                                                                                                                    t1aeG_1_argbuf_d[0],
                                                                                                                                                                                                                    lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_4_argbuf_d[0],
                                                                                                                                                                                                                    lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_4_argbuf_d[0]}), lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_4_argbuf_d, lizzieLet17_5QNone_Int_7QNode_Int_8QNode_Int_1_argbuf_d, t1aeG_1_argbuf_d, lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_4_argbuf_d, lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_4_argbuf_d);
  assign {lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_4_argbuf_r,
          lizzieLet17_5QNone_Int_7QNode_Int_8QNode_Int_1_argbuf_r,
          t1aeG_1_argbuf_r,
          lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_4_argbuf_r,
          lizzieLet17_5QNone_Int_7QNode_Int_3QNode_Int_4_argbuf_r} = {5 {(\f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int4_r  && \f''''''''''''_f''''''''''''_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int4_d [0])}};
  
  /* buf (Ty Go) : (lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_5,Go) > (lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_5_argbuf,Go) */
  Go_t lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_5_bufchan_d;
  logic lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_5_bufchan_r;
  assign lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_5_r = ((! lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_5_bufchan_d[0]) || lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_5_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_5_bufchan_d <= 1'd0;
    else
      if (lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_5_r)
        lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_5_bufchan_d <= lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_5_d;
  Go_t lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_5_bufchan_buf;
  assign lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_5_bufchan_r = (! lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_5_bufchan_buf[0]);
  assign lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_5_argbuf_d = (lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_5_bufchan_buf[0] ? lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_5_bufchan_buf :
                                                                    lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_5_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_5_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_5_argbuf_r && lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_5_bufchan_buf[0]))
        lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_5_bufchan_buf <= 1'd0;
      else if (((! lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_5_argbuf_r) && (! lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_5_bufchan_buf[0])))
        lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_5_bufchan_buf <= lizzieLet17_5QNone_Int_7QNode_Int_5QNode_Int_5_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet17_5QNone_Int_7QNode_Int_5QNone_Int,Go) > (lizzieLet17_5QNone_Int_7QNode_Int_5QNone_Int_1_argbuf,Go) */
  Go_t lizzieLet17_5QNone_Int_7QNode_Int_5QNone_Int_bufchan_d;
  logic lizzieLet17_5QNone_Int_7QNode_Int_5QNone_Int_bufchan_r;
  assign lizzieLet17_5QNone_Int_7QNode_Int_5QNone_Int_r = ((! lizzieLet17_5QNone_Int_7QNode_Int_5QNone_Int_bufchan_d[0]) || lizzieLet17_5QNone_Int_7QNode_Int_5QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNone_Int_7QNode_Int_5QNone_Int_bufchan_d <= 1'd0;
    else
      if (lizzieLet17_5QNone_Int_7QNode_Int_5QNone_Int_r)
        lizzieLet17_5QNone_Int_7QNode_Int_5QNone_Int_bufchan_d <= lizzieLet17_5QNone_Int_7QNode_Int_5QNone_Int_d;
  Go_t lizzieLet17_5QNone_Int_7QNode_Int_5QNone_Int_bufchan_buf;
  assign lizzieLet17_5QNone_Int_7QNode_Int_5QNone_Int_bufchan_r = (! lizzieLet17_5QNone_Int_7QNode_Int_5QNone_Int_bufchan_buf[0]);
  assign lizzieLet17_5QNone_Int_7QNode_Int_5QNone_Int_1_argbuf_d = (lizzieLet17_5QNone_Int_7QNode_Int_5QNone_Int_bufchan_buf[0] ? lizzieLet17_5QNone_Int_7QNode_Int_5QNone_Int_bufchan_buf :
                                                                    lizzieLet17_5QNone_Int_7QNode_Int_5QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNone_Int_7QNode_Int_5QNone_Int_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet17_5QNone_Int_7QNode_Int_5QNone_Int_1_argbuf_r && lizzieLet17_5QNone_Int_7QNode_Int_5QNone_Int_bufchan_buf[0]))
        lizzieLet17_5QNone_Int_7QNode_Int_5QNone_Int_bufchan_buf <= 1'd0;
      else if (((! lizzieLet17_5QNone_Int_7QNode_Int_5QNone_Int_1_argbuf_r) && (! lizzieLet17_5QNone_Int_7QNode_Int_5QNone_Int_bufchan_buf[0])))
        lizzieLet17_5QNone_Int_7QNode_Int_5QNone_Int_bufchan_buf <= lizzieLet17_5QNone_Int_7QNode_Int_5QNone_Int_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet17_5QNone_Int_7QNode_Int_5QVal_Int,Go) > [(lizzieLet17_5QNone_Int_7QNode_Int_5QVal_Int_1,Go),
                                                                   (lizzieLet17_5QNone_Int_7QNode_Int_5QVal_Int_2,Go)] */
  logic [1:0] lizzieLet17_5QNone_Int_7QNode_Int_5QVal_Int_emitted;
  logic [1:0] lizzieLet17_5QNone_Int_7QNode_Int_5QVal_Int_done;
  assign lizzieLet17_5QNone_Int_7QNode_Int_5QVal_Int_1_d = (lizzieLet17_5QNone_Int_7QNode_Int_5QVal_Int_d[0] && (! lizzieLet17_5QNone_Int_7QNode_Int_5QVal_Int_emitted[0]));
  assign lizzieLet17_5QNone_Int_7QNode_Int_5QVal_Int_2_d = (lizzieLet17_5QNone_Int_7QNode_Int_5QVal_Int_d[0] && (! lizzieLet17_5QNone_Int_7QNode_Int_5QVal_Int_emitted[1]));
  assign lizzieLet17_5QNone_Int_7QNode_Int_5QVal_Int_done = (lizzieLet17_5QNone_Int_7QNode_Int_5QVal_Int_emitted | ({lizzieLet17_5QNone_Int_7QNode_Int_5QVal_Int_2_d[0],
                                                                                                                     lizzieLet17_5QNone_Int_7QNode_Int_5QVal_Int_1_d[0]} & {lizzieLet17_5QNone_Int_7QNode_Int_5QVal_Int_2_r,
                                                                                                                                                                            lizzieLet17_5QNone_Int_7QNode_Int_5QVal_Int_1_r}));
  assign lizzieLet17_5QNone_Int_7QNode_Int_5QVal_Int_r = (& lizzieLet17_5QNone_Int_7QNode_Int_5QVal_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNone_Int_7QNode_Int_5QVal_Int_emitted <= 2'd0;
    else
      lizzieLet17_5QNone_Int_7QNode_Int_5QVal_Int_emitted <= (lizzieLet17_5QNone_Int_7QNode_Int_5QVal_Int_r ? 2'd0 :
                                                              lizzieLet17_5QNone_Int_7QNode_Int_5QVal_Int_done);
  
  /* dcon (Ty QTree_Int,
      Dcon QError_Int) : [(lizzieLet17_5QNone_Int_7QNode_Int_5QVal_Int_1,Go)] > (lizzieLet17_5QNone_Int_7QNode_Int_5QVal_Int_1QError_Int,QTree_Int) */
  assign lizzieLet17_5QNone_Int_7QNode_Int_5QVal_Int_1QError_Int_d = QError_Int_dc((& {lizzieLet17_5QNone_Int_7QNode_Int_5QVal_Int_1_d[0]}), lizzieLet17_5QNone_Int_7QNode_Int_5QVal_Int_1_d);
  assign {lizzieLet17_5QNone_Int_7QNode_Int_5QVal_Int_1_r} = {1 {(lizzieLet17_5QNone_Int_7QNode_Int_5QVal_Int_1QError_Int_r && lizzieLet17_5QNone_Int_7QNode_Int_5QVal_Int_1QError_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (lizzieLet17_5QNone_Int_7QNode_Int_5QVal_Int_1QError_Int,QTree_Int) > (lizzieLet25_1_argbuf,QTree_Int) */
  QTree_Int_t lizzieLet17_5QNone_Int_7QNode_Int_5QVal_Int_1QError_Int_bufchan_d;
  logic lizzieLet17_5QNone_Int_7QNode_Int_5QVal_Int_1QError_Int_bufchan_r;
  assign lizzieLet17_5QNone_Int_7QNode_Int_5QVal_Int_1QError_Int_r = ((! lizzieLet17_5QNone_Int_7QNode_Int_5QVal_Int_1QError_Int_bufchan_d[0]) || lizzieLet17_5QNone_Int_7QNode_Int_5QVal_Int_1QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNone_Int_7QNode_Int_5QVal_Int_1QError_Int_bufchan_d <= {66'd0,
                                                                            1'd0};
    else
      if (lizzieLet17_5QNone_Int_7QNode_Int_5QVal_Int_1QError_Int_r)
        lizzieLet17_5QNone_Int_7QNode_Int_5QVal_Int_1QError_Int_bufchan_d <= lizzieLet17_5QNone_Int_7QNode_Int_5QVal_Int_1QError_Int_d;
  QTree_Int_t lizzieLet17_5QNone_Int_7QNode_Int_5QVal_Int_1QError_Int_bufchan_buf;
  assign lizzieLet17_5QNone_Int_7QNode_Int_5QVal_Int_1QError_Int_bufchan_r = (! lizzieLet17_5QNone_Int_7QNode_Int_5QVal_Int_1QError_Int_bufchan_buf[0]);
  assign lizzieLet25_1_argbuf_d = (lizzieLet17_5QNone_Int_7QNode_Int_5QVal_Int_1QError_Int_bufchan_buf[0] ? lizzieLet17_5QNone_Int_7QNode_Int_5QVal_Int_1QError_Int_bufchan_buf :
                                   lizzieLet17_5QNone_Int_7QNode_Int_5QVal_Int_1QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNone_Int_7QNode_Int_5QVal_Int_1QError_Int_bufchan_buf <= {66'd0,
                                                                              1'd0};
    else
      if ((lizzieLet25_1_argbuf_r && lizzieLet17_5QNone_Int_7QNode_Int_5QVal_Int_1QError_Int_bufchan_buf[0]))
        lizzieLet17_5QNone_Int_7QNode_Int_5QVal_Int_1QError_Int_bufchan_buf <= {66'd0,
                                                                                1'd0};
      else if (((! lizzieLet25_1_argbuf_r) && (! lizzieLet17_5QNone_Int_7QNode_Int_5QVal_Int_1QError_Int_bufchan_buf[0])))
        lizzieLet17_5QNone_Int_7QNode_Int_5QVal_Int_1QError_Int_bufchan_buf <= lizzieLet17_5QNone_Int_7QNode_Int_5QVal_Int_1QError_Int_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet17_5QNone_Int_7QNode_Int_5QVal_Int_2,Go) > (lizzieLet17_5QNone_Int_7QNode_Int_5QVal_Int_2_argbuf,Go) */
  Go_t lizzieLet17_5QNone_Int_7QNode_Int_5QVal_Int_2_bufchan_d;
  logic lizzieLet17_5QNone_Int_7QNode_Int_5QVal_Int_2_bufchan_r;
  assign lizzieLet17_5QNone_Int_7QNode_Int_5QVal_Int_2_r = ((! lizzieLet17_5QNone_Int_7QNode_Int_5QVal_Int_2_bufchan_d[0]) || lizzieLet17_5QNone_Int_7QNode_Int_5QVal_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNone_Int_7QNode_Int_5QVal_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet17_5QNone_Int_7QNode_Int_5QVal_Int_2_r)
        lizzieLet17_5QNone_Int_7QNode_Int_5QVal_Int_2_bufchan_d <= lizzieLet17_5QNone_Int_7QNode_Int_5QVal_Int_2_d;
  Go_t lizzieLet17_5QNone_Int_7QNode_Int_5QVal_Int_2_bufchan_buf;
  assign lizzieLet17_5QNone_Int_7QNode_Int_5QVal_Int_2_bufchan_r = (! lizzieLet17_5QNone_Int_7QNode_Int_5QVal_Int_2_bufchan_buf[0]);
  assign lizzieLet17_5QNone_Int_7QNode_Int_5QVal_Int_2_argbuf_d = (lizzieLet17_5QNone_Int_7QNode_Int_5QVal_Int_2_bufchan_buf[0] ? lizzieLet17_5QNone_Int_7QNode_Int_5QVal_Int_2_bufchan_buf :
                                                                   lizzieLet17_5QNone_Int_7QNode_Int_5QVal_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNone_Int_7QNode_Int_5QVal_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet17_5QNone_Int_7QNode_Int_5QVal_Int_2_argbuf_r && lizzieLet17_5QNone_Int_7QNode_Int_5QVal_Int_2_bufchan_buf[0]))
        lizzieLet17_5QNone_Int_7QNode_Int_5QVal_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet17_5QNone_Int_7QNode_Int_5QVal_Int_2_argbuf_r) && (! lizzieLet17_5QNone_Int_7QNode_Int_5QVal_Int_2_bufchan_buf[0])))
        lizzieLet17_5QNone_Int_7QNode_Int_5QVal_Int_2_bufchan_buf <= lizzieLet17_5QNone_Int_7QNode_Int_5QVal_Int_2_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty MyDTInt_Bool) : (lizzieLet17_5QNone_Int_7QNode_Int_6,QTree_Int) (lizzieLet17_5QNone_Int_6QNode_Int,MyDTInt_Bool) > [(_132,MyDTInt_Bool),
                                                                                                                              (_131,MyDTInt_Bool),
                                                                                                                              (lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int,MyDTInt_Bool),
                                                                                                                              (_130,MyDTInt_Bool)] */
  logic [3:0] lizzieLet17_5QNone_Int_6QNode_Int_onehotd;
  always_comb
    if ((lizzieLet17_5QNone_Int_7QNode_Int_6_d[0] && lizzieLet17_5QNone_Int_6QNode_Int_d[0]))
      unique case (lizzieLet17_5QNone_Int_7QNode_Int_6_d[2:1])
        2'd0: lizzieLet17_5QNone_Int_6QNode_Int_onehotd = 4'd1;
        2'd1: lizzieLet17_5QNone_Int_6QNode_Int_onehotd = 4'd2;
        2'd2: lizzieLet17_5QNone_Int_6QNode_Int_onehotd = 4'd4;
        2'd3: lizzieLet17_5QNone_Int_6QNode_Int_onehotd = 4'd8;
        default: lizzieLet17_5QNone_Int_6QNode_Int_onehotd = 4'd0;
      endcase
    else lizzieLet17_5QNone_Int_6QNode_Int_onehotd = 4'd0;
  assign _132_d = lizzieLet17_5QNone_Int_6QNode_Int_onehotd[0];
  assign _131_d = lizzieLet17_5QNone_Int_6QNode_Int_onehotd[1];
  assign lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_d = lizzieLet17_5QNone_Int_6QNode_Int_onehotd[2];
  assign _130_d = lizzieLet17_5QNone_Int_6QNode_Int_onehotd[3];
  assign lizzieLet17_5QNone_Int_6QNode_Int_r = (| (lizzieLet17_5QNone_Int_6QNode_Int_onehotd & {_130_r,
                                                                                                lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_r,
                                                                                                _131_r,
                                                                                                _132_r}));
  assign lizzieLet17_5QNone_Int_7QNode_Int_6_r = lizzieLet17_5QNone_Int_6QNode_Int_r;
  
  /* fork (Ty MyDTInt_Bool) : (lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int,MyDTInt_Bool) > [(lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_1,MyDTInt_Bool),
                                                                                        (lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_2,MyDTInt_Bool),
                                                                                        (lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_3,MyDTInt_Bool),
                                                                                        (lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_4,MyDTInt_Bool)] */
  logic [3:0] lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_emitted;
  logic [3:0] lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_done;
  assign lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_1_d = (lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_d[0] && (! lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_emitted[0]));
  assign lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_2_d = (lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_d[0] && (! lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_emitted[1]));
  assign lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_3_d = (lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_d[0] && (! lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_emitted[2]));
  assign lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_4_d = (lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_d[0] && (! lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_emitted[3]));
  assign lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_done = (lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_emitted | ({lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_4_d[0],
                                                                                                                       lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_3_d[0],
                                                                                                                       lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_2_d[0],
                                                                                                                       lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_1_d[0]} & {lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_4_r,
                                                                                                                                                                               lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_3_r,
                                                                                                                                                                               lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_2_r,
                                                                                                                                                                               lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_1_r}));
  assign lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_r = (& lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_emitted <= 4'd0;
    else
      lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_emitted <= (lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_r ? 4'd0 :
                                                               lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_done);
  
  /* buf (Ty MyDTInt_Bool) : (lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_1,MyDTInt_Bool) > (lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_1_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_1_bufchan_d;
  logic lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_1_bufchan_r;
  assign lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_1_r = ((! lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_1_bufchan_d[0]) || lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_1_bufchan_d <= 1'd0;
    else
      if (lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_1_r)
        lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_1_bufchan_d <= lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_1_d;
  MyDTInt_Bool_t lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_1_bufchan_buf;
  assign lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_1_bufchan_r = (! lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_1_bufchan_buf[0]);
  assign lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_1_argbuf_d = (lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_1_bufchan_buf[0] ? lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_1_bufchan_buf :
                                                                    lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_1_argbuf_r && lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_1_bufchan_buf[0]))
        lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_1_argbuf_r) && (! lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_1_bufchan_buf[0])))
        lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_1_bufchan_buf <= lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_1_bufchan_d;
  
  /* buf (Ty MyDTInt_Bool) : (lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_2,MyDTInt_Bool) > (lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_2_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_2_bufchan_d;
  logic lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_2_bufchan_r;
  assign lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_2_r = ((! lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_2_bufchan_d[0]) || lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_2_r)
        lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_2_bufchan_d <= lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_2_d;
  MyDTInt_Bool_t lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_2_bufchan_buf;
  assign lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_2_bufchan_r = (! lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_2_bufchan_buf[0]);
  assign lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_2_argbuf_d = (lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_2_bufchan_buf[0] ? lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_2_bufchan_buf :
                                                                    lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_2_argbuf_r && lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_2_bufchan_buf[0]))
        lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_2_argbuf_r) && (! lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_2_bufchan_buf[0])))
        lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_2_bufchan_buf <= lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_2_bufchan_d;
  
  /* buf (Ty MyDTInt_Bool) : (lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_3,MyDTInt_Bool) > (lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_3_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_3_bufchan_d;
  logic lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_3_bufchan_r;
  assign lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_3_r = ((! lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_3_bufchan_d[0]) || lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_3_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_3_bufchan_d <= 1'd0;
    else
      if (lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_3_r)
        lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_3_bufchan_d <= lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_3_d;
  MyDTInt_Bool_t lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_3_bufchan_buf;
  assign lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_3_bufchan_r = (! lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_3_bufchan_buf[0]);
  assign lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_3_argbuf_d = (lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_3_bufchan_buf[0] ? lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_3_bufchan_buf :
                                                                    lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_3_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_3_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_3_argbuf_r && lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_3_bufchan_buf[0]))
        lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_3_bufchan_buf <= 1'd0;
      else if (((! lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_3_argbuf_r) && (! lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_3_bufchan_buf[0])))
        lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_3_bufchan_buf <= lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_3_bufchan_d;
  
  /* buf (Ty MyDTInt_Bool) : (lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_4,MyDTInt_Bool) > (lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_4_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_4_bufchan_d;
  logic lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_4_bufchan_r;
  assign lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_4_r = ((! lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_4_bufchan_d[0]) || lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_4_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_4_bufchan_d <= 1'd0;
    else
      if (lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_4_r)
        lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_4_bufchan_d <= lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_4_d;
  MyDTInt_Bool_t lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_4_bufchan_buf;
  assign lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_4_bufchan_r = (! lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_4_bufchan_buf[0]);
  assign lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_4_argbuf_d = (lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_4_bufchan_buf[0] ? lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_4_bufchan_buf :
                                                                    lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_4_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_4_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_4_argbuf_r && lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_4_bufchan_buf[0]))
        lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_4_bufchan_buf <= 1'd0;
      else if (((! lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_4_argbuf_r) && (! lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_4_bufchan_buf[0])))
        lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_4_bufchan_buf <= lizzieLet17_5QNone_Int_7QNode_Int_6QNode_Int_4_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_QTree_Int) : (lizzieLet17_5QNone_Int_7QNode_Int_7,QTree_Int) (lizzieLet17_5QNone_Int_8QNode_Int,Pointer_QTree_Int) > [(lizzieLet17_5QNone_Int_7QNode_Int_7QNone_Int,Pointer_QTree_Int),
                                                                                                                                        (_129,Pointer_QTree_Int),
                                                                                                                                        (_128,Pointer_QTree_Int),
                                                                                                                                        (_127,Pointer_QTree_Int)] */
  logic [3:0] lizzieLet17_5QNone_Int_8QNode_Int_onehotd;
  always_comb
    if ((lizzieLet17_5QNone_Int_7QNode_Int_7_d[0] && lizzieLet17_5QNone_Int_8QNode_Int_d[0]))
      unique case (lizzieLet17_5QNone_Int_7QNode_Int_7_d[2:1])
        2'd0: lizzieLet17_5QNone_Int_8QNode_Int_onehotd = 4'd1;
        2'd1: lizzieLet17_5QNone_Int_8QNode_Int_onehotd = 4'd2;
        2'd2: lizzieLet17_5QNone_Int_8QNode_Int_onehotd = 4'd4;
        2'd3: lizzieLet17_5QNone_Int_8QNode_Int_onehotd = 4'd8;
        default: lizzieLet17_5QNone_Int_8QNode_Int_onehotd = 4'd0;
      endcase
    else lizzieLet17_5QNone_Int_8QNode_Int_onehotd = 4'd0;
  assign lizzieLet17_5QNone_Int_7QNode_Int_7QNone_Int_d = {lizzieLet17_5QNone_Int_8QNode_Int_d[16:1],
                                                           lizzieLet17_5QNone_Int_8QNode_Int_onehotd[0]};
  assign _129_d = {lizzieLet17_5QNone_Int_8QNode_Int_d[16:1],
                   lizzieLet17_5QNone_Int_8QNode_Int_onehotd[1]};
  assign _128_d = {lizzieLet17_5QNone_Int_8QNode_Int_d[16:1],
                   lizzieLet17_5QNone_Int_8QNode_Int_onehotd[2]};
  assign _127_d = {lizzieLet17_5QNone_Int_8QNode_Int_d[16:1],
                   lizzieLet17_5QNone_Int_8QNode_Int_onehotd[3]};
  assign lizzieLet17_5QNone_Int_8QNode_Int_r = (| (lizzieLet17_5QNone_Int_8QNode_Int_onehotd & {_127_r,
                                                                                                _128_r,
                                                                                                _129_r,
                                                                                                lizzieLet17_5QNone_Int_7QNode_Int_7QNone_Int_r}));
  assign lizzieLet17_5QNone_Int_7QNode_Int_7_r = lizzieLet17_5QNone_Int_8QNode_Int_r;
  
  /* buf (Ty Pointer_QTree_Int) : (lizzieLet17_5QNone_Int_7QNode_Int_7QNone_Int,Pointer_QTree_Int) > (lizzieLet17_5QNone_Int_7QNode_Int_7QNone_Int_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t lizzieLet17_5QNone_Int_7QNode_Int_7QNone_Int_bufchan_d;
  logic lizzieLet17_5QNone_Int_7QNode_Int_7QNone_Int_bufchan_r;
  assign lizzieLet17_5QNone_Int_7QNode_Int_7QNone_Int_r = ((! lizzieLet17_5QNone_Int_7QNode_Int_7QNone_Int_bufchan_d[0]) || lizzieLet17_5QNone_Int_7QNode_Int_7QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNone_Int_7QNode_Int_7QNone_Int_bufchan_d <= {16'd0,
                                                                 1'd0};
    else
      if (lizzieLet17_5QNone_Int_7QNode_Int_7QNone_Int_r)
        lizzieLet17_5QNone_Int_7QNode_Int_7QNone_Int_bufchan_d <= lizzieLet17_5QNone_Int_7QNode_Int_7QNone_Int_d;
  Pointer_QTree_Int_t lizzieLet17_5QNone_Int_7QNode_Int_7QNone_Int_bufchan_buf;
  assign lizzieLet17_5QNone_Int_7QNode_Int_7QNone_Int_bufchan_r = (! lizzieLet17_5QNone_Int_7QNode_Int_7QNone_Int_bufchan_buf[0]);
  assign lizzieLet17_5QNone_Int_7QNode_Int_7QNone_Int_1_argbuf_d = (lizzieLet17_5QNone_Int_7QNode_Int_7QNone_Int_bufchan_buf[0] ? lizzieLet17_5QNone_Int_7QNode_Int_7QNone_Int_bufchan_buf :
                                                                    lizzieLet17_5QNone_Int_7QNode_Int_7QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNone_Int_7QNode_Int_7QNone_Int_bufchan_buf <= {16'd0,
                                                                   1'd0};
    else
      if ((lizzieLet17_5QNone_Int_7QNode_Int_7QNone_Int_1_argbuf_r && lizzieLet17_5QNone_Int_7QNode_Int_7QNone_Int_bufchan_buf[0]))
        lizzieLet17_5QNone_Int_7QNode_Int_7QNone_Int_bufchan_buf <= {16'd0,
                                                                     1'd0};
      else if (((! lizzieLet17_5QNone_Int_7QNode_Int_7QNone_Int_1_argbuf_r) && (! lizzieLet17_5QNone_Int_7QNode_Int_7QNone_Int_bufchan_buf[0])))
        lizzieLet17_5QNone_Int_7QNode_Int_7QNone_Int_bufchan_buf <= lizzieLet17_5QNone_Int_7QNode_Int_7QNone_Int_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_QTree_Int) : (lizzieLet17_5QNone_Int_7QNode_Int_8,QTree_Int) (q1aeB_destruct,Pointer_QTree_Int) > [(_126,Pointer_QTree_Int),
                                                                                                                     (_125,Pointer_QTree_Int),
                                                                                                                     (lizzieLet17_5QNone_Int_7QNode_Int_8QNode_Int,Pointer_QTree_Int),
                                                                                                                     (_124,Pointer_QTree_Int)] */
  logic [3:0] q1aeB_destruct_onehotd;
  always_comb
    if ((lizzieLet17_5QNone_Int_7QNode_Int_8_d[0] && q1aeB_destruct_d[0]))
      unique case (lizzieLet17_5QNone_Int_7QNode_Int_8_d[2:1])
        2'd0: q1aeB_destruct_onehotd = 4'd1;
        2'd1: q1aeB_destruct_onehotd = 4'd2;
        2'd2: q1aeB_destruct_onehotd = 4'd4;
        2'd3: q1aeB_destruct_onehotd = 4'd8;
        default: q1aeB_destruct_onehotd = 4'd0;
      endcase
    else q1aeB_destruct_onehotd = 4'd0;
  assign _126_d = {q1aeB_destruct_d[16:1],
                   q1aeB_destruct_onehotd[0]};
  assign _125_d = {q1aeB_destruct_d[16:1],
                   q1aeB_destruct_onehotd[1]};
  assign lizzieLet17_5QNone_Int_7QNode_Int_8QNode_Int_d = {q1aeB_destruct_d[16:1],
                                                           q1aeB_destruct_onehotd[2]};
  assign _124_d = {q1aeB_destruct_d[16:1],
                   q1aeB_destruct_onehotd[3]};
  assign q1aeB_destruct_r = (| (q1aeB_destruct_onehotd & {_124_r,
                                                          lizzieLet17_5QNone_Int_7QNode_Int_8QNode_Int_r,
                                                          _125_r,
                                                          _126_r}));
  assign lizzieLet17_5QNone_Int_7QNode_Int_8_r = q1aeB_destruct_r;
  
  /* buf (Ty Pointer_QTree_Int) : (lizzieLet17_5QNone_Int_7QNode_Int_8QNode_Int,Pointer_QTree_Int) > (lizzieLet17_5QNone_Int_7QNode_Int_8QNode_Int_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t lizzieLet17_5QNone_Int_7QNode_Int_8QNode_Int_bufchan_d;
  logic lizzieLet17_5QNone_Int_7QNode_Int_8QNode_Int_bufchan_r;
  assign lizzieLet17_5QNone_Int_7QNode_Int_8QNode_Int_r = ((! lizzieLet17_5QNone_Int_7QNode_Int_8QNode_Int_bufchan_d[0]) || lizzieLet17_5QNone_Int_7QNode_Int_8QNode_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNone_Int_7QNode_Int_8QNode_Int_bufchan_d <= {16'd0,
                                                                 1'd0};
    else
      if (lizzieLet17_5QNone_Int_7QNode_Int_8QNode_Int_r)
        lizzieLet17_5QNone_Int_7QNode_Int_8QNode_Int_bufchan_d <= lizzieLet17_5QNone_Int_7QNode_Int_8QNode_Int_d;
  Pointer_QTree_Int_t lizzieLet17_5QNone_Int_7QNode_Int_8QNode_Int_bufchan_buf;
  assign lizzieLet17_5QNone_Int_7QNode_Int_8QNode_Int_bufchan_r = (! lizzieLet17_5QNone_Int_7QNode_Int_8QNode_Int_bufchan_buf[0]);
  assign lizzieLet17_5QNone_Int_7QNode_Int_8QNode_Int_1_argbuf_d = (lizzieLet17_5QNone_Int_7QNode_Int_8QNode_Int_bufchan_buf[0] ? lizzieLet17_5QNone_Int_7QNode_Int_8QNode_Int_bufchan_buf :
                                                                    lizzieLet17_5QNone_Int_7QNode_Int_8QNode_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNone_Int_7QNode_Int_8QNode_Int_bufchan_buf <= {16'd0,
                                                                   1'd0};
    else
      if ((lizzieLet17_5QNone_Int_7QNode_Int_8QNode_Int_1_argbuf_r && lizzieLet17_5QNone_Int_7QNode_Int_8QNode_Int_bufchan_buf[0]))
        lizzieLet17_5QNone_Int_7QNode_Int_8QNode_Int_bufchan_buf <= {16'd0,
                                                                     1'd0};
      else if (((! lizzieLet17_5QNone_Int_7QNode_Int_8QNode_Int_1_argbuf_r) && (! lizzieLet17_5QNone_Int_7QNode_Int_8QNode_Int_bufchan_buf[0])))
        lizzieLet17_5QNone_Int_7QNode_Int_8QNode_Int_bufchan_buf <= lizzieLet17_5QNone_Int_7QNode_Int_8QNode_Int_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_QTree_Int) : (lizzieLet17_5QNone_Int_7QNode_Int_9,QTree_Int) (q2aeC_destruct,Pointer_QTree_Int) > [(_123,Pointer_QTree_Int),
                                                                                                                     (_122,Pointer_QTree_Int),
                                                                                                                     (lizzieLet17_5QNone_Int_7QNode_Int_9QNode_Int,Pointer_QTree_Int),
                                                                                                                     (_121,Pointer_QTree_Int)] */
  logic [3:0] q2aeC_destruct_onehotd;
  always_comb
    if ((lizzieLet17_5QNone_Int_7QNode_Int_9_d[0] && q2aeC_destruct_d[0]))
      unique case (lizzieLet17_5QNone_Int_7QNode_Int_9_d[2:1])
        2'd0: q2aeC_destruct_onehotd = 4'd1;
        2'd1: q2aeC_destruct_onehotd = 4'd2;
        2'd2: q2aeC_destruct_onehotd = 4'd4;
        2'd3: q2aeC_destruct_onehotd = 4'd8;
        default: q2aeC_destruct_onehotd = 4'd0;
      endcase
    else q2aeC_destruct_onehotd = 4'd0;
  assign _123_d = {q2aeC_destruct_d[16:1],
                   q2aeC_destruct_onehotd[0]};
  assign _122_d = {q2aeC_destruct_d[16:1],
                   q2aeC_destruct_onehotd[1]};
  assign lizzieLet17_5QNone_Int_7QNode_Int_9QNode_Int_d = {q2aeC_destruct_d[16:1],
                                                           q2aeC_destruct_onehotd[2]};
  assign _121_d = {q2aeC_destruct_d[16:1],
                   q2aeC_destruct_onehotd[3]};
  assign q2aeC_destruct_r = (| (q2aeC_destruct_onehotd & {_121_r,
                                                          lizzieLet17_5QNone_Int_7QNode_Int_9QNode_Int_r,
                                                          _122_r,
                                                          _123_r}));
  assign lizzieLet17_5QNone_Int_7QNode_Int_9_r = q2aeC_destruct_r;
  
  /* buf (Ty Pointer_QTree_Int) : (lizzieLet17_5QNone_Int_7QNode_Int_9QNode_Int,Pointer_QTree_Int) > (lizzieLet17_5QNone_Int_7QNode_Int_9QNode_Int_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t lizzieLet17_5QNone_Int_7QNode_Int_9QNode_Int_bufchan_d;
  logic lizzieLet17_5QNone_Int_7QNode_Int_9QNode_Int_bufchan_r;
  assign lizzieLet17_5QNone_Int_7QNode_Int_9QNode_Int_r = ((! lizzieLet17_5QNone_Int_7QNode_Int_9QNode_Int_bufchan_d[0]) || lizzieLet17_5QNone_Int_7QNode_Int_9QNode_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNone_Int_7QNode_Int_9QNode_Int_bufchan_d <= {16'd0,
                                                                 1'd0};
    else
      if (lizzieLet17_5QNone_Int_7QNode_Int_9QNode_Int_r)
        lizzieLet17_5QNone_Int_7QNode_Int_9QNode_Int_bufchan_d <= lizzieLet17_5QNone_Int_7QNode_Int_9QNode_Int_d;
  Pointer_QTree_Int_t lizzieLet17_5QNone_Int_7QNode_Int_9QNode_Int_bufchan_buf;
  assign lizzieLet17_5QNone_Int_7QNode_Int_9QNode_Int_bufchan_r = (! lizzieLet17_5QNone_Int_7QNode_Int_9QNode_Int_bufchan_buf[0]);
  assign lizzieLet17_5QNone_Int_7QNode_Int_9QNode_Int_1_argbuf_d = (lizzieLet17_5QNone_Int_7QNode_Int_9QNode_Int_bufchan_buf[0] ? lizzieLet17_5QNone_Int_7QNode_Int_9QNode_Int_bufchan_buf :
                                                                    lizzieLet17_5QNone_Int_7QNode_Int_9QNode_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNone_Int_7QNode_Int_9QNode_Int_bufchan_buf <= {16'd0,
                                                                   1'd0};
    else
      if ((lizzieLet17_5QNone_Int_7QNode_Int_9QNode_Int_1_argbuf_r && lizzieLet17_5QNone_Int_7QNode_Int_9QNode_Int_bufchan_buf[0]))
        lizzieLet17_5QNone_Int_7QNode_Int_9QNode_Int_bufchan_buf <= {16'd0,
                                                                     1'd0};
      else if (((! lizzieLet17_5QNone_Int_7QNode_Int_9QNode_Int_1_argbuf_r) && (! lizzieLet17_5QNone_Int_7QNode_Int_9QNode_Int_bufchan_buf[0])))
        lizzieLet17_5QNone_Int_7QNode_Int_9QNode_Int_bufchan_buf <= lizzieLet17_5QNone_Int_7QNode_Int_9QNode_Int_bufchan_d;
  
  /* fork (Ty QTree_Int) : (lizzieLet17_5QNone_Int_7QVal_Int,QTree_Int) > [(lizzieLet17_5QNone_Int_7QVal_Int_1,QTree_Int),
                                                                      (lizzieLet17_5QNone_Int_7QVal_Int_2,QTree_Int),
                                                                      (lizzieLet17_5QNone_Int_7QVal_Int_3,QTree_Int),
                                                                      (lizzieLet17_5QNone_Int_7QVal_Int_4,QTree_Int),
                                                                      (lizzieLet17_5QNone_Int_7QVal_Int_5,QTree_Int),
                                                                      (lizzieLet17_5QNone_Int_7QVal_Int_6,QTree_Int),
                                                                      (lizzieLet17_5QNone_Int_7QVal_Int_7,QTree_Int),
                                                                      (lizzieLet17_5QNone_Int_7QVal_Int_8,QTree_Int)] */
  logic [7:0] lizzieLet17_5QNone_Int_7QVal_Int_emitted;
  logic [7:0] lizzieLet17_5QNone_Int_7QVal_Int_done;
  assign lizzieLet17_5QNone_Int_7QVal_Int_1_d = {lizzieLet17_5QNone_Int_7QVal_Int_d[66:1],
                                                 (lizzieLet17_5QNone_Int_7QVal_Int_d[0] && (! lizzieLet17_5QNone_Int_7QVal_Int_emitted[0]))};
  assign lizzieLet17_5QNone_Int_7QVal_Int_2_d = {lizzieLet17_5QNone_Int_7QVal_Int_d[66:1],
                                                 (lizzieLet17_5QNone_Int_7QVal_Int_d[0] && (! lizzieLet17_5QNone_Int_7QVal_Int_emitted[1]))};
  assign lizzieLet17_5QNone_Int_7QVal_Int_3_d = {lizzieLet17_5QNone_Int_7QVal_Int_d[66:1],
                                                 (lizzieLet17_5QNone_Int_7QVal_Int_d[0] && (! lizzieLet17_5QNone_Int_7QVal_Int_emitted[2]))};
  assign lizzieLet17_5QNone_Int_7QVal_Int_4_d = {lizzieLet17_5QNone_Int_7QVal_Int_d[66:1],
                                                 (lizzieLet17_5QNone_Int_7QVal_Int_d[0] && (! lizzieLet17_5QNone_Int_7QVal_Int_emitted[3]))};
  assign lizzieLet17_5QNone_Int_7QVal_Int_5_d = {lizzieLet17_5QNone_Int_7QVal_Int_d[66:1],
                                                 (lizzieLet17_5QNone_Int_7QVal_Int_d[0] && (! lizzieLet17_5QNone_Int_7QVal_Int_emitted[4]))};
  assign lizzieLet17_5QNone_Int_7QVal_Int_6_d = {lizzieLet17_5QNone_Int_7QVal_Int_d[66:1],
                                                 (lizzieLet17_5QNone_Int_7QVal_Int_d[0] && (! lizzieLet17_5QNone_Int_7QVal_Int_emitted[5]))};
  assign lizzieLet17_5QNone_Int_7QVal_Int_7_d = {lizzieLet17_5QNone_Int_7QVal_Int_d[66:1],
                                                 (lizzieLet17_5QNone_Int_7QVal_Int_d[0] && (! lizzieLet17_5QNone_Int_7QVal_Int_emitted[6]))};
  assign lizzieLet17_5QNone_Int_7QVal_Int_8_d = {lizzieLet17_5QNone_Int_7QVal_Int_d[66:1],
                                                 (lizzieLet17_5QNone_Int_7QVal_Int_d[0] && (! lizzieLet17_5QNone_Int_7QVal_Int_emitted[7]))};
  assign lizzieLet17_5QNone_Int_7QVal_Int_done = (lizzieLet17_5QNone_Int_7QVal_Int_emitted | ({lizzieLet17_5QNone_Int_7QVal_Int_8_d[0],
                                                                                               lizzieLet17_5QNone_Int_7QVal_Int_7_d[0],
                                                                                               lizzieLet17_5QNone_Int_7QVal_Int_6_d[0],
                                                                                               lizzieLet17_5QNone_Int_7QVal_Int_5_d[0],
                                                                                               lizzieLet17_5QNone_Int_7QVal_Int_4_d[0],
                                                                                               lizzieLet17_5QNone_Int_7QVal_Int_3_d[0],
                                                                                               lizzieLet17_5QNone_Int_7QVal_Int_2_d[0],
                                                                                               lizzieLet17_5QNone_Int_7QVal_Int_1_d[0]} & {lizzieLet17_5QNone_Int_7QVal_Int_8_r,
                                                                                                                                           lizzieLet17_5QNone_Int_7QVal_Int_7_r,
                                                                                                                                           lizzieLet17_5QNone_Int_7QVal_Int_6_r,
                                                                                                                                           lizzieLet17_5QNone_Int_7QVal_Int_5_r,
                                                                                                                                           lizzieLet17_5QNone_Int_7QVal_Int_4_r,
                                                                                                                                           lizzieLet17_5QNone_Int_7QVal_Int_3_r,
                                                                                                                                           lizzieLet17_5QNone_Int_7QVal_Int_2_r,
                                                                                                                                           lizzieLet17_5QNone_Int_7QVal_Int_1_r}));
  assign lizzieLet17_5QNone_Int_7QVal_Int_r = (& lizzieLet17_5QNone_Int_7QVal_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNone_Int_7QVal_Int_emitted <= 8'd0;
    else
      lizzieLet17_5QNone_Int_7QVal_Int_emitted <= (lizzieLet17_5QNone_Int_7QVal_Int_r ? 8'd0 :
                                                   lizzieLet17_5QNone_Int_7QVal_Int_done);
  
  /* destruct (Ty QTree_Int,
          Dcon QVal_Int) : (lizzieLet17_5QNone_Int_7QVal_Int_1QVal_Int,QTree_Int) > [(vaew_destruct,Int)] */
  assign vaew_destruct_d = {lizzieLet17_5QNone_Int_7QVal_Int_1QVal_Int_d[34:3],
                            lizzieLet17_5QNone_Int_7QVal_Int_1QVal_Int_d[0]};
  assign lizzieLet17_5QNone_Int_7QVal_Int_1QVal_Int_r = vaew_destruct_r;
  
  /* demux (Ty QTree_Int,
       Ty QTree_Int) : (lizzieLet17_5QNone_Int_7QVal_Int_2,QTree_Int) (lizzieLet17_5QNone_Int_7QVal_Int_1,QTree_Int) > [(_120,QTree_Int),
                                                                                                                        (lizzieLet17_5QNone_Int_7QVal_Int_1QVal_Int,QTree_Int),
                                                                                                                        (_119,QTree_Int),
                                                                                                                        (_118,QTree_Int)] */
  logic [3:0] lizzieLet17_5QNone_Int_7QVal_Int_1_onehotd;
  always_comb
    if ((lizzieLet17_5QNone_Int_7QVal_Int_2_d[0] && lizzieLet17_5QNone_Int_7QVal_Int_1_d[0]))
      unique case (lizzieLet17_5QNone_Int_7QVal_Int_2_d[2:1])
        2'd0: lizzieLet17_5QNone_Int_7QVal_Int_1_onehotd = 4'd1;
        2'd1: lizzieLet17_5QNone_Int_7QVal_Int_1_onehotd = 4'd2;
        2'd2: lizzieLet17_5QNone_Int_7QVal_Int_1_onehotd = 4'd4;
        2'd3: lizzieLet17_5QNone_Int_7QVal_Int_1_onehotd = 4'd8;
        default: lizzieLet17_5QNone_Int_7QVal_Int_1_onehotd = 4'd0;
      endcase
    else lizzieLet17_5QNone_Int_7QVal_Int_1_onehotd = 4'd0;
  assign _120_d = {lizzieLet17_5QNone_Int_7QVal_Int_1_d[66:1],
                   lizzieLet17_5QNone_Int_7QVal_Int_1_onehotd[0]};
  assign lizzieLet17_5QNone_Int_7QVal_Int_1QVal_Int_d = {lizzieLet17_5QNone_Int_7QVal_Int_1_d[66:1],
                                                         lizzieLet17_5QNone_Int_7QVal_Int_1_onehotd[1]};
  assign _119_d = {lizzieLet17_5QNone_Int_7QVal_Int_1_d[66:1],
                   lizzieLet17_5QNone_Int_7QVal_Int_1_onehotd[2]};
  assign _118_d = {lizzieLet17_5QNone_Int_7QVal_Int_1_d[66:1],
                   lizzieLet17_5QNone_Int_7QVal_Int_1_onehotd[3]};
  assign lizzieLet17_5QNone_Int_7QVal_Int_1_r = (| (lizzieLet17_5QNone_Int_7QVal_Int_1_onehotd & {_118_r,
                                                                                                  _119_r,
                                                                                                  lizzieLet17_5QNone_Int_7QVal_Int_1QVal_Int_r,
                                                                                                  _120_r}));
  assign lizzieLet17_5QNone_Int_7QVal_Int_2_r = lizzieLet17_5QNone_Int_7QVal_Int_1_r;
  
  /* demux (Ty QTree_Int,
       Ty MyDTInt_Int_Int) : (lizzieLet17_5QNone_Int_7QVal_Int_3,QTree_Int) (lizzieLet17_5QNone_Int_3QVal_Int,MyDTInt_Int_Int) > [(_117,MyDTInt_Int_Int),
                                                                                                                                  (lizzieLet17_5QNone_Int_7QVal_Int_3QVal_Int,MyDTInt_Int_Int),
                                                                                                                                  (_116,MyDTInt_Int_Int),
                                                                                                                                  (_115,MyDTInt_Int_Int)] */
  logic [3:0] lizzieLet17_5QNone_Int_3QVal_Int_onehotd;
  always_comb
    if ((lizzieLet17_5QNone_Int_7QVal_Int_3_d[0] && lizzieLet17_5QNone_Int_3QVal_Int_d[0]))
      unique case (lizzieLet17_5QNone_Int_7QVal_Int_3_d[2:1])
        2'd0: lizzieLet17_5QNone_Int_3QVal_Int_onehotd = 4'd1;
        2'd1: lizzieLet17_5QNone_Int_3QVal_Int_onehotd = 4'd2;
        2'd2: lizzieLet17_5QNone_Int_3QVal_Int_onehotd = 4'd4;
        2'd3: lizzieLet17_5QNone_Int_3QVal_Int_onehotd = 4'd8;
        default: lizzieLet17_5QNone_Int_3QVal_Int_onehotd = 4'd0;
      endcase
    else lizzieLet17_5QNone_Int_3QVal_Int_onehotd = 4'd0;
  assign _117_d = lizzieLet17_5QNone_Int_3QVal_Int_onehotd[0];
  assign lizzieLet17_5QNone_Int_7QVal_Int_3QVal_Int_d = lizzieLet17_5QNone_Int_3QVal_Int_onehotd[1];
  assign _116_d = lizzieLet17_5QNone_Int_3QVal_Int_onehotd[2];
  assign _115_d = lizzieLet17_5QNone_Int_3QVal_Int_onehotd[3];
  assign lizzieLet17_5QNone_Int_3QVal_Int_r = (| (lizzieLet17_5QNone_Int_3QVal_Int_onehotd & {_115_r,
                                                                                              _116_r,
                                                                                              lizzieLet17_5QNone_Int_7QVal_Int_3QVal_Int_r,
                                                                                              _117_r}));
  assign lizzieLet17_5QNone_Int_7QVal_Int_3_r = lizzieLet17_5QNone_Int_3QVal_Int_r;
  
  /* fork (Ty MyDTInt_Int_Int) : (lizzieLet17_5QNone_Int_7QVal_Int_3QVal_Int,MyDTInt_Int_Int) > [(lizzieLet17_5QNone_Int_7QVal_Int_3QVal_Int_1,MyDTInt_Int_Int),
                                                                                            (lizzieLet17_5QNone_Int_7QVal_Int_3QVal_Int_2,MyDTInt_Int_Int)] */
  logic [1:0] lizzieLet17_5QNone_Int_7QVal_Int_3QVal_Int_emitted;
  logic [1:0] lizzieLet17_5QNone_Int_7QVal_Int_3QVal_Int_done;
  assign lizzieLet17_5QNone_Int_7QVal_Int_3QVal_Int_1_d = (lizzieLet17_5QNone_Int_7QVal_Int_3QVal_Int_d[0] && (! lizzieLet17_5QNone_Int_7QVal_Int_3QVal_Int_emitted[0]));
  assign lizzieLet17_5QNone_Int_7QVal_Int_3QVal_Int_2_d = (lizzieLet17_5QNone_Int_7QVal_Int_3QVal_Int_d[0] && (! lizzieLet17_5QNone_Int_7QVal_Int_3QVal_Int_emitted[1]));
  assign lizzieLet17_5QNone_Int_7QVal_Int_3QVal_Int_done = (lizzieLet17_5QNone_Int_7QVal_Int_3QVal_Int_emitted | ({lizzieLet17_5QNone_Int_7QVal_Int_3QVal_Int_2_d[0],
                                                                                                                   lizzieLet17_5QNone_Int_7QVal_Int_3QVal_Int_1_d[0]} & {lizzieLet17_5QNone_Int_7QVal_Int_3QVal_Int_2_r,
                                                                                                                                                                         lizzieLet17_5QNone_Int_7QVal_Int_3QVal_Int_1_r}));
  assign lizzieLet17_5QNone_Int_7QVal_Int_3QVal_Int_r = (& lizzieLet17_5QNone_Int_7QVal_Int_3QVal_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNone_Int_7QVal_Int_3QVal_Int_emitted <= 2'd0;
    else
      lizzieLet17_5QNone_Int_7QVal_Int_3QVal_Int_emitted <= (lizzieLet17_5QNone_Int_7QVal_Int_3QVal_Int_r ? 2'd0 :
                                                             lizzieLet17_5QNone_Int_7QVal_Int_3QVal_Int_done);
  
  /* buf (Ty MyDTInt_Int_Int) : (lizzieLet17_5QNone_Int_7QVal_Int_3QVal_Int_1,MyDTInt_Int_Int) > (lizzieLet17_5QNone_Int_7QVal_Int_3QVal_Int_1_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t lizzieLet17_5QNone_Int_7QVal_Int_3QVal_Int_1_bufchan_d;
  logic lizzieLet17_5QNone_Int_7QVal_Int_3QVal_Int_1_bufchan_r;
  assign lizzieLet17_5QNone_Int_7QVal_Int_3QVal_Int_1_r = ((! lizzieLet17_5QNone_Int_7QVal_Int_3QVal_Int_1_bufchan_d[0]) || lizzieLet17_5QNone_Int_7QVal_Int_3QVal_Int_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNone_Int_7QVal_Int_3QVal_Int_1_bufchan_d <= 1'd0;
    else
      if (lizzieLet17_5QNone_Int_7QVal_Int_3QVal_Int_1_r)
        lizzieLet17_5QNone_Int_7QVal_Int_3QVal_Int_1_bufchan_d <= lizzieLet17_5QNone_Int_7QVal_Int_3QVal_Int_1_d;
  MyDTInt_Int_Int_t lizzieLet17_5QNone_Int_7QVal_Int_3QVal_Int_1_bufchan_buf;
  assign lizzieLet17_5QNone_Int_7QVal_Int_3QVal_Int_1_bufchan_r = (! lizzieLet17_5QNone_Int_7QVal_Int_3QVal_Int_1_bufchan_buf[0]);
  assign lizzieLet17_5QNone_Int_7QVal_Int_3QVal_Int_1_argbuf_d = (lizzieLet17_5QNone_Int_7QVal_Int_3QVal_Int_1_bufchan_buf[0] ? lizzieLet17_5QNone_Int_7QVal_Int_3QVal_Int_1_bufchan_buf :
                                                                  lizzieLet17_5QNone_Int_7QVal_Int_3QVal_Int_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNone_Int_7QVal_Int_3QVal_Int_1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet17_5QNone_Int_7QVal_Int_3QVal_Int_1_argbuf_r && lizzieLet17_5QNone_Int_7QVal_Int_3QVal_Int_1_bufchan_buf[0]))
        lizzieLet17_5QNone_Int_7QVal_Int_3QVal_Int_1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet17_5QNone_Int_7QVal_Int_3QVal_Int_1_argbuf_r) && (! lizzieLet17_5QNone_Int_7QVal_Int_3QVal_Int_1_bufchan_buf[0])))
        lizzieLet17_5QNone_Int_7QVal_Int_3QVal_Int_1_bufchan_buf <= lizzieLet17_5QNone_Int_7QVal_Int_3QVal_Int_1_bufchan_d;
  
  /* dcon (Ty TupMyDTInt_Int_Int___Int___Int,
      Dcon TupMyDTInt_Int_Int___Int___Int) : [(lizzieLet17_5QNone_Int_7QVal_Int_3QVal_Int_1_argbuf,MyDTInt_Int_Int),
                                              (lizzieLet17_5QNone_Int_7QVal_Int_8QVal_Int_1_argbuf,Int),
                                              (vaew_1_argbuf,Int)] > (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1,TupMyDTInt_Int_Int___Int___Int) */
  assign applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_d = TupMyDTInt_Int_Int___Int___Int_dc((& {lizzieLet17_5QNone_Int_7QVal_Int_3QVal_Int_1_argbuf_d[0],
                                                                                                        lizzieLet17_5QNone_Int_7QVal_Int_8QVal_Int_1_argbuf_d[0],
                                                                                                        vaew_1_argbuf_d[0]}), lizzieLet17_5QNone_Int_7QVal_Int_3QVal_Int_1_argbuf_d, lizzieLet17_5QNone_Int_7QVal_Int_8QVal_Int_1_argbuf_d, vaew_1_argbuf_d);
  assign {lizzieLet17_5QNone_Int_7QVal_Int_3QVal_Int_1_argbuf_r,
          lizzieLet17_5QNone_Int_7QVal_Int_8QVal_Int_1_argbuf_r,
          vaew_1_argbuf_r} = {3 {(applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_r && applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_d[0])}};
  
  /* demux (Ty QTree_Int,
       Ty Pointer_CTf_f_Int) : (lizzieLet17_5QNone_Int_7QVal_Int_4,QTree_Int) (lizzieLet17_5QNone_Int_4QVal_Int,Pointer_CTf_f_Int) > [(lizzieLet17_5QNone_Int_7QVal_Int_4QNone_Int,Pointer_CTf_f_Int),
                                                                                                                                      (lizzieLet17_5QNone_Int_7QVal_Int_4QVal_Int,Pointer_CTf_f_Int),
                                                                                                                                      (lizzieLet17_5QNone_Int_7QVal_Int_4QNode_Int,Pointer_CTf_f_Int),
                                                                                                                                      (lizzieLet17_5QNone_Int_7QVal_Int_4QError_Int,Pointer_CTf_f_Int)] */
  logic [3:0] lizzieLet17_5QNone_Int_4QVal_Int_onehotd;
  always_comb
    if ((lizzieLet17_5QNone_Int_7QVal_Int_4_d[0] && lizzieLet17_5QNone_Int_4QVal_Int_d[0]))
      unique case (lizzieLet17_5QNone_Int_7QVal_Int_4_d[2:1])
        2'd0: lizzieLet17_5QNone_Int_4QVal_Int_onehotd = 4'd1;
        2'd1: lizzieLet17_5QNone_Int_4QVal_Int_onehotd = 4'd2;
        2'd2: lizzieLet17_5QNone_Int_4QVal_Int_onehotd = 4'd4;
        2'd3: lizzieLet17_5QNone_Int_4QVal_Int_onehotd = 4'd8;
        default: lizzieLet17_5QNone_Int_4QVal_Int_onehotd = 4'd0;
      endcase
    else lizzieLet17_5QNone_Int_4QVal_Int_onehotd = 4'd0;
  assign lizzieLet17_5QNone_Int_7QVal_Int_4QNone_Int_d = {lizzieLet17_5QNone_Int_4QVal_Int_d[16:1],
                                                          lizzieLet17_5QNone_Int_4QVal_Int_onehotd[0]};
  assign lizzieLet17_5QNone_Int_7QVal_Int_4QVal_Int_d = {lizzieLet17_5QNone_Int_4QVal_Int_d[16:1],
                                                         lizzieLet17_5QNone_Int_4QVal_Int_onehotd[1]};
  assign lizzieLet17_5QNone_Int_7QVal_Int_4QNode_Int_d = {lizzieLet17_5QNone_Int_4QVal_Int_d[16:1],
                                                          lizzieLet17_5QNone_Int_4QVal_Int_onehotd[2]};
  assign lizzieLet17_5QNone_Int_7QVal_Int_4QError_Int_d = {lizzieLet17_5QNone_Int_4QVal_Int_d[16:1],
                                                           lizzieLet17_5QNone_Int_4QVal_Int_onehotd[3]};
  assign lizzieLet17_5QNone_Int_4QVal_Int_r = (| (lizzieLet17_5QNone_Int_4QVal_Int_onehotd & {lizzieLet17_5QNone_Int_7QVal_Int_4QError_Int_r,
                                                                                              lizzieLet17_5QNone_Int_7QVal_Int_4QNode_Int_r,
                                                                                              lizzieLet17_5QNone_Int_7QVal_Int_4QVal_Int_r,
                                                                                              lizzieLet17_5QNone_Int_7QVal_Int_4QNone_Int_r}));
  assign lizzieLet17_5QNone_Int_7QVal_Int_4_r = lizzieLet17_5QNone_Int_4QVal_Int_r;
  
  /* buf (Ty Pointer_CTf_f_Int) : (lizzieLet17_5QNone_Int_7QVal_Int_4QError_Int,Pointer_CTf_f_Int) > (lizzieLet17_5QNone_Int_7QVal_Int_4QError_Int_1_argbuf,Pointer_CTf_f_Int) */
  Pointer_CTf_f_Int_t lizzieLet17_5QNone_Int_7QVal_Int_4QError_Int_bufchan_d;
  logic lizzieLet17_5QNone_Int_7QVal_Int_4QError_Int_bufchan_r;
  assign lizzieLet17_5QNone_Int_7QVal_Int_4QError_Int_r = ((! lizzieLet17_5QNone_Int_7QVal_Int_4QError_Int_bufchan_d[0]) || lizzieLet17_5QNone_Int_7QVal_Int_4QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNone_Int_7QVal_Int_4QError_Int_bufchan_d <= {16'd0,
                                                                 1'd0};
    else
      if (lizzieLet17_5QNone_Int_7QVal_Int_4QError_Int_r)
        lizzieLet17_5QNone_Int_7QVal_Int_4QError_Int_bufchan_d <= lizzieLet17_5QNone_Int_7QVal_Int_4QError_Int_d;
  Pointer_CTf_f_Int_t lizzieLet17_5QNone_Int_7QVal_Int_4QError_Int_bufchan_buf;
  assign lizzieLet17_5QNone_Int_7QVal_Int_4QError_Int_bufchan_r = (! lizzieLet17_5QNone_Int_7QVal_Int_4QError_Int_bufchan_buf[0]);
  assign lizzieLet17_5QNone_Int_7QVal_Int_4QError_Int_1_argbuf_d = (lizzieLet17_5QNone_Int_7QVal_Int_4QError_Int_bufchan_buf[0] ? lizzieLet17_5QNone_Int_7QVal_Int_4QError_Int_bufchan_buf :
                                                                    lizzieLet17_5QNone_Int_7QVal_Int_4QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNone_Int_7QVal_Int_4QError_Int_bufchan_buf <= {16'd0,
                                                                   1'd0};
    else
      if ((lizzieLet17_5QNone_Int_7QVal_Int_4QError_Int_1_argbuf_r && lizzieLet17_5QNone_Int_7QVal_Int_4QError_Int_bufchan_buf[0]))
        lizzieLet17_5QNone_Int_7QVal_Int_4QError_Int_bufchan_buf <= {16'd0,
                                                                     1'd0};
      else if (((! lizzieLet17_5QNone_Int_7QVal_Int_4QError_Int_1_argbuf_r) && (! lizzieLet17_5QNone_Int_7QVal_Int_4QError_Int_bufchan_buf[0])))
        lizzieLet17_5QNone_Int_7QVal_Int_4QError_Int_bufchan_buf <= lizzieLet17_5QNone_Int_7QVal_Int_4QError_Int_bufchan_d;
  
  /* buf (Ty Pointer_CTf_f_Int) : (lizzieLet17_5QNone_Int_7QVal_Int_4QNode_Int,Pointer_CTf_f_Int) > (lizzieLet17_5QNone_Int_7QVal_Int_4QNode_Int_1_argbuf,Pointer_CTf_f_Int) */
  Pointer_CTf_f_Int_t lizzieLet17_5QNone_Int_7QVal_Int_4QNode_Int_bufchan_d;
  logic lizzieLet17_5QNone_Int_7QVal_Int_4QNode_Int_bufchan_r;
  assign lizzieLet17_5QNone_Int_7QVal_Int_4QNode_Int_r = ((! lizzieLet17_5QNone_Int_7QVal_Int_4QNode_Int_bufchan_d[0]) || lizzieLet17_5QNone_Int_7QVal_Int_4QNode_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNone_Int_7QVal_Int_4QNode_Int_bufchan_d <= {16'd0,
                                                                1'd0};
    else
      if (lizzieLet17_5QNone_Int_7QVal_Int_4QNode_Int_r)
        lizzieLet17_5QNone_Int_7QVal_Int_4QNode_Int_bufchan_d <= lizzieLet17_5QNone_Int_7QVal_Int_4QNode_Int_d;
  Pointer_CTf_f_Int_t lizzieLet17_5QNone_Int_7QVal_Int_4QNode_Int_bufchan_buf;
  assign lizzieLet17_5QNone_Int_7QVal_Int_4QNode_Int_bufchan_r = (! lizzieLet17_5QNone_Int_7QVal_Int_4QNode_Int_bufchan_buf[0]);
  assign lizzieLet17_5QNone_Int_7QVal_Int_4QNode_Int_1_argbuf_d = (lizzieLet17_5QNone_Int_7QVal_Int_4QNode_Int_bufchan_buf[0] ? lizzieLet17_5QNone_Int_7QVal_Int_4QNode_Int_bufchan_buf :
                                                                   lizzieLet17_5QNone_Int_7QVal_Int_4QNode_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNone_Int_7QVal_Int_4QNode_Int_bufchan_buf <= {16'd0,
                                                                  1'd0};
    else
      if ((lizzieLet17_5QNone_Int_7QVal_Int_4QNode_Int_1_argbuf_r && lizzieLet17_5QNone_Int_7QVal_Int_4QNode_Int_bufchan_buf[0]))
        lizzieLet17_5QNone_Int_7QVal_Int_4QNode_Int_bufchan_buf <= {16'd0,
                                                                    1'd0};
      else if (((! lizzieLet17_5QNone_Int_7QVal_Int_4QNode_Int_1_argbuf_r) && (! lizzieLet17_5QNone_Int_7QVal_Int_4QNode_Int_bufchan_buf[0])))
        lizzieLet17_5QNone_Int_7QVal_Int_4QNode_Int_bufchan_buf <= lizzieLet17_5QNone_Int_7QVal_Int_4QNode_Int_bufchan_d;
  
  /* buf (Ty Pointer_CTf_f_Int) : (lizzieLet17_5QNone_Int_7QVal_Int_4QNone_Int,Pointer_CTf_f_Int) > (lizzieLet17_5QNone_Int_7QVal_Int_4QNone_Int_1_argbuf,Pointer_CTf_f_Int) */
  Pointer_CTf_f_Int_t lizzieLet17_5QNone_Int_7QVal_Int_4QNone_Int_bufchan_d;
  logic lizzieLet17_5QNone_Int_7QVal_Int_4QNone_Int_bufchan_r;
  assign lizzieLet17_5QNone_Int_7QVal_Int_4QNone_Int_r = ((! lizzieLet17_5QNone_Int_7QVal_Int_4QNone_Int_bufchan_d[0]) || lizzieLet17_5QNone_Int_7QVal_Int_4QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNone_Int_7QVal_Int_4QNone_Int_bufchan_d <= {16'd0,
                                                                1'd0};
    else
      if (lizzieLet17_5QNone_Int_7QVal_Int_4QNone_Int_r)
        lizzieLet17_5QNone_Int_7QVal_Int_4QNone_Int_bufchan_d <= lizzieLet17_5QNone_Int_7QVal_Int_4QNone_Int_d;
  Pointer_CTf_f_Int_t lizzieLet17_5QNone_Int_7QVal_Int_4QNone_Int_bufchan_buf;
  assign lizzieLet17_5QNone_Int_7QVal_Int_4QNone_Int_bufchan_r = (! lizzieLet17_5QNone_Int_7QVal_Int_4QNone_Int_bufchan_buf[0]);
  assign lizzieLet17_5QNone_Int_7QVal_Int_4QNone_Int_1_argbuf_d = (lizzieLet17_5QNone_Int_7QVal_Int_4QNone_Int_bufchan_buf[0] ? lizzieLet17_5QNone_Int_7QVal_Int_4QNone_Int_bufchan_buf :
                                                                   lizzieLet17_5QNone_Int_7QVal_Int_4QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNone_Int_7QVal_Int_4QNone_Int_bufchan_buf <= {16'd0,
                                                                  1'd0};
    else
      if ((lizzieLet17_5QNone_Int_7QVal_Int_4QNone_Int_1_argbuf_r && lizzieLet17_5QNone_Int_7QVal_Int_4QNone_Int_bufchan_buf[0]))
        lizzieLet17_5QNone_Int_7QVal_Int_4QNone_Int_bufchan_buf <= {16'd0,
                                                                    1'd0};
      else if (((! lizzieLet17_5QNone_Int_7QVal_Int_4QNone_Int_1_argbuf_r) && (! lizzieLet17_5QNone_Int_7QVal_Int_4QNone_Int_bufchan_buf[0])))
        lizzieLet17_5QNone_Int_7QVal_Int_4QNone_Int_bufchan_buf <= lizzieLet17_5QNone_Int_7QVal_Int_4QNone_Int_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Go) : (lizzieLet17_5QNone_Int_7QVal_Int_5,QTree_Int) (lizzieLet17_5QNone_Int_5QVal_Int,Go) > [(lizzieLet17_5QNone_Int_7QVal_Int_5QNone_Int,Go),
                                                                                                        (lizzieLet17_5QNone_Int_7QVal_Int_5QVal_Int,Go),
                                                                                                        (lizzieLet17_5QNone_Int_7QVal_Int_5QNode_Int,Go),
                                                                                                        (lizzieLet17_5QNone_Int_7QVal_Int_5QError_Int,Go)] */
  logic [3:0] lizzieLet17_5QNone_Int_5QVal_Int_onehotd;
  always_comb
    if ((lizzieLet17_5QNone_Int_7QVal_Int_5_d[0] && lizzieLet17_5QNone_Int_5QVal_Int_d[0]))
      unique case (lizzieLet17_5QNone_Int_7QVal_Int_5_d[2:1])
        2'd0: lizzieLet17_5QNone_Int_5QVal_Int_onehotd = 4'd1;
        2'd1: lizzieLet17_5QNone_Int_5QVal_Int_onehotd = 4'd2;
        2'd2: lizzieLet17_5QNone_Int_5QVal_Int_onehotd = 4'd4;
        2'd3: lizzieLet17_5QNone_Int_5QVal_Int_onehotd = 4'd8;
        default: lizzieLet17_5QNone_Int_5QVal_Int_onehotd = 4'd0;
      endcase
    else lizzieLet17_5QNone_Int_5QVal_Int_onehotd = 4'd0;
  assign lizzieLet17_5QNone_Int_7QVal_Int_5QNone_Int_d = lizzieLet17_5QNone_Int_5QVal_Int_onehotd[0];
  assign lizzieLet17_5QNone_Int_7QVal_Int_5QVal_Int_d = lizzieLet17_5QNone_Int_5QVal_Int_onehotd[1];
  assign lizzieLet17_5QNone_Int_7QVal_Int_5QNode_Int_d = lizzieLet17_5QNone_Int_5QVal_Int_onehotd[2];
  assign lizzieLet17_5QNone_Int_7QVal_Int_5QError_Int_d = lizzieLet17_5QNone_Int_5QVal_Int_onehotd[3];
  assign lizzieLet17_5QNone_Int_5QVal_Int_r = (| (lizzieLet17_5QNone_Int_5QVal_Int_onehotd & {lizzieLet17_5QNone_Int_7QVal_Int_5QError_Int_r,
                                                                                              lizzieLet17_5QNone_Int_7QVal_Int_5QNode_Int_r,
                                                                                              lizzieLet17_5QNone_Int_7QVal_Int_5QVal_Int_r,
                                                                                              lizzieLet17_5QNone_Int_7QVal_Int_5QNone_Int_r}));
  assign lizzieLet17_5QNone_Int_7QVal_Int_5_r = lizzieLet17_5QNone_Int_5QVal_Int_r;
  
  /* fork (Ty Go) : (lizzieLet17_5QNone_Int_7QVal_Int_5QError_Int,Go) > [(lizzieLet17_5QNone_Int_7QVal_Int_5QError_Int_1,Go),
                                                                    (lizzieLet17_5QNone_Int_7QVal_Int_5QError_Int_2,Go)] */
  logic [1:0] lizzieLet17_5QNone_Int_7QVal_Int_5QError_Int_emitted;
  logic [1:0] lizzieLet17_5QNone_Int_7QVal_Int_5QError_Int_done;
  assign lizzieLet17_5QNone_Int_7QVal_Int_5QError_Int_1_d = (lizzieLet17_5QNone_Int_7QVal_Int_5QError_Int_d[0] && (! lizzieLet17_5QNone_Int_7QVal_Int_5QError_Int_emitted[0]));
  assign lizzieLet17_5QNone_Int_7QVal_Int_5QError_Int_2_d = (lizzieLet17_5QNone_Int_7QVal_Int_5QError_Int_d[0] && (! lizzieLet17_5QNone_Int_7QVal_Int_5QError_Int_emitted[1]));
  assign lizzieLet17_5QNone_Int_7QVal_Int_5QError_Int_done = (lizzieLet17_5QNone_Int_7QVal_Int_5QError_Int_emitted | ({lizzieLet17_5QNone_Int_7QVal_Int_5QError_Int_2_d[0],
                                                                                                                       lizzieLet17_5QNone_Int_7QVal_Int_5QError_Int_1_d[0]} & {lizzieLet17_5QNone_Int_7QVal_Int_5QError_Int_2_r,
                                                                                                                                                                               lizzieLet17_5QNone_Int_7QVal_Int_5QError_Int_1_r}));
  assign lizzieLet17_5QNone_Int_7QVal_Int_5QError_Int_r = (& lizzieLet17_5QNone_Int_7QVal_Int_5QError_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNone_Int_7QVal_Int_5QError_Int_emitted <= 2'd0;
    else
      lizzieLet17_5QNone_Int_7QVal_Int_5QError_Int_emitted <= (lizzieLet17_5QNone_Int_7QVal_Int_5QError_Int_r ? 2'd0 :
                                                               lizzieLet17_5QNone_Int_7QVal_Int_5QError_Int_done);
  
  /* dcon (Ty QTree_Int,
      Dcon QError_Int) : [(lizzieLet17_5QNone_Int_7QVal_Int_5QError_Int_1,Go)] > (lizzieLet17_5QNone_Int_7QVal_Int_5QError_Int_1QError_Int,QTree_Int) */
  assign lizzieLet17_5QNone_Int_7QVal_Int_5QError_Int_1QError_Int_d = QError_Int_dc((& {lizzieLet17_5QNone_Int_7QVal_Int_5QError_Int_1_d[0]}), lizzieLet17_5QNone_Int_7QVal_Int_5QError_Int_1_d);
  assign {lizzieLet17_5QNone_Int_7QVal_Int_5QError_Int_1_r} = {1 {(lizzieLet17_5QNone_Int_7QVal_Int_5QError_Int_1QError_Int_r && lizzieLet17_5QNone_Int_7QVal_Int_5QError_Int_1QError_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (lizzieLet17_5QNone_Int_7QVal_Int_5QError_Int_1QError_Int,QTree_Int) > (lizzieLet23_1_argbuf,QTree_Int) */
  QTree_Int_t lizzieLet17_5QNone_Int_7QVal_Int_5QError_Int_1QError_Int_bufchan_d;
  logic lizzieLet17_5QNone_Int_7QVal_Int_5QError_Int_1QError_Int_bufchan_r;
  assign lizzieLet17_5QNone_Int_7QVal_Int_5QError_Int_1QError_Int_r = ((! lizzieLet17_5QNone_Int_7QVal_Int_5QError_Int_1QError_Int_bufchan_d[0]) || lizzieLet17_5QNone_Int_7QVal_Int_5QError_Int_1QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNone_Int_7QVal_Int_5QError_Int_1QError_Int_bufchan_d <= {66'd0,
                                                                             1'd0};
    else
      if (lizzieLet17_5QNone_Int_7QVal_Int_5QError_Int_1QError_Int_r)
        lizzieLet17_5QNone_Int_7QVal_Int_5QError_Int_1QError_Int_bufchan_d <= lizzieLet17_5QNone_Int_7QVal_Int_5QError_Int_1QError_Int_d;
  QTree_Int_t lizzieLet17_5QNone_Int_7QVal_Int_5QError_Int_1QError_Int_bufchan_buf;
  assign lizzieLet17_5QNone_Int_7QVal_Int_5QError_Int_1QError_Int_bufchan_r = (! lizzieLet17_5QNone_Int_7QVal_Int_5QError_Int_1QError_Int_bufchan_buf[0]);
  assign lizzieLet23_1_argbuf_d = (lizzieLet17_5QNone_Int_7QVal_Int_5QError_Int_1QError_Int_bufchan_buf[0] ? lizzieLet17_5QNone_Int_7QVal_Int_5QError_Int_1QError_Int_bufchan_buf :
                                   lizzieLet17_5QNone_Int_7QVal_Int_5QError_Int_1QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNone_Int_7QVal_Int_5QError_Int_1QError_Int_bufchan_buf <= {66'd0,
                                                                               1'd0};
    else
      if ((lizzieLet23_1_argbuf_r && lizzieLet17_5QNone_Int_7QVal_Int_5QError_Int_1QError_Int_bufchan_buf[0]))
        lizzieLet17_5QNone_Int_7QVal_Int_5QError_Int_1QError_Int_bufchan_buf <= {66'd0,
                                                                                 1'd0};
      else if (((! lizzieLet23_1_argbuf_r) && (! lizzieLet17_5QNone_Int_7QVal_Int_5QError_Int_1QError_Int_bufchan_buf[0])))
        lizzieLet17_5QNone_Int_7QVal_Int_5QError_Int_1QError_Int_bufchan_buf <= lizzieLet17_5QNone_Int_7QVal_Int_5QError_Int_1QError_Int_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet17_5QNone_Int_7QVal_Int_5QError_Int_2,Go) > (lizzieLet17_5QNone_Int_7QVal_Int_5QError_Int_2_argbuf,Go) */
  Go_t lizzieLet17_5QNone_Int_7QVal_Int_5QError_Int_2_bufchan_d;
  logic lizzieLet17_5QNone_Int_7QVal_Int_5QError_Int_2_bufchan_r;
  assign lizzieLet17_5QNone_Int_7QVal_Int_5QError_Int_2_r = ((! lizzieLet17_5QNone_Int_7QVal_Int_5QError_Int_2_bufchan_d[0]) || lizzieLet17_5QNone_Int_7QVal_Int_5QError_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNone_Int_7QVal_Int_5QError_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet17_5QNone_Int_7QVal_Int_5QError_Int_2_r)
        lizzieLet17_5QNone_Int_7QVal_Int_5QError_Int_2_bufchan_d <= lizzieLet17_5QNone_Int_7QVal_Int_5QError_Int_2_d;
  Go_t lizzieLet17_5QNone_Int_7QVal_Int_5QError_Int_2_bufchan_buf;
  assign lizzieLet17_5QNone_Int_7QVal_Int_5QError_Int_2_bufchan_r = (! lizzieLet17_5QNone_Int_7QVal_Int_5QError_Int_2_bufchan_buf[0]);
  assign lizzieLet17_5QNone_Int_7QVal_Int_5QError_Int_2_argbuf_d = (lizzieLet17_5QNone_Int_7QVal_Int_5QError_Int_2_bufchan_buf[0] ? lizzieLet17_5QNone_Int_7QVal_Int_5QError_Int_2_bufchan_buf :
                                                                    lizzieLet17_5QNone_Int_7QVal_Int_5QError_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNone_Int_7QVal_Int_5QError_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet17_5QNone_Int_7QVal_Int_5QError_Int_2_argbuf_r && lizzieLet17_5QNone_Int_7QVal_Int_5QError_Int_2_bufchan_buf[0]))
        lizzieLet17_5QNone_Int_7QVal_Int_5QError_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet17_5QNone_Int_7QVal_Int_5QError_Int_2_argbuf_r) && (! lizzieLet17_5QNone_Int_7QVal_Int_5QError_Int_2_bufchan_buf[0])))
        lizzieLet17_5QNone_Int_7QVal_Int_5QError_Int_2_bufchan_buf <= lizzieLet17_5QNone_Int_7QVal_Int_5QError_Int_2_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet17_5QNone_Int_7QVal_Int_5QNode_Int,Go) > [(lizzieLet17_5QNone_Int_7QVal_Int_5QNode_Int_1,Go),
                                                                   (lizzieLet17_5QNone_Int_7QVal_Int_5QNode_Int_2,Go)] */
  logic [1:0] lizzieLet17_5QNone_Int_7QVal_Int_5QNode_Int_emitted;
  logic [1:0] lizzieLet17_5QNone_Int_7QVal_Int_5QNode_Int_done;
  assign lizzieLet17_5QNone_Int_7QVal_Int_5QNode_Int_1_d = (lizzieLet17_5QNone_Int_7QVal_Int_5QNode_Int_d[0] && (! lizzieLet17_5QNone_Int_7QVal_Int_5QNode_Int_emitted[0]));
  assign lizzieLet17_5QNone_Int_7QVal_Int_5QNode_Int_2_d = (lizzieLet17_5QNone_Int_7QVal_Int_5QNode_Int_d[0] && (! lizzieLet17_5QNone_Int_7QVal_Int_5QNode_Int_emitted[1]));
  assign lizzieLet17_5QNone_Int_7QVal_Int_5QNode_Int_done = (lizzieLet17_5QNone_Int_7QVal_Int_5QNode_Int_emitted | ({lizzieLet17_5QNone_Int_7QVal_Int_5QNode_Int_2_d[0],
                                                                                                                     lizzieLet17_5QNone_Int_7QVal_Int_5QNode_Int_1_d[0]} & {lizzieLet17_5QNone_Int_7QVal_Int_5QNode_Int_2_r,
                                                                                                                                                                            lizzieLet17_5QNone_Int_7QVal_Int_5QNode_Int_1_r}));
  assign lizzieLet17_5QNone_Int_7QVal_Int_5QNode_Int_r = (& lizzieLet17_5QNone_Int_7QVal_Int_5QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNone_Int_7QVal_Int_5QNode_Int_emitted <= 2'd0;
    else
      lizzieLet17_5QNone_Int_7QVal_Int_5QNode_Int_emitted <= (lizzieLet17_5QNone_Int_7QVal_Int_5QNode_Int_r ? 2'd0 :
                                                              lizzieLet17_5QNone_Int_7QVal_Int_5QNode_Int_done);
  
  /* dcon (Ty QTree_Int,
      Dcon QError_Int) : [(lizzieLet17_5QNone_Int_7QVal_Int_5QNode_Int_1,Go)] > (lizzieLet17_5QNone_Int_7QVal_Int_5QNode_Int_1QError_Int,QTree_Int) */
  assign lizzieLet17_5QNone_Int_7QVal_Int_5QNode_Int_1QError_Int_d = QError_Int_dc((& {lizzieLet17_5QNone_Int_7QVal_Int_5QNode_Int_1_d[0]}), lizzieLet17_5QNone_Int_7QVal_Int_5QNode_Int_1_d);
  assign {lizzieLet17_5QNone_Int_7QVal_Int_5QNode_Int_1_r} = {1 {(lizzieLet17_5QNone_Int_7QVal_Int_5QNode_Int_1QError_Int_r && lizzieLet17_5QNone_Int_7QVal_Int_5QNode_Int_1QError_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (lizzieLet17_5QNone_Int_7QVal_Int_5QNode_Int_1QError_Int,QTree_Int) > (lizzieLet22_1_argbuf,QTree_Int) */
  QTree_Int_t lizzieLet17_5QNone_Int_7QVal_Int_5QNode_Int_1QError_Int_bufchan_d;
  logic lizzieLet17_5QNone_Int_7QVal_Int_5QNode_Int_1QError_Int_bufchan_r;
  assign lizzieLet17_5QNone_Int_7QVal_Int_5QNode_Int_1QError_Int_r = ((! lizzieLet17_5QNone_Int_7QVal_Int_5QNode_Int_1QError_Int_bufchan_d[0]) || lizzieLet17_5QNone_Int_7QVal_Int_5QNode_Int_1QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNone_Int_7QVal_Int_5QNode_Int_1QError_Int_bufchan_d <= {66'd0,
                                                                            1'd0};
    else
      if (lizzieLet17_5QNone_Int_7QVal_Int_5QNode_Int_1QError_Int_r)
        lizzieLet17_5QNone_Int_7QVal_Int_5QNode_Int_1QError_Int_bufchan_d <= lizzieLet17_5QNone_Int_7QVal_Int_5QNode_Int_1QError_Int_d;
  QTree_Int_t lizzieLet17_5QNone_Int_7QVal_Int_5QNode_Int_1QError_Int_bufchan_buf;
  assign lizzieLet17_5QNone_Int_7QVal_Int_5QNode_Int_1QError_Int_bufchan_r = (! lizzieLet17_5QNone_Int_7QVal_Int_5QNode_Int_1QError_Int_bufchan_buf[0]);
  assign lizzieLet22_1_argbuf_d = (lizzieLet17_5QNone_Int_7QVal_Int_5QNode_Int_1QError_Int_bufchan_buf[0] ? lizzieLet17_5QNone_Int_7QVal_Int_5QNode_Int_1QError_Int_bufchan_buf :
                                   lizzieLet17_5QNone_Int_7QVal_Int_5QNode_Int_1QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNone_Int_7QVal_Int_5QNode_Int_1QError_Int_bufchan_buf <= {66'd0,
                                                                              1'd0};
    else
      if ((lizzieLet22_1_argbuf_r && lizzieLet17_5QNone_Int_7QVal_Int_5QNode_Int_1QError_Int_bufchan_buf[0]))
        lizzieLet17_5QNone_Int_7QVal_Int_5QNode_Int_1QError_Int_bufchan_buf <= {66'd0,
                                                                                1'd0};
      else if (((! lizzieLet22_1_argbuf_r) && (! lizzieLet17_5QNone_Int_7QVal_Int_5QNode_Int_1QError_Int_bufchan_buf[0])))
        lizzieLet17_5QNone_Int_7QVal_Int_5QNode_Int_1QError_Int_bufchan_buf <= lizzieLet17_5QNone_Int_7QVal_Int_5QNode_Int_1QError_Int_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet17_5QNone_Int_7QVal_Int_5QNode_Int_2,Go) > (lizzieLet17_5QNone_Int_7QVal_Int_5QNode_Int_2_argbuf,Go) */
  Go_t lizzieLet17_5QNone_Int_7QVal_Int_5QNode_Int_2_bufchan_d;
  logic lizzieLet17_5QNone_Int_7QVal_Int_5QNode_Int_2_bufchan_r;
  assign lizzieLet17_5QNone_Int_7QVal_Int_5QNode_Int_2_r = ((! lizzieLet17_5QNone_Int_7QVal_Int_5QNode_Int_2_bufchan_d[0]) || lizzieLet17_5QNone_Int_7QVal_Int_5QNode_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNone_Int_7QVal_Int_5QNode_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet17_5QNone_Int_7QVal_Int_5QNode_Int_2_r)
        lizzieLet17_5QNone_Int_7QVal_Int_5QNode_Int_2_bufchan_d <= lizzieLet17_5QNone_Int_7QVal_Int_5QNode_Int_2_d;
  Go_t lizzieLet17_5QNone_Int_7QVal_Int_5QNode_Int_2_bufchan_buf;
  assign lizzieLet17_5QNone_Int_7QVal_Int_5QNode_Int_2_bufchan_r = (! lizzieLet17_5QNone_Int_7QVal_Int_5QNode_Int_2_bufchan_buf[0]);
  assign lizzieLet17_5QNone_Int_7QVal_Int_5QNode_Int_2_argbuf_d = (lizzieLet17_5QNone_Int_7QVal_Int_5QNode_Int_2_bufchan_buf[0] ? lizzieLet17_5QNone_Int_7QVal_Int_5QNode_Int_2_bufchan_buf :
                                                                   lizzieLet17_5QNone_Int_7QVal_Int_5QNode_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNone_Int_7QVal_Int_5QNode_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet17_5QNone_Int_7QVal_Int_5QNode_Int_2_argbuf_r && lizzieLet17_5QNone_Int_7QVal_Int_5QNode_Int_2_bufchan_buf[0]))
        lizzieLet17_5QNone_Int_7QVal_Int_5QNode_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet17_5QNone_Int_7QVal_Int_5QNode_Int_2_argbuf_r) && (! lizzieLet17_5QNone_Int_7QVal_Int_5QNode_Int_2_bufchan_buf[0])))
        lizzieLet17_5QNone_Int_7QVal_Int_5QNode_Int_2_bufchan_buf <= lizzieLet17_5QNone_Int_7QVal_Int_5QNode_Int_2_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet17_5QNone_Int_7QVal_Int_5QNone_Int,Go) > (lizzieLet17_5QNone_Int_7QVal_Int_5QNone_Int_1_argbuf,Go) */
  Go_t lizzieLet17_5QNone_Int_7QVal_Int_5QNone_Int_bufchan_d;
  logic lizzieLet17_5QNone_Int_7QVal_Int_5QNone_Int_bufchan_r;
  assign lizzieLet17_5QNone_Int_7QVal_Int_5QNone_Int_r = ((! lizzieLet17_5QNone_Int_7QVal_Int_5QNone_Int_bufchan_d[0]) || lizzieLet17_5QNone_Int_7QVal_Int_5QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNone_Int_7QVal_Int_5QNone_Int_bufchan_d <= 1'd0;
    else
      if (lizzieLet17_5QNone_Int_7QVal_Int_5QNone_Int_r)
        lizzieLet17_5QNone_Int_7QVal_Int_5QNone_Int_bufchan_d <= lizzieLet17_5QNone_Int_7QVal_Int_5QNone_Int_d;
  Go_t lizzieLet17_5QNone_Int_7QVal_Int_5QNone_Int_bufchan_buf;
  assign lizzieLet17_5QNone_Int_7QVal_Int_5QNone_Int_bufchan_r = (! lizzieLet17_5QNone_Int_7QVal_Int_5QNone_Int_bufchan_buf[0]);
  assign lizzieLet17_5QNone_Int_7QVal_Int_5QNone_Int_1_argbuf_d = (lizzieLet17_5QNone_Int_7QVal_Int_5QNone_Int_bufchan_buf[0] ? lizzieLet17_5QNone_Int_7QVal_Int_5QNone_Int_bufchan_buf :
                                                                   lizzieLet17_5QNone_Int_7QVal_Int_5QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNone_Int_7QVal_Int_5QNone_Int_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet17_5QNone_Int_7QVal_Int_5QNone_Int_1_argbuf_r && lizzieLet17_5QNone_Int_7QVal_Int_5QNone_Int_bufchan_buf[0]))
        lizzieLet17_5QNone_Int_7QVal_Int_5QNone_Int_bufchan_buf <= 1'd0;
      else if (((! lizzieLet17_5QNone_Int_7QVal_Int_5QNone_Int_1_argbuf_r) && (! lizzieLet17_5QNone_Int_7QVal_Int_5QNone_Int_bufchan_buf[0])))
        lizzieLet17_5QNone_Int_7QVal_Int_5QNone_Int_bufchan_buf <= lizzieLet17_5QNone_Int_7QVal_Int_5QNone_Int_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet17_5QNone_Int_7QVal_Int_5QVal_Int,Go) > [(lizzieLet17_5QNone_Int_7QVal_Int_5QVal_Int_1,Go),
                                                                  (lizzieLet17_5QNone_Int_7QVal_Int_5QVal_Int_2,Go)] */
  logic [1:0] lizzieLet17_5QNone_Int_7QVal_Int_5QVal_Int_emitted;
  logic [1:0] lizzieLet17_5QNone_Int_7QVal_Int_5QVal_Int_done;
  assign lizzieLet17_5QNone_Int_7QVal_Int_5QVal_Int_1_d = (lizzieLet17_5QNone_Int_7QVal_Int_5QVal_Int_d[0] && (! lizzieLet17_5QNone_Int_7QVal_Int_5QVal_Int_emitted[0]));
  assign lizzieLet17_5QNone_Int_7QVal_Int_5QVal_Int_2_d = (lizzieLet17_5QNone_Int_7QVal_Int_5QVal_Int_d[0] && (! lizzieLet17_5QNone_Int_7QVal_Int_5QVal_Int_emitted[1]));
  assign lizzieLet17_5QNone_Int_7QVal_Int_5QVal_Int_done = (lizzieLet17_5QNone_Int_7QVal_Int_5QVal_Int_emitted | ({lizzieLet17_5QNone_Int_7QVal_Int_5QVal_Int_2_d[0],
                                                                                                                   lizzieLet17_5QNone_Int_7QVal_Int_5QVal_Int_1_d[0]} & {lizzieLet17_5QNone_Int_7QVal_Int_5QVal_Int_2_r,
                                                                                                                                                                         lizzieLet17_5QNone_Int_7QVal_Int_5QVal_Int_1_r}));
  assign lizzieLet17_5QNone_Int_7QVal_Int_5QVal_Int_r = (& lizzieLet17_5QNone_Int_7QVal_Int_5QVal_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNone_Int_7QVal_Int_5QVal_Int_emitted <= 2'd0;
    else
      lizzieLet17_5QNone_Int_7QVal_Int_5QVal_Int_emitted <= (lizzieLet17_5QNone_Int_7QVal_Int_5QVal_Int_r ? 2'd0 :
                                                             lizzieLet17_5QNone_Int_7QVal_Int_5QVal_Int_done);
  
  /* buf (Ty Go) : (lizzieLet17_5QNone_Int_7QVal_Int_5QVal_Int_1,Go) > (lizzieLet17_5QNone_Int_7QVal_Int_5QVal_Int_1_argbuf,Go) */
  Go_t lizzieLet17_5QNone_Int_7QVal_Int_5QVal_Int_1_bufchan_d;
  logic lizzieLet17_5QNone_Int_7QVal_Int_5QVal_Int_1_bufchan_r;
  assign lizzieLet17_5QNone_Int_7QVal_Int_5QVal_Int_1_r = ((! lizzieLet17_5QNone_Int_7QVal_Int_5QVal_Int_1_bufchan_d[0]) || lizzieLet17_5QNone_Int_7QVal_Int_5QVal_Int_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNone_Int_7QVal_Int_5QVal_Int_1_bufchan_d <= 1'd0;
    else
      if (lizzieLet17_5QNone_Int_7QVal_Int_5QVal_Int_1_r)
        lizzieLet17_5QNone_Int_7QVal_Int_5QVal_Int_1_bufchan_d <= lizzieLet17_5QNone_Int_7QVal_Int_5QVal_Int_1_d;
  Go_t lizzieLet17_5QNone_Int_7QVal_Int_5QVal_Int_1_bufchan_buf;
  assign lizzieLet17_5QNone_Int_7QVal_Int_5QVal_Int_1_bufchan_r = (! lizzieLet17_5QNone_Int_7QVal_Int_5QVal_Int_1_bufchan_buf[0]);
  assign lizzieLet17_5QNone_Int_7QVal_Int_5QVal_Int_1_argbuf_d = (lizzieLet17_5QNone_Int_7QVal_Int_5QVal_Int_1_bufchan_buf[0] ? lizzieLet17_5QNone_Int_7QVal_Int_5QVal_Int_1_bufchan_buf :
                                                                  lizzieLet17_5QNone_Int_7QVal_Int_5QVal_Int_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNone_Int_7QVal_Int_5QVal_Int_1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet17_5QNone_Int_7QVal_Int_5QVal_Int_1_argbuf_r && lizzieLet17_5QNone_Int_7QVal_Int_5QVal_Int_1_bufchan_buf[0]))
        lizzieLet17_5QNone_Int_7QVal_Int_5QVal_Int_1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet17_5QNone_Int_7QVal_Int_5QVal_Int_1_argbuf_r) && (! lizzieLet17_5QNone_Int_7QVal_Int_5QVal_Int_1_bufchan_buf[0])))
        lizzieLet17_5QNone_Int_7QVal_Int_5QVal_Int_1_bufchan_buf <= lizzieLet17_5QNone_Int_7QVal_Int_5QVal_Int_1_bufchan_d;
  
  /* dcon (Ty TupGo___MyDTInt_Bool___Int,
      Dcon TupGo___MyDTInt_Bool___Int) : [(lizzieLet17_5QNone_Int_7QVal_Int_5QVal_Int_1_argbuf,Go),
                                          (lizzieLet17_5QNone_Int_7QVal_Int_6QVal_Int_1_argbuf,MyDTInt_Bool),
                                          (es_1_1_1_argbuf,Int)] > (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1,TupGo___MyDTInt_Bool___Int) */
  assign applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_d = TupGo___MyDTInt_Bool___Int_dc((& {lizzieLet17_5QNone_Int_7QVal_Int_5QVal_Int_1_argbuf_d[0],
                                                                                             lizzieLet17_5QNone_Int_7QVal_Int_6QVal_Int_1_argbuf_d[0],
                                                                                             es_1_1_1_argbuf_d[0]}), lizzieLet17_5QNone_Int_7QVal_Int_5QVal_Int_1_argbuf_d, lizzieLet17_5QNone_Int_7QVal_Int_6QVal_Int_1_argbuf_d, es_1_1_1_argbuf_d);
  assign {lizzieLet17_5QNone_Int_7QVal_Int_5QVal_Int_1_argbuf_r,
          lizzieLet17_5QNone_Int_7QVal_Int_6QVal_Int_1_argbuf_r,
          es_1_1_1_argbuf_r} = {3 {(applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_r && applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_d[0])}};
  
  /* demux (Ty QTree_Int,
       Ty MyDTInt_Bool) : (lizzieLet17_5QNone_Int_7QVal_Int_6,QTree_Int) (lizzieLet17_5QNone_Int_6QVal_Int,MyDTInt_Bool) > [(_114,MyDTInt_Bool),
                                                                                                                            (lizzieLet17_5QNone_Int_7QVal_Int_6QVal_Int,MyDTInt_Bool),
                                                                                                                            (_113,MyDTInt_Bool),
                                                                                                                            (_112,MyDTInt_Bool)] */
  logic [3:0] lizzieLet17_5QNone_Int_6QVal_Int_onehotd;
  always_comb
    if ((lizzieLet17_5QNone_Int_7QVal_Int_6_d[0] && lizzieLet17_5QNone_Int_6QVal_Int_d[0]))
      unique case (lizzieLet17_5QNone_Int_7QVal_Int_6_d[2:1])
        2'd0: lizzieLet17_5QNone_Int_6QVal_Int_onehotd = 4'd1;
        2'd1: lizzieLet17_5QNone_Int_6QVal_Int_onehotd = 4'd2;
        2'd2: lizzieLet17_5QNone_Int_6QVal_Int_onehotd = 4'd4;
        2'd3: lizzieLet17_5QNone_Int_6QVal_Int_onehotd = 4'd8;
        default: lizzieLet17_5QNone_Int_6QVal_Int_onehotd = 4'd0;
      endcase
    else lizzieLet17_5QNone_Int_6QVal_Int_onehotd = 4'd0;
  assign _114_d = lizzieLet17_5QNone_Int_6QVal_Int_onehotd[0];
  assign lizzieLet17_5QNone_Int_7QVal_Int_6QVal_Int_d = lizzieLet17_5QNone_Int_6QVal_Int_onehotd[1];
  assign _113_d = lizzieLet17_5QNone_Int_6QVal_Int_onehotd[2];
  assign _112_d = lizzieLet17_5QNone_Int_6QVal_Int_onehotd[3];
  assign lizzieLet17_5QNone_Int_6QVal_Int_r = (| (lizzieLet17_5QNone_Int_6QVal_Int_onehotd & {_112_r,
                                                                                              _113_r,
                                                                                              lizzieLet17_5QNone_Int_7QVal_Int_6QVal_Int_r,
                                                                                              _114_r}));
  assign lizzieLet17_5QNone_Int_7QVal_Int_6_r = lizzieLet17_5QNone_Int_6QVal_Int_r;
  
  /* buf (Ty MyDTInt_Bool) : (lizzieLet17_5QNone_Int_7QVal_Int_6QVal_Int,MyDTInt_Bool) > (lizzieLet17_5QNone_Int_7QVal_Int_6QVal_Int_1_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t lizzieLet17_5QNone_Int_7QVal_Int_6QVal_Int_bufchan_d;
  logic lizzieLet17_5QNone_Int_7QVal_Int_6QVal_Int_bufchan_r;
  assign lizzieLet17_5QNone_Int_7QVal_Int_6QVal_Int_r = ((! lizzieLet17_5QNone_Int_7QVal_Int_6QVal_Int_bufchan_d[0]) || lizzieLet17_5QNone_Int_7QVal_Int_6QVal_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNone_Int_7QVal_Int_6QVal_Int_bufchan_d <= 1'd0;
    else
      if (lizzieLet17_5QNone_Int_7QVal_Int_6QVal_Int_r)
        lizzieLet17_5QNone_Int_7QVal_Int_6QVal_Int_bufchan_d <= lizzieLet17_5QNone_Int_7QVal_Int_6QVal_Int_d;
  MyDTInt_Bool_t lizzieLet17_5QNone_Int_7QVal_Int_6QVal_Int_bufchan_buf;
  assign lizzieLet17_5QNone_Int_7QVal_Int_6QVal_Int_bufchan_r = (! lizzieLet17_5QNone_Int_7QVal_Int_6QVal_Int_bufchan_buf[0]);
  assign lizzieLet17_5QNone_Int_7QVal_Int_6QVal_Int_1_argbuf_d = (lizzieLet17_5QNone_Int_7QVal_Int_6QVal_Int_bufchan_buf[0] ? lizzieLet17_5QNone_Int_7QVal_Int_6QVal_Int_bufchan_buf :
                                                                  lizzieLet17_5QNone_Int_7QVal_Int_6QVal_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNone_Int_7QVal_Int_6QVal_Int_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet17_5QNone_Int_7QVal_Int_6QVal_Int_1_argbuf_r && lizzieLet17_5QNone_Int_7QVal_Int_6QVal_Int_bufchan_buf[0]))
        lizzieLet17_5QNone_Int_7QVal_Int_6QVal_Int_bufchan_buf <= 1'd0;
      else if (((! lizzieLet17_5QNone_Int_7QVal_Int_6QVal_Int_1_argbuf_r) && (! lizzieLet17_5QNone_Int_7QVal_Int_6QVal_Int_bufchan_buf[0])))
        lizzieLet17_5QNone_Int_7QVal_Int_6QVal_Int_bufchan_buf <= lizzieLet17_5QNone_Int_7QVal_Int_6QVal_Int_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_QTree_Int) : (lizzieLet17_5QNone_Int_7QVal_Int_7,QTree_Int) (lizzieLet17_5QNone_Int_8QVal_Int,Pointer_QTree_Int) > [(lizzieLet17_5QNone_Int_7QVal_Int_7QNone_Int,Pointer_QTree_Int),
                                                                                                                                      (_111,Pointer_QTree_Int),
                                                                                                                                      (_110,Pointer_QTree_Int),
                                                                                                                                      (_109,Pointer_QTree_Int)] */
  logic [3:0] lizzieLet17_5QNone_Int_8QVal_Int_onehotd;
  always_comb
    if ((lizzieLet17_5QNone_Int_7QVal_Int_7_d[0] && lizzieLet17_5QNone_Int_8QVal_Int_d[0]))
      unique case (lizzieLet17_5QNone_Int_7QVal_Int_7_d[2:1])
        2'd0: lizzieLet17_5QNone_Int_8QVal_Int_onehotd = 4'd1;
        2'd1: lizzieLet17_5QNone_Int_8QVal_Int_onehotd = 4'd2;
        2'd2: lizzieLet17_5QNone_Int_8QVal_Int_onehotd = 4'd4;
        2'd3: lizzieLet17_5QNone_Int_8QVal_Int_onehotd = 4'd8;
        default: lizzieLet17_5QNone_Int_8QVal_Int_onehotd = 4'd0;
      endcase
    else lizzieLet17_5QNone_Int_8QVal_Int_onehotd = 4'd0;
  assign lizzieLet17_5QNone_Int_7QVal_Int_7QNone_Int_d = {lizzieLet17_5QNone_Int_8QVal_Int_d[16:1],
                                                          lizzieLet17_5QNone_Int_8QVal_Int_onehotd[0]};
  assign _111_d = {lizzieLet17_5QNone_Int_8QVal_Int_d[16:1],
                   lizzieLet17_5QNone_Int_8QVal_Int_onehotd[1]};
  assign _110_d = {lizzieLet17_5QNone_Int_8QVal_Int_d[16:1],
                   lizzieLet17_5QNone_Int_8QVal_Int_onehotd[2]};
  assign _109_d = {lizzieLet17_5QNone_Int_8QVal_Int_d[16:1],
                   lizzieLet17_5QNone_Int_8QVal_Int_onehotd[3]};
  assign lizzieLet17_5QNone_Int_8QVal_Int_r = (| (lizzieLet17_5QNone_Int_8QVal_Int_onehotd & {_109_r,
                                                                                              _110_r,
                                                                                              _111_r,
                                                                                              lizzieLet17_5QNone_Int_7QVal_Int_7QNone_Int_r}));
  assign lizzieLet17_5QNone_Int_7QVal_Int_7_r = lizzieLet17_5QNone_Int_8QVal_Int_r;
  
  /* buf (Ty Pointer_QTree_Int) : (lizzieLet17_5QNone_Int_7QVal_Int_7QNone_Int,Pointer_QTree_Int) > (lizzieLet17_5QNone_Int_7QVal_Int_7QNone_Int_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t lizzieLet17_5QNone_Int_7QVal_Int_7QNone_Int_bufchan_d;
  logic lizzieLet17_5QNone_Int_7QVal_Int_7QNone_Int_bufchan_r;
  assign lizzieLet17_5QNone_Int_7QVal_Int_7QNone_Int_r = ((! lizzieLet17_5QNone_Int_7QVal_Int_7QNone_Int_bufchan_d[0]) || lizzieLet17_5QNone_Int_7QVal_Int_7QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNone_Int_7QVal_Int_7QNone_Int_bufchan_d <= {16'd0,
                                                                1'd0};
    else
      if (lizzieLet17_5QNone_Int_7QVal_Int_7QNone_Int_r)
        lizzieLet17_5QNone_Int_7QVal_Int_7QNone_Int_bufchan_d <= lizzieLet17_5QNone_Int_7QVal_Int_7QNone_Int_d;
  Pointer_QTree_Int_t lizzieLet17_5QNone_Int_7QVal_Int_7QNone_Int_bufchan_buf;
  assign lizzieLet17_5QNone_Int_7QVal_Int_7QNone_Int_bufchan_r = (! lizzieLet17_5QNone_Int_7QVal_Int_7QNone_Int_bufchan_buf[0]);
  assign lizzieLet17_5QNone_Int_7QVal_Int_7QNone_Int_1_argbuf_d = (lizzieLet17_5QNone_Int_7QVal_Int_7QNone_Int_bufchan_buf[0] ? lizzieLet17_5QNone_Int_7QVal_Int_7QNone_Int_bufchan_buf :
                                                                   lizzieLet17_5QNone_Int_7QVal_Int_7QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNone_Int_7QVal_Int_7QNone_Int_bufchan_buf <= {16'd0,
                                                                  1'd0};
    else
      if ((lizzieLet17_5QNone_Int_7QVal_Int_7QNone_Int_1_argbuf_r && lizzieLet17_5QNone_Int_7QVal_Int_7QNone_Int_bufchan_buf[0]))
        lizzieLet17_5QNone_Int_7QVal_Int_7QNone_Int_bufchan_buf <= {16'd0,
                                                                    1'd0};
      else if (((! lizzieLet17_5QNone_Int_7QVal_Int_7QNone_Int_1_argbuf_r) && (! lizzieLet17_5QNone_Int_7QVal_Int_7QNone_Int_bufchan_buf[0])))
        lizzieLet17_5QNone_Int_7QVal_Int_7QNone_Int_bufchan_buf <= lizzieLet17_5QNone_Int_7QVal_Int_7QNone_Int_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Int) : (lizzieLet17_5QNone_Int_7QVal_Int_8,QTree_Int) (v1aev_destruct,Int) > [(_108,Int),
                                                                                        (lizzieLet17_5QNone_Int_7QVal_Int_8QVal_Int,Int),
                                                                                        (_107,Int),
                                                                                        (_106,Int)] */
  logic [3:0] v1aev_destruct_onehotd;
  always_comb
    if ((lizzieLet17_5QNone_Int_7QVal_Int_8_d[0] && v1aev_destruct_d[0]))
      unique case (lizzieLet17_5QNone_Int_7QVal_Int_8_d[2:1])
        2'd0: v1aev_destruct_onehotd = 4'd1;
        2'd1: v1aev_destruct_onehotd = 4'd2;
        2'd2: v1aev_destruct_onehotd = 4'd4;
        2'd3: v1aev_destruct_onehotd = 4'd8;
        default: v1aev_destruct_onehotd = 4'd0;
      endcase
    else v1aev_destruct_onehotd = 4'd0;
  assign _108_d = {v1aev_destruct_d[32:1],
                   v1aev_destruct_onehotd[0]};
  assign lizzieLet17_5QNone_Int_7QVal_Int_8QVal_Int_d = {v1aev_destruct_d[32:1],
                                                         v1aev_destruct_onehotd[1]};
  assign _107_d = {v1aev_destruct_d[32:1],
                   v1aev_destruct_onehotd[2]};
  assign _106_d = {v1aev_destruct_d[32:1],
                   v1aev_destruct_onehotd[3]};
  assign v1aev_destruct_r = (| (v1aev_destruct_onehotd & {_106_r,
                                                          _107_r,
                                                          lizzieLet17_5QNone_Int_7QVal_Int_8QVal_Int_r,
                                                          _108_r}));
  assign lizzieLet17_5QNone_Int_7QVal_Int_8_r = v1aev_destruct_r;
  
  /* fork (Ty Int) : (lizzieLet17_5QNone_Int_7QVal_Int_8QVal_Int,Int) > [(lizzieLet17_5QNone_Int_7QVal_Int_8QVal_Int_1,Int),
                                                                    (lizzieLet17_5QNone_Int_7QVal_Int_8QVal_Int_2,Int)] */
  logic [1:0] lizzieLet17_5QNone_Int_7QVal_Int_8QVal_Int_emitted;
  logic [1:0] lizzieLet17_5QNone_Int_7QVal_Int_8QVal_Int_done;
  assign lizzieLet17_5QNone_Int_7QVal_Int_8QVal_Int_1_d = {lizzieLet17_5QNone_Int_7QVal_Int_8QVal_Int_d[32:1],
                                                           (lizzieLet17_5QNone_Int_7QVal_Int_8QVal_Int_d[0] && (! lizzieLet17_5QNone_Int_7QVal_Int_8QVal_Int_emitted[0]))};
  assign lizzieLet17_5QNone_Int_7QVal_Int_8QVal_Int_2_d = {lizzieLet17_5QNone_Int_7QVal_Int_8QVal_Int_d[32:1],
                                                           (lizzieLet17_5QNone_Int_7QVal_Int_8QVal_Int_d[0] && (! lizzieLet17_5QNone_Int_7QVal_Int_8QVal_Int_emitted[1]))};
  assign lizzieLet17_5QNone_Int_7QVal_Int_8QVal_Int_done = (lizzieLet17_5QNone_Int_7QVal_Int_8QVal_Int_emitted | ({lizzieLet17_5QNone_Int_7QVal_Int_8QVal_Int_2_d[0],
                                                                                                                   lizzieLet17_5QNone_Int_7QVal_Int_8QVal_Int_1_d[0]} & {lizzieLet17_5QNone_Int_7QVal_Int_8QVal_Int_2_r,
                                                                                                                                                                         lizzieLet17_5QNone_Int_7QVal_Int_8QVal_Int_1_r}));
  assign lizzieLet17_5QNone_Int_7QVal_Int_8QVal_Int_r = (& lizzieLet17_5QNone_Int_7QVal_Int_8QVal_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNone_Int_7QVal_Int_8QVal_Int_emitted <= 2'd0;
    else
      lizzieLet17_5QNone_Int_7QVal_Int_8QVal_Int_emitted <= (lizzieLet17_5QNone_Int_7QVal_Int_8QVal_Int_r ? 2'd0 :
                                                             lizzieLet17_5QNone_Int_7QVal_Int_8QVal_Int_done);
  
  /* buf (Ty Int) : (lizzieLet17_5QNone_Int_7QVal_Int_8QVal_Int_1,Int) > (lizzieLet17_5QNone_Int_7QVal_Int_8QVal_Int_1_argbuf,Int) */
  Int_t lizzieLet17_5QNone_Int_7QVal_Int_8QVal_Int_1_bufchan_d;
  logic lizzieLet17_5QNone_Int_7QVal_Int_8QVal_Int_1_bufchan_r;
  assign lizzieLet17_5QNone_Int_7QVal_Int_8QVal_Int_1_r = ((! lizzieLet17_5QNone_Int_7QVal_Int_8QVal_Int_1_bufchan_d[0]) || lizzieLet17_5QNone_Int_7QVal_Int_8QVal_Int_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNone_Int_7QVal_Int_8QVal_Int_1_bufchan_d <= {32'd0,
                                                                 1'd0};
    else
      if (lizzieLet17_5QNone_Int_7QVal_Int_8QVal_Int_1_r)
        lizzieLet17_5QNone_Int_7QVal_Int_8QVal_Int_1_bufchan_d <= lizzieLet17_5QNone_Int_7QVal_Int_8QVal_Int_1_d;
  Int_t lizzieLet17_5QNone_Int_7QVal_Int_8QVal_Int_1_bufchan_buf;
  assign lizzieLet17_5QNone_Int_7QVal_Int_8QVal_Int_1_bufchan_r = (! lizzieLet17_5QNone_Int_7QVal_Int_8QVal_Int_1_bufchan_buf[0]);
  assign lizzieLet17_5QNone_Int_7QVal_Int_8QVal_Int_1_argbuf_d = (lizzieLet17_5QNone_Int_7QVal_Int_8QVal_Int_1_bufchan_buf[0] ? lizzieLet17_5QNone_Int_7QVal_Int_8QVal_Int_1_bufchan_buf :
                                                                  lizzieLet17_5QNone_Int_7QVal_Int_8QVal_Int_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNone_Int_7QVal_Int_8QVal_Int_1_bufchan_buf <= {32'd0,
                                                                   1'd0};
    else
      if ((lizzieLet17_5QNone_Int_7QVal_Int_8QVal_Int_1_argbuf_r && lizzieLet17_5QNone_Int_7QVal_Int_8QVal_Int_1_bufchan_buf[0]))
        lizzieLet17_5QNone_Int_7QVal_Int_8QVal_Int_1_bufchan_buf <= {32'd0,
                                                                     1'd0};
      else if (((! lizzieLet17_5QNone_Int_7QVal_Int_8QVal_Int_1_argbuf_r) && (! lizzieLet17_5QNone_Int_7QVal_Int_8QVal_Int_1_bufchan_buf[0])))
        lizzieLet17_5QNone_Int_7QVal_Int_8QVal_Int_1_bufchan_buf <= lizzieLet17_5QNone_Int_7QVal_Int_8QVal_Int_1_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_QTree_Int) : (lizzieLet17_5QNone_Int_8,QTree_Int) (lizzieLet17_8QNone_Int,Pointer_QTree_Int) > [(_105,Pointer_QTree_Int),
                                                                                                                  (lizzieLet17_5QNone_Int_8QVal_Int,Pointer_QTree_Int),
                                                                                                                  (lizzieLet17_5QNone_Int_8QNode_Int,Pointer_QTree_Int),
                                                                                                                  (_104,Pointer_QTree_Int)] */
  logic [3:0] lizzieLet17_8QNone_Int_onehotd;
  always_comb
    if ((lizzieLet17_5QNone_Int_8_d[0] && lizzieLet17_8QNone_Int_d[0]))
      unique case (lizzieLet17_5QNone_Int_8_d[2:1])
        2'd0: lizzieLet17_8QNone_Int_onehotd = 4'd1;
        2'd1: lizzieLet17_8QNone_Int_onehotd = 4'd2;
        2'd2: lizzieLet17_8QNone_Int_onehotd = 4'd4;
        2'd3: lizzieLet17_8QNone_Int_onehotd = 4'd8;
        default: lizzieLet17_8QNone_Int_onehotd = 4'd0;
      endcase
    else lizzieLet17_8QNone_Int_onehotd = 4'd0;
  assign _105_d = {lizzieLet17_8QNone_Int_d[16:1],
                   lizzieLet17_8QNone_Int_onehotd[0]};
  assign lizzieLet17_5QNone_Int_8QVal_Int_d = {lizzieLet17_8QNone_Int_d[16:1],
                                               lizzieLet17_8QNone_Int_onehotd[1]};
  assign lizzieLet17_5QNone_Int_8QNode_Int_d = {lizzieLet17_8QNone_Int_d[16:1],
                                                lizzieLet17_8QNone_Int_onehotd[2]};
  assign _104_d = {lizzieLet17_8QNone_Int_d[16:1],
                   lizzieLet17_8QNone_Int_onehotd[3]};
  assign lizzieLet17_8QNone_Int_r = (| (lizzieLet17_8QNone_Int_onehotd & {_104_r,
                                                                          lizzieLet17_5QNone_Int_8QNode_Int_r,
                                                                          lizzieLet17_5QNone_Int_8QVal_Int_r,
                                                                          _105_r}));
  assign lizzieLet17_5QNone_Int_8_r = lizzieLet17_8QNone_Int_r;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_QTree_Int) : (lizzieLet17_5QNone_Int_9,QTree_Int) (lizzieLet17_9QNone_Int,Pointer_QTree_Int) > [(lizzieLet17_5QNone_Int_9QNone_Int,Pointer_QTree_Int),
                                                                                                                  (_103,Pointer_QTree_Int),
                                                                                                                  (_102,Pointer_QTree_Int),
                                                                                                                  (_101,Pointer_QTree_Int)] */
  logic [3:0] lizzieLet17_9QNone_Int_onehotd;
  always_comb
    if ((lizzieLet17_5QNone_Int_9_d[0] && lizzieLet17_9QNone_Int_d[0]))
      unique case (lizzieLet17_5QNone_Int_9_d[2:1])
        2'd0: lizzieLet17_9QNone_Int_onehotd = 4'd1;
        2'd1: lizzieLet17_9QNone_Int_onehotd = 4'd2;
        2'd2: lizzieLet17_9QNone_Int_onehotd = 4'd4;
        2'd3: lizzieLet17_9QNone_Int_onehotd = 4'd8;
        default: lizzieLet17_9QNone_Int_onehotd = 4'd0;
      endcase
    else lizzieLet17_9QNone_Int_onehotd = 4'd0;
  assign lizzieLet17_5QNone_Int_9QNone_Int_d = {lizzieLet17_9QNone_Int_d[16:1],
                                                lizzieLet17_9QNone_Int_onehotd[0]};
  assign _103_d = {lizzieLet17_9QNone_Int_d[16:1],
                   lizzieLet17_9QNone_Int_onehotd[1]};
  assign _102_d = {lizzieLet17_9QNone_Int_d[16:1],
                   lizzieLet17_9QNone_Int_onehotd[2]};
  assign _101_d = {lizzieLet17_9QNone_Int_d[16:1],
                   lizzieLet17_9QNone_Int_onehotd[3]};
  assign lizzieLet17_9QNone_Int_r = (| (lizzieLet17_9QNone_Int_onehotd & {_101_r,
                                                                          _102_r,
                                                                          _103_r,
                                                                          lizzieLet17_5QNone_Int_9QNone_Int_r}));
  assign lizzieLet17_5QNone_Int_9_r = lizzieLet17_9QNone_Int_r;
  
  /* buf (Ty Pointer_QTree_Int) : (lizzieLet17_5QNone_Int_9QNone_Int,Pointer_QTree_Int) > (lizzieLet17_5QNone_Int_9QNone_Int_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t lizzieLet17_5QNone_Int_9QNone_Int_bufchan_d;
  logic lizzieLet17_5QNone_Int_9QNone_Int_bufchan_r;
  assign lizzieLet17_5QNone_Int_9QNone_Int_r = ((! lizzieLet17_5QNone_Int_9QNone_Int_bufchan_d[0]) || lizzieLet17_5QNone_Int_9QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNone_Int_9QNone_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet17_5QNone_Int_9QNone_Int_r)
        lizzieLet17_5QNone_Int_9QNone_Int_bufchan_d <= lizzieLet17_5QNone_Int_9QNone_Int_d;
  Pointer_QTree_Int_t lizzieLet17_5QNone_Int_9QNone_Int_bufchan_buf;
  assign lizzieLet17_5QNone_Int_9QNone_Int_bufchan_r = (! lizzieLet17_5QNone_Int_9QNone_Int_bufchan_buf[0]);
  assign lizzieLet17_5QNone_Int_9QNone_Int_1_argbuf_d = (lizzieLet17_5QNone_Int_9QNone_Int_bufchan_buf[0] ? lizzieLet17_5QNone_Int_9QNone_Int_bufchan_buf :
                                                         lizzieLet17_5QNone_Int_9QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QNone_Int_9QNone_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet17_5QNone_Int_9QNone_Int_1_argbuf_r && lizzieLet17_5QNone_Int_9QNone_Int_bufchan_buf[0]))
        lizzieLet17_5QNone_Int_9QNone_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet17_5QNone_Int_9QNone_Int_1_argbuf_r) && (! lizzieLet17_5QNone_Int_9QNone_Int_bufchan_buf[0])))
        lizzieLet17_5QNone_Int_9QNone_Int_bufchan_buf <= lizzieLet17_5QNone_Int_9QNone_Int_bufchan_d;
  
  /* fork (Ty QTree_Int) : (lizzieLet17_5QVal_Int,QTree_Int) > [(lizzieLet17_5QVal_Int_1,QTree_Int),
                                                           (lizzieLet17_5QVal_Int_2,QTree_Int),
                                                           (lizzieLet17_5QVal_Int_3,QTree_Int),
                                                           (lizzieLet17_5QVal_Int_4,QTree_Int),
                                                           (lizzieLet17_5QVal_Int_5,QTree_Int),
                                                           (lizzieLet17_5QVal_Int_6,QTree_Int),
                                                           (lizzieLet17_5QVal_Int_7,QTree_Int),
                                                           (lizzieLet17_5QVal_Int_8,QTree_Int),
                                                           (lizzieLet17_5QVal_Int_9,QTree_Int),
                                                           (lizzieLet17_5QVal_Int_10,QTree_Int)] */
  logic [9:0] lizzieLet17_5QVal_Int_emitted;
  logic [9:0] lizzieLet17_5QVal_Int_done;
  assign lizzieLet17_5QVal_Int_1_d = {lizzieLet17_5QVal_Int_d[66:1],
                                      (lizzieLet17_5QVal_Int_d[0] && (! lizzieLet17_5QVal_Int_emitted[0]))};
  assign lizzieLet17_5QVal_Int_2_d = {lizzieLet17_5QVal_Int_d[66:1],
                                      (lizzieLet17_5QVal_Int_d[0] && (! lizzieLet17_5QVal_Int_emitted[1]))};
  assign lizzieLet17_5QVal_Int_3_d = {lizzieLet17_5QVal_Int_d[66:1],
                                      (lizzieLet17_5QVal_Int_d[0] && (! lizzieLet17_5QVal_Int_emitted[2]))};
  assign lizzieLet17_5QVal_Int_4_d = {lizzieLet17_5QVal_Int_d[66:1],
                                      (lizzieLet17_5QVal_Int_d[0] && (! lizzieLet17_5QVal_Int_emitted[3]))};
  assign lizzieLet17_5QVal_Int_5_d = {lizzieLet17_5QVal_Int_d[66:1],
                                      (lizzieLet17_5QVal_Int_d[0] && (! lizzieLet17_5QVal_Int_emitted[4]))};
  assign lizzieLet17_5QVal_Int_6_d = {lizzieLet17_5QVal_Int_d[66:1],
                                      (lizzieLet17_5QVal_Int_d[0] && (! lizzieLet17_5QVal_Int_emitted[5]))};
  assign lizzieLet17_5QVal_Int_7_d = {lizzieLet17_5QVal_Int_d[66:1],
                                      (lizzieLet17_5QVal_Int_d[0] && (! lizzieLet17_5QVal_Int_emitted[6]))};
  assign lizzieLet17_5QVal_Int_8_d = {lizzieLet17_5QVal_Int_d[66:1],
                                      (lizzieLet17_5QVal_Int_d[0] && (! lizzieLet17_5QVal_Int_emitted[7]))};
  assign lizzieLet17_5QVal_Int_9_d = {lizzieLet17_5QVal_Int_d[66:1],
                                      (lizzieLet17_5QVal_Int_d[0] && (! lizzieLet17_5QVal_Int_emitted[8]))};
  assign lizzieLet17_5QVal_Int_10_d = {lizzieLet17_5QVal_Int_d[66:1],
                                       (lizzieLet17_5QVal_Int_d[0] && (! lizzieLet17_5QVal_Int_emitted[9]))};
  assign lizzieLet17_5QVal_Int_done = (lizzieLet17_5QVal_Int_emitted | ({lizzieLet17_5QVal_Int_10_d[0],
                                                                         lizzieLet17_5QVal_Int_9_d[0],
                                                                         lizzieLet17_5QVal_Int_8_d[0],
                                                                         lizzieLet17_5QVal_Int_7_d[0],
                                                                         lizzieLet17_5QVal_Int_6_d[0],
                                                                         lizzieLet17_5QVal_Int_5_d[0],
                                                                         lizzieLet17_5QVal_Int_4_d[0],
                                                                         lizzieLet17_5QVal_Int_3_d[0],
                                                                         lizzieLet17_5QVal_Int_2_d[0],
                                                                         lizzieLet17_5QVal_Int_1_d[0]} & {lizzieLet17_5QVal_Int_10_r,
                                                                                                          lizzieLet17_5QVal_Int_9_r,
                                                                                                          lizzieLet17_5QVal_Int_8_r,
                                                                                                          lizzieLet17_5QVal_Int_7_r,
                                                                                                          lizzieLet17_5QVal_Int_6_r,
                                                                                                          lizzieLet17_5QVal_Int_5_r,
                                                                                                          lizzieLet17_5QVal_Int_4_r,
                                                                                                          lizzieLet17_5QVal_Int_3_r,
                                                                                                          lizzieLet17_5QVal_Int_2_r,
                                                                                                          lizzieLet17_5QVal_Int_1_r}));
  assign lizzieLet17_5QVal_Int_r = (& lizzieLet17_5QVal_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet17_5QVal_Int_emitted <= 10'd0;
    else
      lizzieLet17_5QVal_Int_emitted <= (lizzieLet17_5QVal_Int_r ? 10'd0 :
                                        lizzieLet17_5QVal_Int_done);
  
  /* demux (Ty QTree_Int,
       Ty Int) : (lizzieLet17_5QVal_Int_10,QTree_Int) (v1aeK_destruct,Int) > [(lizzieLet17_5QVal_Int_10QNone_Int,Int),
                                                                              (lizzieLet17_5QVal_Int_10QVal_Int,Int),
                                                                              (_100,Int),
                                                                              (_99,Int)] */
  logic [3:0] v1aeK_destruct_onehotd;
  always_comb
    if ((lizzieLet17_5QVal_Int_10_d[0] && v1aeK_destruct_d[0]))
      unique case (lizzieLet17_5QVal_Int_10_d[2:1])
        2'd0: v1aeK_destruct_onehotd = 4'd1;
        2'd1: v1aeK_destruct_onehotd = 4'd2;
        2'd2: v1aeK_destruct_onehotd = 4'd4;
        2'd3: v1aeK_destruct_onehotd = 4'd8;
        default: v1aeK_destruct_onehotd = 4'd0;
      endcase
    else v1aeK_destruct_onehotd = 4'd0;
  assign lizzieLet17_5QVal_Int_10QNone_Int_d = {v1aeK_destruct_d[32:1],
                                                v1aeK_destruct_onehotd[0]};
  assign lizzieLet17_5QVal_Int_10QVal_Int_d = {v1aeK_destruct_d[32:1],
                                               v1aeK_destruct_onehotd[1]};
  assign _100_d = {v1aeK_destruct_d[32:1],
                   v1aeK_destruct_onehotd[2]};
  assign _99_d = {v1aeK_destruct_d[32:1], v1aeK_destruct_onehotd[3]};
  assign v1aeK_destruct_r = (| (v1aeK_destruct_onehotd & {_99_r,
                                                          _100_r,
                                                          lizzieLet17_5QVal_Int_10QVal_Int_r,
                                                          lizzieLet17_5QVal_Int_10QNone_Int_r}));
  assign lizzieLet17_5QVal_Int_10_r = v1aeK_destruct_r;
  
  /* fork (Ty Int) : (lizzieLet17_5QVal_Int_10QVal_Int,Int) > [(lizzieLet17_5QVal_Int_10QVal_Int_1,Int),
                                                          (lizzieLet17_5QVal_Int_10QVal_Int_2,Int)] */
  logic [1:0] lizzieLet17_5QVal_Int_10QVal_Int_emitted;
  logic [1:0] lizzieLet17_5QVal_Int_10QVal_Int_done;
  assign lizzieLet17_5QVal_Int_10QVal_Int_1_d = {lizzieLet17_5QVal_Int_10QVal_Int_d[32:1],
                                                 (lizzieLet17_5QVal_Int_10QVal_Int_d[0] && (! lizzieLet17_5QVal_Int_10QVal_Int_emitted[0]))};
  assign lizzieLet17_5QVal_Int_10QVal_Int_2_d = {lizzieLet17_5QVal_Int_10QVal_Int_d[32:1],
                                                 (lizzieLet17_5QVal_Int_10QVal_Int_d[0] && (! lizzieLet17_5QVal_Int_10QVal_Int_emitted[1]))};
  assign lizzieLet17_5QVal_Int_10QVal_Int_done = (lizzieLet17_5QVal_Int_10QVal_Int_emitted | ({lizzieLet17_5QVal_Int_10QVal_Int_2_d[0],
                                                                                               lizzieLet17_5QVal_Int_10QVal_Int_1_d[0]} & {lizzieLet17_5QVal_Int_10QVal_Int_2_r,
                                                                                                                                           lizzieLet17_5QVal_Int_10QVal_Int_1_r}));
  assign lizzieLet17_5QVal_Int_10QVal_Int_r = (& lizzieLet17_5QVal_Int_10QVal_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QVal_Int_10QVal_Int_emitted <= 2'd0;
    else
      lizzieLet17_5QVal_Int_10QVal_Int_emitted <= (lizzieLet17_5QVal_Int_10QVal_Int_r ? 2'd0 :
                                                   lizzieLet17_5QVal_Int_10QVal_Int_done);
  
  /* buf (Ty Int) : (lizzieLet17_5QVal_Int_10QVal_Int_1,Int) > (lizzieLet17_5QVal_Int_10QVal_Int_1_argbuf,Int) */
  Int_t lizzieLet17_5QVal_Int_10QVal_Int_1_bufchan_d;
  logic lizzieLet17_5QVal_Int_10QVal_Int_1_bufchan_r;
  assign lizzieLet17_5QVal_Int_10QVal_Int_1_r = ((! lizzieLet17_5QVal_Int_10QVal_Int_1_bufchan_d[0]) || lizzieLet17_5QVal_Int_10QVal_Int_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QVal_Int_10QVal_Int_1_bufchan_d <= {32'd0, 1'd0};
    else
      if (lizzieLet17_5QVal_Int_10QVal_Int_1_r)
        lizzieLet17_5QVal_Int_10QVal_Int_1_bufchan_d <= lizzieLet17_5QVal_Int_10QVal_Int_1_d;
  Int_t lizzieLet17_5QVal_Int_10QVal_Int_1_bufchan_buf;
  assign lizzieLet17_5QVal_Int_10QVal_Int_1_bufchan_r = (! lizzieLet17_5QVal_Int_10QVal_Int_1_bufchan_buf[0]);
  assign lizzieLet17_5QVal_Int_10QVal_Int_1_argbuf_d = (lizzieLet17_5QVal_Int_10QVal_Int_1_bufchan_buf[0] ? lizzieLet17_5QVal_Int_10QVal_Int_1_bufchan_buf :
                                                        lizzieLet17_5QVal_Int_10QVal_Int_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QVal_Int_10QVal_Int_1_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((lizzieLet17_5QVal_Int_10QVal_Int_1_argbuf_r && lizzieLet17_5QVal_Int_10QVal_Int_1_bufchan_buf[0]))
        lizzieLet17_5QVal_Int_10QVal_Int_1_bufchan_buf <= {32'd0, 1'd0};
      else if (((! lizzieLet17_5QVal_Int_10QVal_Int_1_argbuf_r) && (! lizzieLet17_5QVal_Int_10QVal_Int_1_bufchan_buf[0])))
        lizzieLet17_5QVal_Int_10QVal_Int_1_bufchan_buf <= lizzieLet17_5QVal_Int_10QVal_Int_1_bufchan_d;
  
  /* destruct (Ty QTree_Int,
          Dcon QVal_Int) : (lizzieLet17_5QVal_Int_1QVal_Int,QTree_Int) > [(vaeQ_destruct,Int)] */
  assign vaeQ_destruct_d = {lizzieLet17_5QVal_Int_1QVal_Int_d[34:3],
                            lizzieLet17_5QVal_Int_1QVal_Int_d[0]};
  assign lizzieLet17_5QVal_Int_1QVal_Int_r = vaeQ_destruct_r;
  
  /* demux (Ty QTree_Int,
       Ty QTree_Int) : (lizzieLet17_5QVal_Int_2,QTree_Int) (lizzieLet17_5QVal_Int_1,QTree_Int) > [(_98,QTree_Int),
                                                                                                  (lizzieLet17_5QVal_Int_1QVal_Int,QTree_Int),
                                                                                                  (_97,QTree_Int),
                                                                                                  (_96,QTree_Int)] */
  logic [3:0] lizzieLet17_5QVal_Int_1_onehotd;
  always_comb
    if ((lizzieLet17_5QVal_Int_2_d[0] && lizzieLet17_5QVal_Int_1_d[0]))
      unique case (lizzieLet17_5QVal_Int_2_d[2:1])
        2'd0: lizzieLet17_5QVal_Int_1_onehotd = 4'd1;
        2'd1: lizzieLet17_5QVal_Int_1_onehotd = 4'd2;
        2'd2: lizzieLet17_5QVal_Int_1_onehotd = 4'd4;
        2'd3: lizzieLet17_5QVal_Int_1_onehotd = 4'd8;
        default: lizzieLet17_5QVal_Int_1_onehotd = 4'd0;
      endcase
    else lizzieLet17_5QVal_Int_1_onehotd = 4'd0;
  assign _98_d = {lizzieLet17_5QVal_Int_1_d[66:1],
                  lizzieLet17_5QVal_Int_1_onehotd[0]};
  assign lizzieLet17_5QVal_Int_1QVal_Int_d = {lizzieLet17_5QVal_Int_1_d[66:1],
                                              lizzieLet17_5QVal_Int_1_onehotd[1]};
  assign _97_d = {lizzieLet17_5QVal_Int_1_d[66:1],
                  lizzieLet17_5QVal_Int_1_onehotd[2]};
  assign _96_d = {lizzieLet17_5QVal_Int_1_d[66:1],
                  lizzieLet17_5QVal_Int_1_onehotd[3]};
  assign lizzieLet17_5QVal_Int_1_r = (| (lizzieLet17_5QVal_Int_1_onehotd & {_96_r,
                                                                            _97_r,
                                                                            lizzieLet17_5QVal_Int_1QVal_Int_r,
                                                                            _98_r}));
  assign lizzieLet17_5QVal_Int_2_r = lizzieLet17_5QVal_Int_1_r;
  
  /* demux (Ty QTree_Int,
       Ty MyDTInt_Int_Int) : (lizzieLet17_5QVal_Int_3,QTree_Int) (lizzieLet17_10QVal_Int,MyDTInt_Int_Int) > [(lizzieLet17_5QVal_Int_3QNone_Int,MyDTInt_Int_Int),
                                                                                                             (lizzieLet17_5QVal_Int_3QVal_Int,MyDTInt_Int_Int),
                                                                                                             (_95,MyDTInt_Int_Int),
                                                                                                             (_94,MyDTInt_Int_Int)] */
  logic [3:0] lizzieLet17_10QVal_Int_onehotd;
  always_comb
    if ((lizzieLet17_5QVal_Int_3_d[0] && lizzieLet17_10QVal_Int_d[0]))
      unique case (lizzieLet17_5QVal_Int_3_d[2:1])
        2'd0: lizzieLet17_10QVal_Int_onehotd = 4'd1;
        2'd1: lizzieLet17_10QVal_Int_onehotd = 4'd2;
        2'd2: lizzieLet17_10QVal_Int_onehotd = 4'd4;
        2'd3: lizzieLet17_10QVal_Int_onehotd = 4'd8;
        default: lizzieLet17_10QVal_Int_onehotd = 4'd0;
      endcase
    else lizzieLet17_10QVal_Int_onehotd = 4'd0;
  assign lizzieLet17_5QVal_Int_3QNone_Int_d = lizzieLet17_10QVal_Int_onehotd[0];
  assign lizzieLet17_5QVal_Int_3QVal_Int_d = lizzieLet17_10QVal_Int_onehotd[1];
  assign _95_d = lizzieLet17_10QVal_Int_onehotd[2];
  assign _94_d = lizzieLet17_10QVal_Int_onehotd[3];
  assign lizzieLet17_10QVal_Int_r = (| (lizzieLet17_10QVal_Int_onehotd & {_94_r,
                                                                          _95_r,
                                                                          lizzieLet17_5QVal_Int_3QVal_Int_r,
                                                                          lizzieLet17_5QVal_Int_3QNone_Int_r}));
  assign lizzieLet17_5QVal_Int_3_r = lizzieLet17_10QVal_Int_r;
  
  /* fork (Ty MyDTInt_Int_Int) : (lizzieLet17_5QVal_Int_3QVal_Int,MyDTInt_Int_Int) > [(lizzieLet17_5QVal_Int_3QVal_Int_1,MyDTInt_Int_Int),
                                                                                 (lizzieLet17_5QVal_Int_3QVal_Int_2,MyDTInt_Int_Int)] */
  logic [1:0] lizzieLet17_5QVal_Int_3QVal_Int_emitted;
  logic [1:0] lizzieLet17_5QVal_Int_3QVal_Int_done;
  assign lizzieLet17_5QVal_Int_3QVal_Int_1_d = (lizzieLet17_5QVal_Int_3QVal_Int_d[0] && (! lizzieLet17_5QVal_Int_3QVal_Int_emitted[0]));
  assign lizzieLet17_5QVal_Int_3QVal_Int_2_d = (lizzieLet17_5QVal_Int_3QVal_Int_d[0] && (! lizzieLet17_5QVal_Int_3QVal_Int_emitted[1]));
  assign lizzieLet17_5QVal_Int_3QVal_Int_done = (lizzieLet17_5QVal_Int_3QVal_Int_emitted | ({lizzieLet17_5QVal_Int_3QVal_Int_2_d[0],
                                                                                             lizzieLet17_5QVal_Int_3QVal_Int_1_d[0]} & {lizzieLet17_5QVal_Int_3QVal_Int_2_r,
                                                                                                                                        lizzieLet17_5QVal_Int_3QVal_Int_1_r}));
  assign lizzieLet17_5QVal_Int_3QVal_Int_r = (& lizzieLet17_5QVal_Int_3QVal_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QVal_Int_3QVal_Int_emitted <= 2'd0;
    else
      lizzieLet17_5QVal_Int_3QVal_Int_emitted <= (lizzieLet17_5QVal_Int_3QVal_Int_r ? 2'd0 :
                                                  lizzieLet17_5QVal_Int_3QVal_Int_done);
  
  /* buf (Ty MyDTInt_Int_Int) : (lizzieLet17_5QVal_Int_3QVal_Int_1,MyDTInt_Int_Int) > (lizzieLet17_5QVal_Int_3QVal_Int_1_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t lizzieLet17_5QVal_Int_3QVal_Int_1_bufchan_d;
  logic lizzieLet17_5QVal_Int_3QVal_Int_1_bufchan_r;
  assign lizzieLet17_5QVal_Int_3QVal_Int_1_r = ((! lizzieLet17_5QVal_Int_3QVal_Int_1_bufchan_d[0]) || lizzieLet17_5QVal_Int_3QVal_Int_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QVal_Int_3QVal_Int_1_bufchan_d <= 1'd0;
    else
      if (lizzieLet17_5QVal_Int_3QVal_Int_1_r)
        lizzieLet17_5QVal_Int_3QVal_Int_1_bufchan_d <= lizzieLet17_5QVal_Int_3QVal_Int_1_d;
  MyDTInt_Int_Int_t lizzieLet17_5QVal_Int_3QVal_Int_1_bufchan_buf;
  assign lizzieLet17_5QVal_Int_3QVal_Int_1_bufchan_r = (! lizzieLet17_5QVal_Int_3QVal_Int_1_bufchan_buf[0]);
  assign lizzieLet17_5QVal_Int_3QVal_Int_1_argbuf_d = (lizzieLet17_5QVal_Int_3QVal_Int_1_bufchan_buf[0] ? lizzieLet17_5QVal_Int_3QVal_Int_1_bufchan_buf :
                                                       lizzieLet17_5QVal_Int_3QVal_Int_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QVal_Int_3QVal_Int_1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet17_5QVal_Int_3QVal_Int_1_argbuf_r && lizzieLet17_5QVal_Int_3QVal_Int_1_bufchan_buf[0]))
        lizzieLet17_5QVal_Int_3QVal_Int_1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet17_5QVal_Int_3QVal_Int_1_argbuf_r) && (! lizzieLet17_5QVal_Int_3QVal_Int_1_bufchan_buf[0])))
        lizzieLet17_5QVal_Int_3QVal_Int_1_bufchan_buf <= lizzieLet17_5QVal_Int_3QVal_Int_1_bufchan_d;
  
  /* dcon (Ty TupMyDTInt_Int_Int___Int___Int,
      Dcon TupMyDTInt_Int_Int___Int___Int) : [(lizzieLet17_5QVal_Int_3QVal_Int_1_argbuf,MyDTInt_Int_Int),
                                              (lizzieLet17_5QVal_Int_10QVal_Int_1_argbuf,Int),
                                              (vaeQ_1_argbuf,Int)] > (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int7,TupMyDTInt_Int_Int___Int___Int) */
  assign applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int7_d = TupMyDTInt_Int_Int___Int___Int_dc((& {lizzieLet17_5QVal_Int_3QVal_Int_1_argbuf_d[0],
                                                                                                       lizzieLet17_5QVal_Int_10QVal_Int_1_argbuf_d[0],
                                                                                                       vaeQ_1_argbuf_d[0]}), lizzieLet17_5QVal_Int_3QVal_Int_1_argbuf_d, lizzieLet17_5QVal_Int_10QVal_Int_1_argbuf_d, vaeQ_1_argbuf_d);
  assign {lizzieLet17_5QVal_Int_3QVal_Int_1_argbuf_r,
          lizzieLet17_5QVal_Int_10QVal_Int_1_argbuf_r,
          vaeQ_1_argbuf_r} = {3 {(applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int7_r && applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int7_d[0])}};
  
  /* demux (Ty QTree_Int,
       Ty Pointer_CTf_f_Int) : (lizzieLet17_5QVal_Int_4,QTree_Int) (lizzieLet17_11QVal_Int,Pointer_CTf_f_Int) > [(lizzieLet17_5QVal_Int_4QNone_Int,Pointer_CTf_f_Int),
                                                                                                                 (lizzieLet17_5QVal_Int_4QVal_Int,Pointer_CTf_f_Int),
                                                                                                                 (lizzieLet17_5QVal_Int_4QNode_Int,Pointer_CTf_f_Int),
                                                                                                                 (lizzieLet17_5QVal_Int_4QError_Int,Pointer_CTf_f_Int)] */
  logic [3:0] lizzieLet17_11QVal_Int_onehotd;
  always_comb
    if ((lizzieLet17_5QVal_Int_4_d[0] && lizzieLet17_11QVal_Int_d[0]))
      unique case (lizzieLet17_5QVal_Int_4_d[2:1])
        2'd0: lizzieLet17_11QVal_Int_onehotd = 4'd1;
        2'd1: lizzieLet17_11QVal_Int_onehotd = 4'd2;
        2'd2: lizzieLet17_11QVal_Int_onehotd = 4'd4;
        2'd3: lizzieLet17_11QVal_Int_onehotd = 4'd8;
        default: lizzieLet17_11QVal_Int_onehotd = 4'd0;
      endcase
    else lizzieLet17_11QVal_Int_onehotd = 4'd0;
  assign lizzieLet17_5QVal_Int_4QNone_Int_d = {lizzieLet17_11QVal_Int_d[16:1],
                                               lizzieLet17_11QVal_Int_onehotd[0]};
  assign lizzieLet17_5QVal_Int_4QVal_Int_d = {lizzieLet17_11QVal_Int_d[16:1],
                                              lizzieLet17_11QVal_Int_onehotd[1]};
  assign lizzieLet17_5QVal_Int_4QNode_Int_d = {lizzieLet17_11QVal_Int_d[16:1],
                                               lizzieLet17_11QVal_Int_onehotd[2]};
  assign lizzieLet17_5QVal_Int_4QError_Int_d = {lizzieLet17_11QVal_Int_d[16:1],
                                                lizzieLet17_11QVal_Int_onehotd[3]};
  assign lizzieLet17_11QVal_Int_r = (| (lizzieLet17_11QVal_Int_onehotd & {lizzieLet17_5QVal_Int_4QError_Int_r,
                                                                          lizzieLet17_5QVal_Int_4QNode_Int_r,
                                                                          lizzieLet17_5QVal_Int_4QVal_Int_r,
                                                                          lizzieLet17_5QVal_Int_4QNone_Int_r}));
  assign lizzieLet17_5QVal_Int_4_r = lizzieLet17_11QVal_Int_r;
  
  /* buf (Ty Pointer_CTf_f_Int) : (lizzieLet17_5QVal_Int_4QError_Int,Pointer_CTf_f_Int) > (lizzieLet17_5QVal_Int_4QError_Int_1_argbuf,Pointer_CTf_f_Int) */
  Pointer_CTf_f_Int_t lizzieLet17_5QVal_Int_4QError_Int_bufchan_d;
  logic lizzieLet17_5QVal_Int_4QError_Int_bufchan_r;
  assign lizzieLet17_5QVal_Int_4QError_Int_r = ((! lizzieLet17_5QVal_Int_4QError_Int_bufchan_d[0]) || lizzieLet17_5QVal_Int_4QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QVal_Int_4QError_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet17_5QVal_Int_4QError_Int_r)
        lizzieLet17_5QVal_Int_4QError_Int_bufchan_d <= lizzieLet17_5QVal_Int_4QError_Int_d;
  Pointer_CTf_f_Int_t lizzieLet17_5QVal_Int_4QError_Int_bufchan_buf;
  assign lizzieLet17_5QVal_Int_4QError_Int_bufchan_r = (! lizzieLet17_5QVal_Int_4QError_Int_bufchan_buf[0]);
  assign lizzieLet17_5QVal_Int_4QError_Int_1_argbuf_d = (lizzieLet17_5QVal_Int_4QError_Int_bufchan_buf[0] ? lizzieLet17_5QVal_Int_4QError_Int_bufchan_buf :
                                                         lizzieLet17_5QVal_Int_4QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QVal_Int_4QError_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet17_5QVal_Int_4QError_Int_1_argbuf_r && lizzieLet17_5QVal_Int_4QError_Int_bufchan_buf[0]))
        lizzieLet17_5QVal_Int_4QError_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet17_5QVal_Int_4QError_Int_1_argbuf_r) && (! lizzieLet17_5QVal_Int_4QError_Int_bufchan_buf[0])))
        lizzieLet17_5QVal_Int_4QError_Int_bufchan_buf <= lizzieLet17_5QVal_Int_4QError_Int_bufchan_d;
  
  /* buf (Ty Pointer_CTf_f_Int) : (lizzieLet17_5QVal_Int_4QNode_Int,Pointer_CTf_f_Int) > (lizzieLet17_5QVal_Int_4QNode_Int_1_argbuf,Pointer_CTf_f_Int) */
  Pointer_CTf_f_Int_t lizzieLet17_5QVal_Int_4QNode_Int_bufchan_d;
  logic lizzieLet17_5QVal_Int_4QNode_Int_bufchan_r;
  assign lizzieLet17_5QVal_Int_4QNode_Int_r = ((! lizzieLet17_5QVal_Int_4QNode_Int_bufchan_d[0]) || lizzieLet17_5QVal_Int_4QNode_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QVal_Int_4QNode_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet17_5QVal_Int_4QNode_Int_r)
        lizzieLet17_5QVal_Int_4QNode_Int_bufchan_d <= lizzieLet17_5QVal_Int_4QNode_Int_d;
  Pointer_CTf_f_Int_t lizzieLet17_5QVal_Int_4QNode_Int_bufchan_buf;
  assign lizzieLet17_5QVal_Int_4QNode_Int_bufchan_r = (! lizzieLet17_5QVal_Int_4QNode_Int_bufchan_buf[0]);
  assign lizzieLet17_5QVal_Int_4QNode_Int_1_argbuf_d = (lizzieLet17_5QVal_Int_4QNode_Int_bufchan_buf[0] ? lizzieLet17_5QVal_Int_4QNode_Int_bufchan_buf :
                                                        lizzieLet17_5QVal_Int_4QNode_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QVal_Int_4QNode_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet17_5QVal_Int_4QNode_Int_1_argbuf_r && lizzieLet17_5QVal_Int_4QNode_Int_bufchan_buf[0]))
        lizzieLet17_5QVal_Int_4QNode_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet17_5QVal_Int_4QNode_Int_1_argbuf_r) && (! lizzieLet17_5QVal_Int_4QNode_Int_bufchan_buf[0])))
        lizzieLet17_5QVal_Int_4QNode_Int_bufchan_buf <= lizzieLet17_5QVal_Int_4QNode_Int_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Go) : (lizzieLet17_5QVal_Int_5,QTree_Int) (lizzieLet17_3QVal_Int,Go) > [(lizzieLet17_5QVal_Int_5QNone_Int,Go),
                                                                                  (lizzieLet17_5QVal_Int_5QVal_Int,Go),
                                                                                  (lizzieLet17_5QVal_Int_5QNode_Int,Go),
                                                                                  (lizzieLet17_5QVal_Int_5QError_Int,Go)] */
  logic [3:0] lizzieLet17_3QVal_Int_onehotd;
  always_comb
    if ((lizzieLet17_5QVal_Int_5_d[0] && lizzieLet17_3QVal_Int_d[0]))
      unique case (lizzieLet17_5QVal_Int_5_d[2:1])
        2'd0: lizzieLet17_3QVal_Int_onehotd = 4'd1;
        2'd1: lizzieLet17_3QVal_Int_onehotd = 4'd2;
        2'd2: lizzieLet17_3QVal_Int_onehotd = 4'd4;
        2'd3: lizzieLet17_3QVal_Int_onehotd = 4'd8;
        default: lizzieLet17_3QVal_Int_onehotd = 4'd0;
      endcase
    else lizzieLet17_3QVal_Int_onehotd = 4'd0;
  assign lizzieLet17_5QVal_Int_5QNone_Int_d = lizzieLet17_3QVal_Int_onehotd[0];
  assign lizzieLet17_5QVal_Int_5QVal_Int_d = lizzieLet17_3QVal_Int_onehotd[1];
  assign lizzieLet17_5QVal_Int_5QNode_Int_d = lizzieLet17_3QVal_Int_onehotd[2];
  assign lizzieLet17_5QVal_Int_5QError_Int_d = lizzieLet17_3QVal_Int_onehotd[3];
  assign lizzieLet17_3QVal_Int_r = (| (lizzieLet17_3QVal_Int_onehotd & {lizzieLet17_5QVal_Int_5QError_Int_r,
                                                                        lizzieLet17_5QVal_Int_5QNode_Int_r,
                                                                        lizzieLet17_5QVal_Int_5QVal_Int_r,
                                                                        lizzieLet17_5QVal_Int_5QNone_Int_r}));
  assign lizzieLet17_5QVal_Int_5_r = lizzieLet17_3QVal_Int_r;
  
  /* fork (Ty Go) : (lizzieLet17_5QVal_Int_5QError_Int,Go) > [(lizzieLet17_5QVal_Int_5QError_Int_1,Go),
                                                         (lizzieLet17_5QVal_Int_5QError_Int_2,Go)] */
  logic [1:0] lizzieLet17_5QVal_Int_5QError_Int_emitted;
  logic [1:0] lizzieLet17_5QVal_Int_5QError_Int_done;
  assign lizzieLet17_5QVal_Int_5QError_Int_1_d = (lizzieLet17_5QVal_Int_5QError_Int_d[0] && (! lizzieLet17_5QVal_Int_5QError_Int_emitted[0]));
  assign lizzieLet17_5QVal_Int_5QError_Int_2_d = (lizzieLet17_5QVal_Int_5QError_Int_d[0] && (! lizzieLet17_5QVal_Int_5QError_Int_emitted[1]));
  assign lizzieLet17_5QVal_Int_5QError_Int_done = (lizzieLet17_5QVal_Int_5QError_Int_emitted | ({lizzieLet17_5QVal_Int_5QError_Int_2_d[0],
                                                                                                 lizzieLet17_5QVal_Int_5QError_Int_1_d[0]} & {lizzieLet17_5QVal_Int_5QError_Int_2_r,
                                                                                                                                              lizzieLet17_5QVal_Int_5QError_Int_1_r}));
  assign lizzieLet17_5QVal_Int_5QError_Int_r = (& lizzieLet17_5QVal_Int_5QError_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QVal_Int_5QError_Int_emitted <= 2'd0;
    else
      lizzieLet17_5QVal_Int_5QError_Int_emitted <= (lizzieLet17_5QVal_Int_5QError_Int_r ? 2'd0 :
                                                    lizzieLet17_5QVal_Int_5QError_Int_done);
  
  /* dcon (Ty QTree_Int,
      Dcon QError_Int) : [(lizzieLet17_5QVal_Int_5QError_Int_1,Go)] > (lizzieLet17_5QVal_Int_5QError_Int_1QError_Int,QTree_Int) */
  assign lizzieLet17_5QVal_Int_5QError_Int_1QError_Int_d = QError_Int_dc((& {lizzieLet17_5QVal_Int_5QError_Int_1_d[0]}), lizzieLet17_5QVal_Int_5QError_Int_1_d);
  assign {lizzieLet17_5QVal_Int_5QError_Int_1_r} = {1 {(lizzieLet17_5QVal_Int_5QError_Int_1QError_Int_r && lizzieLet17_5QVal_Int_5QError_Int_1QError_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (lizzieLet17_5QVal_Int_5QError_Int_1QError_Int,QTree_Int) > (lizzieLet42_1_argbuf,QTree_Int) */
  QTree_Int_t lizzieLet17_5QVal_Int_5QError_Int_1QError_Int_bufchan_d;
  logic lizzieLet17_5QVal_Int_5QError_Int_1QError_Int_bufchan_r;
  assign lizzieLet17_5QVal_Int_5QError_Int_1QError_Int_r = ((! lizzieLet17_5QVal_Int_5QError_Int_1QError_Int_bufchan_d[0]) || lizzieLet17_5QVal_Int_5QError_Int_1QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QVal_Int_5QError_Int_1QError_Int_bufchan_d <= {66'd0,
                                                                  1'd0};
    else
      if (lizzieLet17_5QVal_Int_5QError_Int_1QError_Int_r)
        lizzieLet17_5QVal_Int_5QError_Int_1QError_Int_bufchan_d <= lizzieLet17_5QVal_Int_5QError_Int_1QError_Int_d;
  QTree_Int_t lizzieLet17_5QVal_Int_5QError_Int_1QError_Int_bufchan_buf;
  assign lizzieLet17_5QVal_Int_5QError_Int_1QError_Int_bufchan_r = (! lizzieLet17_5QVal_Int_5QError_Int_1QError_Int_bufchan_buf[0]);
  assign lizzieLet42_1_argbuf_d = (lizzieLet17_5QVal_Int_5QError_Int_1QError_Int_bufchan_buf[0] ? lizzieLet17_5QVal_Int_5QError_Int_1QError_Int_bufchan_buf :
                                   lizzieLet17_5QVal_Int_5QError_Int_1QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QVal_Int_5QError_Int_1QError_Int_bufchan_buf <= {66'd0,
                                                                    1'd0};
    else
      if ((lizzieLet42_1_argbuf_r && lizzieLet17_5QVal_Int_5QError_Int_1QError_Int_bufchan_buf[0]))
        lizzieLet17_5QVal_Int_5QError_Int_1QError_Int_bufchan_buf <= {66'd0,
                                                                      1'd0};
      else if (((! lizzieLet42_1_argbuf_r) && (! lizzieLet17_5QVal_Int_5QError_Int_1QError_Int_bufchan_buf[0])))
        lizzieLet17_5QVal_Int_5QError_Int_1QError_Int_bufchan_buf <= lizzieLet17_5QVal_Int_5QError_Int_1QError_Int_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet17_5QVal_Int_5QError_Int_2,Go) > (lizzieLet17_5QVal_Int_5QError_Int_2_argbuf,Go) */
  Go_t lizzieLet17_5QVal_Int_5QError_Int_2_bufchan_d;
  logic lizzieLet17_5QVal_Int_5QError_Int_2_bufchan_r;
  assign lizzieLet17_5QVal_Int_5QError_Int_2_r = ((! lizzieLet17_5QVal_Int_5QError_Int_2_bufchan_d[0]) || lizzieLet17_5QVal_Int_5QError_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QVal_Int_5QError_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet17_5QVal_Int_5QError_Int_2_r)
        lizzieLet17_5QVal_Int_5QError_Int_2_bufchan_d <= lizzieLet17_5QVal_Int_5QError_Int_2_d;
  Go_t lizzieLet17_5QVal_Int_5QError_Int_2_bufchan_buf;
  assign lizzieLet17_5QVal_Int_5QError_Int_2_bufchan_r = (! lizzieLet17_5QVal_Int_5QError_Int_2_bufchan_buf[0]);
  assign lizzieLet17_5QVal_Int_5QError_Int_2_argbuf_d = (lizzieLet17_5QVal_Int_5QError_Int_2_bufchan_buf[0] ? lizzieLet17_5QVal_Int_5QError_Int_2_bufchan_buf :
                                                         lizzieLet17_5QVal_Int_5QError_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QVal_Int_5QError_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet17_5QVal_Int_5QError_Int_2_argbuf_r && lizzieLet17_5QVal_Int_5QError_Int_2_bufchan_buf[0]))
        lizzieLet17_5QVal_Int_5QError_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet17_5QVal_Int_5QError_Int_2_argbuf_r) && (! lizzieLet17_5QVal_Int_5QError_Int_2_bufchan_buf[0])))
        lizzieLet17_5QVal_Int_5QError_Int_2_bufchan_buf <= lizzieLet17_5QVal_Int_5QError_Int_2_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet17_5QVal_Int_5QNode_Int,Go) > [(lizzieLet17_5QVal_Int_5QNode_Int_1,Go),
                                                        (lizzieLet17_5QVal_Int_5QNode_Int_2,Go)] */
  logic [1:0] lizzieLet17_5QVal_Int_5QNode_Int_emitted;
  logic [1:0] lizzieLet17_5QVal_Int_5QNode_Int_done;
  assign lizzieLet17_5QVal_Int_5QNode_Int_1_d = (lizzieLet17_5QVal_Int_5QNode_Int_d[0] && (! lizzieLet17_5QVal_Int_5QNode_Int_emitted[0]));
  assign lizzieLet17_5QVal_Int_5QNode_Int_2_d = (lizzieLet17_5QVal_Int_5QNode_Int_d[0] && (! lizzieLet17_5QVal_Int_5QNode_Int_emitted[1]));
  assign lizzieLet17_5QVal_Int_5QNode_Int_done = (lizzieLet17_5QVal_Int_5QNode_Int_emitted | ({lizzieLet17_5QVal_Int_5QNode_Int_2_d[0],
                                                                                               lizzieLet17_5QVal_Int_5QNode_Int_1_d[0]} & {lizzieLet17_5QVal_Int_5QNode_Int_2_r,
                                                                                                                                           lizzieLet17_5QVal_Int_5QNode_Int_1_r}));
  assign lizzieLet17_5QVal_Int_5QNode_Int_r = (& lizzieLet17_5QVal_Int_5QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QVal_Int_5QNode_Int_emitted <= 2'd0;
    else
      lizzieLet17_5QVal_Int_5QNode_Int_emitted <= (lizzieLet17_5QVal_Int_5QNode_Int_r ? 2'd0 :
                                                   lizzieLet17_5QVal_Int_5QNode_Int_done);
  
  /* dcon (Ty QTree_Int,
      Dcon QError_Int) : [(lizzieLet17_5QVal_Int_5QNode_Int_1,Go)] > (lizzieLet17_5QVal_Int_5QNode_Int_1QError_Int,QTree_Int) */
  assign lizzieLet17_5QVal_Int_5QNode_Int_1QError_Int_d = QError_Int_dc((& {lizzieLet17_5QVal_Int_5QNode_Int_1_d[0]}), lizzieLet17_5QVal_Int_5QNode_Int_1_d);
  assign {lizzieLet17_5QVal_Int_5QNode_Int_1_r} = {1 {(lizzieLet17_5QVal_Int_5QNode_Int_1QError_Int_r && lizzieLet17_5QVal_Int_5QNode_Int_1QError_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (lizzieLet17_5QVal_Int_5QNode_Int_1QError_Int,QTree_Int) > (lizzieLet41_1_argbuf,QTree_Int) */
  QTree_Int_t lizzieLet17_5QVal_Int_5QNode_Int_1QError_Int_bufchan_d;
  logic lizzieLet17_5QVal_Int_5QNode_Int_1QError_Int_bufchan_r;
  assign lizzieLet17_5QVal_Int_5QNode_Int_1QError_Int_r = ((! lizzieLet17_5QVal_Int_5QNode_Int_1QError_Int_bufchan_d[0]) || lizzieLet17_5QVal_Int_5QNode_Int_1QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QVal_Int_5QNode_Int_1QError_Int_bufchan_d <= {66'd0,
                                                                 1'd0};
    else
      if (lizzieLet17_5QVal_Int_5QNode_Int_1QError_Int_r)
        lizzieLet17_5QVal_Int_5QNode_Int_1QError_Int_bufchan_d <= lizzieLet17_5QVal_Int_5QNode_Int_1QError_Int_d;
  QTree_Int_t lizzieLet17_5QVal_Int_5QNode_Int_1QError_Int_bufchan_buf;
  assign lizzieLet17_5QVal_Int_5QNode_Int_1QError_Int_bufchan_r = (! lizzieLet17_5QVal_Int_5QNode_Int_1QError_Int_bufchan_buf[0]);
  assign lizzieLet41_1_argbuf_d = (lizzieLet17_5QVal_Int_5QNode_Int_1QError_Int_bufchan_buf[0] ? lizzieLet17_5QVal_Int_5QNode_Int_1QError_Int_bufchan_buf :
                                   lizzieLet17_5QVal_Int_5QNode_Int_1QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QVal_Int_5QNode_Int_1QError_Int_bufchan_buf <= {66'd0,
                                                                   1'd0};
    else
      if ((lizzieLet41_1_argbuf_r && lizzieLet17_5QVal_Int_5QNode_Int_1QError_Int_bufchan_buf[0]))
        lizzieLet17_5QVal_Int_5QNode_Int_1QError_Int_bufchan_buf <= {66'd0,
                                                                     1'd0};
      else if (((! lizzieLet41_1_argbuf_r) && (! lizzieLet17_5QVal_Int_5QNode_Int_1QError_Int_bufchan_buf[0])))
        lizzieLet17_5QVal_Int_5QNode_Int_1QError_Int_bufchan_buf <= lizzieLet17_5QVal_Int_5QNode_Int_1QError_Int_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet17_5QVal_Int_5QNode_Int_2,Go) > (lizzieLet17_5QVal_Int_5QNode_Int_2_argbuf,Go) */
  Go_t lizzieLet17_5QVal_Int_5QNode_Int_2_bufchan_d;
  logic lizzieLet17_5QVal_Int_5QNode_Int_2_bufchan_r;
  assign lizzieLet17_5QVal_Int_5QNode_Int_2_r = ((! lizzieLet17_5QVal_Int_5QNode_Int_2_bufchan_d[0]) || lizzieLet17_5QVal_Int_5QNode_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QVal_Int_5QNode_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet17_5QVal_Int_5QNode_Int_2_r)
        lizzieLet17_5QVal_Int_5QNode_Int_2_bufchan_d <= lizzieLet17_5QVal_Int_5QNode_Int_2_d;
  Go_t lizzieLet17_5QVal_Int_5QNode_Int_2_bufchan_buf;
  assign lizzieLet17_5QVal_Int_5QNode_Int_2_bufchan_r = (! lizzieLet17_5QVal_Int_5QNode_Int_2_bufchan_buf[0]);
  assign lizzieLet17_5QVal_Int_5QNode_Int_2_argbuf_d = (lizzieLet17_5QVal_Int_5QNode_Int_2_bufchan_buf[0] ? lizzieLet17_5QVal_Int_5QNode_Int_2_bufchan_buf :
                                                        lizzieLet17_5QVal_Int_5QNode_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QVal_Int_5QNode_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet17_5QVal_Int_5QNode_Int_2_argbuf_r && lizzieLet17_5QVal_Int_5QNode_Int_2_bufchan_buf[0]))
        lizzieLet17_5QVal_Int_5QNode_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet17_5QVal_Int_5QNode_Int_2_argbuf_r) && (! lizzieLet17_5QVal_Int_5QNode_Int_2_bufchan_buf[0])))
        lizzieLet17_5QVal_Int_5QNode_Int_2_bufchan_buf <= lizzieLet17_5QVal_Int_5QNode_Int_2_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet17_5QVal_Int_5QVal_Int,Go) > [(lizzieLet17_5QVal_Int_5QVal_Int_1,Go),
                                                       (lizzieLet17_5QVal_Int_5QVal_Int_2,Go)] */
  logic [1:0] lizzieLet17_5QVal_Int_5QVal_Int_emitted;
  logic [1:0] lizzieLet17_5QVal_Int_5QVal_Int_done;
  assign lizzieLet17_5QVal_Int_5QVal_Int_1_d = (lizzieLet17_5QVal_Int_5QVal_Int_d[0] && (! lizzieLet17_5QVal_Int_5QVal_Int_emitted[0]));
  assign lizzieLet17_5QVal_Int_5QVal_Int_2_d = (lizzieLet17_5QVal_Int_5QVal_Int_d[0] && (! lizzieLet17_5QVal_Int_5QVal_Int_emitted[1]));
  assign lizzieLet17_5QVal_Int_5QVal_Int_done = (lizzieLet17_5QVal_Int_5QVal_Int_emitted | ({lizzieLet17_5QVal_Int_5QVal_Int_2_d[0],
                                                                                             lizzieLet17_5QVal_Int_5QVal_Int_1_d[0]} & {lizzieLet17_5QVal_Int_5QVal_Int_2_r,
                                                                                                                                        lizzieLet17_5QVal_Int_5QVal_Int_1_r}));
  assign lizzieLet17_5QVal_Int_5QVal_Int_r = (& lizzieLet17_5QVal_Int_5QVal_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QVal_Int_5QVal_Int_emitted <= 2'd0;
    else
      lizzieLet17_5QVal_Int_5QVal_Int_emitted <= (lizzieLet17_5QVal_Int_5QVal_Int_r ? 2'd0 :
                                                  lizzieLet17_5QVal_Int_5QVal_Int_done);
  
  /* buf (Ty Go) : (lizzieLet17_5QVal_Int_5QVal_Int_1,Go) > (lizzieLet17_5QVal_Int_5QVal_Int_1_argbuf,Go) */
  Go_t lizzieLet17_5QVal_Int_5QVal_Int_1_bufchan_d;
  logic lizzieLet17_5QVal_Int_5QVal_Int_1_bufchan_r;
  assign lizzieLet17_5QVal_Int_5QVal_Int_1_r = ((! lizzieLet17_5QVal_Int_5QVal_Int_1_bufchan_d[0]) || lizzieLet17_5QVal_Int_5QVal_Int_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QVal_Int_5QVal_Int_1_bufchan_d <= 1'd0;
    else
      if (lizzieLet17_5QVal_Int_5QVal_Int_1_r)
        lizzieLet17_5QVal_Int_5QVal_Int_1_bufchan_d <= lizzieLet17_5QVal_Int_5QVal_Int_1_d;
  Go_t lizzieLet17_5QVal_Int_5QVal_Int_1_bufchan_buf;
  assign lizzieLet17_5QVal_Int_5QVal_Int_1_bufchan_r = (! lizzieLet17_5QVal_Int_5QVal_Int_1_bufchan_buf[0]);
  assign lizzieLet17_5QVal_Int_5QVal_Int_1_argbuf_d = (lizzieLet17_5QVal_Int_5QVal_Int_1_bufchan_buf[0] ? lizzieLet17_5QVal_Int_5QVal_Int_1_bufchan_buf :
                                                       lizzieLet17_5QVal_Int_5QVal_Int_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QVal_Int_5QVal_Int_1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet17_5QVal_Int_5QVal_Int_1_argbuf_r && lizzieLet17_5QVal_Int_5QVal_Int_1_bufchan_buf[0]))
        lizzieLet17_5QVal_Int_5QVal_Int_1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet17_5QVal_Int_5QVal_Int_1_argbuf_r) && (! lizzieLet17_5QVal_Int_5QVal_Int_1_bufchan_buf[0])))
        lizzieLet17_5QVal_Int_5QVal_Int_1_bufchan_buf <= lizzieLet17_5QVal_Int_5QVal_Int_1_bufchan_d;
  
  /* dcon (Ty TupGo___MyDTInt_Bool___Int,
      Dcon TupGo___MyDTInt_Bool___Int) : [(lizzieLet17_5QVal_Int_5QVal_Int_1_argbuf,Go),
                                          (lizzieLet17_5QVal_Int_6QVal_Int_1_argbuf,MyDTInt_Bool),
                                          (es_13_1_argbuf,Int)] > (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int4,TupGo___MyDTInt_Bool___Int) */
  assign applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int4_d = TupGo___MyDTInt_Bool___Int_dc((& {lizzieLet17_5QVal_Int_5QVal_Int_1_argbuf_d[0],
                                                                                            lizzieLet17_5QVal_Int_6QVal_Int_1_argbuf_d[0],
                                                                                            es_13_1_argbuf_d[0]}), lizzieLet17_5QVal_Int_5QVal_Int_1_argbuf_d, lizzieLet17_5QVal_Int_6QVal_Int_1_argbuf_d, es_13_1_argbuf_d);
  assign {lizzieLet17_5QVal_Int_5QVal_Int_1_argbuf_r,
          lizzieLet17_5QVal_Int_6QVal_Int_1_argbuf_r,
          es_13_1_argbuf_r} = {3 {(applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int4_r && applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int4_d[0])}};
  
  /* demux (Ty QTree_Int,
       Ty MyDTInt_Bool) : (lizzieLet17_5QVal_Int_6,QTree_Int) (lizzieLet17_4QVal_Int,MyDTInt_Bool) > [(lizzieLet17_5QVal_Int_6QNone_Int,MyDTInt_Bool),
                                                                                                      (lizzieLet17_5QVal_Int_6QVal_Int,MyDTInt_Bool),
                                                                                                      (_93,MyDTInt_Bool),
                                                                                                      (_92,MyDTInt_Bool)] */
  logic [3:0] lizzieLet17_4QVal_Int_onehotd;
  always_comb
    if ((lizzieLet17_5QVal_Int_6_d[0] && lizzieLet17_4QVal_Int_d[0]))
      unique case (lizzieLet17_5QVal_Int_6_d[2:1])
        2'd0: lizzieLet17_4QVal_Int_onehotd = 4'd1;
        2'd1: lizzieLet17_4QVal_Int_onehotd = 4'd2;
        2'd2: lizzieLet17_4QVal_Int_onehotd = 4'd4;
        2'd3: lizzieLet17_4QVal_Int_onehotd = 4'd8;
        default: lizzieLet17_4QVal_Int_onehotd = 4'd0;
      endcase
    else lizzieLet17_4QVal_Int_onehotd = 4'd0;
  assign lizzieLet17_5QVal_Int_6QNone_Int_d = lizzieLet17_4QVal_Int_onehotd[0];
  assign lizzieLet17_5QVal_Int_6QVal_Int_d = lizzieLet17_4QVal_Int_onehotd[1];
  assign _93_d = lizzieLet17_4QVal_Int_onehotd[2];
  assign _92_d = lizzieLet17_4QVal_Int_onehotd[3];
  assign lizzieLet17_4QVal_Int_r = (| (lizzieLet17_4QVal_Int_onehotd & {_92_r,
                                                                        _93_r,
                                                                        lizzieLet17_5QVal_Int_6QVal_Int_r,
                                                                        lizzieLet17_5QVal_Int_6QNone_Int_r}));
  assign lizzieLet17_5QVal_Int_6_r = lizzieLet17_4QVal_Int_r;
  
  /* fork (Ty MyDTInt_Bool) : (lizzieLet17_5QVal_Int_6QVal_Int,MyDTInt_Bool) > [(lizzieLet17_5QVal_Int_6QVal_Int_1,MyDTInt_Bool),
                                                                           (lizzieLet17_5QVal_Int_6QVal_Int_2,MyDTInt_Bool)] */
  logic [1:0] lizzieLet17_5QVal_Int_6QVal_Int_emitted;
  logic [1:0] lizzieLet17_5QVal_Int_6QVal_Int_done;
  assign lizzieLet17_5QVal_Int_6QVal_Int_1_d = (lizzieLet17_5QVal_Int_6QVal_Int_d[0] && (! lizzieLet17_5QVal_Int_6QVal_Int_emitted[0]));
  assign lizzieLet17_5QVal_Int_6QVal_Int_2_d = (lizzieLet17_5QVal_Int_6QVal_Int_d[0] && (! lizzieLet17_5QVal_Int_6QVal_Int_emitted[1]));
  assign lizzieLet17_5QVal_Int_6QVal_Int_done = (lizzieLet17_5QVal_Int_6QVal_Int_emitted | ({lizzieLet17_5QVal_Int_6QVal_Int_2_d[0],
                                                                                             lizzieLet17_5QVal_Int_6QVal_Int_1_d[0]} & {lizzieLet17_5QVal_Int_6QVal_Int_2_r,
                                                                                                                                        lizzieLet17_5QVal_Int_6QVal_Int_1_r}));
  assign lizzieLet17_5QVal_Int_6QVal_Int_r = (& lizzieLet17_5QVal_Int_6QVal_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QVal_Int_6QVal_Int_emitted <= 2'd0;
    else
      lizzieLet17_5QVal_Int_6QVal_Int_emitted <= (lizzieLet17_5QVal_Int_6QVal_Int_r ? 2'd0 :
                                                  lizzieLet17_5QVal_Int_6QVal_Int_done);
  
  /* buf (Ty MyDTInt_Bool) : (lizzieLet17_5QVal_Int_6QVal_Int_1,MyDTInt_Bool) > (lizzieLet17_5QVal_Int_6QVal_Int_1_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t lizzieLet17_5QVal_Int_6QVal_Int_1_bufchan_d;
  logic lizzieLet17_5QVal_Int_6QVal_Int_1_bufchan_r;
  assign lizzieLet17_5QVal_Int_6QVal_Int_1_r = ((! lizzieLet17_5QVal_Int_6QVal_Int_1_bufchan_d[0]) || lizzieLet17_5QVal_Int_6QVal_Int_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QVal_Int_6QVal_Int_1_bufchan_d <= 1'd0;
    else
      if (lizzieLet17_5QVal_Int_6QVal_Int_1_r)
        lizzieLet17_5QVal_Int_6QVal_Int_1_bufchan_d <= lizzieLet17_5QVal_Int_6QVal_Int_1_d;
  MyDTInt_Bool_t lizzieLet17_5QVal_Int_6QVal_Int_1_bufchan_buf;
  assign lizzieLet17_5QVal_Int_6QVal_Int_1_bufchan_r = (! lizzieLet17_5QVal_Int_6QVal_Int_1_bufchan_buf[0]);
  assign lizzieLet17_5QVal_Int_6QVal_Int_1_argbuf_d = (lizzieLet17_5QVal_Int_6QVal_Int_1_bufchan_buf[0] ? lizzieLet17_5QVal_Int_6QVal_Int_1_bufchan_buf :
                                                       lizzieLet17_5QVal_Int_6QVal_Int_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QVal_Int_6QVal_Int_1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet17_5QVal_Int_6QVal_Int_1_argbuf_r && lizzieLet17_5QVal_Int_6QVal_Int_1_bufchan_buf[0]))
        lizzieLet17_5QVal_Int_6QVal_Int_1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet17_5QVal_Int_6QVal_Int_1_argbuf_r) && (! lizzieLet17_5QVal_Int_6QVal_Int_1_bufchan_buf[0])))
        lizzieLet17_5QVal_Int_6QVal_Int_1_bufchan_buf <= lizzieLet17_5QVal_Int_6QVal_Int_1_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty QTree_Int) : (lizzieLet17_5QVal_Int_7,QTree_Int) (lizzieLet17_6QVal_Int,QTree_Int) > [(lizzieLet17_5QVal_Int_7QNone_Int,QTree_Int),
                                                                                                (lizzieLet17_5QVal_Int_7QVal_Int,QTree_Int),
                                                                                                (_91,QTree_Int),
                                                                                                (_90,QTree_Int)] */
  logic [3:0] lizzieLet17_6QVal_Int_onehotd;
  always_comb
    if ((lizzieLet17_5QVal_Int_7_d[0] && lizzieLet17_6QVal_Int_d[0]))
      unique case (lizzieLet17_5QVal_Int_7_d[2:1])
        2'd0: lizzieLet17_6QVal_Int_onehotd = 4'd1;
        2'd1: lizzieLet17_6QVal_Int_onehotd = 4'd2;
        2'd2: lizzieLet17_6QVal_Int_onehotd = 4'd4;
        2'd3: lizzieLet17_6QVal_Int_onehotd = 4'd8;
        default: lizzieLet17_6QVal_Int_onehotd = 4'd0;
      endcase
    else lizzieLet17_6QVal_Int_onehotd = 4'd0;
  assign lizzieLet17_5QVal_Int_7QNone_Int_d = {lizzieLet17_6QVal_Int_d[66:1],
                                               lizzieLet17_6QVal_Int_onehotd[0]};
  assign lizzieLet17_5QVal_Int_7QVal_Int_d = {lizzieLet17_6QVal_Int_d[66:1],
                                              lizzieLet17_6QVal_Int_onehotd[1]};
  assign _91_d = {lizzieLet17_6QVal_Int_d[66:1],
                  lizzieLet17_6QVal_Int_onehotd[2]};
  assign _90_d = {lizzieLet17_6QVal_Int_d[66:1],
                  lizzieLet17_6QVal_Int_onehotd[3]};
  assign lizzieLet17_6QVal_Int_r = (| (lizzieLet17_6QVal_Int_onehotd & {_90_r,
                                                                        _91_r,
                                                                        lizzieLet17_5QVal_Int_7QVal_Int_r,
                                                                        lizzieLet17_5QVal_Int_7QNone_Int_r}));
  assign lizzieLet17_5QVal_Int_7_r = lizzieLet17_6QVal_Int_r;
  
  /* fork (Ty QTree_Int) : (lizzieLet17_5QVal_Int_7QNone_Int,QTree_Int) > [(lizzieLet17_5QVal_Int_7QNone_Int_1,QTree_Int),
                                                                      (lizzieLet17_5QVal_Int_7QNone_Int_2,QTree_Int),
                                                                      (lizzieLet17_5QVal_Int_7QNone_Int_3,QTree_Int),
                                                                      (lizzieLet17_5QVal_Int_7QNone_Int_4,QTree_Int),
                                                                      (lizzieLet17_5QVal_Int_7QNone_Int_5,QTree_Int),
                                                                      (lizzieLet17_5QVal_Int_7QNone_Int_6,QTree_Int),
                                                                      (lizzieLet17_5QVal_Int_7QNone_Int_7,QTree_Int),
                                                                      (lizzieLet17_5QVal_Int_7QNone_Int_8,QTree_Int)] */
  logic [7:0] lizzieLet17_5QVal_Int_7QNone_Int_emitted;
  logic [7:0] lizzieLet17_5QVal_Int_7QNone_Int_done;
  assign lizzieLet17_5QVal_Int_7QNone_Int_1_d = {lizzieLet17_5QVal_Int_7QNone_Int_d[66:1],
                                                 (lizzieLet17_5QVal_Int_7QNone_Int_d[0] && (! lizzieLet17_5QVal_Int_7QNone_Int_emitted[0]))};
  assign lizzieLet17_5QVal_Int_7QNone_Int_2_d = {lizzieLet17_5QVal_Int_7QNone_Int_d[66:1],
                                                 (lizzieLet17_5QVal_Int_7QNone_Int_d[0] && (! lizzieLet17_5QVal_Int_7QNone_Int_emitted[1]))};
  assign lizzieLet17_5QVal_Int_7QNone_Int_3_d = {lizzieLet17_5QVal_Int_7QNone_Int_d[66:1],
                                                 (lizzieLet17_5QVal_Int_7QNone_Int_d[0] && (! lizzieLet17_5QVal_Int_7QNone_Int_emitted[2]))};
  assign lizzieLet17_5QVal_Int_7QNone_Int_4_d = {lizzieLet17_5QVal_Int_7QNone_Int_d[66:1],
                                                 (lizzieLet17_5QVal_Int_7QNone_Int_d[0] && (! lizzieLet17_5QVal_Int_7QNone_Int_emitted[3]))};
  assign lizzieLet17_5QVal_Int_7QNone_Int_5_d = {lizzieLet17_5QVal_Int_7QNone_Int_d[66:1],
                                                 (lizzieLet17_5QVal_Int_7QNone_Int_d[0] && (! lizzieLet17_5QVal_Int_7QNone_Int_emitted[4]))};
  assign lizzieLet17_5QVal_Int_7QNone_Int_6_d = {lizzieLet17_5QVal_Int_7QNone_Int_d[66:1],
                                                 (lizzieLet17_5QVal_Int_7QNone_Int_d[0] && (! lizzieLet17_5QVal_Int_7QNone_Int_emitted[5]))};
  assign lizzieLet17_5QVal_Int_7QNone_Int_7_d = {lizzieLet17_5QVal_Int_7QNone_Int_d[66:1],
                                                 (lizzieLet17_5QVal_Int_7QNone_Int_d[0] && (! lizzieLet17_5QVal_Int_7QNone_Int_emitted[6]))};
  assign lizzieLet17_5QVal_Int_7QNone_Int_8_d = {lizzieLet17_5QVal_Int_7QNone_Int_d[66:1],
                                                 (lizzieLet17_5QVal_Int_7QNone_Int_d[0] && (! lizzieLet17_5QVal_Int_7QNone_Int_emitted[7]))};
  assign lizzieLet17_5QVal_Int_7QNone_Int_done = (lizzieLet17_5QVal_Int_7QNone_Int_emitted | ({lizzieLet17_5QVal_Int_7QNone_Int_8_d[0],
                                                                                               lizzieLet17_5QVal_Int_7QNone_Int_7_d[0],
                                                                                               lizzieLet17_5QVal_Int_7QNone_Int_6_d[0],
                                                                                               lizzieLet17_5QVal_Int_7QNone_Int_5_d[0],
                                                                                               lizzieLet17_5QVal_Int_7QNone_Int_4_d[0],
                                                                                               lizzieLet17_5QVal_Int_7QNone_Int_3_d[0],
                                                                                               lizzieLet17_5QVal_Int_7QNone_Int_2_d[0],
                                                                                               lizzieLet17_5QVal_Int_7QNone_Int_1_d[0]} & {lizzieLet17_5QVal_Int_7QNone_Int_8_r,
                                                                                                                                           lizzieLet17_5QVal_Int_7QNone_Int_7_r,
                                                                                                                                           lizzieLet17_5QVal_Int_7QNone_Int_6_r,
                                                                                                                                           lizzieLet17_5QVal_Int_7QNone_Int_5_r,
                                                                                                                                           lizzieLet17_5QVal_Int_7QNone_Int_4_r,
                                                                                                                                           lizzieLet17_5QVal_Int_7QNone_Int_3_r,
                                                                                                                                           lizzieLet17_5QVal_Int_7QNone_Int_2_r,
                                                                                                                                           lizzieLet17_5QVal_Int_7QNone_Int_1_r}));
  assign lizzieLet17_5QVal_Int_7QNone_Int_r = (& lizzieLet17_5QVal_Int_7QNone_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QVal_Int_7QNone_Int_emitted <= 8'd0;
    else
      lizzieLet17_5QVal_Int_7QNone_Int_emitted <= (lizzieLet17_5QVal_Int_7QNone_Int_r ? 8'd0 :
                                                   lizzieLet17_5QVal_Int_7QNone_Int_done);
  
  /* destruct (Ty QTree_Int,
          Dcon QVal_Int) : (lizzieLet17_5QVal_Int_7QNone_Int_1QVal_Int,QTree_Int) > [(vaeL_destruct,Int)] */
  assign vaeL_destruct_d = {lizzieLet17_5QVal_Int_7QNone_Int_1QVal_Int_d[34:3],
                            lizzieLet17_5QVal_Int_7QNone_Int_1QVal_Int_d[0]};
  assign lizzieLet17_5QVal_Int_7QNone_Int_1QVal_Int_r = vaeL_destruct_r;
  
  /* demux (Ty QTree_Int,
       Ty QTree_Int) : (lizzieLet17_5QVal_Int_7QNone_Int_2,QTree_Int) (lizzieLet17_5QVal_Int_7QNone_Int_1,QTree_Int) > [(_89,QTree_Int),
                                                                                                                        (lizzieLet17_5QVal_Int_7QNone_Int_1QVal_Int,QTree_Int),
                                                                                                                        (_88,QTree_Int),
                                                                                                                        (_87,QTree_Int)] */
  logic [3:0] lizzieLet17_5QVal_Int_7QNone_Int_1_onehotd;
  always_comb
    if ((lizzieLet17_5QVal_Int_7QNone_Int_2_d[0] && lizzieLet17_5QVal_Int_7QNone_Int_1_d[0]))
      unique case (lizzieLet17_5QVal_Int_7QNone_Int_2_d[2:1])
        2'd0: lizzieLet17_5QVal_Int_7QNone_Int_1_onehotd = 4'd1;
        2'd1: lizzieLet17_5QVal_Int_7QNone_Int_1_onehotd = 4'd2;
        2'd2: lizzieLet17_5QVal_Int_7QNone_Int_1_onehotd = 4'd4;
        2'd3: lizzieLet17_5QVal_Int_7QNone_Int_1_onehotd = 4'd8;
        default: lizzieLet17_5QVal_Int_7QNone_Int_1_onehotd = 4'd0;
      endcase
    else lizzieLet17_5QVal_Int_7QNone_Int_1_onehotd = 4'd0;
  assign _89_d = {lizzieLet17_5QVal_Int_7QNone_Int_1_d[66:1],
                  lizzieLet17_5QVal_Int_7QNone_Int_1_onehotd[0]};
  assign lizzieLet17_5QVal_Int_7QNone_Int_1QVal_Int_d = {lizzieLet17_5QVal_Int_7QNone_Int_1_d[66:1],
                                                         lizzieLet17_5QVal_Int_7QNone_Int_1_onehotd[1]};
  assign _88_d = {lizzieLet17_5QVal_Int_7QNone_Int_1_d[66:1],
                  lizzieLet17_5QVal_Int_7QNone_Int_1_onehotd[2]};
  assign _87_d = {lizzieLet17_5QVal_Int_7QNone_Int_1_d[66:1],
                  lizzieLet17_5QVal_Int_7QNone_Int_1_onehotd[3]};
  assign lizzieLet17_5QVal_Int_7QNone_Int_1_r = (| (lizzieLet17_5QVal_Int_7QNone_Int_1_onehotd & {_87_r,
                                                                                                  _88_r,
                                                                                                  lizzieLet17_5QVal_Int_7QNone_Int_1QVal_Int_r,
                                                                                                  _89_r}));
  assign lizzieLet17_5QVal_Int_7QNone_Int_2_r = lizzieLet17_5QVal_Int_7QNone_Int_1_r;
  
  /* demux (Ty QTree_Int,
       Ty Int) : (lizzieLet17_5QVal_Int_7QNone_Int_3,QTree_Int) (lizzieLet17_5QVal_Int_10QNone_Int,Int) > [(_86,Int),
                                                                                                           (lizzieLet17_5QVal_Int_7QNone_Int_3QVal_Int,Int),
                                                                                                           (_85,Int),
                                                                                                           (_84,Int)] */
  logic [3:0] lizzieLet17_5QVal_Int_10QNone_Int_onehotd;
  always_comb
    if ((lizzieLet17_5QVal_Int_7QNone_Int_3_d[0] && lizzieLet17_5QVal_Int_10QNone_Int_d[0]))
      unique case (lizzieLet17_5QVal_Int_7QNone_Int_3_d[2:1])
        2'd0: lizzieLet17_5QVal_Int_10QNone_Int_onehotd = 4'd1;
        2'd1: lizzieLet17_5QVal_Int_10QNone_Int_onehotd = 4'd2;
        2'd2: lizzieLet17_5QVal_Int_10QNone_Int_onehotd = 4'd4;
        2'd3: lizzieLet17_5QVal_Int_10QNone_Int_onehotd = 4'd8;
        default: lizzieLet17_5QVal_Int_10QNone_Int_onehotd = 4'd0;
      endcase
    else lizzieLet17_5QVal_Int_10QNone_Int_onehotd = 4'd0;
  assign _86_d = {lizzieLet17_5QVal_Int_10QNone_Int_d[32:1],
                  lizzieLet17_5QVal_Int_10QNone_Int_onehotd[0]};
  assign lizzieLet17_5QVal_Int_7QNone_Int_3QVal_Int_d = {lizzieLet17_5QVal_Int_10QNone_Int_d[32:1],
                                                         lizzieLet17_5QVal_Int_10QNone_Int_onehotd[1]};
  assign _85_d = {lizzieLet17_5QVal_Int_10QNone_Int_d[32:1],
                  lizzieLet17_5QVal_Int_10QNone_Int_onehotd[2]};
  assign _84_d = {lizzieLet17_5QVal_Int_10QNone_Int_d[32:1],
                  lizzieLet17_5QVal_Int_10QNone_Int_onehotd[3]};
  assign lizzieLet17_5QVal_Int_10QNone_Int_r = (| (lizzieLet17_5QVal_Int_10QNone_Int_onehotd & {_84_r,
                                                                                                _85_r,
                                                                                                lizzieLet17_5QVal_Int_7QNone_Int_3QVal_Int_r,
                                                                                                _86_r}));
  assign lizzieLet17_5QVal_Int_7QNone_Int_3_r = lizzieLet17_5QVal_Int_10QNone_Int_r;
  
  /* fork (Ty Int) : (lizzieLet17_5QVal_Int_7QNone_Int_3QVal_Int,Int) > [(lizzieLet17_5QVal_Int_7QNone_Int_3QVal_Int_1,Int),
                                                                    (lizzieLet17_5QVal_Int_7QNone_Int_3QVal_Int_2,Int)] */
  logic [1:0] lizzieLet17_5QVal_Int_7QNone_Int_3QVal_Int_emitted;
  logic [1:0] lizzieLet17_5QVal_Int_7QNone_Int_3QVal_Int_done;
  assign lizzieLet17_5QVal_Int_7QNone_Int_3QVal_Int_1_d = {lizzieLet17_5QVal_Int_7QNone_Int_3QVal_Int_d[32:1],
                                                           (lizzieLet17_5QVal_Int_7QNone_Int_3QVal_Int_d[0] && (! lizzieLet17_5QVal_Int_7QNone_Int_3QVal_Int_emitted[0]))};
  assign lizzieLet17_5QVal_Int_7QNone_Int_3QVal_Int_2_d = {lizzieLet17_5QVal_Int_7QNone_Int_3QVal_Int_d[32:1],
                                                           (lizzieLet17_5QVal_Int_7QNone_Int_3QVal_Int_d[0] && (! lizzieLet17_5QVal_Int_7QNone_Int_3QVal_Int_emitted[1]))};
  assign lizzieLet17_5QVal_Int_7QNone_Int_3QVal_Int_done = (lizzieLet17_5QVal_Int_7QNone_Int_3QVal_Int_emitted | ({lizzieLet17_5QVal_Int_7QNone_Int_3QVal_Int_2_d[0],
                                                                                                                   lizzieLet17_5QVal_Int_7QNone_Int_3QVal_Int_1_d[0]} & {lizzieLet17_5QVal_Int_7QNone_Int_3QVal_Int_2_r,
                                                                                                                                                                         lizzieLet17_5QVal_Int_7QNone_Int_3QVal_Int_1_r}));
  assign lizzieLet17_5QVal_Int_7QNone_Int_3QVal_Int_r = (& lizzieLet17_5QVal_Int_7QNone_Int_3QVal_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QVal_Int_7QNone_Int_3QVal_Int_emitted <= 2'd0;
    else
      lizzieLet17_5QVal_Int_7QNone_Int_3QVal_Int_emitted <= (lizzieLet17_5QVal_Int_7QNone_Int_3QVal_Int_r ? 2'd0 :
                                                             lizzieLet17_5QVal_Int_7QNone_Int_3QVal_Int_done);
  
  /* buf (Ty Int) : (lizzieLet17_5QVal_Int_7QNone_Int_3QVal_Int_1,Int) > (lizzieLet17_5QVal_Int_7QNone_Int_3QVal_Int_1_argbuf,Int) */
  Int_t lizzieLet17_5QVal_Int_7QNone_Int_3QVal_Int_1_bufchan_d;
  logic lizzieLet17_5QVal_Int_7QNone_Int_3QVal_Int_1_bufchan_r;
  assign lizzieLet17_5QVal_Int_7QNone_Int_3QVal_Int_1_r = ((! lizzieLet17_5QVal_Int_7QNone_Int_3QVal_Int_1_bufchan_d[0]) || lizzieLet17_5QVal_Int_7QNone_Int_3QVal_Int_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QVal_Int_7QNone_Int_3QVal_Int_1_bufchan_d <= {32'd0,
                                                                 1'd0};
    else
      if (lizzieLet17_5QVal_Int_7QNone_Int_3QVal_Int_1_r)
        lizzieLet17_5QVal_Int_7QNone_Int_3QVal_Int_1_bufchan_d <= lizzieLet17_5QVal_Int_7QNone_Int_3QVal_Int_1_d;
  Int_t lizzieLet17_5QVal_Int_7QNone_Int_3QVal_Int_1_bufchan_buf;
  assign lizzieLet17_5QVal_Int_7QNone_Int_3QVal_Int_1_bufchan_r = (! lizzieLet17_5QVal_Int_7QNone_Int_3QVal_Int_1_bufchan_buf[0]);
  assign lizzieLet17_5QVal_Int_7QNone_Int_3QVal_Int_1_argbuf_d = (lizzieLet17_5QVal_Int_7QNone_Int_3QVal_Int_1_bufchan_buf[0] ? lizzieLet17_5QVal_Int_7QNone_Int_3QVal_Int_1_bufchan_buf :
                                                                  lizzieLet17_5QVal_Int_7QNone_Int_3QVal_Int_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QVal_Int_7QNone_Int_3QVal_Int_1_bufchan_buf <= {32'd0,
                                                                   1'd0};
    else
      if ((lizzieLet17_5QVal_Int_7QNone_Int_3QVal_Int_1_argbuf_r && lizzieLet17_5QVal_Int_7QNone_Int_3QVal_Int_1_bufchan_buf[0]))
        lizzieLet17_5QVal_Int_7QNone_Int_3QVal_Int_1_bufchan_buf <= {32'd0,
                                                                     1'd0};
      else if (((! lizzieLet17_5QVal_Int_7QNone_Int_3QVal_Int_1_argbuf_r) && (! lizzieLet17_5QVal_Int_7QNone_Int_3QVal_Int_1_bufchan_buf[0])))
        lizzieLet17_5QVal_Int_7QNone_Int_3QVal_Int_1_bufchan_buf <= lizzieLet17_5QVal_Int_7QNone_Int_3QVal_Int_1_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty MyDTInt_Int_Int) : (lizzieLet17_5QVal_Int_7QNone_Int_4,QTree_Int) (lizzieLet17_5QVal_Int_3QNone_Int,MyDTInt_Int_Int) > [(_83,MyDTInt_Int_Int),
                                                                                                                                  (lizzieLet17_5QVal_Int_7QNone_Int_4QVal_Int,MyDTInt_Int_Int),
                                                                                                                                  (_82,MyDTInt_Int_Int),
                                                                                                                                  (_81,MyDTInt_Int_Int)] */
  logic [3:0] lizzieLet17_5QVal_Int_3QNone_Int_onehotd;
  always_comb
    if ((lizzieLet17_5QVal_Int_7QNone_Int_4_d[0] && lizzieLet17_5QVal_Int_3QNone_Int_d[0]))
      unique case (lizzieLet17_5QVal_Int_7QNone_Int_4_d[2:1])
        2'd0: lizzieLet17_5QVal_Int_3QNone_Int_onehotd = 4'd1;
        2'd1: lizzieLet17_5QVal_Int_3QNone_Int_onehotd = 4'd2;
        2'd2: lizzieLet17_5QVal_Int_3QNone_Int_onehotd = 4'd4;
        2'd3: lizzieLet17_5QVal_Int_3QNone_Int_onehotd = 4'd8;
        default: lizzieLet17_5QVal_Int_3QNone_Int_onehotd = 4'd0;
      endcase
    else lizzieLet17_5QVal_Int_3QNone_Int_onehotd = 4'd0;
  assign _83_d = lizzieLet17_5QVal_Int_3QNone_Int_onehotd[0];
  assign lizzieLet17_5QVal_Int_7QNone_Int_4QVal_Int_d = lizzieLet17_5QVal_Int_3QNone_Int_onehotd[1];
  assign _82_d = lizzieLet17_5QVal_Int_3QNone_Int_onehotd[2];
  assign _81_d = lizzieLet17_5QVal_Int_3QNone_Int_onehotd[3];
  assign lizzieLet17_5QVal_Int_3QNone_Int_r = (| (lizzieLet17_5QVal_Int_3QNone_Int_onehotd & {_81_r,
                                                                                              _82_r,
                                                                                              lizzieLet17_5QVal_Int_7QNone_Int_4QVal_Int_r,
                                                                                              _83_r}));
  assign lizzieLet17_5QVal_Int_7QNone_Int_4_r = lizzieLet17_5QVal_Int_3QNone_Int_r;
  
  /* fork (Ty MyDTInt_Int_Int) : (lizzieLet17_5QVal_Int_7QNone_Int_4QVal_Int,MyDTInt_Int_Int) > [(lizzieLet17_5QVal_Int_7QNone_Int_4QVal_Int_1,MyDTInt_Int_Int),
                                                                                            (lizzieLet17_5QVal_Int_7QNone_Int_4QVal_Int_2,MyDTInt_Int_Int)] */
  logic [1:0] lizzieLet17_5QVal_Int_7QNone_Int_4QVal_Int_emitted;
  logic [1:0] lizzieLet17_5QVal_Int_7QNone_Int_4QVal_Int_done;
  assign lizzieLet17_5QVal_Int_7QNone_Int_4QVal_Int_1_d = (lizzieLet17_5QVal_Int_7QNone_Int_4QVal_Int_d[0] && (! lizzieLet17_5QVal_Int_7QNone_Int_4QVal_Int_emitted[0]));
  assign lizzieLet17_5QVal_Int_7QNone_Int_4QVal_Int_2_d = (lizzieLet17_5QVal_Int_7QNone_Int_4QVal_Int_d[0] && (! lizzieLet17_5QVal_Int_7QNone_Int_4QVal_Int_emitted[1]));
  assign lizzieLet17_5QVal_Int_7QNone_Int_4QVal_Int_done = (lizzieLet17_5QVal_Int_7QNone_Int_4QVal_Int_emitted | ({lizzieLet17_5QVal_Int_7QNone_Int_4QVal_Int_2_d[0],
                                                                                                                   lizzieLet17_5QVal_Int_7QNone_Int_4QVal_Int_1_d[0]} & {lizzieLet17_5QVal_Int_7QNone_Int_4QVal_Int_2_r,
                                                                                                                                                                         lizzieLet17_5QVal_Int_7QNone_Int_4QVal_Int_1_r}));
  assign lizzieLet17_5QVal_Int_7QNone_Int_4QVal_Int_r = (& lizzieLet17_5QVal_Int_7QNone_Int_4QVal_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QVal_Int_7QNone_Int_4QVal_Int_emitted <= 2'd0;
    else
      lizzieLet17_5QVal_Int_7QNone_Int_4QVal_Int_emitted <= (lizzieLet17_5QVal_Int_7QNone_Int_4QVal_Int_r ? 2'd0 :
                                                             lizzieLet17_5QVal_Int_7QNone_Int_4QVal_Int_done);
  
  /* buf (Ty MyDTInt_Int_Int) : (lizzieLet17_5QVal_Int_7QNone_Int_4QVal_Int_1,MyDTInt_Int_Int) > (lizzieLet17_5QVal_Int_7QNone_Int_4QVal_Int_1_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t lizzieLet17_5QVal_Int_7QNone_Int_4QVal_Int_1_bufchan_d;
  logic lizzieLet17_5QVal_Int_7QNone_Int_4QVal_Int_1_bufchan_r;
  assign lizzieLet17_5QVal_Int_7QNone_Int_4QVal_Int_1_r = ((! lizzieLet17_5QVal_Int_7QNone_Int_4QVal_Int_1_bufchan_d[0]) || lizzieLet17_5QVal_Int_7QNone_Int_4QVal_Int_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QVal_Int_7QNone_Int_4QVal_Int_1_bufchan_d <= 1'd0;
    else
      if (lizzieLet17_5QVal_Int_7QNone_Int_4QVal_Int_1_r)
        lizzieLet17_5QVal_Int_7QNone_Int_4QVal_Int_1_bufchan_d <= lizzieLet17_5QVal_Int_7QNone_Int_4QVal_Int_1_d;
  MyDTInt_Int_Int_t lizzieLet17_5QVal_Int_7QNone_Int_4QVal_Int_1_bufchan_buf;
  assign lizzieLet17_5QVal_Int_7QNone_Int_4QVal_Int_1_bufchan_r = (! lizzieLet17_5QVal_Int_7QNone_Int_4QVal_Int_1_bufchan_buf[0]);
  assign lizzieLet17_5QVal_Int_7QNone_Int_4QVal_Int_1_argbuf_d = (lizzieLet17_5QVal_Int_7QNone_Int_4QVal_Int_1_bufchan_buf[0] ? lizzieLet17_5QVal_Int_7QNone_Int_4QVal_Int_1_bufchan_buf :
                                                                  lizzieLet17_5QVal_Int_7QNone_Int_4QVal_Int_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QVal_Int_7QNone_Int_4QVal_Int_1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet17_5QVal_Int_7QNone_Int_4QVal_Int_1_argbuf_r && lizzieLet17_5QVal_Int_7QNone_Int_4QVal_Int_1_bufchan_buf[0]))
        lizzieLet17_5QVal_Int_7QNone_Int_4QVal_Int_1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet17_5QVal_Int_7QNone_Int_4QVal_Int_1_argbuf_r) && (! lizzieLet17_5QVal_Int_7QNone_Int_4QVal_Int_1_bufchan_buf[0])))
        lizzieLet17_5QVal_Int_7QNone_Int_4QVal_Int_1_bufchan_buf <= lizzieLet17_5QVal_Int_7QNone_Int_4QVal_Int_1_bufchan_d;
  
  /* dcon (Ty TupMyDTInt_Int_Int___Int___Int,
      Dcon TupMyDTInt_Int_Int___Int___Int) : [(lizzieLet17_5QVal_Int_7QNone_Int_4QVal_Int_1_argbuf,MyDTInt_Int_Int),
                                              (lizzieLet17_5QVal_Int_7QNone_Int_3QVal_Int_1_argbuf,Int),
                                              (vaeL_1_argbuf,Int)] > (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int5,TupMyDTInt_Int_Int___Int___Int) */
  assign applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int5_d = TupMyDTInt_Int_Int___Int___Int_dc((& {lizzieLet17_5QVal_Int_7QNone_Int_4QVal_Int_1_argbuf_d[0],
                                                                                                       lizzieLet17_5QVal_Int_7QNone_Int_3QVal_Int_1_argbuf_d[0],
                                                                                                       vaeL_1_argbuf_d[0]}), lizzieLet17_5QVal_Int_7QNone_Int_4QVal_Int_1_argbuf_d, lizzieLet17_5QVal_Int_7QNone_Int_3QVal_Int_1_argbuf_d, vaeL_1_argbuf_d);
  assign {lizzieLet17_5QVal_Int_7QNone_Int_4QVal_Int_1_argbuf_r,
          lizzieLet17_5QVal_Int_7QNone_Int_3QVal_Int_1_argbuf_r,
          vaeL_1_argbuf_r} = {3 {(applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int5_r && applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int5_d[0])}};
  
  /* demux (Ty QTree_Int,
       Ty Pointer_CTf_f_Int) : (lizzieLet17_5QVal_Int_7QNone_Int_5,QTree_Int) (lizzieLet17_5QVal_Int_4QNone_Int,Pointer_CTf_f_Int) > [(lizzieLet17_5QVal_Int_7QNone_Int_5QNone_Int,Pointer_CTf_f_Int),
                                                                                                                                      (lizzieLet17_5QVal_Int_7QNone_Int_5QVal_Int,Pointer_CTf_f_Int),
                                                                                                                                      (lizzieLet17_5QVal_Int_7QNone_Int_5QNode_Int,Pointer_CTf_f_Int),
                                                                                                                                      (lizzieLet17_5QVal_Int_7QNone_Int_5QError_Int,Pointer_CTf_f_Int)] */
  logic [3:0] lizzieLet17_5QVal_Int_4QNone_Int_onehotd;
  always_comb
    if ((lizzieLet17_5QVal_Int_7QNone_Int_5_d[0] && lizzieLet17_5QVal_Int_4QNone_Int_d[0]))
      unique case (lizzieLet17_5QVal_Int_7QNone_Int_5_d[2:1])
        2'd0: lizzieLet17_5QVal_Int_4QNone_Int_onehotd = 4'd1;
        2'd1: lizzieLet17_5QVal_Int_4QNone_Int_onehotd = 4'd2;
        2'd2: lizzieLet17_5QVal_Int_4QNone_Int_onehotd = 4'd4;
        2'd3: lizzieLet17_5QVal_Int_4QNone_Int_onehotd = 4'd8;
        default: lizzieLet17_5QVal_Int_4QNone_Int_onehotd = 4'd0;
      endcase
    else lizzieLet17_5QVal_Int_4QNone_Int_onehotd = 4'd0;
  assign lizzieLet17_5QVal_Int_7QNone_Int_5QNone_Int_d = {lizzieLet17_5QVal_Int_4QNone_Int_d[16:1],
                                                          lizzieLet17_5QVal_Int_4QNone_Int_onehotd[0]};
  assign lizzieLet17_5QVal_Int_7QNone_Int_5QVal_Int_d = {lizzieLet17_5QVal_Int_4QNone_Int_d[16:1],
                                                         lizzieLet17_5QVal_Int_4QNone_Int_onehotd[1]};
  assign lizzieLet17_5QVal_Int_7QNone_Int_5QNode_Int_d = {lizzieLet17_5QVal_Int_4QNone_Int_d[16:1],
                                                          lizzieLet17_5QVal_Int_4QNone_Int_onehotd[2]};
  assign lizzieLet17_5QVal_Int_7QNone_Int_5QError_Int_d = {lizzieLet17_5QVal_Int_4QNone_Int_d[16:1],
                                                           lizzieLet17_5QVal_Int_4QNone_Int_onehotd[3]};
  assign lizzieLet17_5QVal_Int_4QNone_Int_r = (| (lizzieLet17_5QVal_Int_4QNone_Int_onehotd & {lizzieLet17_5QVal_Int_7QNone_Int_5QError_Int_r,
                                                                                              lizzieLet17_5QVal_Int_7QNone_Int_5QNode_Int_r,
                                                                                              lizzieLet17_5QVal_Int_7QNone_Int_5QVal_Int_r,
                                                                                              lizzieLet17_5QVal_Int_7QNone_Int_5QNone_Int_r}));
  assign lizzieLet17_5QVal_Int_7QNone_Int_5_r = lizzieLet17_5QVal_Int_4QNone_Int_r;
  
  /* buf (Ty Pointer_CTf_f_Int) : (lizzieLet17_5QVal_Int_7QNone_Int_5QError_Int,Pointer_CTf_f_Int) > (lizzieLet17_5QVal_Int_7QNone_Int_5QError_Int_1_argbuf,Pointer_CTf_f_Int) */
  Pointer_CTf_f_Int_t lizzieLet17_5QVal_Int_7QNone_Int_5QError_Int_bufchan_d;
  logic lizzieLet17_5QVal_Int_7QNone_Int_5QError_Int_bufchan_r;
  assign lizzieLet17_5QVal_Int_7QNone_Int_5QError_Int_r = ((! lizzieLet17_5QVal_Int_7QNone_Int_5QError_Int_bufchan_d[0]) || lizzieLet17_5QVal_Int_7QNone_Int_5QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QVal_Int_7QNone_Int_5QError_Int_bufchan_d <= {16'd0,
                                                                 1'd0};
    else
      if (lizzieLet17_5QVal_Int_7QNone_Int_5QError_Int_r)
        lizzieLet17_5QVal_Int_7QNone_Int_5QError_Int_bufchan_d <= lizzieLet17_5QVal_Int_7QNone_Int_5QError_Int_d;
  Pointer_CTf_f_Int_t lizzieLet17_5QVal_Int_7QNone_Int_5QError_Int_bufchan_buf;
  assign lizzieLet17_5QVal_Int_7QNone_Int_5QError_Int_bufchan_r = (! lizzieLet17_5QVal_Int_7QNone_Int_5QError_Int_bufchan_buf[0]);
  assign lizzieLet17_5QVal_Int_7QNone_Int_5QError_Int_1_argbuf_d = (lizzieLet17_5QVal_Int_7QNone_Int_5QError_Int_bufchan_buf[0] ? lizzieLet17_5QVal_Int_7QNone_Int_5QError_Int_bufchan_buf :
                                                                    lizzieLet17_5QVal_Int_7QNone_Int_5QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QVal_Int_7QNone_Int_5QError_Int_bufchan_buf <= {16'd0,
                                                                   1'd0};
    else
      if ((lizzieLet17_5QVal_Int_7QNone_Int_5QError_Int_1_argbuf_r && lizzieLet17_5QVal_Int_7QNone_Int_5QError_Int_bufchan_buf[0]))
        lizzieLet17_5QVal_Int_7QNone_Int_5QError_Int_bufchan_buf <= {16'd0,
                                                                     1'd0};
      else if (((! lizzieLet17_5QVal_Int_7QNone_Int_5QError_Int_1_argbuf_r) && (! lizzieLet17_5QVal_Int_7QNone_Int_5QError_Int_bufchan_buf[0])))
        lizzieLet17_5QVal_Int_7QNone_Int_5QError_Int_bufchan_buf <= lizzieLet17_5QVal_Int_7QNone_Int_5QError_Int_bufchan_d;
  
  /* buf (Ty Pointer_CTf_f_Int) : (lizzieLet17_5QVal_Int_7QNone_Int_5QNode_Int,Pointer_CTf_f_Int) > (lizzieLet17_5QVal_Int_7QNone_Int_5QNode_Int_1_argbuf,Pointer_CTf_f_Int) */
  Pointer_CTf_f_Int_t lizzieLet17_5QVal_Int_7QNone_Int_5QNode_Int_bufchan_d;
  logic lizzieLet17_5QVal_Int_7QNone_Int_5QNode_Int_bufchan_r;
  assign lizzieLet17_5QVal_Int_7QNone_Int_5QNode_Int_r = ((! lizzieLet17_5QVal_Int_7QNone_Int_5QNode_Int_bufchan_d[0]) || lizzieLet17_5QVal_Int_7QNone_Int_5QNode_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QVal_Int_7QNone_Int_5QNode_Int_bufchan_d <= {16'd0,
                                                                1'd0};
    else
      if (lizzieLet17_5QVal_Int_7QNone_Int_5QNode_Int_r)
        lizzieLet17_5QVal_Int_7QNone_Int_5QNode_Int_bufchan_d <= lizzieLet17_5QVal_Int_7QNone_Int_5QNode_Int_d;
  Pointer_CTf_f_Int_t lizzieLet17_5QVal_Int_7QNone_Int_5QNode_Int_bufchan_buf;
  assign lizzieLet17_5QVal_Int_7QNone_Int_5QNode_Int_bufchan_r = (! lizzieLet17_5QVal_Int_7QNone_Int_5QNode_Int_bufchan_buf[0]);
  assign lizzieLet17_5QVal_Int_7QNone_Int_5QNode_Int_1_argbuf_d = (lizzieLet17_5QVal_Int_7QNone_Int_5QNode_Int_bufchan_buf[0] ? lizzieLet17_5QVal_Int_7QNone_Int_5QNode_Int_bufchan_buf :
                                                                   lizzieLet17_5QVal_Int_7QNone_Int_5QNode_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QVal_Int_7QNone_Int_5QNode_Int_bufchan_buf <= {16'd0,
                                                                  1'd0};
    else
      if ((lizzieLet17_5QVal_Int_7QNone_Int_5QNode_Int_1_argbuf_r && lizzieLet17_5QVal_Int_7QNone_Int_5QNode_Int_bufchan_buf[0]))
        lizzieLet17_5QVal_Int_7QNone_Int_5QNode_Int_bufchan_buf <= {16'd0,
                                                                    1'd0};
      else if (((! lizzieLet17_5QVal_Int_7QNone_Int_5QNode_Int_1_argbuf_r) && (! lizzieLet17_5QVal_Int_7QNone_Int_5QNode_Int_bufchan_buf[0])))
        lizzieLet17_5QVal_Int_7QNone_Int_5QNode_Int_bufchan_buf <= lizzieLet17_5QVal_Int_7QNone_Int_5QNode_Int_bufchan_d;
  
  /* buf (Ty Pointer_CTf_f_Int) : (lizzieLet17_5QVal_Int_7QNone_Int_5QNone_Int,Pointer_CTf_f_Int) > (lizzieLet17_5QVal_Int_7QNone_Int_5QNone_Int_1_argbuf,Pointer_CTf_f_Int) */
  Pointer_CTf_f_Int_t lizzieLet17_5QVal_Int_7QNone_Int_5QNone_Int_bufchan_d;
  logic lizzieLet17_5QVal_Int_7QNone_Int_5QNone_Int_bufchan_r;
  assign lizzieLet17_5QVal_Int_7QNone_Int_5QNone_Int_r = ((! lizzieLet17_5QVal_Int_7QNone_Int_5QNone_Int_bufchan_d[0]) || lizzieLet17_5QVal_Int_7QNone_Int_5QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QVal_Int_7QNone_Int_5QNone_Int_bufchan_d <= {16'd0,
                                                                1'd0};
    else
      if (lizzieLet17_5QVal_Int_7QNone_Int_5QNone_Int_r)
        lizzieLet17_5QVal_Int_7QNone_Int_5QNone_Int_bufchan_d <= lizzieLet17_5QVal_Int_7QNone_Int_5QNone_Int_d;
  Pointer_CTf_f_Int_t lizzieLet17_5QVal_Int_7QNone_Int_5QNone_Int_bufchan_buf;
  assign lizzieLet17_5QVal_Int_7QNone_Int_5QNone_Int_bufchan_r = (! lizzieLet17_5QVal_Int_7QNone_Int_5QNone_Int_bufchan_buf[0]);
  assign lizzieLet17_5QVal_Int_7QNone_Int_5QNone_Int_1_argbuf_d = (lizzieLet17_5QVal_Int_7QNone_Int_5QNone_Int_bufchan_buf[0] ? lizzieLet17_5QVal_Int_7QNone_Int_5QNone_Int_bufchan_buf :
                                                                   lizzieLet17_5QVal_Int_7QNone_Int_5QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QVal_Int_7QNone_Int_5QNone_Int_bufchan_buf <= {16'd0,
                                                                  1'd0};
    else
      if ((lizzieLet17_5QVal_Int_7QNone_Int_5QNone_Int_1_argbuf_r && lizzieLet17_5QVal_Int_7QNone_Int_5QNone_Int_bufchan_buf[0]))
        lizzieLet17_5QVal_Int_7QNone_Int_5QNone_Int_bufchan_buf <= {16'd0,
                                                                    1'd0};
      else if (((! lizzieLet17_5QVal_Int_7QNone_Int_5QNone_Int_1_argbuf_r) && (! lizzieLet17_5QVal_Int_7QNone_Int_5QNone_Int_bufchan_buf[0])))
        lizzieLet17_5QVal_Int_7QNone_Int_5QNone_Int_bufchan_buf <= lizzieLet17_5QVal_Int_7QNone_Int_5QNone_Int_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Go) : (lizzieLet17_5QVal_Int_7QNone_Int_6,QTree_Int) (lizzieLet17_5QVal_Int_5QNone_Int,Go) > [(lizzieLet17_5QVal_Int_7QNone_Int_6QNone_Int,Go),
                                                                                                        (lizzieLet17_5QVal_Int_7QNone_Int_6QVal_Int,Go),
                                                                                                        (lizzieLet17_5QVal_Int_7QNone_Int_6QNode_Int,Go),
                                                                                                        (lizzieLet17_5QVal_Int_7QNone_Int_6QError_Int,Go)] */
  logic [3:0] lizzieLet17_5QVal_Int_5QNone_Int_onehotd;
  always_comb
    if ((lizzieLet17_5QVal_Int_7QNone_Int_6_d[0] && lizzieLet17_5QVal_Int_5QNone_Int_d[0]))
      unique case (lizzieLet17_5QVal_Int_7QNone_Int_6_d[2:1])
        2'd0: lizzieLet17_5QVal_Int_5QNone_Int_onehotd = 4'd1;
        2'd1: lizzieLet17_5QVal_Int_5QNone_Int_onehotd = 4'd2;
        2'd2: lizzieLet17_5QVal_Int_5QNone_Int_onehotd = 4'd4;
        2'd3: lizzieLet17_5QVal_Int_5QNone_Int_onehotd = 4'd8;
        default: lizzieLet17_5QVal_Int_5QNone_Int_onehotd = 4'd0;
      endcase
    else lizzieLet17_5QVal_Int_5QNone_Int_onehotd = 4'd0;
  assign lizzieLet17_5QVal_Int_7QNone_Int_6QNone_Int_d = lizzieLet17_5QVal_Int_5QNone_Int_onehotd[0];
  assign lizzieLet17_5QVal_Int_7QNone_Int_6QVal_Int_d = lizzieLet17_5QVal_Int_5QNone_Int_onehotd[1];
  assign lizzieLet17_5QVal_Int_7QNone_Int_6QNode_Int_d = lizzieLet17_5QVal_Int_5QNone_Int_onehotd[2];
  assign lizzieLet17_5QVal_Int_7QNone_Int_6QError_Int_d = lizzieLet17_5QVal_Int_5QNone_Int_onehotd[3];
  assign lizzieLet17_5QVal_Int_5QNone_Int_r = (| (lizzieLet17_5QVal_Int_5QNone_Int_onehotd & {lizzieLet17_5QVal_Int_7QNone_Int_6QError_Int_r,
                                                                                              lizzieLet17_5QVal_Int_7QNone_Int_6QNode_Int_r,
                                                                                              lizzieLet17_5QVal_Int_7QNone_Int_6QVal_Int_r,
                                                                                              lizzieLet17_5QVal_Int_7QNone_Int_6QNone_Int_r}));
  assign lizzieLet17_5QVal_Int_7QNone_Int_6_r = lizzieLet17_5QVal_Int_5QNone_Int_r;
  
  /* fork (Ty Go) : (lizzieLet17_5QVal_Int_7QNone_Int_6QError_Int,Go) > [(lizzieLet17_5QVal_Int_7QNone_Int_6QError_Int_1,Go),
                                                                    (lizzieLet17_5QVal_Int_7QNone_Int_6QError_Int_2,Go)] */
  logic [1:0] lizzieLet17_5QVal_Int_7QNone_Int_6QError_Int_emitted;
  logic [1:0] lizzieLet17_5QVal_Int_7QNone_Int_6QError_Int_done;
  assign lizzieLet17_5QVal_Int_7QNone_Int_6QError_Int_1_d = (lizzieLet17_5QVal_Int_7QNone_Int_6QError_Int_d[0] && (! lizzieLet17_5QVal_Int_7QNone_Int_6QError_Int_emitted[0]));
  assign lizzieLet17_5QVal_Int_7QNone_Int_6QError_Int_2_d = (lizzieLet17_5QVal_Int_7QNone_Int_6QError_Int_d[0] && (! lizzieLet17_5QVal_Int_7QNone_Int_6QError_Int_emitted[1]));
  assign lizzieLet17_5QVal_Int_7QNone_Int_6QError_Int_done = (lizzieLet17_5QVal_Int_7QNone_Int_6QError_Int_emitted | ({lizzieLet17_5QVal_Int_7QNone_Int_6QError_Int_2_d[0],
                                                                                                                       lizzieLet17_5QVal_Int_7QNone_Int_6QError_Int_1_d[0]} & {lizzieLet17_5QVal_Int_7QNone_Int_6QError_Int_2_r,
                                                                                                                                                                               lizzieLet17_5QVal_Int_7QNone_Int_6QError_Int_1_r}));
  assign lizzieLet17_5QVal_Int_7QNone_Int_6QError_Int_r = (& lizzieLet17_5QVal_Int_7QNone_Int_6QError_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QVal_Int_7QNone_Int_6QError_Int_emitted <= 2'd0;
    else
      lizzieLet17_5QVal_Int_7QNone_Int_6QError_Int_emitted <= (lizzieLet17_5QVal_Int_7QNone_Int_6QError_Int_r ? 2'd0 :
                                                               lizzieLet17_5QVal_Int_7QNone_Int_6QError_Int_done);
  
  /* dcon (Ty QTree_Int,
      Dcon QError_Int) : [(lizzieLet17_5QVal_Int_7QNone_Int_6QError_Int_1,Go)] > (lizzieLet17_5QVal_Int_7QNone_Int_6QError_Int_1QError_Int,QTree_Int) */
  assign lizzieLet17_5QVal_Int_7QNone_Int_6QError_Int_1QError_Int_d = QError_Int_dc((& {lizzieLet17_5QVal_Int_7QNone_Int_6QError_Int_1_d[0]}), lizzieLet17_5QVal_Int_7QNone_Int_6QError_Int_1_d);
  assign {lizzieLet17_5QVal_Int_7QNone_Int_6QError_Int_1_r} = {1 {(lizzieLet17_5QVal_Int_7QNone_Int_6QError_Int_1QError_Int_r && lizzieLet17_5QVal_Int_7QNone_Int_6QError_Int_1QError_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (lizzieLet17_5QVal_Int_7QNone_Int_6QError_Int_1QError_Int,QTree_Int) > (lizzieLet34_1_argbuf,QTree_Int) */
  QTree_Int_t lizzieLet17_5QVal_Int_7QNone_Int_6QError_Int_1QError_Int_bufchan_d;
  logic lizzieLet17_5QVal_Int_7QNone_Int_6QError_Int_1QError_Int_bufchan_r;
  assign lizzieLet17_5QVal_Int_7QNone_Int_6QError_Int_1QError_Int_r = ((! lizzieLet17_5QVal_Int_7QNone_Int_6QError_Int_1QError_Int_bufchan_d[0]) || lizzieLet17_5QVal_Int_7QNone_Int_6QError_Int_1QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QVal_Int_7QNone_Int_6QError_Int_1QError_Int_bufchan_d <= {66'd0,
                                                                             1'd0};
    else
      if (lizzieLet17_5QVal_Int_7QNone_Int_6QError_Int_1QError_Int_r)
        lizzieLet17_5QVal_Int_7QNone_Int_6QError_Int_1QError_Int_bufchan_d <= lizzieLet17_5QVal_Int_7QNone_Int_6QError_Int_1QError_Int_d;
  QTree_Int_t lizzieLet17_5QVal_Int_7QNone_Int_6QError_Int_1QError_Int_bufchan_buf;
  assign lizzieLet17_5QVal_Int_7QNone_Int_6QError_Int_1QError_Int_bufchan_r = (! lizzieLet17_5QVal_Int_7QNone_Int_6QError_Int_1QError_Int_bufchan_buf[0]);
  assign lizzieLet34_1_argbuf_d = (lizzieLet17_5QVal_Int_7QNone_Int_6QError_Int_1QError_Int_bufchan_buf[0] ? lizzieLet17_5QVal_Int_7QNone_Int_6QError_Int_1QError_Int_bufchan_buf :
                                   lizzieLet17_5QVal_Int_7QNone_Int_6QError_Int_1QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QVal_Int_7QNone_Int_6QError_Int_1QError_Int_bufchan_buf <= {66'd0,
                                                                               1'd0};
    else
      if ((lizzieLet34_1_argbuf_r && lizzieLet17_5QVal_Int_7QNone_Int_6QError_Int_1QError_Int_bufchan_buf[0]))
        lizzieLet17_5QVal_Int_7QNone_Int_6QError_Int_1QError_Int_bufchan_buf <= {66'd0,
                                                                                 1'd0};
      else if (((! lizzieLet34_1_argbuf_r) && (! lizzieLet17_5QVal_Int_7QNone_Int_6QError_Int_1QError_Int_bufchan_buf[0])))
        lizzieLet17_5QVal_Int_7QNone_Int_6QError_Int_1QError_Int_bufchan_buf <= lizzieLet17_5QVal_Int_7QNone_Int_6QError_Int_1QError_Int_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet17_5QVal_Int_7QNone_Int_6QError_Int_2,Go) > (lizzieLet17_5QVal_Int_7QNone_Int_6QError_Int_2_argbuf,Go) */
  Go_t lizzieLet17_5QVal_Int_7QNone_Int_6QError_Int_2_bufchan_d;
  logic lizzieLet17_5QVal_Int_7QNone_Int_6QError_Int_2_bufchan_r;
  assign lizzieLet17_5QVal_Int_7QNone_Int_6QError_Int_2_r = ((! lizzieLet17_5QVal_Int_7QNone_Int_6QError_Int_2_bufchan_d[0]) || lizzieLet17_5QVal_Int_7QNone_Int_6QError_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QVal_Int_7QNone_Int_6QError_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet17_5QVal_Int_7QNone_Int_6QError_Int_2_r)
        lizzieLet17_5QVal_Int_7QNone_Int_6QError_Int_2_bufchan_d <= lizzieLet17_5QVal_Int_7QNone_Int_6QError_Int_2_d;
  Go_t lizzieLet17_5QVal_Int_7QNone_Int_6QError_Int_2_bufchan_buf;
  assign lizzieLet17_5QVal_Int_7QNone_Int_6QError_Int_2_bufchan_r = (! lizzieLet17_5QVal_Int_7QNone_Int_6QError_Int_2_bufchan_buf[0]);
  assign lizzieLet17_5QVal_Int_7QNone_Int_6QError_Int_2_argbuf_d = (lizzieLet17_5QVal_Int_7QNone_Int_6QError_Int_2_bufchan_buf[0] ? lizzieLet17_5QVal_Int_7QNone_Int_6QError_Int_2_bufchan_buf :
                                                                    lizzieLet17_5QVal_Int_7QNone_Int_6QError_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QVal_Int_7QNone_Int_6QError_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet17_5QVal_Int_7QNone_Int_6QError_Int_2_argbuf_r && lizzieLet17_5QVal_Int_7QNone_Int_6QError_Int_2_bufchan_buf[0]))
        lizzieLet17_5QVal_Int_7QNone_Int_6QError_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet17_5QVal_Int_7QNone_Int_6QError_Int_2_argbuf_r) && (! lizzieLet17_5QVal_Int_7QNone_Int_6QError_Int_2_bufchan_buf[0])))
        lizzieLet17_5QVal_Int_7QNone_Int_6QError_Int_2_bufchan_buf <= lizzieLet17_5QVal_Int_7QNone_Int_6QError_Int_2_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet17_5QVal_Int_7QNone_Int_6QNode_Int,Go) > [(lizzieLet17_5QVal_Int_7QNone_Int_6QNode_Int_1,Go),
                                                                   (lizzieLet17_5QVal_Int_7QNone_Int_6QNode_Int_2,Go)] */
  logic [1:0] lizzieLet17_5QVal_Int_7QNone_Int_6QNode_Int_emitted;
  logic [1:0] lizzieLet17_5QVal_Int_7QNone_Int_6QNode_Int_done;
  assign lizzieLet17_5QVal_Int_7QNone_Int_6QNode_Int_1_d = (lizzieLet17_5QVal_Int_7QNone_Int_6QNode_Int_d[0] && (! lizzieLet17_5QVal_Int_7QNone_Int_6QNode_Int_emitted[0]));
  assign lizzieLet17_5QVal_Int_7QNone_Int_6QNode_Int_2_d = (lizzieLet17_5QVal_Int_7QNone_Int_6QNode_Int_d[0] && (! lizzieLet17_5QVal_Int_7QNone_Int_6QNode_Int_emitted[1]));
  assign lizzieLet17_5QVal_Int_7QNone_Int_6QNode_Int_done = (lizzieLet17_5QVal_Int_7QNone_Int_6QNode_Int_emitted | ({lizzieLet17_5QVal_Int_7QNone_Int_6QNode_Int_2_d[0],
                                                                                                                     lizzieLet17_5QVal_Int_7QNone_Int_6QNode_Int_1_d[0]} & {lizzieLet17_5QVal_Int_7QNone_Int_6QNode_Int_2_r,
                                                                                                                                                                            lizzieLet17_5QVal_Int_7QNone_Int_6QNode_Int_1_r}));
  assign lizzieLet17_5QVal_Int_7QNone_Int_6QNode_Int_r = (& lizzieLet17_5QVal_Int_7QNone_Int_6QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QVal_Int_7QNone_Int_6QNode_Int_emitted <= 2'd0;
    else
      lizzieLet17_5QVal_Int_7QNone_Int_6QNode_Int_emitted <= (lizzieLet17_5QVal_Int_7QNone_Int_6QNode_Int_r ? 2'd0 :
                                                              lizzieLet17_5QVal_Int_7QNone_Int_6QNode_Int_done);
  
  /* dcon (Ty QTree_Int,
      Dcon QError_Int) : [(lizzieLet17_5QVal_Int_7QNone_Int_6QNode_Int_1,Go)] > (lizzieLet17_5QVal_Int_7QNone_Int_6QNode_Int_1QError_Int,QTree_Int) */
  assign lizzieLet17_5QVal_Int_7QNone_Int_6QNode_Int_1QError_Int_d = QError_Int_dc((& {lizzieLet17_5QVal_Int_7QNone_Int_6QNode_Int_1_d[0]}), lizzieLet17_5QVal_Int_7QNone_Int_6QNode_Int_1_d);
  assign {lizzieLet17_5QVal_Int_7QNone_Int_6QNode_Int_1_r} = {1 {(lizzieLet17_5QVal_Int_7QNone_Int_6QNode_Int_1QError_Int_r && lizzieLet17_5QVal_Int_7QNone_Int_6QNode_Int_1QError_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (lizzieLet17_5QVal_Int_7QNone_Int_6QNode_Int_1QError_Int,QTree_Int) > (lizzieLet33_1_argbuf,QTree_Int) */
  QTree_Int_t lizzieLet17_5QVal_Int_7QNone_Int_6QNode_Int_1QError_Int_bufchan_d;
  logic lizzieLet17_5QVal_Int_7QNone_Int_6QNode_Int_1QError_Int_bufchan_r;
  assign lizzieLet17_5QVal_Int_7QNone_Int_6QNode_Int_1QError_Int_r = ((! lizzieLet17_5QVal_Int_7QNone_Int_6QNode_Int_1QError_Int_bufchan_d[0]) || lizzieLet17_5QVal_Int_7QNone_Int_6QNode_Int_1QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QVal_Int_7QNone_Int_6QNode_Int_1QError_Int_bufchan_d <= {66'd0,
                                                                            1'd0};
    else
      if (lizzieLet17_5QVal_Int_7QNone_Int_6QNode_Int_1QError_Int_r)
        lizzieLet17_5QVal_Int_7QNone_Int_6QNode_Int_1QError_Int_bufchan_d <= lizzieLet17_5QVal_Int_7QNone_Int_6QNode_Int_1QError_Int_d;
  QTree_Int_t lizzieLet17_5QVal_Int_7QNone_Int_6QNode_Int_1QError_Int_bufchan_buf;
  assign lizzieLet17_5QVal_Int_7QNone_Int_6QNode_Int_1QError_Int_bufchan_r = (! lizzieLet17_5QVal_Int_7QNone_Int_6QNode_Int_1QError_Int_bufchan_buf[0]);
  assign lizzieLet33_1_argbuf_d = (lizzieLet17_5QVal_Int_7QNone_Int_6QNode_Int_1QError_Int_bufchan_buf[0] ? lizzieLet17_5QVal_Int_7QNone_Int_6QNode_Int_1QError_Int_bufchan_buf :
                                   lizzieLet17_5QVal_Int_7QNone_Int_6QNode_Int_1QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QVal_Int_7QNone_Int_6QNode_Int_1QError_Int_bufchan_buf <= {66'd0,
                                                                              1'd0};
    else
      if ((lizzieLet33_1_argbuf_r && lizzieLet17_5QVal_Int_7QNone_Int_6QNode_Int_1QError_Int_bufchan_buf[0]))
        lizzieLet17_5QVal_Int_7QNone_Int_6QNode_Int_1QError_Int_bufchan_buf <= {66'd0,
                                                                                1'd0};
      else if (((! lizzieLet33_1_argbuf_r) && (! lizzieLet17_5QVal_Int_7QNone_Int_6QNode_Int_1QError_Int_bufchan_buf[0])))
        lizzieLet17_5QVal_Int_7QNone_Int_6QNode_Int_1QError_Int_bufchan_buf <= lizzieLet17_5QVal_Int_7QNone_Int_6QNode_Int_1QError_Int_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet17_5QVal_Int_7QNone_Int_6QNode_Int_2,Go) > (lizzieLet17_5QVal_Int_7QNone_Int_6QNode_Int_2_argbuf,Go) */
  Go_t lizzieLet17_5QVal_Int_7QNone_Int_6QNode_Int_2_bufchan_d;
  logic lizzieLet17_5QVal_Int_7QNone_Int_6QNode_Int_2_bufchan_r;
  assign lizzieLet17_5QVal_Int_7QNone_Int_6QNode_Int_2_r = ((! lizzieLet17_5QVal_Int_7QNone_Int_6QNode_Int_2_bufchan_d[0]) || lizzieLet17_5QVal_Int_7QNone_Int_6QNode_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QVal_Int_7QNone_Int_6QNode_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet17_5QVal_Int_7QNone_Int_6QNode_Int_2_r)
        lizzieLet17_5QVal_Int_7QNone_Int_6QNode_Int_2_bufchan_d <= lizzieLet17_5QVal_Int_7QNone_Int_6QNode_Int_2_d;
  Go_t lizzieLet17_5QVal_Int_7QNone_Int_6QNode_Int_2_bufchan_buf;
  assign lizzieLet17_5QVal_Int_7QNone_Int_6QNode_Int_2_bufchan_r = (! lizzieLet17_5QVal_Int_7QNone_Int_6QNode_Int_2_bufchan_buf[0]);
  assign lizzieLet17_5QVal_Int_7QNone_Int_6QNode_Int_2_argbuf_d = (lizzieLet17_5QVal_Int_7QNone_Int_6QNode_Int_2_bufchan_buf[0] ? lizzieLet17_5QVal_Int_7QNone_Int_6QNode_Int_2_bufchan_buf :
                                                                   lizzieLet17_5QVal_Int_7QNone_Int_6QNode_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QVal_Int_7QNone_Int_6QNode_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet17_5QVal_Int_7QNone_Int_6QNode_Int_2_argbuf_r && lizzieLet17_5QVal_Int_7QNone_Int_6QNode_Int_2_bufchan_buf[0]))
        lizzieLet17_5QVal_Int_7QNone_Int_6QNode_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet17_5QVal_Int_7QNone_Int_6QNode_Int_2_argbuf_r) && (! lizzieLet17_5QVal_Int_7QNone_Int_6QNode_Int_2_bufchan_buf[0])))
        lizzieLet17_5QVal_Int_7QNone_Int_6QNode_Int_2_bufchan_buf <= lizzieLet17_5QVal_Int_7QNone_Int_6QNode_Int_2_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet17_5QVal_Int_7QNone_Int_6QNone_Int,Go) > (lizzieLet17_5QVal_Int_7QNone_Int_6QNone_Int_1_argbuf,Go) */
  Go_t lizzieLet17_5QVal_Int_7QNone_Int_6QNone_Int_bufchan_d;
  logic lizzieLet17_5QVal_Int_7QNone_Int_6QNone_Int_bufchan_r;
  assign lizzieLet17_5QVal_Int_7QNone_Int_6QNone_Int_r = ((! lizzieLet17_5QVal_Int_7QNone_Int_6QNone_Int_bufchan_d[0]) || lizzieLet17_5QVal_Int_7QNone_Int_6QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QVal_Int_7QNone_Int_6QNone_Int_bufchan_d <= 1'd0;
    else
      if (lizzieLet17_5QVal_Int_7QNone_Int_6QNone_Int_r)
        lizzieLet17_5QVal_Int_7QNone_Int_6QNone_Int_bufchan_d <= lizzieLet17_5QVal_Int_7QNone_Int_6QNone_Int_d;
  Go_t lizzieLet17_5QVal_Int_7QNone_Int_6QNone_Int_bufchan_buf;
  assign lizzieLet17_5QVal_Int_7QNone_Int_6QNone_Int_bufchan_r = (! lizzieLet17_5QVal_Int_7QNone_Int_6QNone_Int_bufchan_buf[0]);
  assign lizzieLet17_5QVal_Int_7QNone_Int_6QNone_Int_1_argbuf_d = (lizzieLet17_5QVal_Int_7QNone_Int_6QNone_Int_bufchan_buf[0] ? lizzieLet17_5QVal_Int_7QNone_Int_6QNone_Int_bufchan_buf :
                                                                   lizzieLet17_5QVal_Int_7QNone_Int_6QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QVal_Int_7QNone_Int_6QNone_Int_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet17_5QVal_Int_7QNone_Int_6QNone_Int_1_argbuf_r && lizzieLet17_5QVal_Int_7QNone_Int_6QNone_Int_bufchan_buf[0]))
        lizzieLet17_5QVal_Int_7QNone_Int_6QNone_Int_bufchan_buf <= 1'd0;
      else if (((! lizzieLet17_5QVal_Int_7QNone_Int_6QNone_Int_1_argbuf_r) && (! lizzieLet17_5QVal_Int_7QNone_Int_6QNone_Int_bufchan_buf[0])))
        lizzieLet17_5QVal_Int_7QNone_Int_6QNone_Int_bufchan_buf <= lizzieLet17_5QVal_Int_7QNone_Int_6QNone_Int_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet17_5QVal_Int_7QNone_Int_6QVal_Int,Go) > [(lizzieLet17_5QVal_Int_7QNone_Int_6QVal_Int_1,Go),
                                                                  (lizzieLet17_5QVal_Int_7QNone_Int_6QVal_Int_2,Go)] */
  logic [1:0] lizzieLet17_5QVal_Int_7QNone_Int_6QVal_Int_emitted;
  logic [1:0] lizzieLet17_5QVal_Int_7QNone_Int_6QVal_Int_done;
  assign lizzieLet17_5QVal_Int_7QNone_Int_6QVal_Int_1_d = (lizzieLet17_5QVal_Int_7QNone_Int_6QVal_Int_d[0] && (! lizzieLet17_5QVal_Int_7QNone_Int_6QVal_Int_emitted[0]));
  assign lizzieLet17_5QVal_Int_7QNone_Int_6QVal_Int_2_d = (lizzieLet17_5QVal_Int_7QNone_Int_6QVal_Int_d[0] && (! lizzieLet17_5QVal_Int_7QNone_Int_6QVal_Int_emitted[1]));
  assign lizzieLet17_5QVal_Int_7QNone_Int_6QVal_Int_done = (lizzieLet17_5QVal_Int_7QNone_Int_6QVal_Int_emitted | ({lizzieLet17_5QVal_Int_7QNone_Int_6QVal_Int_2_d[0],
                                                                                                                   lizzieLet17_5QVal_Int_7QNone_Int_6QVal_Int_1_d[0]} & {lizzieLet17_5QVal_Int_7QNone_Int_6QVal_Int_2_r,
                                                                                                                                                                         lizzieLet17_5QVal_Int_7QNone_Int_6QVal_Int_1_r}));
  assign lizzieLet17_5QVal_Int_7QNone_Int_6QVal_Int_r = (& lizzieLet17_5QVal_Int_7QNone_Int_6QVal_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QVal_Int_7QNone_Int_6QVal_Int_emitted <= 2'd0;
    else
      lizzieLet17_5QVal_Int_7QNone_Int_6QVal_Int_emitted <= (lizzieLet17_5QVal_Int_7QNone_Int_6QVal_Int_r ? 2'd0 :
                                                             lizzieLet17_5QVal_Int_7QNone_Int_6QVal_Int_done);
  
  /* buf (Ty Go) : (lizzieLet17_5QVal_Int_7QNone_Int_6QVal_Int_1,Go) > (lizzieLet17_5QVal_Int_7QNone_Int_6QVal_Int_1_argbuf,Go) */
  Go_t lizzieLet17_5QVal_Int_7QNone_Int_6QVal_Int_1_bufchan_d;
  logic lizzieLet17_5QVal_Int_7QNone_Int_6QVal_Int_1_bufchan_r;
  assign lizzieLet17_5QVal_Int_7QNone_Int_6QVal_Int_1_r = ((! lizzieLet17_5QVal_Int_7QNone_Int_6QVal_Int_1_bufchan_d[0]) || lizzieLet17_5QVal_Int_7QNone_Int_6QVal_Int_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QVal_Int_7QNone_Int_6QVal_Int_1_bufchan_d <= 1'd0;
    else
      if (lizzieLet17_5QVal_Int_7QNone_Int_6QVal_Int_1_r)
        lizzieLet17_5QVal_Int_7QNone_Int_6QVal_Int_1_bufchan_d <= lizzieLet17_5QVal_Int_7QNone_Int_6QVal_Int_1_d;
  Go_t lizzieLet17_5QVal_Int_7QNone_Int_6QVal_Int_1_bufchan_buf;
  assign lizzieLet17_5QVal_Int_7QNone_Int_6QVal_Int_1_bufchan_r = (! lizzieLet17_5QVal_Int_7QNone_Int_6QVal_Int_1_bufchan_buf[0]);
  assign lizzieLet17_5QVal_Int_7QNone_Int_6QVal_Int_1_argbuf_d = (lizzieLet17_5QVal_Int_7QNone_Int_6QVal_Int_1_bufchan_buf[0] ? lizzieLet17_5QVal_Int_7QNone_Int_6QVal_Int_1_bufchan_buf :
                                                                  lizzieLet17_5QVal_Int_7QNone_Int_6QVal_Int_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QVal_Int_7QNone_Int_6QVal_Int_1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet17_5QVal_Int_7QNone_Int_6QVal_Int_1_argbuf_r && lizzieLet17_5QVal_Int_7QNone_Int_6QVal_Int_1_bufchan_buf[0]))
        lizzieLet17_5QVal_Int_7QNone_Int_6QVal_Int_1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet17_5QVal_Int_7QNone_Int_6QVal_Int_1_argbuf_r) && (! lizzieLet17_5QVal_Int_7QNone_Int_6QVal_Int_1_bufchan_buf[0])))
        lizzieLet17_5QVal_Int_7QNone_Int_6QVal_Int_1_bufchan_buf <= lizzieLet17_5QVal_Int_7QNone_Int_6QVal_Int_1_bufchan_d;
  
  /* dcon (Ty TupGo___MyDTInt_Bool___Int,
      Dcon TupGo___MyDTInt_Bool___Int) : [(lizzieLet17_5QVal_Int_7QNone_Int_6QVal_Int_1_argbuf,Go),
                                          (lizzieLet17_5QVal_Int_7QNone_Int_7QVal_Int_1_argbuf,MyDTInt_Bool),
                                          (es_9_1_argbuf,Int)] > (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int3,TupGo___MyDTInt_Bool___Int) */
  assign applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int3_d = TupGo___MyDTInt_Bool___Int_dc((& {lizzieLet17_5QVal_Int_7QNone_Int_6QVal_Int_1_argbuf_d[0],
                                                                                            lizzieLet17_5QVal_Int_7QNone_Int_7QVal_Int_1_argbuf_d[0],
                                                                                            es_9_1_argbuf_d[0]}), lizzieLet17_5QVal_Int_7QNone_Int_6QVal_Int_1_argbuf_d, lizzieLet17_5QVal_Int_7QNone_Int_7QVal_Int_1_argbuf_d, es_9_1_argbuf_d);
  assign {lizzieLet17_5QVal_Int_7QNone_Int_6QVal_Int_1_argbuf_r,
          lizzieLet17_5QVal_Int_7QNone_Int_7QVal_Int_1_argbuf_r,
          es_9_1_argbuf_r} = {3 {(applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int3_r && applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int3_d[0])}};
  
  /* demux (Ty QTree_Int,
       Ty MyDTInt_Bool) : (lizzieLet17_5QVal_Int_7QNone_Int_7,QTree_Int) (lizzieLet17_5QVal_Int_6QNone_Int,MyDTInt_Bool) > [(_80,MyDTInt_Bool),
                                                                                                                            (lizzieLet17_5QVal_Int_7QNone_Int_7QVal_Int,MyDTInt_Bool),
                                                                                                                            (_79,MyDTInt_Bool),
                                                                                                                            (_78,MyDTInt_Bool)] */
  logic [3:0] lizzieLet17_5QVal_Int_6QNone_Int_onehotd;
  always_comb
    if ((lizzieLet17_5QVal_Int_7QNone_Int_7_d[0] && lizzieLet17_5QVal_Int_6QNone_Int_d[0]))
      unique case (lizzieLet17_5QVal_Int_7QNone_Int_7_d[2:1])
        2'd0: lizzieLet17_5QVal_Int_6QNone_Int_onehotd = 4'd1;
        2'd1: lizzieLet17_5QVal_Int_6QNone_Int_onehotd = 4'd2;
        2'd2: lizzieLet17_5QVal_Int_6QNone_Int_onehotd = 4'd4;
        2'd3: lizzieLet17_5QVal_Int_6QNone_Int_onehotd = 4'd8;
        default: lizzieLet17_5QVal_Int_6QNone_Int_onehotd = 4'd0;
      endcase
    else lizzieLet17_5QVal_Int_6QNone_Int_onehotd = 4'd0;
  assign _80_d = lizzieLet17_5QVal_Int_6QNone_Int_onehotd[0];
  assign lizzieLet17_5QVal_Int_7QNone_Int_7QVal_Int_d = lizzieLet17_5QVal_Int_6QNone_Int_onehotd[1];
  assign _79_d = lizzieLet17_5QVal_Int_6QNone_Int_onehotd[2];
  assign _78_d = lizzieLet17_5QVal_Int_6QNone_Int_onehotd[3];
  assign lizzieLet17_5QVal_Int_6QNone_Int_r = (| (lizzieLet17_5QVal_Int_6QNone_Int_onehotd & {_78_r,
                                                                                              _79_r,
                                                                                              lizzieLet17_5QVal_Int_7QNone_Int_7QVal_Int_r,
                                                                                              _80_r}));
  assign lizzieLet17_5QVal_Int_7QNone_Int_7_r = lizzieLet17_5QVal_Int_6QNone_Int_r;
  
  /* buf (Ty MyDTInt_Bool) : (lizzieLet17_5QVal_Int_7QNone_Int_7QVal_Int,MyDTInt_Bool) > (lizzieLet17_5QVal_Int_7QNone_Int_7QVal_Int_1_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t lizzieLet17_5QVal_Int_7QNone_Int_7QVal_Int_bufchan_d;
  logic lizzieLet17_5QVal_Int_7QNone_Int_7QVal_Int_bufchan_r;
  assign lizzieLet17_5QVal_Int_7QNone_Int_7QVal_Int_r = ((! lizzieLet17_5QVal_Int_7QNone_Int_7QVal_Int_bufchan_d[0]) || lizzieLet17_5QVal_Int_7QNone_Int_7QVal_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QVal_Int_7QNone_Int_7QVal_Int_bufchan_d <= 1'd0;
    else
      if (lizzieLet17_5QVal_Int_7QNone_Int_7QVal_Int_r)
        lizzieLet17_5QVal_Int_7QNone_Int_7QVal_Int_bufchan_d <= lizzieLet17_5QVal_Int_7QNone_Int_7QVal_Int_d;
  MyDTInt_Bool_t lizzieLet17_5QVal_Int_7QNone_Int_7QVal_Int_bufchan_buf;
  assign lizzieLet17_5QVal_Int_7QNone_Int_7QVal_Int_bufchan_r = (! lizzieLet17_5QVal_Int_7QNone_Int_7QVal_Int_bufchan_buf[0]);
  assign lizzieLet17_5QVal_Int_7QNone_Int_7QVal_Int_1_argbuf_d = (lizzieLet17_5QVal_Int_7QNone_Int_7QVal_Int_bufchan_buf[0] ? lizzieLet17_5QVal_Int_7QNone_Int_7QVal_Int_bufchan_buf :
                                                                  lizzieLet17_5QVal_Int_7QNone_Int_7QVal_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QVal_Int_7QNone_Int_7QVal_Int_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet17_5QVal_Int_7QNone_Int_7QVal_Int_1_argbuf_r && lizzieLet17_5QVal_Int_7QNone_Int_7QVal_Int_bufchan_buf[0]))
        lizzieLet17_5QVal_Int_7QNone_Int_7QVal_Int_bufchan_buf <= 1'd0;
      else if (((! lizzieLet17_5QVal_Int_7QNone_Int_7QVal_Int_1_argbuf_r) && (! lizzieLet17_5QVal_Int_7QNone_Int_7QVal_Int_bufchan_buf[0])))
        lizzieLet17_5QVal_Int_7QNone_Int_7QVal_Int_bufchan_buf <= lizzieLet17_5QVal_Int_7QNone_Int_7QVal_Int_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_QTree_Int) : (lizzieLet17_5QVal_Int_7QNone_Int_8,QTree_Int) (lizzieLet17_5QVal_Int_8QNone_Int,Pointer_QTree_Int) > [(lizzieLet17_5QVal_Int_7QNone_Int_8QNone_Int,Pointer_QTree_Int),
                                                                                                                                      (_77,Pointer_QTree_Int),
                                                                                                                                      (_76,Pointer_QTree_Int),
                                                                                                                                      (_75,Pointer_QTree_Int)] */
  logic [3:0] lizzieLet17_5QVal_Int_8QNone_Int_onehotd;
  always_comb
    if ((lizzieLet17_5QVal_Int_7QNone_Int_8_d[0] && lizzieLet17_5QVal_Int_8QNone_Int_d[0]))
      unique case (lizzieLet17_5QVal_Int_7QNone_Int_8_d[2:1])
        2'd0: lizzieLet17_5QVal_Int_8QNone_Int_onehotd = 4'd1;
        2'd1: lizzieLet17_5QVal_Int_8QNone_Int_onehotd = 4'd2;
        2'd2: lizzieLet17_5QVal_Int_8QNone_Int_onehotd = 4'd4;
        2'd3: lizzieLet17_5QVal_Int_8QNone_Int_onehotd = 4'd8;
        default: lizzieLet17_5QVal_Int_8QNone_Int_onehotd = 4'd0;
      endcase
    else lizzieLet17_5QVal_Int_8QNone_Int_onehotd = 4'd0;
  assign lizzieLet17_5QVal_Int_7QNone_Int_8QNone_Int_d = {lizzieLet17_5QVal_Int_8QNone_Int_d[16:1],
                                                          lizzieLet17_5QVal_Int_8QNone_Int_onehotd[0]};
  assign _77_d = {lizzieLet17_5QVal_Int_8QNone_Int_d[16:1],
                  lizzieLet17_5QVal_Int_8QNone_Int_onehotd[1]};
  assign _76_d = {lizzieLet17_5QVal_Int_8QNone_Int_d[16:1],
                  lizzieLet17_5QVal_Int_8QNone_Int_onehotd[2]};
  assign _75_d = {lizzieLet17_5QVal_Int_8QNone_Int_d[16:1],
                  lizzieLet17_5QVal_Int_8QNone_Int_onehotd[3]};
  assign lizzieLet17_5QVal_Int_8QNone_Int_r = (| (lizzieLet17_5QVal_Int_8QNone_Int_onehotd & {_75_r,
                                                                                              _76_r,
                                                                                              _77_r,
                                                                                              lizzieLet17_5QVal_Int_7QNone_Int_8QNone_Int_r}));
  assign lizzieLet17_5QVal_Int_7QNone_Int_8_r = lizzieLet17_5QVal_Int_8QNone_Int_r;
  
  /* buf (Ty Pointer_QTree_Int) : (lizzieLet17_5QVal_Int_7QNone_Int_8QNone_Int,Pointer_QTree_Int) > (lizzieLet17_5QVal_Int_7QNone_Int_8QNone_Int_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t lizzieLet17_5QVal_Int_7QNone_Int_8QNone_Int_bufchan_d;
  logic lizzieLet17_5QVal_Int_7QNone_Int_8QNone_Int_bufchan_r;
  assign lizzieLet17_5QVal_Int_7QNone_Int_8QNone_Int_r = ((! lizzieLet17_5QVal_Int_7QNone_Int_8QNone_Int_bufchan_d[0]) || lizzieLet17_5QVal_Int_7QNone_Int_8QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QVal_Int_7QNone_Int_8QNone_Int_bufchan_d <= {16'd0,
                                                                1'd0};
    else
      if (lizzieLet17_5QVal_Int_7QNone_Int_8QNone_Int_r)
        lizzieLet17_5QVal_Int_7QNone_Int_8QNone_Int_bufchan_d <= lizzieLet17_5QVal_Int_7QNone_Int_8QNone_Int_d;
  Pointer_QTree_Int_t lizzieLet17_5QVal_Int_7QNone_Int_8QNone_Int_bufchan_buf;
  assign lizzieLet17_5QVal_Int_7QNone_Int_8QNone_Int_bufchan_r = (! lizzieLet17_5QVal_Int_7QNone_Int_8QNone_Int_bufchan_buf[0]);
  assign lizzieLet17_5QVal_Int_7QNone_Int_8QNone_Int_1_argbuf_d = (lizzieLet17_5QVal_Int_7QNone_Int_8QNone_Int_bufchan_buf[0] ? lizzieLet17_5QVal_Int_7QNone_Int_8QNone_Int_bufchan_buf :
                                                                   lizzieLet17_5QVal_Int_7QNone_Int_8QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_5QVal_Int_7QNone_Int_8QNone_Int_bufchan_buf <= {16'd0,
                                                                  1'd0};
    else
      if ((lizzieLet17_5QVal_Int_7QNone_Int_8QNone_Int_1_argbuf_r && lizzieLet17_5QVal_Int_7QNone_Int_8QNone_Int_bufchan_buf[0]))
        lizzieLet17_5QVal_Int_7QNone_Int_8QNone_Int_bufchan_buf <= {16'd0,
                                                                    1'd0};
      else if (((! lizzieLet17_5QVal_Int_7QNone_Int_8QNone_Int_1_argbuf_r) && (! lizzieLet17_5QVal_Int_7QNone_Int_8QNone_Int_bufchan_buf[0])))
        lizzieLet17_5QVal_Int_7QNone_Int_8QNone_Int_bufchan_buf <= lizzieLet17_5QVal_Int_7QNone_Int_8QNone_Int_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_QTree_Int) : (lizzieLet17_5QVal_Int_8,QTree_Int) (lizzieLet17_7QVal_Int,Pointer_QTree_Int) > [(lizzieLet17_5QVal_Int_8QNone_Int,Pointer_QTree_Int),
                                                                                                                (_74,Pointer_QTree_Int),
                                                                                                                (_73,Pointer_QTree_Int),
                                                                                                                (_72,Pointer_QTree_Int)] */
  logic [3:0] lizzieLet17_7QVal_Int_onehotd;
  always_comb
    if ((lizzieLet17_5QVal_Int_8_d[0] && lizzieLet17_7QVal_Int_d[0]))
      unique case (lizzieLet17_5QVal_Int_8_d[2:1])
        2'd0: lizzieLet17_7QVal_Int_onehotd = 4'd1;
        2'd1: lizzieLet17_7QVal_Int_onehotd = 4'd2;
        2'd2: lizzieLet17_7QVal_Int_onehotd = 4'd4;
        2'd3: lizzieLet17_7QVal_Int_onehotd = 4'd8;
        default: lizzieLet17_7QVal_Int_onehotd = 4'd0;
      endcase
    else lizzieLet17_7QVal_Int_onehotd = 4'd0;
  assign lizzieLet17_5QVal_Int_8QNone_Int_d = {lizzieLet17_7QVal_Int_d[16:1],
                                               lizzieLet17_7QVal_Int_onehotd[0]};
  assign _74_d = {lizzieLet17_7QVal_Int_d[16:1],
                  lizzieLet17_7QVal_Int_onehotd[1]};
  assign _73_d = {lizzieLet17_7QVal_Int_d[16:1],
                  lizzieLet17_7QVal_Int_onehotd[2]};
  assign _72_d = {lizzieLet17_7QVal_Int_d[16:1],
                  lizzieLet17_7QVal_Int_onehotd[3]};
  assign lizzieLet17_7QVal_Int_r = (| (lizzieLet17_7QVal_Int_onehotd & {_72_r,
                                                                        _73_r,
                                                                        _74_r,
                                                                        lizzieLet17_5QVal_Int_8QNone_Int_r}));
  assign lizzieLet17_5QVal_Int_8_r = lizzieLet17_7QVal_Int_r;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_QTree_Int) : (lizzieLet17_5QVal_Int_9,QTree_Int) (lizzieLet17_9QVal_Int,Pointer_QTree_Int) > [(_71,Pointer_QTree_Int),
                                                                                                                (lizzieLet17_5QVal_Int_9QVal_Int,Pointer_QTree_Int),
                                                                                                                (_70,Pointer_QTree_Int),
                                                                                                                (_69,Pointer_QTree_Int)] */
  logic [3:0] lizzieLet17_9QVal_Int_onehotd;
  always_comb
    if ((lizzieLet17_5QVal_Int_9_d[0] && lizzieLet17_9QVal_Int_d[0]))
      unique case (lizzieLet17_5QVal_Int_9_d[2:1])
        2'd0: lizzieLet17_9QVal_Int_onehotd = 4'd1;
        2'd1: lizzieLet17_9QVal_Int_onehotd = 4'd2;
        2'd2: lizzieLet17_9QVal_Int_onehotd = 4'd4;
        2'd3: lizzieLet17_9QVal_Int_onehotd = 4'd8;
        default: lizzieLet17_9QVal_Int_onehotd = 4'd0;
      endcase
    else lizzieLet17_9QVal_Int_onehotd = 4'd0;
  assign _71_d = {lizzieLet17_9QVal_Int_d[16:1],
                  lizzieLet17_9QVal_Int_onehotd[0]};
  assign lizzieLet17_5QVal_Int_9QVal_Int_d = {lizzieLet17_9QVal_Int_d[16:1],
                                              lizzieLet17_9QVal_Int_onehotd[1]};
  assign _70_d = {lizzieLet17_9QVal_Int_d[16:1],
                  lizzieLet17_9QVal_Int_onehotd[2]};
  assign _69_d = {lizzieLet17_9QVal_Int_d[16:1],
                  lizzieLet17_9QVal_Int_onehotd[3]};
  assign lizzieLet17_9QVal_Int_r = (| (lizzieLet17_9QVal_Int_onehotd & {_69_r,
                                                                        _70_r,
                                                                        lizzieLet17_5QVal_Int_9QVal_Int_r,
                                                                        _71_r}));
  assign lizzieLet17_5QVal_Int_9_r = lizzieLet17_9QVal_Int_r;
  
  /* demux (Ty QTree_Int,
       Ty QTree_Int) : (lizzieLet17_6,QTree_Int) (readPointer_QTree_Intm3aes_1_argbuf_rwb,QTree_Int) > [(lizzieLet17_6QNone_Int,QTree_Int),
                                                                                                        (lizzieLet17_6QVal_Int,QTree_Int),
                                                                                                        (lizzieLet17_6QNode_Int,QTree_Int),
                                                                                                        (_68,QTree_Int)] */
  logic [3:0] readPointer_QTree_Intm3aes_1_argbuf_rwb_onehotd;
  always_comb
    if ((lizzieLet17_6_d[0] && readPointer_QTree_Intm3aes_1_argbuf_rwb_d[0]))
      unique case (lizzieLet17_6_d[2:1])
        2'd0: readPointer_QTree_Intm3aes_1_argbuf_rwb_onehotd = 4'd1;
        2'd1: readPointer_QTree_Intm3aes_1_argbuf_rwb_onehotd = 4'd2;
        2'd2: readPointer_QTree_Intm3aes_1_argbuf_rwb_onehotd = 4'd4;
        2'd3: readPointer_QTree_Intm3aes_1_argbuf_rwb_onehotd = 4'd8;
        default: readPointer_QTree_Intm3aes_1_argbuf_rwb_onehotd = 4'd0;
      endcase
    else readPointer_QTree_Intm3aes_1_argbuf_rwb_onehotd = 4'd0;
  assign lizzieLet17_6QNone_Int_d = {readPointer_QTree_Intm3aes_1_argbuf_rwb_d[66:1],
                                     readPointer_QTree_Intm3aes_1_argbuf_rwb_onehotd[0]};
  assign lizzieLet17_6QVal_Int_d = {readPointer_QTree_Intm3aes_1_argbuf_rwb_d[66:1],
                                    readPointer_QTree_Intm3aes_1_argbuf_rwb_onehotd[1]};
  assign lizzieLet17_6QNode_Int_d = {readPointer_QTree_Intm3aes_1_argbuf_rwb_d[66:1],
                                     readPointer_QTree_Intm3aes_1_argbuf_rwb_onehotd[2]};
  assign _68_d = {readPointer_QTree_Intm3aes_1_argbuf_rwb_d[66:1],
                  readPointer_QTree_Intm3aes_1_argbuf_rwb_onehotd[3]};
  assign readPointer_QTree_Intm3aes_1_argbuf_rwb_r = (| (readPointer_QTree_Intm3aes_1_argbuf_rwb_onehotd & {_68_r,
                                                                                                            lizzieLet17_6QNode_Int_r,
                                                                                                            lizzieLet17_6QVal_Int_r,
                                                                                                            lizzieLet17_6QNone_Int_r}));
  assign lizzieLet17_6_r = readPointer_QTree_Intm3aes_1_argbuf_rwb_r;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_QTree_Int) : (lizzieLet17_7,QTree_Int) (m1aeq_2,Pointer_QTree_Int) > [(_67,Pointer_QTree_Int),
                                                                                        (lizzieLet17_7QVal_Int,Pointer_QTree_Int),
                                                                                        (lizzieLet17_7QNode_Int,Pointer_QTree_Int),
                                                                                        (_66,Pointer_QTree_Int)] */
  logic [3:0] m1aeq_2_onehotd;
  always_comb
    if ((lizzieLet17_7_d[0] && m1aeq_2_d[0]))
      unique case (lizzieLet17_7_d[2:1])
        2'd0: m1aeq_2_onehotd = 4'd1;
        2'd1: m1aeq_2_onehotd = 4'd2;
        2'd2: m1aeq_2_onehotd = 4'd4;
        2'd3: m1aeq_2_onehotd = 4'd8;
        default: m1aeq_2_onehotd = 4'd0;
      endcase
    else m1aeq_2_onehotd = 4'd0;
  assign _67_d = {m1aeq_2_d[16:1], m1aeq_2_onehotd[0]};
  assign lizzieLet17_7QVal_Int_d = {m1aeq_2_d[16:1],
                                    m1aeq_2_onehotd[1]};
  assign lizzieLet17_7QNode_Int_d = {m1aeq_2_d[16:1],
                                     m1aeq_2_onehotd[2]};
  assign _66_d = {m1aeq_2_d[16:1], m1aeq_2_onehotd[3]};
  assign m1aeq_2_r = (| (m1aeq_2_onehotd & {_66_r,
                                            lizzieLet17_7QNode_Int_r,
                                            lizzieLet17_7QVal_Int_r,
                                            _67_r}));
  assign lizzieLet17_7_r = m1aeq_2_r;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_QTree_Int) : (lizzieLet17_8,QTree_Int) (m2aer_2,Pointer_QTree_Int) > [(lizzieLet17_8QNone_Int,Pointer_QTree_Int),
                                                                                        (_65,Pointer_QTree_Int),
                                                                                        (_64,Pointer_QTree_Int),
                                                                                        (_63,Pointer_QTree_Int)] */
  logic [3:0] m2aer_2_onehotd;
  always_comb
    if ((lizzieLet17_8_d[0] && m2aer_2_d[0]))
      unique case (lizzieLet17_8_d[2:1])
        2'd0: m2aer_2_onehotd = 4'd1;
        2'd1: m2aer_2_onehotd = 4'd2;
        2'd2: m2aer_2_onehotd = 4'd4;
        2'd3: m2aer_2_onehotd = 4'd8;
        default: m2aer_2_onehotd = 4'd0;
      endcase
    else m2aer_2_onehotd = 4'd0;
  assign lizzieLet17_8QNone_Int_d = {m2aer_2_d[16:1],
                                     m2aer_2_onehotd[0]};
  assign _65_d = {m2aer_2_d[16:1], m2aer_2_onehotd[1]};
  assign _64_d = {m2aer_2_d[16:1], m2aer_2_onehotd[2]};
  assign _63_d = {m2aer_2_d[16:1], m2aer_2_onehotd[3]};
  assign m2aer_2_r = (| (m2aer_2_onehotd & {_63_r,
                                            _64_r,
                                            _65_r,
                                            lizzieLet17_8QNone_Int_r}));
  assign lizzieLet17_8_r = m2aer_2_r;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_QTree_Int) : (lizzieLet17_9,QTree_Int) (m3aes_2,Pointer_QTree_Int) > [(lizzieLet17_9QNone_Int,Pointer_QTree_Int),
                                                                                        (lizzieLet17_9QVal_Int,Pointer_QTree_Int),
                                                                                        (_62,Pointer_QTree_Int),
                                                                                        (_61,Pointer_QTree_Int)] */
  logic [3:0] m3aes_2_onehotd;
  always_comb
    if ((lizzieLet17_9_d[0] && m3aes_2_d[0]))
      unique case (lizzieLet17_9_d[2:1])
        2'd0: m3aes_2_onehotd = 4'd1;
        2'd1: m3aes_2_onehotd = 4'd2;
        2'd2: m3aes_2_onehotd = 4'd4;
        2'd3: m3aes_2_onehotd = 4'd8;
        default: m3aes_2_onehotd = 4'd0;
      endcase
    else m3aes_2_onehotd = 4'd0;
  assign lizzieLet17_9QNone_Int_d = {m3aes_2_d[16:1],
                                     m3aes_2_onehotd[0]};
  assign lizzieLet17_9QVal_Int_d = {m3aes_2_d[16:1],
                                    m3aes_2_onehotd[1]};
  assign _62_d = {m3aes_2_d[16:1], m3aes_2_onehotd[2]};
  assign _61_d = {m3aes_2_d[16:1], m3aes_2_onehotd[3]};
  assign m3aes_2_r = (| (m3aes_2_onehotd & {_61_r,
                                            _62_r,
                                            lizzieLet17_9QVal_Int_r,
                                            lizzieLet17_9QNone_Int_r}));
  assign lizzieLet17_9_r = m3aes_2_r;
  
  /* buf (Ty Bool) : (lizzieLet1_1wild1Xv_1_Eq,Bool) > (lizzieLet2_1_argbuf,Bool) */
  Bool_t lizzieLet1_1wild1Xv_1_Eq_bufchan_d;
  logic lizzieLet1_1wild1Xv_1_Eq_bufchan_r;
  assign lizzieLet1_1wild1Xv_1_Eq_r = ((! lizzieLet1_1wild1Xv_1_Eq_bufchan_d[0]) || lizzieLet1_1wild1Xv_1_Eq_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet1_1wild1Xv_1_Eq_bufchan_d <= {1'd0, 1'd0};
    else
      if (lizzieLet1_1wild1Xv_1_Eq_r)
        lizzieLet1_1wild1Xv_1_Eq_bufchan_d <= lizzieLet1_1wild1Xv_1_Eq_d;
  Bool_t lizzieLet1_1wild1Xv_1_Eq_bufchan_buf;
  assign lizzieLet1_1wild1Xv_1_Eq_bufchan_r = (! lizzieLet1_1wild1Xv_1_Eq_bufchan_buf[0]);
  assign lizzieLet2_1_argbuf_d = (lizzieLet1_1wild1Xv_1_Eq_bufchan_buf[0] ? lizzieLet1_1wild1Xv_1_Eq_bufchan_buf :
                                  lizzieLet1_1wild1Xv_1_Eq_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet1_1wild1Xv_1_Eq_bufchan_buf <= {1'd0, 1'd0};
    else
      if ((lizzieLet2_1_argbuf_r && lizzieLet1_1wild1Xv_1_Eq_bufchan_buf[0]))
        lizzieLet1_1wild1Xv_1_Eq_bufchan_buf <= {1'd0, 1'd0};
      else if (((! lizzieLet2_1_argbuf_r) && (! lizzieLet1_1wild1Xv_1_Eq_bufchan_buf[0])))
        lizzieLet1_1wild1Xv_1_Eq_bufchan_buf <= lizzieLet1_1wild1Xv_1_Eq_bufchan_d;
  
  /* demux (Ty MyBool,
       Ty Go) : (lizzieLet3_1,MyBool) (arg0_1Dcon_isZ_3I#_3,Go) > [(lizzieLet3_1MyFalse,Go),
                                                                   (lizzieLet3_1MyTrue,Go)] */
  logic [1:0] \arg0_1Dcon_isZ_3I#_3_onehotd ;
  always_comb
    if ((lizzieLet3_1_d[0] && \arg0_1Dcon_isZ_3I#_3_d [0]))
      unique case (lizzieLet3_1_d[1:1])
        1'd0: \arg0_1Dcon_isZ_3I#_3_onehotd  = 2'd1;
        1'd1: \arg0_1Dcon_isZ_3I#_3_onehotd  = 2'd2;
        default: \arg0_1Dcon_isZ_3I#_3_onehotd  = 2'd0;
      endcase
    else \arg0_1Dcon_isZ_3I#_3_onehotd  = 2'd0;
  assign lizzieLet3_1MyFalse_d = \arg0_1Dcon_isZ_3I#_3_onehotd [0];
  assign lizzieLet3_1MyTrue_d = \arg0_1Dcon_isZ_3I#_3_onehotd [1];
  assign \arg0_1Dcon_isZ_3I#_3_r  = (| (\arg0_1Dcon_isZ_3I#_3_onehotd  & {lizzieLet3_1MyTrue_r,
                                                                          lizzieLet3_1MyFalse_r}));
  assign lizzieLet3_1_r = \arg0_1Dcon_isZ_3I#_3_r ;
  
  /* dcon (Ty MyBool,
      Dcon MyFalse) : [(lizzieLet3_1MyFalse,Go)] > (lizzieLet3_1MyFalse_1MyFalse,MyBool) */
  assign lizzieLet3_1MyFalse_1MyFalse_d = MyFalse_dc((& {lizzieLet3_1MyFalse_d[0]}), lizzieLet3_1MyFalse_d);
  assign {lizzieLet3_1MyFalse_r} = {1 {(lizzieLet3_1MyFalse_1MyFalse_r && lizzieLet3_1MyFalse_1MyFalse_d[0])}};
  
  /* dcon (Ty MyBool,
      Dcon MyTrue) : [(lizzieLet3_1MyTrue,Go)] > (lizzieLet3_1MyTrue_1MyTrue,MyBool) */
  assign lizzieLet3_1MyTrue_1MyTrue_d = MyTrue_dc((& {lizzieLet3_1MyTrue_d[0]}), lizzieLet3_1MyTrue_d);
  assign {lizzieLet3_1MyTrue_r} = {1 {(lizzieLet3_1MyTrue_1MyTrue_r && lizzieLet3_1MyTrue_1MyTrue_d[0])}};
  
  /* mux (Ty MyBool,
     Ty MyBool) : (lizzieLet3_2,MyBool) [(lizzieLet3_1MyFalse_1MyFalse,MyBool),
                                         (lizzieLet3_1MyTrue_1MyTrue,MyBool)] > (lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux,MyBool) */
  logic [1:0] lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux;
  logic [1:0] lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_onehot;
  always_comb
    unique case (lizzieLet3_2_d[1:1])
      1'd0:
        {lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_onehot,
         lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux} = {2'd1,
                                                                            lizzieLet3_1MyFalse_1MyFalse_d};
      1'd1:
        {lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_onehot,
         lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux} = {2'd2,
                                                                            lizzieLet3_1MyTrue_1MyTrue_d};
      default:
        {lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_onehot,
         lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux} = {2'd0,
                                                                            {1'd0, 1'd0}};
    endcase
  assign lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_d = {lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux[1:1],
                                                                         (lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux[0] && lizzieLet3_2_d[0])};
  assign lizzieLet3_2_r = (lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_d[0] && lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_r);
  assign {lizzieLet3_1MyTrue_1MyTrue_r,
          lizzieLet3_1MyFalse_1MyFalse_r} = (lizzieLet3_2_r ? lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_onehot :
                                             2'd0);
  
  /* destruct (Ty QTree_Int,
          Dcon QNode_Int) : (lizzieLet4_1QNode_Int,QTree_Int) > [(q1a8r_destruct,Pointer_QTree_Int),
                                                                 (q2a8s_destruct,Pointer_QTree_Int),
                                                                 (q3a8t_destruct,Pointer_QTree_Int),
                                                                 (q4a8u_destruct,Pointer_QTree_Int)] */
  logic [3:0] lizzieLet4_1QNode_Int_emitted;
  logic [3:0] lizzieLet4_1QNode_Int_done;
  assign q1a8r_destruct_d = {lizzieLet4_1QNode_Int_d[18:3],
                             (lizzieLet4_1QNode_Int_d[0] && (! lizzieLet4_1QNode_Int_emitted[0]))};
  assign q2a8s_destruct_d = {lizzieLet4_1QNode_Int_d[34:19],
                             (lizzieLet4_1QNode_Int_d[0] && (! lizzieLet4_1QNode_Int_emitted[1]))};
  assign q3a8t_destruct_d = {lizzieLet4_1QNode_Int_d[50:35],
                             (lizzieLet4_1QNode_Int_d[0] && (! lizzieLet4_1QNode_Int_emitted[2]))};
  assign q4a8u_destruct_d = {lizzieLet4_1QNode_Int_d[66:51],
                             (lizzieLet4_1QNode_Int_d[0] && (! lizzieLet4_1QNode_Int_emitted[3]))};
  assign lizzieLet4_1QNode_Int_done = (lizzieLet4_1QNode_Int_emitted | ({q4a8u_destruct_d[0],
                                                                         q3a8t_destruct_d[0],
                                                                         q2a8s_destruct_d[0],
                                                                         q1a8r_destruct_d[0]} & {q4a8u_destruct_r,
                                                                                                 q3a8t_destruct_r,
                                                                                                 q2a8s_destruct_r,
                                                                                                 q1a8r_destruct_r}));
  assign lizzieLet4_1QNode_Int_r = (& lizzieLet4_1QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_1QNode_Int_emitted <= 4'd0;
    else
      lizzieLet4_1QNode_Int_emitted <= (lizzieLet4_1QNode_Int_r ? 4'd0 :
                                        lizzieLet4_1QNode_Int_done);
  
  /* demux (Ty QTree_Int,
       Ty QTree_Int) : (lizzieLet4_2,QTree_Int) (lizzieLet4_1,QTree_Int) > [(_60,QTree_Int),
                                                                            (_59,QTree_Int),
                                                                            (lizzieLet4_1QNode_Int,QTree_Int),
                                                                            (_58,QTree_Int)] */
  logic [3:0] lizzieLet4_1_onehotd;
  always_comb
    if ((lizzieLet4_2_d[0] && lizzieLet4_1_d[0]))
      unique case (lizzieLet4_2_d[2:1])
        2'd0: lizzieLet4_1_onehotd = 4'd1;
        2'd1: lizzieLet4_1_onehotd = 4'd2;
        2'd2: lizzieLet4_1_onehotd = 4'd4;
        2'd3: lizzieLet4_1_onehotd = 4'd8;
        default: lizzieLet4_1_onehotd = 4'd0;
      endcase
    else lizzieLet4_1_onehotd = 4'd0;
  assign _60_d = {lizzieLet4_1_d[66:1], lizzieLet4_1_onehotd[0]};
  assign _59_d = {lizzieLet4_1_d[66:1], lizzieLet4_1_onehotd[1]};
  assign lizzieLet4_1QNode_Int_d = {lizzieLet4_1_d[66:1],
                                    lizzieLet4_1_onehotd[2]};
  assign _58_d = {lizzieLet4_1_d[66:1], lizzieLet4_1_onehotd[3]};
  assign lizzieLet4_1_r = (| (lizzieLet4_1_onehotd & {_58_r,
                                                      lizzieLet4_1QNode_Int_r,
                                                      _59_r,
                                                      _60_r}));
  assign lizzieLet4_2_r = lizzieLet4_1_r;
  
  /* demux (Ty QTree_Int,
       Ty Go) : (lizzieLet4_3,QTree_Int) (go_8_goMux_data,Go) > [(lizzieLet4_3QNone_Int,Go),
                                                                 (lizzieLet4_3QVal_Int,Go),
                                                                 (lizzieLet4_3QNode_Int,Go),
                                                                 (lizzieLet4_3QError_Int,Go)] */
  logic [3:0] go_8_goMux_data_onehotd;
  always_comb
    if ((lizzieLet4_3_d[0] && go_8_goMux_data_d[0]))
      unique case (lizzieLet4_3_d[2:1])
        2'd0: go_8_goMux_data_onehotd = 4'd1;
        2'd1: go_8_goMux_data_onehotd = 4'd2;
        2'd2: go_8_goMux_data_onehotd = 4'd4;
        2'd3: go_8_goMux_data_onehotd = 4'd8;
        default: go_8_goMux_data_onehotd = 4'd0;
      endcase
    else go_8_goMux_data_onehotd = 4'd0;
  assign lizzieLet4_3QNone_Int_d = go_8_goMux_data_onehotd[0];
  assign lizzieLet4_3QVal_Int_d = go_8_goMux_data_onehotd[1];
  assign lizzieLet4_3QNode_Int_d = go_8_goMux_data_onehotd[2];
  assign lizzieLet4_3QError_Int_d = go_8_goMux_data_onehotd[3];
  assign go_8_goMux_data_r = (| (go_8_goMux_data_onehotd & {lizzieLet4_3QError_Int_r,
                                                            lizzieLet4_3QNode_Int_r,
                                                            lizzieLet4_3QVal_Int_r,
                                                            lizzieLet4_3QNone_Int_r}));
  assign lizzieLet4_3_r = go_8_goMux_data_r;
  
  /* fork (Ty Go) : (lizzieLet4_3QError_Int,Go) > [(lizzieLet4_3QError_Int_1,Go),
                                              (lizzieLet4_3QError_Int_2,Go)] */
  logic [1:0] lizzieLet4_3QError_Int_emitted;
  logic [1:0] lizzieLet4_3QError_Int_done;
  assign lizzieLet4_3QError_Int_1_d = (lizzieLet4_3QError_Int_d[0] && (! lizzieLet4_3QError_Int_emitted[0]));
  assign lizzieLet4_3QError_Int_2_d = (lizzieLet4_3QError_Int_d[0] && (! lizzieLet4_3QError_Int_emitted[1]));
  assign lizzieLet4_3QError_Int_done = (lizzieLet4_3QError_Int_emitted | ({lizzieLet4_3QError_Int_2_d[0],
                                                                           lizzieLet4_3QError_Int_1_d[0]} & {lizzieLet4_3QError_Int_2_r,
                                                                                                             lizzieLet4_3QError_Int_1_r}));
  assign lizzieLet4_3QError_Int_r = (& lizzieLet4_3QError_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3QError_Int_emitted <= 2'd0;
    else
      lizzieLet4_3QError_Int_emitted <= (lizzieLet4_3QError_Int_r ? 2'd0 :
                                         lizzieLet4_3QError_Int_done);
  
  /* buf (Ty Go) : (lizzieLet4_3QError_Int_1,Go) > (lizzieLet4_3QError_Int_1_argbuf,Go) */
  Go_t lizzieLet4_3QError_Int_1_bufchan_d;
  logic lizzieLet4_3QError_Int_1_bufchan_r;
  assign lizzieLet4_3QError_Int_1_r = ((! lizzieLet4_3QError_Int_1_bufchan_d[0]) || lizzieLet4_3QError_Int_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3QError_Int_1_bufchan_d <= 1'd0;
    else
      if (lizzieLet4_3QError_Int_1_r)
        lizzieLet4_3QError_Int_1_bufchan_d <= lizzieLet4_3QError_Int_1_d;
  Go_t lizzieLet4_3QError_Int_1_bufchan_buf;
  assign lizzieLet4_3QError_Int_1_bufchan_r = (! lizzieLet4_3QError_Int_1_bufchan_buf[0]);
  assign lizzieLet4_3QError_Int_1_argbuf_d = (lizzieLet4_3QError_Int_1_bufchan_buf[0] ? lizzieLet4_3QError_Int_1_bufchan_buf :
                                              lizzieLet4_3QError_Int_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3QError_Int_1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet4_3QError_Int_1_argbuf_r && lizzieLet4_3QError_Int_1_bufchan_buf[0]))
        lizzieLet4_3QError_Int_1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet4_3QError_Int_1_argbuf_r) && (! lizzieLet4_3QError_Int_1_bufchan_buf[0])))
        lizzieLet4_3QError_Int_1_bufchan_buf <= lizzieLet4_3QError_Int_1_bufchan_d;
  
  /* const (Ty Int#,
       Lit 0) : (lizzieLet4_3QError_Int_1_argbuf,Go) > (lizzieLet4_3QError_Int_1_argbuf_0,Int#) */
  assign lizzieLet4_3QError_Int_1_argbuf_0_d = {32'd0,
                                                lizzieLet4_3QError_Int_1_argbuf_d[0]};
  assign lizzieLet4_3QError_Int_1_argbuf_r = lizzieLet4_3QError_Int_1_argbuf_0_r;
  
  /* buf (Ty Int#) : (lizzieLet4_3QError_Int_1_argbuf_0,Int#) > (lizzieLet37_1_1_argbuf,Int#) */
  \Int#_t  lizzieLet4_3QError_Int_1_argbuf_0_bufchan_d;
  logic lizzieLet4_3QError_Int_1_argbuf_0_bufchan_r;
  assign lizzieLet4_3QError_Int_1_argbuf_0_r = ((! lizzieLet4_3QError_Int_1_argbuf_0_bufchan_d[0]) || lizzieLet4_3QError_Int_1_argbuf_0_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_3QError_Int_1_argbuf_0_bufchan_d <= {32'd0, 1'd0};
    else
      if (lizzieLet4_3QError_Int_1_argbuf_0_r)
        lizzieLet4_3QError_Int_1_argbuf_0_bufchan_d <= lizzieLet4_3QError_Int_1_argbuf_0_d;
  \Int#_t  lizzieLet4_3QError_Int_1_argbuf_0_bufchan_buf;
  assign lizzieLet4_3QError_Int_1_argbuf_0_bufchan_r = (! lizzieLet4_3QError_Int_1_argbuf_0_bufchan_buf[0]);
  assign lizzieLet37_1_1_argbuf_d = (lizzieLet4_3QError_Int_1_argbuf_0_bufchan_buf[0] ? lizzieLet4_3QError_Int_1_argbuf_0_bufchan_buf :
                                     lizzieLet4_3QError_Int_1_argbuf_0_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_3QError_Int_1_argbuf_0_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((lizzieLet37_1_1_argbuf_r && lizzieLet4_3QError_Int_1_argbuf_0_bufchan_buf[0]))
        lizzieLet4_3QError_Int_1_argbuf_0_bufchan_buf <= {32'd0, 1'd0};
      else if (((! lizzieLet37_1_1_argbuf_r) && (! lizzieLet4_3QError_Int_1_argbuf_0_bufchan_buf[0])))
        lizzieLet4_3QError_Int_1_argbuf_0_bufchan_buf <= lizzieLet4_3QError_Int_1_argbuf_0_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet4_3QError_Int_2,Go) > (lizzieLet4_3QError_Int_2_argbuf,Go) */
  Go_t lizzieLet4_3QError_Int_2_bufchan_d;
  logic lizzieLet4_3QError_Int_2_bufchan_r;
  assign lizzieLet4_3QError_Int_2_r = ((! lizzieLet4_3QError_Int_2_bufchan_d[0]) || lizzieLet4_3QError_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3QError_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet4_3QError_Int_2_r)
        lizzieLet4_3QError_Int_2_bufchan_d <= lizzieLet4_3QError_Int_2_d;
  Go_t lizzieLet4_3QError_Int_2_bufchan_buf;
  assign lizzieLet4_3QError_Int_2_bufchan_r = (! lizzieLet4_3QError_Int_2_bufchan_buf[0]);
  assign lizzieLet4_3QError_Int_2_argbuf_d = (lizzieLet4_3QError_Int_2_bufchan_buf[0] ? lizzieLet4_3QError_Int_2_bufchan_buf :
                                              lizzieLet4_3QError_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3QError_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet4_3QError_Int_2_argbuf_r && lizzieLet4_3QError_Int_2_bufchan_buf[0]))
        lizzieLet4_3QError_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet4_3QError_Int_2_argbuf_r) && (! lizzieLet4_3QError_Int_2_bufchan_buf[0])))
        lizzieLet4_3QError_Int_2_bufchan_buf <= lizzieLet4_3QError_Int_2_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet4_3QNode_Int,Go) > (lizzieLet4_3QNode_Int_1_argbuf,Go) */
  Go_t lizzieLet4_3QNode_Int_bufchan_d;
  logic lizzieLet4_3QNode_Int_bufchan_r;
  assign lizzieLet4_3QNode_Int_r = ((! lizzieLet4_3QNode_Int_bufchan_d[0]) || lizzieLet4_3QNode_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3QNode_Int_bufchan_d <= 1'd0;
    else
      if (lizzieLet4_3QNode_Int_r)
        lizzieLet4_3QNode_Int_bufchan_d <= lizzieLet4_3QNode_Int_d;
  Go_t lizzieLet4_3QNode_Int_bufchan_buf;
  assign lizzieLet4_3QNode_Int_bufchan_r = (! lizzieLet4_3QNode_Int_bufchan_buf[0]);
  assign lizzieLet4_3QNode_Int_1_argbuf_d = (lizzieLet4_3QNode_Int_bufchan_buf[0] ? lizzieLet4_3QNode_Int_bufchan_buf :
                                             lizzieLet4_3QNode_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3QNode_Int_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet4_3QNode_Int_1_argbuf_r && lizzieLet4_3QNode_Int_bufchan_buf[0]))
        lizzieLet4_3QNode_Int_bufchan_buf <= 1'd0;
      else if (((! lizzieLet4_3QNode_Int_1_argbuf_r) && (! lizzieLet4_3QNode_Int_bufchan_buf[0])))
        lizzieLet4_3QNode_Int_bufchan_buf <= lizzieLet4_3QNode_Int_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet4_3QNone_Int,Go) > [(lizzieLet4_3QNone_Int_1,Go),
                                             (lizzieLet4_3QNone_Int_2,Go)] */
  logic [1:0] lizzieLet4_3QNone_Int_emitted;
  logic [1:0] lizzieLet4_3QNone_Int_done;
  assign lizzieLet4_3QNone_Int_1_d = (lizzieLet4_3QNone_Int_d[0] && (! lizzieLet4_3QNone_Int_emitted[0]));
  assign lizzieLet4_3QNone_Int_2_d = (lizzieLet4_3QNone_Int_d[0] && (! lizzieLet4_3QNone_Int_emitted[1]));
  assign lizzieLet4_3QNone_Int_done = (lizzieLet4_3QNone_Int_emitted | ({lizzieLet4_3QNone_Int_2_d[0],
                                                                         lizzieLet4_3QNone_Int_1_d[0]} & {lizzieLet4_3QNone_Int_2_r,
                                                                                                          lizzieLet4_3QNone_Int_1_r}));
  assign lizzieLet4_3QNone_Int_r = (& lizzieLet4_3QNone_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3QNone_Int_emitted <= 2'd0;
    else
      lizzieLet4_3QNone_Int_emitted <= (lizzieLet4_3QNone_Int_r ? 2'd0 :
                                        lizzieLet4_3QNone_Int_done);
  
  /* buf (Ty Go) : (lizzieLet4_3QNone_Int_1,Go) > (lizzieLet4_3QNone_Int_1_argbuf,Go) */
  Go_t lizzieLet4_3QNone_Int_1_bufchan_d;
  logic lizzieLet4_3QNone_Int_1_bufchan_r;
  assign lizzieLet4_3QNone_Int_1_r = ((! lizzieLet4_3QNone_Int_1_bufchan_d[0]) || lizzieLet4_3QNone_Int_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3QNone_Int_1_bufchan_d <= 1'd0;
    else
      if (lizzieLet4_3QNone_Int_1_r)
        lizzieLet4_3QNone_Int_1_bufchan_d <= lizzieLet4_3QNone_Int_1_d;
  Go_t lizzieLet4_3QNone_Int_1_bufchan_buf;
  assign lizzieLet4_3QNone_Int_1_bufchan_r = (! lizzieLet4_3QNone_Int_1_bufchan_buf[0]);
  assign lizzieLet4_3QNone_Int_1_argbuf_d = (lizzieLet4_3QNone_Int_1_bufchan_buf[0] ? lizzieLet4_3QNone_Int_1_bufchan_buf :
                                             lizzieLet4_3QNone_Int_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3QNone_Int_1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet4_3QNone_Int_1_argbuf_r && lizzieLet4_3QNone_Int_1_bufchan_buf[0]))
        lizzieLet4_3QNone_Int_1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet4_3QNone_Int_1_argbuf_r) && (! lizzieLet4_3QNone_Int_1_bufchan_buf[0])))
        lizzieLet4_3QNone_Int_1_bufchan_buf <= lizzieLet4_3QNone_Int_1_bufchan_d;
  
  /* const (Ty Int#,
       Lit 0) : (lizzieLet4_3QNone_Int_1_argbuf,Go) > (lizzieLet4_3QNone_Int_1_argbuf_0,Int#) */
  assign lizzieLet4_3QNone_Int_1_argbuf_0_d = {32'd0,
                                               lizzieLet4_3QNone_Int_1_argbuf_d[0]};
  assign lizzieLet4_3QNone_Int_1_argbuf_r = lizzieLet4_3QNone_Int_1_argbuf_0_r;
  
  /* buf (Ty Int#) : (lizzieLet4_3QNone_Int_1_argbuf_0,Int#) > (lizzieLet37_1_argbuf,Int#) */
  \Int#_t  lizzieLet4_3QNone_Int_1_argbuf_0_bufchan_d;
  logic lizzieLet4_3QNone_Int_1_argbuf_0_bufchan_r;
  assign lizzieLet4_3QNone_Int_1_argbuf_0_r = ((! lizzieLet4_3QNone_Int_1_argbuf_0_bufchan_d[0]) || lizzieLet4_3QNone_Int_1_argbuf_0_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_3QNone_Int_1_argbuf_0_bufchan_d <= {32'd0, 1'd0};
    else
      if (lizzieLet4_3QNone_Int_1_argbuf_0_r)
        lizzieLet4_3QNone_Int_1_argbuf_0_bufchan_d <= lizzieLet4_3QNone_Int_1_argbuf_0_d;
  \Int#_t  lizzieLet4_3QNone_Int_1_argbuf_0_bufchan_buf;
  assign lizzieLet4_3QNone_Int_1_argbuf_0_bufchan_r = (! lizzieLet4_3QNone_Int_1_argbuf_0_bufchan_buf[0]);
  assign lizzieLet37_1_argbuf_d = (lizzieLet4_3QNone_Int_1_argbuf_0_bufchan_buf[0] ? lizzieLet4_3QNone_Int_1_argbuf_0_bufchan_buf :
                                   lizzieLet4_3QNone_Int_1_argbuf_0_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_3QNone_Int_1_argbuf_0_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((lizzieLet37_1_argbuf_r && lizzieLet4_3QNone_Int_1_argbuf_0_bufchan_buf[0]))
        lizzieLet4_3QNone_Int_1_argbuf_0_bufchan_buf <= {32'd0, 1'd0};
      else if (((! lizzieLet37_1_argbuf_r) && (! lizzieLet4_3QNone_Int_1_argbuf_0_bufchan_buf[0])))
        lizzieLet4_3QNone_Int_1_argbuf_0_bufchan_buf <= lizzieLet4_3QNone_Int_1_argbuf_0_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet4_3QNone_Int_2,Go) > (lizzieLet4_3QNone_Int_2_argbuf,Go) */
  Go_t lizzieLet4_3QNone_Int_2_bufchan_d;
  logic lizzieLet4_3QNone_Int_2_bufchan_r;
  assign lizzieLet4_3QNone_Int_2_r = ((! lizzieLet4_3QNone_Int_2_bufchan_d[0]) || lizzieLet4_3QNone_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3QNone_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet4_3QNone_Int_2_r)
        lizzieLet4_3QNone_Int_2_bufchan_d <= lizzieLet4_3QNone_Int_2_d;
  Go_t lizzieLet4_3QNone_Int_2_bufchan_buf;
  assign lizzieLet4_3QNone_Int_2_bufchan_r = (! lizzieLet4_3QNone_Int_2_bufchan_buf[0]);
  assign lizzieLet4_3QNone_Int_2_argbuf_d = (lizzieLet4_3QNone_Int_2_bufchan_buf[0] ? lizzieLet4_3QNone_Int_2_bufchan_buf :
                                             lizzieLet4_3QNone_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3QNone_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet4_3QNone_Int_2_argbuf_r && lizzieLet4_3QNone_Int_2_bufchan_buf[0]))
        lizzieLet4_3QNone_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet4_3QNone_Int_2_argbuf_r) && (! lizzieLet4_3QNone_Int_2_bufchan_buf[0])))
        lizzieLet4_3QNone_Int_2_bufchan_buf <= lizzieLet4_3QNone_Int_2_bufchan_d;
  
  /* mergectrl (Ty C4,Ty Go) : [(lizzieLet4_3QNone_Int_2_argbuf,Go),
                           (lizzieLet58_3Lcall_$wnnz0_1_argbuf,Go),
                           (lizzieLet4_3QVal_Int_2_argbuf,Go),
                           (lizzieLet4_3QError_Int_2_argbuf,Go)] > (go_13_goMux_choice,C4) (go_13_goMux_data,Go) */
  logic [3:0] lizzieLet4_3QNone_Int_2_argbuf_select_d;
  assign lizzieLet4_3QNone_Int_2_argbuf_select_d = ((| lizzieLet4_3QNone_Int_2_argbuf_select_q) ? lizzieLet4_3QNone_Int_2_argbuf_select_q :
                                                    (lizzieLet4_3QNone_Int_2_argbuf_d[0] ? 4'd1 :
                                                     (lizzieLet58_3Lcall_$wnnz0_1_argbuf_d[0] ? 4'd2 :
                                                      (lizzieLet4_3QVal_Int_2_argbuf_d[0] ? 4'd4 :
                                                       (lizzieLet4_3QError_Int_2_argbuf_d[0] ? 4'd8 :
                                                        4'd0)))));
  logic [3:0] lizzieLet4_3QNone_Int_2_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_3QNone_Int_2_argbuf_select_q <= 4'd0;
    else
      lizzieLet4_3QNone_Int_2_argbuf_select_q <= (lizzieLet4_3QNone_Int_2_argbuf_done ? 4'd0 :
                                                  lizzieLet4_3QNone_Int_2_argbuf_select_d);
  logic [1:0] lizzieLet4_3QNone_Int_2_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3QNone_Int_2_argbuf_emit_q <= 2'd0;
    else
      lizzieLet4_3QNone_Int_2_argbuf_emit_q <= (lizzieLet4_3QNone_Int_2_argbuf_done ? 2'd0 :
                                                lizzieLet4_3QNone_Int_2_argbuf_emit_d);
  logic [1:0] lizzieLet4_3QNone_Int_2_argbuf_emit_d;
  assign lizzieLet4_3QNone_Int_2_argbuf_emit_d = (lizzieLet4_3QNone_Int_2_argbuf_emit_q | ({go_13_goMux_choice_d[0],
                                                                                            go_13_goMux_data_d[0]} & {go_13_goMux_choice_r,
                                                                                                                      go_13_goMux_data_r}));
  logic lizzieLet4_3QNone_Int_2_argbuf_done;
  assign lizzieLet4_3QNone_Int_2_argbuf_done = (& lizzieLet4_3QNone_Int_2_argbuf_emit_d);
  assign {lizzieLet4_3QError_Int_2_argbuf_r,
          lizzieLet4_3QVal_Int_2_argbuf_r,
          lizzieLet58_3Lcall_$wnnz0_1_argbuf_r,
          lizzieLet4_3QNone_Int_2_argbuf_r} = (lizzieLet4_3QNone_Int_2_argbuf_done ? lizzieLet4_3QNone_Int_2_argbuf_select_d :
                                               4'd0);
  assign go_13_goMux_data_d = ((lizzieLet4_3QNone_Int_2_argbuf_select_d[0] && (! lizzieLet4_3QNone_Int_2_argbuf_emit_q[0])) ? lizzieLet4_3QNone_Int_2_argbuf_d :
                               ((lizzieLet4_3QNone_Int_2_argbuf_select_d[1] && (! lizzieLet4_3QNone_Int_2_argbuf_emit_q[0])) ? lizzieLet58_3Lcall_$wnnz0_1_argbuf_d :
                                ((lizzieLet4_3QNone_Int_2_argbuf_select_d[2] && (! lizzieLet4_3QNone_Int_2_argbuf_emit_q[0])) ? lizzieLet4_3QVal_Int_2_argbuf_d :
                                 ((lizzieLet4_3QNone_Int_2_argbuf_select_d[3] && (! lizzieLet4_3QNone_Int_2_argbuf_emit_q[0])) ? lizzieLet4_3QError_Int_2_argbuf_d :
                                  1'd0))));
  assign go_13_goMux_choice_d = ((lizzieLet4_3QNone_Int_2_argbuf_select_d[0] && (! lizzieLet4_3QNone_Int_2_argbuf_emit_q[1])) ? C1_4_dc(1'd1) :
                                 ((lizzieLet4_3QNone_Int_2_argbuf_select_d[1] && (! lizzieLet4_3QNone_Int_2_argbuf_emit_q[1])) ? C2_4_dc(1'd1) :
                                  ((lizzieLet4_3QNone_Int_2_argbuf_select_d[2] && (! lizzieLet4_3QNone_Int_2_argbuf_emit_q[1])) ? C3_4_dc(1'd1) :
                                   ((lizzieLet4_3QNone_Int_2_argbuf_select_d[3] && (! lizzieLet4_3QNone_Int_2_argbuf_emit_q[1])) ? C4_4_dc(1'd1) :
                                    {2'd0, 1'd0}))));
  
  /* fork (Ty Go) : (lizzieLet4_3QVal_Int,Go) > [(lizzieLet4_3QVal_Int_1,Go),
                                            (lizzieLet4_3QVal_Int_2,Go)] */
  logic [1:0] lizzieLet4_3QVal_Int_emitted;
  logic [1:0] lizzieLet4_3QVal_Int_done;
  assign lizzieLet4_3QVal_Int_1_d = (lizzieLet4_3QVal_Int_d[0] && (! lizzieLet4_3QVal_Int_emitted[0]));
  assign lizzieLet4_3QVal_Int_2_d = (lizzieLet4_3QVal_Int_d[0] && (! lizzieLet4_3QVal_Int_emitted[1]));
  assign lizzieLet4_3QVal_Int_done = (lizzieLet4_3QVal_Int_emitted | ({lizzieLet4_3QVal_Int_2_d[0],
                                                                       lizzieLet4_3QVal_Int_1_d[0]} & {lizzieLet4_3QVal_Int_2_r,
                                                                                                       lizzieLet4_3QVal_Int_1_r}));
  assign lizzieLet4_3QVal_Int_r = (& lizzieLet4_3QVal_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3QVal_Int_emitted <= 2'd0;
    else
      lizzieLet4_3QVal_Int_emitted <= (lizzieLet4_3QVal_Int_r ? 2'd0 :
                                       lizzieLet4_3QVal_Int_done);
  
  /* buf (Ty Go) : (lizzieLet4_3QVal_Int_1,Go) > (lizzieLet4_3QVal_Int_1_argbuf,Go) */
  Go_t lizzieLet4_3QVal_Int_1_bufchan_d;
  logic lizzieLet4_3QVal_Int_1_bufchan_r;
  assign lizzieLet4_3QVal_Int_1_r = ((! lizzieLet4_3QVal_Int_1_bufchan_d[0]) || lizzieLet4_3QVal_Int_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3QVal_Int_1_bufchan_d <= 1'd0;
    else
      if (lizzieLet4_3QVal_Int_1_r)
        lizzieLet4_3QVal_Int_1_bufchan_d <= lizzieLet4_3QVal_Int_1_d;
  Go_t lizzieLet4_3QVal_Int_1_bufchan_buf;
  assign lizzieLet4_3QVal_Int_1_bufchan_r = (! lizzieLet4_3QVal_Int_1_bufchan_buf[0]);
  assign lizzieLet4_3QVal_Int_1_argbuf_d = (lizzieLet4_3QVal_Int_1_bufchan_buf[0] ? lizzieLet4_3QVal_Int_1_bufchan_buf :
                                            lizzieLet4_3QVal_Int_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3QVal_Int_1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet4_3QVal_Int_1_argbuf_r && lizzieLet4_3QVal_Int_1_bufchan_buf[0]))
        lizzieLet4_3QVal_Int_1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet4_3QVal_Int_1_argbuf_r) && (! lizzieLet4_3QVal_Int_1_bufchan_buf[0])))
        lizzieLet4_3QVal_Int_1_bufchan_buf <= lizzieLet4_3QVal_Int_1_bufchan_d;
  
  /* const (Ty Int#,
       Lit 1) : (lizzieLet4_3QVal_Int_1_argbuf,Go) > (lizzieLet4_3QVal_Int_1_argbuf_1,Int#) */
  assign lizzieLet4_3QVal_Int_1_argbuf_1_d = {32'd1,
                                              lizzieLet4_3QVal_Int_1_argbuf_d[0]};
  assign lizzieLet4_3QVal_Int_1_argbuf_r = lizzieLet4_3QVal_Int_1_argbuf_1_r;
  
  /* buf (Ty Int#) : (lizzieLet4_3QVal_Int_1_argbuf_1,Int#) > (lizzieLet38_1_argbuf,Int#) */
  \Int#_t  lizzieLet4_3QVal_Int_1_argbuf_1_bufchan_d;
  logic lizzieLet4_3QVal_Int_1_argbuf_1_bufchan_r;
  assign lizzieLet4_3QVal_Int_1_argbuf_1_r = ((! lizzieLet4_3QVal_Int_1_argbuf_1_bufchan_d[0]) || lizzieLet4_3QVal_Int_1_argbuf_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_3QVal_Int_1_argbuf_1_bufchan_d <= {32'd0, 1'd0};
    else
      if (lizzieLet4_3QVal_Int_1_argbuf_1_r)
        lizzieLet4_3QVal_Int_1_argbuf_1_bufchan_d <= lizzieLet4_3QVal_Int_1_argbuf_1_d;
  \Int#_t  lizzieLet4_3QVal_Int_1_argbuf_1_bufchan_buf;
  assign lizzieLet4_3QVal_Int_1_argbuf_1_bufchan_r = (! lizzieLet4_3QVal_Int_1_argbuf_1_bufchan_buf[0]);
  assign lizzieLet38_1_argbuf_d = (lizzieLet4_3QVal_Int_1_argbuf_1_bufchan_buf[0] ? lizzieLet4_3QVal_Int_1_argbuf_1_bufchan_buf :
                                   lizzieLet4_3QVal_Int_1_argbuf_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_3QVal_Int_1_argbuf_1_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((lizzieLet38_1_argbuf_r && lizzieLet4_3QVal_Int_1_argbuf_1_bufchan_buf[0]))
        lizzieLet4_3QVal_Int_1_argbuf_1_bufchan_buf <= {32'd0, 1'd0};
      else if (((! lizzieLet38_1_argbuf_r) && (! lizzieLet4_3QVal_Int_1_argbuf_1_bufchan_buf[0])))
        lizzieLet4_3QVal_Int_1_argbuf_1_bufchan_buf <= lizzieLet4_3QVal_Int_1_argbuf_1_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet4_3QVal_Int_2,Go) > (lizzieLet4_3QVal_Int_2_argbuf,Go) */
  Go_t lizzieLet4_3QVal_Int_2_bufchan_d;
  logic lizzieLet4_3QVal_Int_2_bufchan_r;
  assign lizzieLet4_3QVal_Int_2_r = ((! lizzieLet4_3QVal_Int_2_bufchan_d[0]) || lizzieLet4_3QVal_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3QVal_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet4_3QVal_Int_2_r)
        lizzieLet4_3QVal_Int_2_bufchan_d <= lizzieLet4_3QVal_Int_2_d;
  Go_t lizzieLet4_3QVal_Int_2_bufchan_buf;
  assign lizzieLet4_3QVal_Int_2_bufchan_r = (! lizzieLet4_3QVal_Int_2_bufchan_buf[0]);
  assign lizzieLet4_3QVal_Int_2_argbuf_d = (lizzieLet4_3QVal_Int_2_bufchan_buf[0] ? lizzieLet4_3QVal_Int_2_bufchan_buf :
                                            lizzieLet4_3QVal_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3QVal_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet4_3QVal_Int_2_argbuf_r && lizzieLet4_3QVal_Int_2_bufchan_buf[0]))
        lizzieLet4_3QVal_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet4_3QVal_Int_2_argbuf_r) && (! lizzieLet4_3QVal_Int_2_bufchan_buf[0])))
        lizzieLet4_3QVal_Int_2_bufchan_buf <= lizzieLet4_3QVal_Int_2_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_CT$wnnz) : (lizzieLet4_4,QTree_Int) (sc_0_goMux_mux,Pointer_CT$wnnz) > [(lizzieLet4_4QNone_Int,Pointer_CT$wnnz),
                                                                                          (lizzieLet4_4QVal_Int,Pointer_CT$wnnz),
                                                                                          (lizzieLet4_4QNode_Int,Pointer_CT$wnnz),
                                                                                          (lizzieLet4_4QError_Int,Pointer_CT$wnnz)] */
  logic [3:0] sc_0_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet4_4_d[0] && sc_0_goMux_mux_d[0]))
      unique case (lizzieLet4_4_d[2:1])
        2'd0: sc_0_goMux_mux_onehotd = 4'd1;
        2'd1: sc_0_goMux_mux_onehotd = 4'd2;
        2'd2: sc_0_goMux_mux_onehotd = 4'd4;
        2'd3: sc_0_goMux_mux_onehotd = 4'd8;
        default: sc_0_goMux_mux_onehotd = 4'd0;
      endcase
    else sc_0_goMux_mux_onehotd = 4'd0;
  assign lizzieLet4_4QNone_Int_d = {sc_0_goMux_mux_d[16:1],
                                    sc_0_goMux_mux_onehotd[0]};
  assign lizzieLet4_4QVal_Int_d = {sc_0_goMux_mux_d[16:1],
                                   sc_0_goMux_mux_onehotd[1]};
  assign lizzieLet4_4QNode_Int_d = {sc_0_goMux_mux_d[16:1],
                                    sc_0_goMux_mux_onehotd[2]};
  assign lizzieLet4_4QError_Int_d = {sc_0_goMux_mux_d[16:1],
                                     sc_0_goMux_mux_onehotd[3]};
  assign sc_0_goMux_mux_r = (| (sc_0_goMux_mux_onehotd & {lizzieLet4_4QError_Int_r,
                                                          lizzieLet4_4QNode_Int_r,
                                                          lizzieLet4_4QVal_Int_r,
                                                          lizzieLet4_4QNone_Int_r}));
  assign lizzieLet4_4_r = sc_0_goMux_mux_r;
  
  /* buf (Ty Pointer_CT$wnnz) : (lizzieLet4_4QError_Int,Pointer_CT$wnnz) > (lizzieLet4_4QError_Int_1_argbuf,Pointer_CT$wnnz) */
  Pointer_CT$wnnz_t lizzieLet4_4QError_Int_bufchan_d;
  logic lizzieLet4_4QError_Int_bufchan_r;
  assign lizzieLet4_4QError_Int_r = ((! lizzieLet4_4QError_Int_bufchan_d[0]) || lizzieLet4_4QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_4QError_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet4_4QError_Int_r)
        lizzieLet4_4QError_Int_bufchan_d <= lizzieLet4_4QError_Int_d;
  Pointer_CT$wnnz_t lizzieLet4_4QError_Int_bufchan_buf;
  assign lizzieLet4_4QError_Int_bufchan_r = (! lizzieLet4_4QError_Int_bufchan_buf[0]);
  assign lizzieLet4_4QError_Int_1_argbuf_d = (lizzieLet4_4QError_Int_bufchan_buf[0] ? lizzieLet4_4QError_Int_bufchan_buf :
                                              lizzieLet4_4QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_4QError_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet4_4QError_Int_1_argbuf_r && lizzieLet4_4QError_Int_bufchan_buf[0]))
        lizzieLet4_4QError_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet4_4QError_Int_1_argbuf_r) && (! lizzieLet4_4QError_Int_bufchan_buf[0])))
        lizzieLet4_4QError_Int_bufchan_buf <= lizzieLet4_4QError_Int_bufchan_d;
  
  /* dcon (Ty CT$wnnz,
      Dcon Lcall_$wnnz3) : [(lizzieLet4_4QNode_Int,Pointer_CT$wnnz),
                            (q4a8u_destruct,Pointer_QTree_Int),
                            (q3a8t_destruct,Pointer_QTree_Int),
                            (q2a8s_destruct,Pointer_QTree_Int)] > (lizzieLet4_4QNode_Int_1q4a8u_1q3a8t_1q2a8s_1Lcall_$wnnz3,CT$wnnz) */
  assign lizzieLet4_4QNode_Int_1q4a8u_1q3a8t_1q2a8s_1Lcall_$wnnz3_d = Lcall_$wnnz3_dc((& {lizzieLet4_4QNode_Int_d[0],
                                                                                          q4a8u_destruct_d[0],
                                                                                          q3a8t_destruct_d[0],
                                                                                          q2a8s_destruct_d[0]}), lizzieLet4_4QNode_Int_d, q4a8u_destruct_d, q3a8t_destruct_d, q2a8s_destruct_d);
  assign {lizzieLet4_4QNode_Int_r,
          q4a8u_destruct_r,
          q3a8t_destruct_r,
          q2a8s_destruct_r} = {4 {(lizzieLet4_4QNode_Int_1q4a8u_1q3a8t_1q2a8s_1Lcall_$wnnz3_r && lizzieLet4_4QNode_Int_1q4a8u_1q3a8t_1q2a8s_1Lcall_$wnnz3_d[0])}};
  
  /* buf (Ty CT$wnnz) : (lizzieLet4_4QNode_Int_1q4a8u_1q3a8t_1q2a8s_1Lcall_$wnnz3,CT$wnnz) > (lizzieLet5_1_argbuf,CT$wnnz) */
  CT$wnnz_t lizzieLet4_4QNode_Int_1q4a8u_1q3a8t_1q2a8s_1Lcall_$wnnz3_bufchan_d;
  logic lizzieLet4_4QNode_Int_1q4a8u_1q3a8t_1q2a8s_1Lcall_$wnnz3_bufchan_r;
  assign lizzieLet4_4QNode_Int_1q4a8u_1q3a8t_1q2a8s_1Lcall_$wnnz3_r = ((! lizzieLet4_4QNode_Int_1q4a8u_1q3a8t_1q2a8s_1Lcall_$wnnz3_bufchan_d[0]) || lizzieLet4_4QNode_Int_1q4a8u_1q3a8t_1q2a8s_1Lcall_$wnnz3_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_4QNode_Int_1q4a8u_1q3a8t_1q2a8s_1Lcall_$wnnz3_bufchan_d <= {115'd0,
                                                                             1'd0};
    else
      if (lizzieLet4_4QNode_Int_1q4a8u_1q3a8t_1q2a8s_1Lcall_$wnnz3_r)
        lizzieLet4_4QNode_Int_1q4a8u_1q3a8t_1q2a8s_1Lcall_$wnnz3_bufchan_d <= lizzieLet4_4QNode_Int_1q4a8u_1q3a8t_1q2a8s_1Lcall_$wnnz3_d;
  CT$wnnz_t lizzieLet4_4QNode_Int_1q4a8u_1q3a8t_1q2a8s_1Lcall_$wnnz3_bufchan_buf;
  assign lizzieLet4_4QNode_Int_1q4a8u_1q3a8t_1q2a8s_1Lcall_$wnnz3_bufchan_r = (! lizzieLet4_4QNode_Int_1q4a8u_1q3a8t_1q2a8s_1Lcall_$wnnz3_bufchan_buf[0]);
  assign lizzieLet5_1_argbuf_d = (lizzieLet4_4QNode_Int_1q4a8u_1q3a8t_1q2a8s_1Lcall_$wnnz3_bufchan_buf[0] ? lizzieLet4_4QNode_Int_1q4a8u_1q3a8t_1q2a8s_1Lcall_$wnnz3_bufchan_buf :
                                  lizzieLet4_4QNode_Int_1q4a8u_1q3a8t_1q2a8s_1Lcall_$wnnz3_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_4QNode_Int_1q4a8u_1q3a8t_1q2a8s_1Lcall_$wnnz3_bufchan_buf <= {115'd0,
                                                                               1'd0};
    else
      if ((lizzieLet5_1_argbuf_r && lizzieLet4_4QNode_Int_1q4a8u_1q3a8t_1q2a8s_1Lcall_$wnnz3_bufchan_buf[0]))
        lizzieLet4_4QNode_Int_1q4a8u_1q3a8t_1q2a8s_1Lcall_$wnnz3_bufchan_buf <= {115'd0,
                                                                                 1'd0};
      else if (((! lizzieLet5_1_argbuf_r) && (! lizzieLet4_4QNode_Int_1q4a8u_1q3a8t_1q2a8s_1Lcall_$wnnz3_bufchan_buf[0])))
        lizzieLet4_4QNode_Int_1q4a8u_1q3a8t_1q2a8s_1Lcall_$wnnz3_bufchan_buf <= lizzieLet4_4QNode_Int_1q4a8u_1q3a8t_1q2a8s_1Lcall_$wnnz3_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz) : (lizzieLet4_4QNone_Int,Pointer_CT$wnnz) > (lizzieLet4_4QNone_Int_1_argbuf,Pointer_CT$wnnz) */
  Pointer_CT$wnnz_t lizzieLet4_4QNone_Int_bufchan_d;
  logic lizzieLet4_4QNone_Int_bufchan_r;
  assign lizzieLet4_4QNone_Int_r = ((! lizzieLet4_4QNone_Int_bufchan_d[0]) || lizzieLet4_4QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_4QNone_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet4_4QNone_Int_r)
        lizzieLet4_4QNone_Int_bufchan_d <= lizzieLet4_4QNone_Int_d;
  Pointer_CT$wnnz_t lizzieLet4_4QNone_Int_bufchan_buf;
  assign lizzieLet4_4QNone_Int_bufchan_r = (! lizzieLet4_4QNone_Int_bufchan_buf[0]);
  assign lizzieLet4_4QNone_Int_1_argbuf_d = (lizzieLet4_4QNone_Int_bufchan_buf[0] ? lizzieLet4_4QNone_Int_bufchan_buf :
                                             lizzieLet4_4QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_4QNone_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet4_4QNone_Int_1_argbuf_r && lizzieLet4_4QNone_Int_bufchan_buf[0]))
        lizzieLet4_4QNone_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet4_4QNone_Int_1_argbuf_r) && (! lizzieLet4_4QNone_Int_bufchan_buf[0])))
        lizzieLet4_4QNone_Int_bufchan_buf <= lizzieLet4_4QNone_Int_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz) : (lizzieLet4_4QVal_Int,Pointer_CT$wnnz) > (lizzieLet4_4QVal_Int_1_argbuf,Pointer_CT$wnnz) */
  Pointer_CT$wnnz_t lizzieLet4_4QVal_Int_bufchan_d;
  logic lizzieLet4_4QVal_Int_bufchan_r;
  assign lizzieLet4_4QVal_Int_r = ((! lizzieLet4_4QVal_Int_bufchan_d[0]) || lizzieLet4_4QVal_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_4QVal_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet4_4QVal_Int_r)
        lizzieLet4_4QVal_Int_bufchan_d <= lizzieLet4_4QVal_Int_d;
  Pointer_CT$wnnz_t lizzieLet4_4QVal_Int_bufchan_buf;
  assign lizzieLet4_4QVal_Int_bufchan_r = (! lizzieLet4_4QVal_Int_bufchan_buf[0]);
  assign lizzieLet4_4QVal_Int_1_argbuf_d = (lizzieLet4_4QVal_Int_bufchan_buf[0] ? lizzieLet4_4QVal_Int_bufchan_buf :
                                            lizzieLet4_4QVal_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_4QVal_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet4_4QVal_Int_1_argbuf_r && lizzieLet4_4QVal_Int_bufchan_buf[0]))
        lizzieLet4_4QVal_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet4_4QVal_Int_1_argbuf_r) && (! lizzieLet4_4QVal_Int_bufchan_buf[0])))
        lizzieLet4_4QVal_Int_bufchan_buf <= lizzieLet4_4QVal_Int_bufchan_d;
  
  /* destruct (Ty CT$wnnz,
          Dcon Lcall_$wnnz0) : (lizzieLet58_1Lcall_$wnnz0,CT$wnnz) > [(wwsmn_4_destruct,Int#),
                                                                      (ww1XmW_2_destruct,Int#),
                                                                      (ww2XmZ_1_destruct,Int#),
                                                                      (sc_0_6_destruct,Pointer_CT$wnnz)] */
  logic [3:0] lizzieLet58_1Lcall_$wnnz0_emitted;
  logic [3:0] lizzieLet58_1Lcall_$wnnz0_done;
  assign wwsmn_4_destruct_d = {lizzieLet58_1Lcall_$wnnz0_d[35:4],
                               (lizzieLet58_1Lcall_$wnnz0_d[0] && (! lizzieLet58_1Lcall_$wnnz0_emitted[0]))};
  assign ww1XmW_2_destruct_d = {lizzieLet58_1Lcall_$wnnz0_d[67:36],
                                (lizzieLet58_1Lcall_$wnnz0_d[0] && (! lizzieLet58_1Lcall_$wnnz0_emitted[1]))};
  assign ww2XmZ_1_destruct_d = {lizzieLet58_1Lcall_$wnnz0_d[99:68],
                                (lizzieLet58_1Lcall_$wnnz0_d[0] && (! lizzieLet58_1Lcall_$wnnz0_emitted[2]))};
  assign sc_0_6_destruct_d = {lizzieLet58_1Lcall_$wnnz0_d[115:100],
                              (lizzieLet58_1Lcall_$wnnz0_d[0] && (! lizzieLet58_1Lcall_$wnnz0_emitted[3]))};
  assign lizzieLet58_1Lcall_$wnnz0_done = (lizzieLet58_1Lcall_$wnnz0_emitted | ({sc_0_6_destruct_d[0],
                                                                                 ww2XmZ_1_destruct_d[0],
                                                                                 ww1XmW_2_destruct_d[0],
                                                                                 wwsmn_4_destruct_d[0]} & {sc_0_6_destruct_r,
                                                                                                           ww2XmZ_1_destruct_r,
                                                                                                           ww1XmW_2_destruct_r,
                                                                                                           wwsmn_4_destruct_r}));
  assign lizzieLet58_1Lcall_$wnnz0_r = (& lizzieLet58_1Lcall_$wnnz0_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet58_1Lcall_$wnnz0_emitted <= 4'd0;
    else
      lizzieLet58_1Lcall_$wnnz0_emitted <= (lizzieLet58_1Lcall_$wnnz0_r ? 4'd0 :
                                            lizzieLet58_1Lcall_$wnnz0_done);
  
  /* destruct (Ty CT$wnnz,
          Dcon Lcall_$wnnz1) : (lizzieLet58_1Lcall_$wnnz1,CT$wnnz) > [(wwsmn_3_destruct,Int#),
                                                                      (ww1XmW_1_destruct,Int#),
                                                                      (sc_0_5_destruct,Pointer_CT$wnnz),
                                                                      (q4a8u_3_destruct,Pointer_QTree_Int)] */
  logic [3:0] lizzieLet58_1Lcall_$wnnz1_emitted;
  logic [3:0] lizzieLet58_1Lcall_$wnnz1_done;
  assign wwsmn_3_destruct_d = {lizzieLet58_1Lcall_$wnnz1_d[35:4],
                               (lizzieLet58_1Lcall_$wnnz1_d[0] && (! lizzieLet58_1Lcall_$wnnz1_emitted[0]))};
  assign ww1XmW_1_destruct_d = {lizzieLet58_1Lcall_$wnnz1_d[67:36],
                                (lizzieLet58_1Lcall_$wnnz1_d[0] && (! lizzieLet58_1Lcall_$wnnz1_emitted[1]))};
  assign sc_0_5_destruct_d = {lizzieLet58_1Lcall_$wnnz1_d[83:68],
                              (lizzieLet58_1Lcall_$wnnz1_d[0] && (! lizzieLet58_1Lcall_$wnnz1_emitted[2]))};
  assign q4a8u_3_destruct_d = {lizzieLet58_1Lcall_$wnnz1_d[99:84],
                               (lizzieLet58_1Lcall_$wnnz1_d[0] && (! lizzieLet58_1Lcall_$wnnz1_emitted[3]))};
  assign lizzieLet58_1Lcall_$wnnz1_done = (lizzieLet58_1Lcall_$wnnz1_emitted | ({q4a8u_3_destruct_d[0],
                                                                                 sc_0_5_destruct_d[0],
                                                                                 ww1XmW_1_destruct_d[0],
                                                                                 wwsmn_3_destruct_d[0]} & {q4a8u_3_destruct_r,
                                                                                                           sc_0_5_destruct_r,
                                                                                                           ww1XmW_1_destruct_r,
                                                                                                           wwsmn_3_destruct_r}));
  assign lizzieLet58_1Lcall_$wnnz1_r = (& lizzieLet58_1Lcall_$wnnz1_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet58_1Lcall_$wnnz1_emitted <= 4'd0;
    else
      lizzieLet58_1Lcall_$wnnz1_emitted <= (lizzieLet58_1Lcall_$wnnz1_r ? 4'd0 :
                                            lizzieLet58_1Lcall_$wnnz1_done);
  
  /* destruct (Ty CT$wnnz,
          Dcon Lcall_$wnnz2) : (lizzieLet58_1Lcall_$wnnz2,CT$wnnz) > [(wwsmn_2_destruct,Int#),
                                                                      (sc_0_4_destruct,Pointer_CT$wnnz),
                                                                      (q4a8u_2_destruct,Pointer_QTree_Int),
                                                                      (q3a8t_2_destruct,Pointer_QTree_Int)] */
  logic [3:0] lizzieLet58_1Lcall_$wnnz2_emitted;
  logic [3:0] lizzieLet58_1Lcall_$wnnz2_done;
  assign wwsmn_2_destruct_d = {lizzieLet58_1Lcall_$wnnz2_d[35:4],
                               (lizzieLet58_1Lcall_$wnnz2_d[0] && (! lizzieLet58_1Lcall_$wnnz2_emitted[0]))};
  assign sc_0_4_destruct_d = {lizzieLet58_1Lcall_$wnnz2_d[51:36],
                              (lizzieLet58_1Lcall_$wnnz2_d[0] && (! lizzieLet58_1Lcall_$wnnz2_emitted[1]))};
  assign q4a8u_2_destruct_d = {lizzieLet58_1Lcall_$wnnz2_d[67:52],
                               (lizzieLet58_1Lcall_$wnnz2_d[0] && (! lizzieLet58_1Lcall_$wnnz2_emitted[2]))};
  assign q3a8t_2_destruct_d = {lizzieLet58_1Lcall_$wnnz2_d[83:68],
                               (lizzieLet58_1Lcall_$wnnz2_d[0] && (! lizzieLet58_1Lcall_$wnnz2_emitted[3]))};
  assign lizzieLet58_1Lcall_$wnnz2_done = (lizzieLet58_1Lcall_$wnnz2_emitted | ({q3a8t_2_destruct_d[0],
                                                                                 q4a8u_2_destruct_d[0],
                                                                                 sc_0_4_destruct_d[0],
                                                                                 wwsmn_2_destruct_d[0]} & {q3a8t_2_destruct_r,
                                                                                                           q4a8u_2_destruct_r,
                                                                                                           sc_0_4_destruct_r,
                                                                                                           wwsmn_2_destruct_r}));
  assign lizzieLet58_1Lcall_$wnnz2_r = (& lizzieLet58_1Lcall_$wnnz2_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet58_1Lcall_$wnnz2_emitted <= 4'd0;
    else
      lizzieLet58_1Lcall_$wnnz2_emitted <= (lizzieLet58_1Lcall_$wnnz2_r ? 4'd0 :
                                            lizzieLet58_1Lcall_$wnnz2_done);
  
  /* destruct (Ty CT$wnnz,
          Dcon Lcall_$wnnz3) : (lizzieLet58_1Lcall_$wnnz3,CT$wnnz) > [(sc_0_3_destruct,Pointer_CT$wnnz),
                                                                      (q4a8u_1_destruct,Pointer_QTree_Int),
                                                                      (q3a8t_1_destruct,Pointer_QTree_Int),
                                                                      (q2a8s_1_destruct,Pointer_QTree_Int)] */
  logic [3:0] lizzieLet58_1Lcall_$wnnz3_emitted;
  logic [3:0] lizzieLet58_1Lcall_$wnnz3_done;
  assign sc_0_3_destruct_d = {lizzieLet58_1Lcall_$wnnz3_d[19:4],
                              (lizzieLet58_1Lcall_$wnnz3_d[0] && (! lizzieLet58_1Lcall_$wnnz3_emitted[0]))};
  assign q4a8u_1_destruct_d = {lizzieLet58_1Lcall_$wnnz3_d[35:20],
                               (lizzieLet58_1Lcall_$wnnz3_d[0] && (! lizzieLet58_1Lcall_$wnnz3_emitted[1]))};
  assign q3a8t_1_destruct_d = {lizzieLet58_1Lcall_$wnnz3_d[51:36],
                               (lizzieLet58_1Lcall_$wnnz3_d[0] && (! lizzieLet58_1Lcall_$wnnz3_emitted[2]))};
  assign q2a8s_1_destruct_d = {lizzieLet58_1Lcall_$wnnz3_d[67:52],
                               (lizzieLet58_1Lcall_$wnnz3_d[0] && (! lizzieLet58_1Lcall_$wnnz3_emitted[3]))};
  assign lizzieLet58_1Lcall_$wnnz3_done = (lizzieLet58_1Lcall_$wnnz3_emitted | ({q2a8s_1_destruct_d[0],
                                                                                 q3a8t_1_destruct_d[0],
                                                                                 q4a8u_1_destruct_d[0],
                                                                                 sc_0_3_destruct_d[0]} & {q2a8s_1_destruct_r,
                                                                                                          q3a8t_1_destruct_r,
                                                                                                          q4a8u_1_destruct_r,
                                                                                                          sc_0_3_destruct_r}));
  assign lizzieLet58_1Lcall_$wnnz3_r = (& lizzieLet58_1Lcall_$wnnz3_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet58_1Lcall_$wnnz3_emitted <= 4'd0;
    else
      lizzieLet58_1Lcall_$wnnz3_emitted <= (lizzieLet58_1Lcall_$wnnz3_r ? 4'd0 :
                                            lizzieLet58_1Lcall_$wnnz3_done);
  
  /* demux (Ty CT$wnnz,
       Ty CT$wnnz) : (lizzieLet58_2,CT$wnnz) (lizzieLet58_1,CT$wnnz) > [(_57,CT$wnnz),
                                                                        (lizzieLet58_1Lcall_$wnnz3,CT$wnnz),
                                                                        (lizzieLet58_1Lcall_$wnnz2,CT$wnnz),
                                                                        (lizzieLet58_1Lcall_$wnnz1,CT$wnnz),
                                                                        (lizzieLet58_1Lcall_$wnnz0,CT$wnnz)] */
  logic [4:0] lizzieLet58_1_onehotd;
  always_comb
    if ((lizzieLet58_2_d[0] && lizzieLet58_1_d[0]))
      unique case (lizzieLet58_2_d[3:1])
        3'd0: lizzieLet58_1_onehotd = 5'd1;
        3'd1: lizzieLet58_1_onehotd = 5'd2;
        3'd2: lizzieLet58_1_onehotd = 5'd4;
        3'd3: lizzieLet58_1_onehotd = 5'd8;
        3'd4: lizzieLet58_1_onehotd = 5'd16;
        default: lizzieLet58_1_onehotd = 5'd0;
      endcase
    else lizzieLet58_1_onehotd = 5'd0;
  assign _57_d = {lizzieLet58_1_d[115:1], lizzieLet58_1_onehotd[0]};
  assign lizzieLet58_1Lcall_$wnnz3_d = {lizzieLet58_1_d[115:1],
                                        lizzieLet58_1_onehotd[1]};
  assign lizzieLet58_1Lcall_$wnnz2_d = {lizzieLet58_1_d[115:1],
                                        lizzieLet58_1_onehotd[2]};
  assign lizzieLet58_1Lcall_$wnnz1_d = {lizzieLet58_1_d[115:1],
                                        lizzieLet58_1_onehotd[3]};
  assign lizzieLet58_1Lcall_$wnnz0_d = {lizzieLet58_1_d[115:1],
                                        lizzieLet58_1_onehotd[4]};
  assign lizzieLet58_1_r = (| (lizzieLet58_1_onehotd & {lizzieLet58_1Lcall_$wnnz0_r,
                                                        lizzieLet58_1Lcall_$wnnz1_r,
                                                        lizzieLet58_1Lcall_$wnnz2_r,
                                                        lizzieLet58_1Lcall_$wnnz3_r,
                                                        _57_r}));
  assign lizzieLet58_2_r = lizzieLet58_1_r;
  
  /* demux (Ty CT$wnnz,
       Ty Go) : (lizzieLet58_3,CT$wnnz) (go_13_goMux_data,Go) > [(_56,Go),
                                                                 (lizzieLet58_3Lcall_$wnnz3,Go),
                                                                 (lizzieLet58_3Lcall_$wnnz2,Go),
                                                                 (lizzieLet58_3Lcall_$wnnz1,Go),
                                                                 (lizzieLet58_3Lcall_$wnnz0,Go)] */
  logic [4:0] go_13_goMux_data_onehotd;
  always_comb
    if ((lizzieLet58_3_d[0] && go_13_goMux_data_d[0]))
      unique case (lizzieLet58_3_d[3:1])
        3'd0: go_13_goMux_data_onehotd = 5'd1;
        3'd1: go_13_goMux_data_onehotd = 5'd2;
        3'd2: go_13_goMux_data_onehotd = 5'd4;
        3'd3: go_13_goMux_data_onehotd = 5'd8;
        3'd4: go_13_goMux_data_onehotd = 5'd16;
        default: go_13_goMux_data_onehotd = 5'd0;
      endcase
    else go_13_goMux_data_onehotd = 5'd0;
  assign _56_d = go_13_goMux_data_onehotd[0];
  assign lizzieLet58_3Lcall_$wnnz3_d = go_13_goMux_data_onehotd[1];
  assign lizzieLet58_3Lcall_$wnnz2_d = go_13_goMux_data_onehotd[2];
  assign lizzieLet58_3Lcall_$wnnz1_d = go_13_goMux_data_onehotd[3];
  assign lizzieLet58_3Lcall_$wnnz0_d = go_13_goMux_data_onehotd[4];
  assign go_13_goMux_data_r = (| (go_13_goMux_data_onehotd & {lizzieLet58_3Lcall_$wnnz0_r,
                                                              lizzieLet58_3Lcall_$wnnz1_r,
                                                              lizzieLet58_3Lcall_$wnnz2_r,
                                                              lizzieLet58_3Lcall_$wnnz3_r,
                                                              _56_r}));
  assign lizzieLet58_3_r = go_13_goMux_data_r;
  
  /* buf (Ty Go) : (lizzieLet58_3Lcall_$wnnz0,Go) > (lizzieLet58_3Lcall_$wnnz0_1_argbuf,Go) */
  Go_t lizzieLet58_3Lcall_$wnnz0_bufchan_d;
  logic lizzieLet58_3Lcall_$wnnz0_bufchan_r;
  assign lizzieLet58_3Lcall_$wnnz0_r = ((! lizzieLet58_3Lcall_$wnnz0_bufchan_d[0]) || lizzieLet58_3Lcall_$wnnz0_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet58_3Lcall_$wnnz0_bufchan_d <= 1'd0;
    else
      if (lizzieLet58_3Lcall_$wnnz0_r)
        lizzieLet58_3Lcall_$wnnz0_bufchan_d <= lizzieLet58_3Lcall_$wnnz0_d;
  Go_t lizzieLet58_3Lcall_$wnnz0_bufchan_buf;
  assign lizzieLet58_3Lcall_$wnnz0_bufchan_r = (! lizzieLet58_3Lcall_$wnnz0_bufchan_buf[0]);
  assign lizzieLet58_3Lcall_$wnnz0_1_argbuf_d = (lizzieLet58_3Lcall_$wnnz0_bufchan_buf[0] ? lizzieLet58_3Lcall_$wnnz0_bufchan_buf :
                                                 lizzieLet58_3Lcall_$wnnz0_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet58_3Lcall_$wnnz0_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet58_3Lcall_$wnnz0_1_argbuf_r && lizzieLet58_3Lcall_$wnnz0_bufchan_buf[0]))
        lizzieLet58_3Lcall_$wnnz0_bufchan_buf <= 1'd0;
      else if (((! lizzieLet58_3Lcall_$wnnz0_1_argbuf_r) && (! lizzieLet58_3Lcall_$wnnz0_bufchan_buf[0])))
        lizzieLet58_3Lcall_$wnnz0_bufchan_buf <= lizzieLet58_3Lcall_$wnnz0_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet58_3Lcall_$wnnz1,Go) > (lizzieLet58_3Lcall_$wnnz1_1_argbuf,Go) */
  Go_t lizzieLet58_3Lcall_$wnnz1_bufchan_d;
  logic lizzieLet58_3Lcall_$wnnz1_bufchan_r;
  assign lizzieLet58_3Lcall_$wnnz1_r = ((! lizzieLet58_3Lcall_$wnnz1_bufchan_d[0]) || lizzieLet58_3Lcall_$wnnz1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet58_3Lcall_$wnnz1_bufchan_d <= 1'd0;
    else
      if (lizzieLet58_3Lcall_$wnnz1_r)
        lizzieLet58_3Lcall_$wnnz1_bufchan_d <= lizzieLet58_3Lcall_$wnnz1_d;
  Go_t lizzieLet58_3Lcall_$wnnz1_bufchan_buf;
  assign lizzieLet58_3Lcall_$wnnz1_bufchan_r = (! lizzieLet58_3Lcall_$wnnz1_bufchan_buf[0]);
  assign lizzieLet58_3Lcall_$wnnz1_1_argbuf_d = (lizzieLet58_3Lcall_$wnnz1_bufchan_buf[0] ? lizzieLet58_3Lcall_$wnnz1_bufchan_buf :
                                                 lizzieLet58_3Lcall_$wnnz1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet58_3Lcall_$wnnz1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet58_3Lcall_$wnnz1_1_argbuf_r && lizzieLet58_3Lcall_$wnnz1_bufchan_buf[0]))
        lizzieLet58_3Lcall_$wnnz1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet58_3Lcall_$wnnz1_1_argbuf_r) && (! lizzieLet58_3Lcall_$wnnz1_bufchan_buf[0])))
        lizzieLet58_3Lcall_$wnnz1_bufchan_buf <= lizzieLet58_3Lcall_$wnnz1_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet58_3Lcall_$wnnz2,Go) > (lizzieLet58_3Lcall_$wnnz2_1_argbuf,Go) */
  Go_t lizzieLet58_3Lcall_$wnnz2_bufchan_d;
  logic lizzieLet58_3Lcall_$wnnz2_bufchan_r;
  assign lizzieLet58_3Lcall_$wnnz2_r = ((! lizzieLet58_3Lcall_$wnnz2_bufchan_d[0]) || lizzieLet58_3Lcall_$wnnz2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet58_3Lcall_$wnnz2_bufchan_d <= 1'd0;
    else
      if (lizzieLet58_3Lcall_$wnnz2_r)
        lizzieLet58_3Lcall_$wnnz2_bufchan_d <= lizzieLet58_3Lcall_$wnnz2_d;
  Go_t lizzieLet58_3Lcall_$wnnz2_bufchan_buf;
  assign lizzieLet58_3Lcall_$wnnz2_bufchan_r = (! lizzieLet58_3Lcall_$wnnz2_bufchan_buf[0]);
  assign lizzieLet58_3Lcall_$wnnz2_1_argbuf_d = (lizzieLet58_3Lcall_$wnnz2_bufchan_buf[0] ? lizzieLet58_3Lcall_$wnnz2_bufchan_buf :
                                                 lizzieLet58_3Lcall_$wnnz2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet58_3Lcall_$wnnz2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet58_3Lcall_$wnnz2_1_argbuf_r && lizzieLet58_3Lcall_$wnnz2_bufchan_buf[0]))
        lizzieLet58_3Lcall_$wnnz2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet58_3Lcall_$wnnz2_1_argbuf_r) && (! lizzieLet58_3Lcall_$wnnz2_bufchan_buf[0])))
        lizzieLet58_3Lcall_$wnnz2_bufchan_buf <= lizzieLet58_3Lcall_$wnnz2_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet58_3Lcall_$wnnz3,Go) > (lizzieLet58_3Lcall_$wnnz3_1_argbuf,Go) */
  Go_t lizzieLet58_3Lcall_$wnnz3_bufchan_d;
  logic lizzieLet58_3Lcall_$wnnz3_bufchan_r;
  assign lizzieLet58_3Lcall_$wnnz3_r = ((! lizzieLet58_3Lcall_$wnnz3_bufchan_d[0]) || lizzieLet58_3Lcall_$wnnz3_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet58_3Lcall_$wnnz3_bufchan_d <= 1'd0;
    else
      if (lizzieLet58_3Lcall_$wnnz3_r)
        lizzieLet58_3Lcall_$wnnz3_bufchan_d <= lizzieLet58_3Lcall_$wnnz3_d;
  Go_t lizzieLet58_3Lcall_$wnnz3_bufchan_buf;
  assign lizzieLet58_3Lcall_$wnnz3_bufchan_r = (! lizzieLet58_3Lcall_$wnnz3_bufchan_buf[0]);
  assign lizzieLet58_3Lcall_$wnnz3_1_argbuf_d = (lizzieLet58_3Lcall_$wnnz3_bufchan_buf[0] ? lizzieLet58_3Lcall_$wnnz3_bufchan_buf :
                                                 lizzieLet58_3Lcall_$wnnz3_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet58_3Lcall_$wnnz3_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet58_3Lcall_$wnnz3_1_argbuf_r && lizzieLet58_3Lcall_$wnnz3_bufchan_buf[0]))
        lizzieLet58_3Lcall_$wnnz3_bufchan_buf <= 1'd0;
      else if (((! lizzieLet58_3Lcall_$wnnz3_1_argbuf_r) && (! lizzieLet58_3Lcall_$wnnz3_bufchan_buf[0])))
        lizzieLet58_3Lcall_$wnnz3_bufchan_buf <= lizzieLet58_3Lcall_$wnnz3_bufchan_d;
  
  /* demux (Ty CT$wnnz,
       Ty Int#) : (lizzieLet58_4,CT$wnnz) (srtarg_0_goMux_mux,Int#) > [(lizzieLet58_4L$wnnzsbos,Int#),
                                                                       (lizzieLet58_4Lcall_$wnnz3,Int#),
                                                                       (lizzieLet58_4Lcall_$wnnz2,Int#),
                                                                       (lizzieLet58_4Lcall_$wnnz1,Int#),
                                                                       (lizzieLet58_4Lcall_$wnnz0,Int#)] */
  logic [4:0] srtarg_0_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet58_4_d[0] && srtarg_0_goMux_mux_d[0]))
      unique case (lizzieLet58_4_d[3:1])
        3'd0: srtarg_0_goMux_mux_onehotd = 5'd1;
        3'd1: srtarg_0_goMux_mux_onehotd = 5'd2;
        3'd2: srtarg_0_goMux_mux_onehotd = 5'd4;
        3'd3: srtarg_0_goMux_mux_onehotd = 5'd8;
        3'd4: srtarg_0_goMux_mux_onehotd = 5'd16;
        default: srtarg_0_goMux_mux_onehotd = 5'd0;
      endcase
    else srtarg_0_goMux_mux_onehotd = 5'd0;
  assign lizzieLet58_4L$wnnzsbos_d = {srtarg_0_goMux_mux_d[32:1],
                                      srtarg_0_goMux_mux_onehotd[0]};
  assign lizzieLet58_4Lcall_$wnnz3_d = {srtarg_0_goMux_mux_d[32:1],
                                        srtarg_0_goMux_mux_onehotd[1]};
  assign lizzieLet58_4Lcall_$wnnz2_d = {srtarg_0_goMux_mux_d[32:1],
                                        srtarg_0_goMux_mux_onehotd[2]};
  assign lizzieLet58_4Lcall_$wnnz1_d = {srtarg_0_goMux_mux_d[32:1],
                                        srtarg_0_goMux_mux_onehotd[3]};
  assign lizzieLet58_4Lcall_$wnnz0_d = {srtarg_0_goMux_mux_d[32:1],
                                        srtarg_0_goMux_mux_onehotd[4]};
  assign srtarg_0_goMux_mux_r = (| (srtarg_0_goMux_mux_onehotd & {lizzieLet58_4Lcall_$wnnz0_r,
                                                                  lizzieLet58_4Lcall_$wnnz1_r,
                                                                  lizzieLet58_4Lcall_$wnnz2_r,
                                                                  lizzieLet58_4Lcall_$wnnz3_r,
                                                                  lizzieLet58_4L$wnnzsbos_r}));
  assign lizzieLet58_4_r = srtarg_0_goMux_mux_r;
  
  /* fork (Ty Int#) : (lizzieLet58_4L$wnnzsbos,Int#) > [(lizzieLet58_4L$wnnzsbos_1_merge_merge_fork_1,Int#),
                                                   (lizzieLet58_4L$wnnzsbos_1_merge_merge_fork_2,Int#)] */
  logic [1:0] lizzieLet58_4L$wnnzsbos_emitted;
  logic [1:0] lizzieLet58_4L$wnnzsbos_done;
  assign lizzieLet58_4L$wnnzsbos_1_merge_merge_fork_1_d = {lizzieLet58_4L$wnnzsbos_d[32:1],
                                                           (lizzieLet58_4L$wnnzsbos_d[0] && (! lizzieLet58_4L$wnnzsbos_emitted[0]))};
  assign lizzieLet58_4L$wnnzsbos_1_merge_merge_fork_2_d = {lizzieLet58_4L$wnnzsbos_d[32:1],
                                                           (lizzieLet58_4L$wnnzsbos_d[0] && (! lizzieLet58_4L$wnnzsbos_emitted[1]))};
  assign lizzieLet58_4L$wnnzsbos_done = (lizzieLet58_4L$wnnzsbos_emitted | ({lizzieLet58_4L$wnnzsbos_1_merge_merge_fork_2_d[0],
                                                                             lizzieLet58_4L$wnnzsbos_1_merge_merge_fork_1_d[0]} & {lizzieLet58_4L$wnnzsbos_1_merge_merge_fork_2_r,
                                                                                                                                   lizzieLet58_4L$wnnzsbos_1_merge_merge_fork_1_r}));
  assign lizzieLet58_4L$wnnzsbos_r = (& lizzieLet58_4L$wnnzsbos_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet58_4L$wnnzsbos_emitted <= 2'd0;
    else
      lizzieLet58_4L$wnnzsbos_emitted <= (lizzieLet58_4L$wnnzsbos_r ? 2'd0 :
                                          lizzieLet58_4L$wnnzsbos_done);
  
  /* togo (Ty Int#) : (lizzieLet58_4L$wnnzsbos_1_merge_merge_fork_1,Int#) > (call_$wnnz_goConst,Go) */
  assign call_$wnnz_goConst_d = lizzieLet58_4L$wnnzsbos_1_merge_merge_fork_1_d[0];
  assign lizzieLet58_4L$wnnzsbos_1_merge_merge_fork_1_r = call_$wnnz_goConst_r;
  
  /* buf (Ty Int#) : (lizzieLet58_4L$wnnzsbos_1_merge_merge_fork_2,Int#) > ($wnnz_resbuf,Int#) */
  \Int#_t  lizzieLet58_4L$wnnzsbos_1_merge_merge_fork_2_bufchan_d;
  logic lizzieLet58_4L$wnnzsbos_1_merge_merge_fork_2_bufchan_r;
  assign lizzieLet58_4L$wnnzsbos_1_merge_merge_fork_2_r = ((! lizzieLet58_4L$wnnzsbos_1_merge_merge_fork_2_bufchan_d[0]) || lizzieLet58_4L$wnnzsbos_1_merge_merge_fork_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet58_4L$wnnzsbos_1_merge_merge_fork_2_bufchan_d <= {32'd0,
                                                                 1'd0};
    else
      if (lizzieLet58_4L$wnnzsbos_1_merge_merge_fork_2_r)
        lizzieLet58_4L$wnnzsbos_1_merge_merge_fork_2_bufchan_d <= lizzieLet58_4L$wnnzsbos_1_merge_merge_fork_2_d;
  \Int#_t  lizzieLet58_4L$wnnzsbos_1_merge_merge_fork_2_bufchan_buf;
  assign lizzieLet58_4L$wnnzsbos_1_merge_merge_fork_2_bufchan_r = (! lizzieLet58_4L$wnnzsbos_1_merge_merge_fork_2_bufchan_buf[0]);
  assign \$wnnz_resbuf_d  = (lizzieLet58_4L$wnnzsbos_1_merge_merge_fork_2_bufchan_buf[0] ? lizzieLet58_4L$wnnzsbos_1_merge_merge_fork_2_bufchan_buf :
                             lizzieLet58_4L$wnnzsbos_1_merge_merge_fork_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet58_4L$wnnzsbos_1_merge_merge_fork_2_bufchan_buf <= {32'd0,
                                                                   1'd0};
    else
      if ((\$wnnz_resbuf_r  && lizzieLet58_4L$wnnzsbos_1_merge_merge_fork_2_bufchan_buf[0]))
        lizzieLet58_4L$wnnzsbos_1_merge_merge_fork_2_bufchan_buf <= {32'd0,
                                                                     1'd0};
      else if (((! \$wnnz_resbuf_r ) && (! lizzieLet58_4L$wnnzsbos_1_merge_merge_fork_2_bufchan_buf[0])))
        lizzieLet58_4L$wnnzsbos_1_merge_merge_fork_2_bufchan_buf <= lizzieLet58_4L$wnnzsbos_1_merge_merge_fork_2_bufchan_d;
  
  /* dcon (Ty CT$wnnz,
      Dcon Lcall_$wnnz2) : [(lizzieLet58_4Lcall_$wnnz3,Int#),
                            (sc_0_3_destruct,Pointer_CT$wnnz),
                            (q4a8u_1_destruct,Pointer_QTree_Int),
                            (q3a8t_1_destruct,Pointer_QTree_Int)] > (lizzieLet58_4Lcall_$wnnz3_1sc_0_3_1q4a8u_1_1q3a8t_1_1Lcall_$wnnz2,CT$wnnz) */
  assign lizzieLet58_4Lcall_$wnnz3_1sc_0_3_1q4a8u_1_1q3a8t_1_1Lcall_$wnnz2_d = Lcall_$wnnz2_dc((& {lizzieLet58_4Lcall_$wnnz3_d[0],
                                                                                                   sc_0_3_destruct_d[0],
                                                                                                   q4a8u_1_destruct_d[0],
                                                                                                   q3a8t_1_destruct_d[0]}), lizzieLet58_4Lcall_$wnnz3_d, sc_0_3_destruct_d, q4a8u_1_destruct_d, q3a8t_1_destruct_d);
  assign {lizzieLet58_4Lcall_$wnnz3_r,
          sc_0_3_destruct_r,
          q4a8u_1_destruct_r,
          q3a8t_1_destruct_r} = {4 {(lizzieLet58_4Lcall_$wnnz3_1sc_0_3_1q4a8u_1_1q3a8t_1_1Lcall_$wnnz2_r && lizzieLet58_4Lcall_$wnnz3_1sc_0_3_1q4a8u_1_1q3a8t_1_1Lcall_$wnnz2_d[0])}};
  
  /* buf (Ty CT$wnnz) : (lizzieLet58_4Lcall_$wnnz3_1sc_0_3_1q4a8u_1_1q3a8t_1_1Lcall_$wnnz2,CT$wnnz) > (lizzieLet59_1_argbuf,CT$wnnz) */
  CT$wnnz_t lizzieLet58_4Lcall_$wnnz3_1sc_0_3_1q4a8u_1_1q3a8t_1_1Lcall_$wnnz2_bufchan_d;
  logic lizzieLet58_4Lcall_$wnnz3_1sc_0_3_1q4a8u_1_1q3a8t_1_1Lcall_$wnnz2_bufchan_r;
  assign lizzieLet58_4Lcall_$wnnz3_1sc_0_3_1q4a8u_1_1q3a8t_1_1Lcall_$wnnz2_r = ((! lizzieLet58_4Lcall_$wnnz3_1sc_0_3_1q4a8u_1_1q3a8t_1_1Lcall_$wnnz2_bufchan_d[0]) || lizzieLet58_4Lcall_$wnnz3_1sc_0_3_1q4a8u_1_1q3a8t_1_1Lcall_$wnnz2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet58_4Lcall_$wnnz3_1sc_0_3_1q4a8u_1_1q3a8t_1_1Lcall_$wnnz2_bufchan_d <= {115'd0,
                                                                                      1'd0};
    else
      if (lizzieLet58_4Lcall_$wnnz3_1sc_0_3_1q4a8u_1_1q3a8t_1_1Lcall_$wnnz2_r)
        lizzieLet58_4Lcall_$wnnz3_1sc_0_3_1q4a8u_1_1q3a8t_1_1Lcall_$wnnz2_bufchan_d <= lizzieLet58_4Lcall_$wnnz3_1sc_0_3_1q4a8u_1_1q3a8t_1_1Lcall_$wnnz2_d;
  CT$wnnz_t lizzieLet58_4Lcall_$wnnz3_1sc_0_3_1q4a8u_1_1q3a8t_1_1Lcall_$wnnz2_bufchan_buf;
  assign lizzieLet58_4Lcall_$wnnz3_1sc_0_3_1q4a8u_1_1q3a8t_1_1Lcall_$wnnz2_bufchan_r = (! lizzieLet58_4Lcall_$wnnz3_1sc_0_3_1q4a8u_1_1q3a8t_1_1Lcall_$wnnz2_bufchan_buf[0]);
  assign lizzieLet59_1_argbuf_d = (lizzieLet58_4Lcall_$wnnz3_1sc_0_3_1q4a8u_1_1q3a8t_1_1Lcall_$wnnz2_bufchan_buf[0] ? lizzieLet58_4Lcall_$wnnz3_1sc_0_3_1q4a8u_1_1q3a8t_1_1Lcall_$wnnz2_bufchan_buf :
                                   lizzieLet58_4Lcall_$wnnz3_1sc_0_3_1q4a8u_1_1q3a8t_1_1Lcall_$wnnz2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet58_4Lcall_$wnnz3_1sc_0_3_1q4a8u_1_1q3a8t_1_1Lcall_$wnnz2_bufchan_buf <= {115'd0,
                                                                                        1'd0};
    else
      if ((lizzieLet59_1_argbuf_r && lizzieLet58_4Lcall_$wnnz3_1sc_0_3_1q4a8u_1_1q3a8t_1_1Lcall_$wnnz2_bufchan_buf[0]))
        lizzieLet58_4Lcall_$wnnz3_1sc_0_3_1q4a8u_1_1q3a8t_1_1Lcall_$wnnz2_bufchan_buf <= {115'd0,
                                                                                          1'd0};
      else if (((! lizzieLet59_1_argbuf_r) && (! lizzieLet58_4Lcall_$wnnz3_1sc_0_3_1q4a8u_1_1q3a8t_1_1Lcall_$wnnz2_bufchan_buf[0])))
        lizzieLet58_4Lcall_$wnnz3_1sc_0_3_1q4a8u_1_1q3a8t_1_1Lcall_$wnnz2_bufchan_buf <= lizzieLet58_4Lcall_$wnnz3_1sc_0_3_1q4a8u_1_1q3a8t_1_1Lcall_$wnnz2_bufchan_d;
  
  /* destruct (Ty CTf''''''''''''_f''''''''''''_Int,
          Dcon Lcall_f''''''''''''_f''''''''''''_Int0) : (lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int0,CTf''''''''''''_f''''''''''''_Int) > [(es_5_2_destruct,Pointer_QTree_Int),
                                                                                                                                                    (es_6_4_destruct,Pointer_QTree_Int),
                                                                                                                                                    (es_7_3_destruct,Pointer_QTree_Int),
                                                                                                                                                    (sc_0_10_destruct,Pointer_CTf''''''''''''_f''''''''''''_Int)] */
  logic [3:0] \lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int0_emitted ;
  logic [3:0] \lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int0_done ;
  assign es_5_2_destruct_d = {\lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int0_d [19:4],
                              (\lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int0_d [0] && (! \lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int0_emitted [0]))};
  assign es_6_4_destruct_d = {\lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int0_d [35:20],
                              (\lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int0_d [0] && (! \lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int0_emitted [1]))};
  assign es_7_3_destruct_d = {\lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int0_d [51:36],
                              (\lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int0_d [0] && (! \lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int0_emitted [2]))};
  assign sc_0_10_destruct_d = {\lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int0_d [67:52],
                               (\lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int0_d [0] && (! \lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int0_emitted [3]))};
  assign \lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int0_done  = (\lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int0_emitted  | ({sc_0_10_destruct_d[0],
                                                                                                                                         es_7_3_destruct_d[0],
                                                                                                                                         es_6_4_destruct_d[0],
                                                                                                                                         es_5_2_destruct_d[0]} & {sc_0_10_destruct_r,
                                                                                                                                                                  es_7_3_destruct_r,
                                                                                                                                                                  es_6_4_destruct_r,
                                                                                                                                                                  es_5_2_destruct_r}));
  assign \lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int0_r  = (& \lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int0_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int0_emitted  <= 4'd0;
    else
      \lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int0_emitted  <= (\lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int0_r  ? 4'd0 :
                                                                        \lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int0_done );
  
  /* destruct (Ty CTf''''''''''''_f''''''''''''_Int,
          Dcon Lcall_f''''''''''''_f''''''''''''_Int1) : (lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int1,CTf''''''''''''_f''''''''''''_Int) > [(es_6_3_destruct,Pointer_QTree_Int),
                                                                                                                                                    (es_7_2_destruct,Pointer_QTree_Int),
                                                                                                                                                    (sc_0_9_destruct,Pointer_CTf''''''''''''_f''''''''''''_Int),
                                                                                                                                                    (q1aft_3_destruct,Pointer_QTree_Int),
                                                                                                                                                    (t1afy_3_destruct,Pointer_QTree_Int),
                                                                                                                                                    (is_zafl_4_destruct,MyDTInt_Bool),
                                                                                                                                                    (op_addafm_4_destruct,MyDTInt_Int_Int)] */
  logic [6:0] \lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int1_emitted ;
  logic [6:0] \lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int1_done ;
  assign es_6_3_destruct_d = {\lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int1_d [19:4],
                              (\lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int1_d [0] && (! \lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int1_emitted [0]))};
  assign es_7_2_destruct_d = {\lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int1_d [35:20],
                              (\lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int1_d [0] && (! \lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int1_emitted [1]))};
  assign sc_0_9_destruct_d = {\lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int1_d [51:36],
                              (\lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int1_d [0] && (! \lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int1_emitted [2]))};
  assign q1aft_3_destruct_d = {\lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int1_d [67:52],
                               (\lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int1_d [0] && (! \lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int1_emitted [3]))};
  assign t1afy_3_destruct_d = {\lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int1_d [83:68],
                               (\lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int1_d [0] && (! \lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int1_emitted [4]))};
  assign is_zafl_4_destruct_d = (\lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int1_d [0] && (! \lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int1_emitted [5]));
  assign op_addafm_4_destruct_d = (\lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int1_d [0] && (! \lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int1_emitted [6]));
  assign \lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int1_done  = (\lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int1_emitted  | ({op_addafm_4_destruct_d[0],
                                                                                                                                         is_zafl_4_destruct_d[0],
                                                                                                                                         t1afy_3_destruct_d[0],
                                                                                                                                         q1aft_3_destruct_d[0],
                                                                                                                                         sc_0_9_destruct_d[0],
                                                                                                                                         es_7_2_destruct_d[0],
                                                                                                                                         es_6_3_destruct_d[0]} & {op_addafm_4_destruct_r,
                                                                                                                                                                  is_zafl_4_destruct_r,
                                                                                                                                                                  t1afy_3_destruct_r,
                                                                                                                                                                  q1aft_3_destruct_r,
                                                                                                                                                                  sc_0_9_destruct_r,
                                                                                                                                                                  es_7_2_destruct_r,
                                                                                                                                                                  es_6_3_destruct_r}));
  assign \lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int1_r  = (& \lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int1_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int1_emitted  <= 7'd0;
    else
      \lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int1_emitted  <= (\lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int1_r  ? 7'd0 :
                                                                        \lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int1_done );
  
  /* destruct (Ty CTf''''''''''''_f''''''''''''_Int,
          Dcon Lcall_f''''''''''''_f''''''''''''_Int2) : (lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int2,CTf''''''''''''_f''''''''''''_Int) > [(es_7_1_destruct,Pointer_QTree_Int),
                                                                                                                                                    (sc_0_8_destruct,Pointer_CTf''''''''''''_f''''''''''''_Int),
                                                                                                                                                    (q1aft_2_destruct,Pointer_QTree_Int),
                                                                                                                                                    (t1afy_2_destruct,Pointer_QTree_Int),
                                                                                                                                                    (is_zafl_3_destruct,MyDTInt_Bool),
                                                                                                                                                    (op_addafm_3_destruct,MyDTInt_Int_Int),
                                                                                                                                                    (q2afu_2_destruct,Pointer_QTree_Int),
                                                                                                                                                    (t2afz_2_destruct,Pointer_QTree_Int)] */
  logic [7:0] \lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int2_emitted ;
  logic [7:0] \lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int2_done ;
  assign es_7_1_destruct_d = {\lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int2_d [19:4],
                              (\lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int2_d [0] && (! \lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int2_emitted [0]))};
  assign sc_0_8_destruct_d = {\lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int2_d [35:20],
                              (\lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int2_d [0] && (! \lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int2_emitted [1]))};
  assign q1aft_2_destruct_d = {\lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int2_d [51:36],
                               (\lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int2_d [0] && (! \lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int2_emitted [2]))};
  assign t1afy_2_destruct_d = {\lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int2_d [67:52],
                               (\lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int2_d [0] && (! \lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int2_emitted [3]))};
  assign is_zafl_3_destruct_d = (\lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int2_d [0] && (! \lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int2_emitted [4]));
  assign op_addafm_3_destruct_d = (\lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int2_d [0] && (! \lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int2_emitted [5]));
  assign q2afu_2_destruct_d = {\lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int2_d [83:68],
                               (\lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int2_d [0] && (! \lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int2_emitted [6]))};
  assign t2afz_2_destruct_d = {\lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int2_d [99:84],
                               (\lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int2_d [0] && (! \lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int2_emitted [7]))};
  assign \lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int2_done  = (\lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int2_emitted  | ({t2afz_2_destruct_d[0],
                                                                                                                                         q2afu_2_destruct_d[0],
                                                                                                                                         op_addafm_3_destruct_d[0],
                                                                                                                                         is_zafl_3_destruct_d[0],
                                                                                                                                         t1afy_2_destruct_d[0],
                                                                                                                                         q1aft_2_destruct_d[0],
                                                                                                                                         sc_0_8_destruct_d[0],
                                                                                                                                         es_7_1_destruct_d[0]} & {t2afz_2_destruct_r,
                                                                                                                                                                  q2afu_2_destruct_r,
                                                                                                                                                                  op_addafm_3_destruct_r,
                                                                                                                                                                  is_zafl_3_destruct_r,
                                                                                                                                                                  t1afy_2_destruct_r,
                                                                                                                                                                  q1aft_2_destruct_r,
                                                                                                                                                                  sc_0_8_destruct_r,
                                                                                                                                                                  es_7_1_destruct_r}));
  assign \lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int2_r  = (& \lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int2_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int2_emitted  <= 8'd0;
    else
      \lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int2_emitted  <= (\lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int2_r  ? 8'd0 :
                                                                        \lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int2_done );
  
  /* destruct (Ty CTf''''''''''''_f''''''''''''_Int,
          Dcon Lcall_f''''''''''''_f''''''''''''_Int3) : (lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int3,CTf''''''''''''_f''''''''''''_Int) > [(sc_0_7_destruct,Pointer_CTf''''''''''''_f''''''''''''_Int),
                                                                                                                                                    (q1aft_1_destruct,Pointer_QTree_Int),
                                                                                                                                                    (t1afy_1_destruct,Pointer_QTree_Int),
                                                                                                                                                    (is_zafl_2_destruct,MyDTInt_Bool),
                                                                                                                                                    (op_addafm_2_destruct,MyDTInt_Int_Int),
                                                                                                                                                    (q2afu_1_destruct,Pointer_QTree_Int),
                                                                                                                                                    (t2afz_1_destruct,Pointer_QTree_Int),
                                                                                                                                                    (q3afv_1_destruct,Pointer_QTree_Int),
                                                                                                                                                    (t3afA_1_destruct,Pointer_QTree_Int)] */
  logic [8:0] \lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int3_emitted ;
  logic [8:0] \lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int3_done ;
  assign sc_0_7_destruct_d = {\lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int3_d [19:4],
                              (\lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int3_d [0] && (! \lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int3_emitted [0]))};
  assign q1aft_1_destruct_d = {\lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int3_d [35:20],
                               (\lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int3_d [0] && (! \lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int3_emitted [1]))};
  assign t1afy_1_destruct_d = {\lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int3_d [51:36],
                               (\lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int3_d [0] && (! \lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int3_emitted [2]))};
  assign is_zafl_2_destruct_d = (\lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int3_d [0] && (! \lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int3_emitted [3]));
  assign op_addafm_2_destruct_d = (\lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int3_d [0] && (! \lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int3_emitted [4]));
  assign q2afu_1_destruct_d = {\lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int3_d [67:52],
                               (\lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int3_d [0] && (! \lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int3_emitted [5]))};
  assign t2afz_1_destruct_d = {\lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int3_d [83:68],
                               (\lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int3_d [0] && (! \lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int3_emitted [6]))};
  assign q3afv_1_destruct_d = {\lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int3_d [99:84],
                               (\lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int3_d [0] && (! \lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int3_emitted [7]))};
  assign t3afA_1_destruct_d = {\lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int3_d [115:100],
                               (\lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int3_d [0] && (! \lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int3_emitted [8]))};
  assign \lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int3_done  = (\lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int3_emitted  | ({t3afA_1_destruct_d[0],
                                                                                                                                         q3afv_1_destruct_d[0],
                                                                                                                                         t2afz_1_destruct_d[0],
                                                                                                                                         q2afu_1_destruct_d[0],
                                                                                                                                         op_addafm_2_destruct_d[0],
                                                                                                                                         is_zafl_2_destruct_d[0],
                                                                                                                                         t1afy_1_destruct_d[0],
                                                                                                                                         q1aft_1_destruct_d[0],
                                                                                                                                         sc_0_7_destruct_d[0]} & {t3afA_1_destruct_r,
                                                                                                                                                                  q3afv_1_destruct_r,
                                                                                                                                                                  t2afz_1_destruct_r,
                                                                                                                                                                  q2afu_1_destruct_r,
                                                                                                                                                                  op_addafm_2_destruct_r,
                                                                                                                                                                  is_zafl_2_destruct_r,
                                                                                                                                                                  t1afy_1_destruct_r,
                                                                                                                                                                  q1aft_1_destruct_r,
                                                                                                                                                                  sc_0_7_destruct_r}));
  assign \lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int3_r  = (& \lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int3_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int3_emitted  <= 9'd0;
    else
      \lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int3_emitted  <= (\lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int3_r  ? 9'd0 :
                                                                        \lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int3_done );
  
  /* demux (Ty CTf''''''''''''_f''''''''''''_Int,
       Ty CTf''''''''''''_f''''''''''''_Int) : (lizzieLet62_2,CTf''''''''''''_f''''''''''''_Int) (lizzieLet62_1,CTf''''''''''''_f''''''''''''_Int) > [(_55,CTf''''''''''''_f''''''''''''_Int),
                                                                                                                                                      (lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int3,CTf''''''''''''_f''''''''''''_Int),
                                                                                                                                                      (lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int2,CTf''''''''''''_f''''''''''''_Int),
                                                                                                                                                      (lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int1,CTf''''''''''''_f''''''''''''_Int),
                                                                                                                                                      (lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int0,CTf''''''''''''_f''''''''''''_Int)] */
  logic [4:0] lizzieLet62_1_onehotd;
  always_comb
    if ((lizzieLet62_2_d[0] && lizzieLet62_1_d[0]))
      unique case (lizzieLet62_2_d[3:1])
        3'd0: lizzieLet62_1_onehotd = 5'd1;
        3'd1: lizzieLet62_1_onehotd = 5'd2;
        3'd2: lizzieLet62_1_onehotd = 5'd4;
        3'd3: lizzieLet62_1_onehotd = 5'd8;
        3'd4: lizzieLet62_1_onehotd = 5'd16;
        default: lizzieLet62_1_onehotd = 5'd0;
      endcase
    else lizzieLet62_1_onehotd = 5'd0;
  assign _55_d = {lizzieLet62_1_d[115:1], lizzieLet62_1_onehotd[0]};
  assign \lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int3_d  = {lizzieLet62_1_d[115:1],
                                                                    lizzieLet62_1_onehotd[1]};
  assign \lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int2_d  = {lizzieLet62_1_d[115:1],
                                                                    lizzieLet62_1_onehotd[2]};
  assign \lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int1_d  = {lizzieLet62_1_d[115:1],
                                                                    lizzieLet62_1_onehotd[3]};
  assign \lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int0_d  = {lizzieLet62_1_d[115:1],
                                                                    lizzieLet62_1_onehotd[4]};
  assign lizzieLet62_1_r = (| (lizzieLet62_1_onehotd & {\lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int0_r ,
                                                        \lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int1_r ,
                                                        \lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int2_r ,
                                                        \lizzieLet62_1Lcall_f''''''''''''_f''''''''''''_Int3_r ,
                                                        _55_r}));
  assign lizzieLet62_2_r = lizzieLet62_1_r;
  
  /* demux (Ty CTf''''''''''''_f''''''''''''_Int,
       Ty Go) : (lizzieLet62_3,CTf''''''''''''_f''''''''''''_Int) (go_14_goMux_data,Go) > [(_54,Go),
                                                                                           (lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int3,Go),
                                                                                           (lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int2,Go),
                                                                                           (lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int1,Go),
                                                                                           (lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int0,Go)] */
  logic [4:0] go_14_goMux_data_onehotd;
  always_comb
    if ((lizzieLet62_3_d[0] && go_14_goMux_data_d[0]))
      unique case (lizzieLet62_3_d[3:1])
        3'd0: go_14_goMux_data_onehotd = 5'd1;
        3'd1: go_14_goMux_data_onehotd = 5'd2;
        3'd2: go_14_goMux_data_onehotd = 5'd4;
        3'd3: go_14_goMux_data_onehotd = 5'd8;
        3'd4: go_14_goMux_data_onehotd = 5'd16;
        default: go_14_goMux_data_onehotd = 5'd0;
      endcase
    else go_14_goMux_data_onehotd = 5'd0;
  assign _54_d = go_14_goMux_data_onehotd[0];
  assign \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int3_d  = go_14_goMux_data_onehotd[1];
  assign \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int2_d  = go_14_goMux_data_onehotd[2];
  assign \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int1_d  = go_14_goMux_data_onehotd[3];
  assign \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int0_d  = go_14_goMux_data_onehotd[4];
  assign go_14_goMux_data_r = (| (go_14_goMux_data_onehotd & {\lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int0_r ,
                                                              \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int1_r ,
                                                              \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int2_r ,
                                                              \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int3_r ,
                                                              _54_r}));
  assign lizzieLet62_3_r = go_14_goMux_data_r;
  
  /* buf (Ty Go) : (lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int0,Go) > (lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int0_1_argbuf,Go) */
  Go_t \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int0_bufchan_d ;
  logic \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int0_bufchan_r ;
  assign \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int0_r  = ((! \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int0_bufchan_d [0]) || \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int0_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int0_bufchan_d  <= 1'd0;
    else
      if (\lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int0_r )
        \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int0_bufchan_d  <= \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int0_d ;
  Go_t \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int0_bufchan_buf ;
  assign \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int0_bufchan_r  = (! \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int0_bufchan_buf [0]);
  assign \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int0_1_argbuf_d  = (\lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int0_bufchan_buf [0] ? \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int0_bufchan_buf  :
                                                                             \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int0_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int0_bufchan_buf  <= 1'd0;
    else
      if ((\lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int0_1_argbuf_r  && \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int0_bufchan_buf [0]))
        \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int0_bufchan_buf  <= 1'd0;
      else if (((! \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int0_1_argbuf_r ) && (! \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int0_bufchan_buf [0])))
        \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int0_bufchan_buf  <= \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int0_bufchan_d ;
  
  /* buf (Ty Go) : (lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int1,Go) > (lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int1_1_argbuf,Go) */
  Go_t \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int1_bufchan_d ;
  logic \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int1_bufchan_r ;
  assign \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int1_r  = ((! \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int1_bufchan_d [0]) || \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int1_bufchan_d  <= 1'd0;
    else
      if (\lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int1_r )
        \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int1_bufchan_d  <= \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int1_d ;
  Go_t \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int1_bufchan_buf ;
  assign \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int1_bufchan_r  = (! \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int1_bufchan_buf [0]);
  assign \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int1_1_argbuf_d  = (\lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int1_bufchan_buf [0] ? \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int1_bufchan_buf  :
                                                                             \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int1_bufchan_buf  <= 1'd0;
    else
      if ((\lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int1_1_argbuf_r  && \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int1_bufchan_buf [0]))
        \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int1_bufchan_buf  <= 1'd0;
      else if (((! \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int1_1_argbuf_r ) && (! \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int1_bufchan_buf [0])))
        \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int1_bufchan_buf  <= \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int1_bufchan_d ;
  
  /* buf (Ty Go) : (lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int2,Go) > (lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int2_1_argbuf,Go) */
  Go_t \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int2_bufchan_d ;
  logic \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int2_bufchan_r ;
  assign \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int2_r  = ((! \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int2_bufchan_d [0]) || \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int2_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int2_bufchan_d  <= 1'd0;
    else
      if (\lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int2_r )
        \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int2_bufchan_d  <= \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int2_d ;
  Go_t \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int2_bufchan_buf ;
  assign \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int2_bufchan_r  = (! \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int2_bufchan_buf [0]);
  assign \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int2_1_argbuf_d  = (\lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int2_bufchan_buf [0] ? \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int2_bufchan_buf  :
                                                                             \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int2_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int2_bufchan_buf  <= 1'd0;
    else
      if ((\lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int2_1_argbuf_r  && \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int2_bufchan_buf [0]))
        \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int2_bufchan_buf  <= 1'd0;
      else if (((! \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int2_1_argbuf_r ) && (! \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int2_bufchan_buf [0])))
        \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int2_bufchan_buf  <= \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int2_bufchan_d ;
  
  /* buf (Ty Go) : (lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int3,Go) > (lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int3_1_argbuf,Go) */
  Go_t \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int3_bufchan_d ;
  logic \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int3_bufchan_r ;
  assign \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int3_r  = ((! \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int3_bufchan_d [0]) || \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int3_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int3_bufchan_d  <= 1'd0;
    else
      if (\lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int3_r )
        \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int3_bufchan_d  <= \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int3_d ;
  Go_t \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int3_bufchan_buf ;
  assign \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int3_bufchan_r  = (! \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int3_bufchan_buf [0]);
  assign \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int3_1_argbuf_d  = (\lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int3_bufchan_buf [0] ? \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int3_bufchan_buf  :
                                                                             \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int3_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int3_bufchan_buf  <= 1'd0;
    else
      if ((\lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int3_1_argbuf_r  && \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int3_bufchan_buf [0]))
        \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int3_bufchan_buf  <= 1'd0;
      else if (((! \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int3_1_argbuf_r ) && (! \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int3_bufchan_buf [0])))
        \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int3_bufchan_buf  <= \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int3_bufchan_d ;
  
  /* demux (Ty CTf''''''''''''_f''''''''''''_Int,
       Ty Pointer_QTree_Int) : (lizzieLet62_4,CTf''''''''''''_f''''''''''''_Int) (srtarg_0_1_goMux_mux,Pointer_QTree_Int) > [(lizzieLet62_4Lf''''''''''''_f''''''''''''_Intsbos,Pointer_QTree_Int),
                                                                                                                             (lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int3,Pointer_QTree_Int),
                                                                                                                             (lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int2,Pointer_QTree_Int),
                                                                                                                             (lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int1,Pointer_QTree_Int),
                                                                                                                             (lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int0,Pointer_QTree_Int)] */
  logic [4:0] srtarg_0_1_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet62_4_d[0] && srtarg_0_1_goMux_mux_d[0]))
      unique case (lizzieLet62_4_d[3:1])
        3'd0: srtarg_0_1_goMux_mux_onehotd = 5'd1;
        3'd1: srtarg_0_1_goMux_mux_onehotd = 5'd2;
        3'd2: srtarg_0_1_goMux_mux_onehotd = 5'd4;
        3'd3: srtarg_0_1_goMux_mux_onehotd = 5'd8;
        3'd4: srtarg_0_1_goMux_mux_onehotd = 5'd16;
        default: srtarg_0_1_goMux_mux_onehotd = 5'd0;
      endcase
    else srtarg_0_1_goMux_mux_onehotd = 5'd0;
  assign \lizzieLet62_4Lf''''''''''''_f''''''''''''_Intsbos_d  = {srtarg_0_1_goMux_mux_d[16:1],
                                                                  srtarg_0_1_goMux_mux_onehotd[0]};
  assign \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int3_d  = {srtarg_0_1_goMux_mux_d[16:1],
                                                                    srtarg_0_1_goMux_mux_onehotd[1]};
  assign \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int2_d  = {srtarg_0_1_goMux_mux_d[16:1],
                                                                    srtarg_0_1_goMux_mux_onehotd[2]};
  assign \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int1_d  = {srtarg_0_1_goMux_mux_d[16:1],
                                                                    srtarg_0_1_goMux_mux_onehotd[3]};
  assign \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int0_d  = {srtarg_0_1_goMux_mux_d[16:1],
                                                                    srtarg_0_1_goMux_mux_onehotd[4]};
  assign srtarg_0_1_goMux_mux_r = (| (srtarg_0_1_goMux_mux_onehotd & {\lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int0_r ,
                                                                      \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int1_r ,
                                                                      \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int2_r ,
                                                                      \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int3_r ,
                                                                      \lizzieLet62_4Lf''''''''''''_f''''''''''''_Intsbos_r }));
  assign lizzieLet62_4_r = srtarg_0_1_goMux_mux_r;
  
  /* dcon (Ty QTree_Int,
      Dcon QNode_Int) : [(lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int0,Pointer_QTree_Int),
                         (es_5_2_destruct,Pointer_QTree_Int),
                         (es_6_4_destruct,Pointer_QTree_Int),
                         (es_7_3_destruct,Pointer_QTree_Int)] > (lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int0_1es_5_2_1es_6_4_1es_7_3_1QNode_Int,QTree_Int) */
  assign \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int0_1es_5_2_1es_6_4_1es_7_3_1QNode_Int_d  = QNode_Int_dc((& {\lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int0_d [0],
                                                                                                                       es_5_2_destruct_d[0],
                                                                                                                       es_6_4_destruct_d[0],
                                                                                                                       es_7_3_destruct_d[0]}), \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int0_d , es_5_2_destruct_d, es_6_4_destruct_d, es_7_3_destruct_d);
  assign {\lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int0_r ,
          es_5_2_destruct_r,
          es_6_4_destruct_r,
          es_7_3_destruct_r} = {4 {(\lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int0_1es_5_2_1es_6_4_1es_7_3_1QNode_Int_r  && \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int0_1es_5_2_1es_6_4_1es_7_3_1QNode_Int_d [0])}};
  
  /* buf (Ty QTree_Int) : (lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int0_1es_5_2_1es_6_4_1es_7_3_1QNode_Int,QTree_Int) > (lizzieLet66_1_argbuf,QTree_Int) */
  QTree_Int_t \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int0_1es_5_2_1es_6_4_1es_7_3_1QNode_Int_bufchan_d ;
  logic \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int0_1es_5_2_1es_6_4_1es_7_3_1QNode_Int_bufchan_r ;
  assign \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int0_1es_5_2_1es_6_4_1es_7_3_1QNode_Int_r  = ((! \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int0_1es_5_2_1es_6_4_1es_7_3_1QNode_Int_bufchan_d [0]) || \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int0_1es_5_2_1es_6_4_1es_7_3_1QNode_Int_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int0_1es_5_2_1es_6_4_1es_7_3_1QNode_Int_bufchan_d  <= {66'd0,
                                                                                                             1'd0};
    else
      if (\lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int0_1es_5_2_1es_6_4_1es_7_3_1QNode_Int_r )
        \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int0_1es_5_2_1es_6_4_1es_7_3_1QNode_Int_bufchan_d  <= \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int0_1es_5_2_1es_6_4_1es_7_3_1QNode_Int_d ;
  QTree_Int_t \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int0_1es_5_2_1es_6_4_1es_7_3_1QNode_Int_bufchan_buf ;
  assign \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int0_1es_5_2_1es_6_4_1es_7_3_1QNode_Int_bufchan_r  = (! \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int0_1es_5_2_1es_6_4_1es_7_3_1QNode_Int_bufchan_buf [0]);
  assign lizzieLet66_1_argbuf_d = (\lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int0_1es_5_2_1es_6_4_1es_7_3_1QNode_Int_bufchan_buf [0] ? \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int0_1es_5_2_1es_6_4_1es_7_3_1QNode_Int_bufchan_buf  :
                                   \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int0_1es_5_2_1es_6_4_1es_7_3_1QNode_Int_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int0_1es_5_2_1es_6_4_1es_7_3_1QNode_Int_bufchan_buf  <= {66'd0,
                                                                                                               1'd0};
    else
      if ((lizzieLet66_1_argbuf_r && \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int0_1es_5_2_1es_6_4_1es_7_3_1QNode_Int_bufchan_buf [0]))
        \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int0_1es_5_2_1es_6_4_1es_7_3_1QNode_Int_bufchan_buf  <= {66'd0,
                                                                                                                 1'd0};
      else if (((! lizzieLet66_1_argbuf_r) && (! \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int0_1es_5_2_1es_6_4_1es_7_3_1QNode_Int_bufchan_buf [0])))
        \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int0_1es_5_2_1es_6_4_1es_7_3_1QNode_Int_bufchan_buf  <= \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int0_1es_5_2_1es_6_4_1es_7_3_1QNode_Int_bufchan_d ;
  
  /* dcon (Ty CTf''''''''''''_f''''''''''''_Int,
      Dcon Lcall_f''''''''''''_f''''''''''''_Int0) : [(lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int1,Pointer_QTree_Int),
                                                      (es_6_3_destruct,Pointer_QTree_Int),
                                                      (es_7_2_destruct,Pointer_QTree_Int),
                                                      (sc_0_9_destruct,Pointer_CTf''''''''''''_f''''''''''''_Int)] > (lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int1_1es_6_3_1es_7_2_1sc_0_9_1Lcall_f''''''''''''_f''''''''''''_Int0,CTf''''''''''''_f''''''''''''_Int) */
  assign \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int1_1es_6_3_1es_7_2_1sc_0_9_1Lcall_f''''''''''''_f''''''''''''_Int0_d  = \Lcall_f''''''''''''_f''''''''''''_Int0_dc ((& {\lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int1_d [0],
                                                                                                                                                                                   es_6_3_destruct_d[0],
                                                                                                                                                                                   es_7_2_destruct_d[0],
                                                                                                                                                                                   sc_0_9_destruct_d[0]}), \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int1_d , es_6_3_destruct_d, es_7_2_destruct_d, sc_0_9_destruct_d);
  assign {\lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int1_r ,
          es_6_3_destruct_r,
          es_7_2_destruct_r,
          sc_0_9_destruct_r} = {4 {(\lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int1_1es_6_3_1es_7_2_1sc_0_9_1Lcall_f''''''''''''_f''''''''''''_Int0_r  && \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int1_1es_6_3_1es_7_2_1sc_0_9_1Lcall_f''''''''''''_f''''''''''''_Int0_d [0])}};
  
  /* buf (Ty CTf''''''''''''_f''''''''''''_Int) : (lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int1_1es_6_3_1es_7_2_1sc_0_9_1Lcall_f''''''''''''_f''''''''''''_Int0,CTf''''''''''''_f''''''''''''_Int) > (lizzieLet65_1_argbuf,CTf''''''''''''_f''''''''''''_Int) */
  \CTf''''''''''''_f''''''''''''_Int_t  \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int1_1es_6_3_1es_7_2_1sc_0_9_1Lcall_f''''''''''''_f''''''''''''_Int0_bufchan_d ;
  logic \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int1_1es_6_3_1es_7_2_1sc_0_9_1Lcall_f''''''''''''_f''''''''''''_Int0_bufchan_r ;
  assign \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int1_1es_6_3_1es_7_2_1sc_0_9_1Lcall_f''''''''''''_f''''''''''''_Int0_r  = ((! \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int1_1es_6_3_1es_7_2_1sc_0_9_1Lcall_f''''''''''''_f''''''''''''_Int0_bufchan_d [0]) || \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int1_1es_6_3_1es_7_2_1sc_0_9_1Lcall_f''''''''''''_f''''''''''''_Int0_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int1_1es_6_3_1es_7_2_1sc_0_9_1Lcall_f''''''''''''_f''''''''''''_Int0_bufchan_d  <= {115'd0,
                                                                                                                                          1'd0};
    else
      if (\lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int1_1es_6_3_1es_7_2_1sc_0_9_1Lcall_f''''''''''''_f''''''''''''_Int0_r )
        \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int1_1es_6_3_1es_7_2_1sc_0_9_1Lcall_f''''''''''''_f''''''''''''_Int0_bufchan_d  <= \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int1_1es_6_3_1es_7_2_1sc_0_9_1Lcall_f''''''''''''_f''''''''''''_Int0_d ;
  \CTf''''''''''''_f''''''''''''_Int_t  \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int1_1es_6_3_1es_7_2_1sc_0_9_1Lcall_f''''''''''''_f''''''''''''_Int0_bufchan_buf ;
  assign \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int1_1es_6_3_1es_7_2_1sc_0_9_1Lcall_f''''''''''''_f''''''''''''_Int0_bufchan_r  = (! \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int1_1es_6_3_1es_7_2_1sc_0_9_1Lcall_f''''''''''''_f''''''''''''_Int0_bufchan_buf [0]);
  assign lizzieLet65_1_argbuf_d = (\lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int1_1es_6_3_1es_7_2_1sc_0_9_1Lcall_f''''''''''''_f''''''''''''_Int0_bufchan_buf [0] ? \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int1_1es_6_3_1es_7_2_1sc_0_9_1Lcall_f''''''''''''_f''''''''''''_Int0_bufchan_buf  :
                                   \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int1_1es_6_3_1es_7_2_1sc_0_9_1Lcall_f''''''''''''_f''''''''''''_Int0_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int1_1es_6_3_1es_7_2_1sc_0_9_1Lcall_f''''''''''''_f''''''''''''_Int0_bufchan_buf  <= {115'd0,
                                                                                                                                            1'd0};
    else
      if ((lizzieLet65_1_argbuf_r && \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int1_1es_6_3_1es_7_2_1sc_0_9_1Lcall_f''''''''''''_f''''''''''''_Int0_bufchan_buf [0]))
        \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int1_1es_6_3_1es_7_2_1sc_0_9_1Lcall_f''''''''''''_f''''''''''''_Int0_bufchan_buf  <= {115'd0,
                                                                                                                                              1'd0};
      else if (((! lizzieLet65_1_argbuf_r) && (! \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int1_1es_6_3_1es_7_2_1sc_0_9_1Lcall_f''''''''''''_f''''''''''''_Int0_bufchan_buf [0])))
        \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int1_1es_6_3_1es_7_2_1sc_0_9_1Lcall_f''''''''''''_f''''''''''''_Int0_bufchan_buf  <= \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int1_1es_6_3_1es_7_2_1sc_0_9_1Lcall_f''''''''''''_f''''''''''''_Int0_bufchan_d ;
  
  /* dcon (Ty CTf''''''''''''_f''''''''''''_Int,
      Dcon Lcall_f''''''''''''_f''''''''''''_Int1) : [(lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int2,Pointer_QTree_Int),
                                                      (es_7_1_destruct,Pointer_QTree_Int),
                                                      (sc_0_8_destruct,Pointer_CTf''''''''''''_f''''''''''''_Int),
                                                      (q1aft_2_destruct,Pointer_QTree_Int),
                                                      (t1afy_2_destruct,Pointer_QTree_Int),
                                                      (is_zafl_3_1,MyDTInt_Bool),
                                                      (op_addafm_3_1,MyDTInt_Int_Int)] > (lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int2_1es_7_1_1sc_0_8_1q1aft_2_1t1afy_2_1is_zafl_3_1op_addafm_3_1Lcall_f''''''''''''_f''''''''''''_Int1,CTf''''''''''''_f''''''''''''_Int) */
  assign \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int2_1es_7_1_1sc_0_8_1q1aft_2_1t1afy_2_1is_zafl_3_1op_addafm_3_1Lcall_f''''''''''''_f''''''''''''_Int1_d  = \Lcall_f''''''''''''_f''''''''''''_Int1_dc ((& {\lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int2_d [0],
                                                                                                                                                                                                                     es_7_1_destruct_d[0],
                                                                                                                                                                                                                     sc_0_8_destruct_d[0],
                                                                                                                                                                                                                     q1aft_2_destruct_d[0],
                                                                                                                                                                                                                     t1afy_2_destruct_d[0],
                                                                                                                                                                                                                     is_zafl_3_1_d[0],
                                                                                                                                                                                                                     op_addafm_3_1_d[0]}), \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int2_d , es_7_1_destruct_d, sc_0_8_destruct_d, q1aft_2_destruct_d, t1afy_2_destruct_d, is_zafl_3_1_d, op_addafm_3_1_d);
  assign {\lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int2_r ,
          es_7_1_destruct_r,
          sc_0_8_destruct_r,
          q1aft_2_destruct_r,
          t1afy_2_destruct_r,
          is_zafl_3_1_r,
          op_addafm_3_1_r} = {7 {(\lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int2_1es_7_1_1sc_0_8_1q1aft_2_1t1afy_2_1is_zafl_3_1op_addafm_3_1Lcall_f''''''''''''_f''''''''''''_Int1_r  && \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int2_1es_7_1_1sc_0_8_1q1aft_2_1t1afy_2_1is_zafl_3_1op_addafm_3_1Lcall_f''''''''''''_f''''''''''''_Int1_d [0])}};
  
  /* buf (Ty CTf''''''''''''_f''''''''''''_Int) : (lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int2_1es_7_1_1sc_0_8_1q1aft_2_1t1afy_2_1is_zafl_3_1op_addafm_3_1Lcall_f''''''''''''_f''''''''''''_Int1,CTf''''''''''''_f''''''''''''_Int) > (lizzieLet64_1_argbuf,CTf''''''''''''_f''''''''''''_Int) */
  \CTf''''''''''''_f''''''''''''_Int_t  \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int2_1es_7_1_1sc_0_8_1q1aft_2_1t1afy_2_1is_zafl_3_1op_addafm_3_1Lcall_f''''''''''''_f''''''''''''_Int1_bufchan_d ;
  logic \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int2_1es_7_1_1sc_0_8_1q1aft_2_1t1afy_2_1is_zafl_3_1op_addafm_3_1Lcall_f''''''''''''_f''''''''''''_Int1_bufchan_r ;
  assign \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int2_1es_7_1_1sc_0_8_1q1aft_2_1t1afy_2_1is_zafl_3_1op_addafm_3_1Lcall_f''''''''''''_f''''''''''''_Int1_r  = ((! \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int2_1es_7_1_1sc_0_8_1q1aft_2_1t1afy_2_1is_zafl_3_1op_addafm_3_1Lcall_f''''''''''''_f''''''''''''_Int1_bufchan_d [0]) || \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int2_1es_7_1_1sc_0_8_1q1aft_2_1t1afy_2_1is_zafl_3_1op_addafm_3_1Lcall_f''''''''''''_f''''''''''''_Int1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int2_1es_7_1_1sc_0_8_1q1aft_2_1t1afy_2_1is_zafl_3_1op_addafm_3_1Lcall_f''''''''''''_f''''''''''''_Int1_bufchan_d  <= {115'd0,
                                                                                                                                                                            1'd0};
    else
      if (\lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int2_1es_7_1_1sc_0_8_1q1aft_2_1t1afy_2_1is_zafl_3_1op_addafm_3_1Lcall_f''''''''''''_f''''''''''''_Int1_r )
        \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int2_1es_7_1_1sc_0_8_1q1aft_2_1t1afy_2_1is_zafl_3_1op_addafm_3_1Lcall_f''''''''''''_f''''''''''''_Int1_bufchan_d  <= \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int2_1es_7_1_1sc_0_8_1q1aft_2_1t1afy_2_1is_zafl_3_1op_addafm_3_1Lcall_f''''''''''''_f''''''''''''_Int1_d ;
  \CTf''''''''''''_f''''''''''''_Int_t  \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int2_1es_7_1_1sc_0_8_1q1aft_2_1t1afy_2_1is_zafl_3_1op_addafm_3_1Lcall_f''''''''''''_f''''''''''''_Int1_bufchan_buf ;
  assign \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int2_1es_7_1_1sc_0_8_1q1aft_2_1t1afy_2_1is_zafl_3_1op_addafm_3_1Lcall_f''''''''''''_f''''''''''''_Int1_bufchan_r  = (! \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int2_1es_7_1_1sc_0_8_1q1aft_2_1t1afy_2_1is_zafl_3_1op_addafm_3_1Lcall_f''''''''''''_f''''''''''''_Int1_bufchan_buf [0]);
  assign lizzieLet64_1_argbuf_d = (\lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int2_1es_7_1_1sc_0_8_1q1aft_2_1t1afy_2_1is_zafl_3_1op_addafm_3_1Lcall_f''''''''''''_f''''''''''''_Int1_bufchan_buf [0] ? \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int2_1es_7_1_1sc_0_8_1q1aft_2_1t1afy_2_1is_zafl_3_1op_addafm_3_1Lcall_f''''''''''''_f''''''''''''_Int1_bufchan_buf  :
                                   \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int2_1es_7_1_1sc_0_8_1q1aft_2_1t1afy_2_1is_zafl_3_1op_addafm_3_1Lcall_f''''''''''''_f''''''''''''_Int1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int2_1es_7_1_1sc_0_8_1q1aft_2_1t1afy_2_1is_zafl_3_1op_addafm_3_1Lcall_f''''''''''''_f''''''''''''_Int1_bufchan_buf  <= {115'd0,
                                                                                                                                                                              1'd0};
    else
      if ((lizzieLet64_1_argbuf_r && \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int2_1es_7_1_1sc_0_8_1q1aft_2_1t1afy_2_1is_zafl_3_1op_addafm_3_1Lcall_f''''''''''''_f''''''''''''_Int1_bufchan_buf [0]))
        \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int2_1es_7_1_1sc_0_8_1q1aft_2_1t1afy_2_1is_zafl_3_1op_addafm_3_1Lcall_f''''''''''''_f''''''''''''_Int1_bufchan_buf  <= {115'd0,
                                                                                                                                                                                1'd0};
      else if (((! lizzieLet64_1_argbuf_r) && (! \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int2_1es_7_1_1sc_0_8_1q1aft_2_1t1afy_2_1is_zafl_3_1op_addafm_3_1Lcall_f''''''''''''_f''''''''''''_Int1_bufchan_buf [0])))
        \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int2_1es_7_1_1sc_0_8_1q1aft_2_1t1afy_2_1is_zafl_3_1op_addafm_3_1Lcall_f''''''''''''_f''''''''''''_Int1_bufchan_buf  <= \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int2_1es_7_1_1sc_0_8_1q1aft_2_1t1afy_2_1is_zafl_3_1op_addafm_3_1Lcall_f''''''''''''_f''''''''''''_Int1_bufchan_d ;
  
  /* dcon (Ty CTf''''''''''''_f''''''''''''_Int,
      Dcon Lcall_f''''''''''''_f''''''''''''_Int2) : [(lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int3,Pointer_QTree_Int),
                                                      (sc_0_7_destruct,Pointer_CTf''''''''''''_f''''''''''''_Int),
                                                      (q1aft_1_destruct,Pointer_QTree_Int),
                                                      (t1afy_1_destruct,Pointer_QTree_Int),
                                                      (is_zafl_2_1,MyDTInt_Bool),
                                                      (op_addafm_2_1,MyDTInt_Int_Int),
                                                      (q2afu_1_destruct,Pointer_QTree_Int),
                                                      (t2afz_1_destruct,Pointer_QTree_Int)] > (lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int3_1sc_0_7_1q1aft_1_1t1afy_1_1is_zafl_2_1op_addafm_2_1q2afu_1_1t2afz_1_1Lcall_f''''''''''''_f''''''''''''_Int2,CTf''''''''''''_f''''''''''''_Int) */
  assign \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int3_1sc_0_7_1q1aft_1_1t1afy_1_1is_zafl_2_1op_addafm_2_1q2afu_1_1t2afz_1_1Lcall_f''''''''''''_f''''''''''''_Int2_d  = \Lcall_f''''''''''''_f''''''''''''_Int2_dc ((& {\lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int3_d [0],
                                                                                                                                                                                                                               sc_0_7_destruct_d[0],
                                                                                                                                                                                                                               q1aft_1_destruct_d[0],
                                                                                                                                                                                                                               t1afy_1_destruct_d[0],
                                                                                                                                                                                                                               is_zafl_2_1_d[0],
                                                                                                                                                                                                                               op_addafm_2_1_d[0],
                                                                                                                                                                                                                               q2afu_1_destruct_d[0],
                                                                                                                                                                                                                               t2afz_1_destruct_d[0]}), \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int3_d , sc_0_7_destruct_d, q1aft_1_destruct_d, t1afy_1_destruct_d, is_zafl_2_1_d, op_addafm_2_1_d, q2afu_1_destruct_d, t2afz_1_destruct_d);
  assign {\lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int3_r ,
          sc_0_7_destruct_r,
          q1aft_1_destruct_r,
          t1afy_1_destruct_r,
          is_zafl_2_1_r,
          op_addafm_2_1_r,
          q2afu_1_destruct_r,
          t2afz_1_destruct_r} = {8 {(\lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int3_1sc_0_7_1q1aft_1_1t1afy_1_1is_zafl_2_1op_addafm_2_1q2afu_1_1t2afz_1_1Lcall_f''''''''''''_f''''''''''''_Int2_r  && \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int3_1sc_0_7_1q1aft_1_1t1afy_1_1is_zafl_2_1op_addafm_2_1q2afu_1_1t2afz_1_1Lcall_f''''''''''''_f''''''''''''_Int2_d [0])}};
  
  /* buf (Ty CTf''''''''''''_f''''''''''''_Int) : (lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int3_1sc_0_7_1q1aft_1_1t1afy_1_1is_zafl_2_1op_addafm_2_1q2afu_1_1t2afz_1_1Lcall_f''''''''''''_f''''''''''''_Int2,CTf''''''''''''_f''''''''''''_Int) > (lizzieLet63_1_argbuf,CTf''''''''''''_f''''''''''''_Int) */
  \CTf''''''''''''_f''''''''''''_Int_t  \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int3_1sc_0_7_1q1aft_1_1t1afy_1_1is_zafl_2_1op_addafm_2_1q2afu_1_1t2afz_1_1Lcall_f''''''''''''_f''''''''''''_Int2_bufchan_d ;
  logic \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int3_1sc_0_7_1q1aft_1_1t1afy_1_1is_zafl_2_1op_addafm_2_1q2afu_1_1t2afz_1_1Lcall_f''''''''''''_f''''''''''''_Int2_bufchan_r ;
  assign \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int3_1sc_0_7_1q1aft_1_1t1afy_1_1is_zafl_2_1op_addafm_2_1q2afu_1_1t2afz_1_1Lcall_f''''''''''''_f''''''''''''_Int2_r  = ((! \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int3_1sc_0_7_1q1aft_1_1t1afy_1_1is_zafl_2_1op_addafm_2_1q2afu_1_1t2afz_1_1Lcall_f''''''''''''_f''''''''''''_Int2_bufchan_d [0]) || \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int3_1sc_0_7_1q1aft_1_1t1afy_1_1is_zafl_2_1op_addafm_2_1q2afu_1_1t2afz_1_1Lcall_f''''''''''''_f''''''''''''_Int2_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int3_1sc_0_7_1q1aft_1_1t1afy_1_1is_zafl_2_1op_addafm_2_1q2afu_1_1t2afz_1_1Lcall_f''''''''''''_f''''''''''''_Int2_bufchan_d  <= {115'd0,
                                                                                                                                                                                      1'd0};
    else
      if (\lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int3_1sc_0_7_1q1aft_1_1t1afy_1_1is_zafl_2_1op_addafm_2_1q2afu_1_1t2afz_1_1Lcall_f''''''''''''_f''''''''''''_Int2_r )
        \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int3_1sc_0_7_1q1aft_1_1t1afy_1_1is_zafl_2_1op_addafm_2_1q2afu_1_1t2afz_1_1Lcall_f''''''''''''_f''''''''''''_Int2_bufchan_d  <= \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int3_1sc_0_7_1q1aft_1_1t1afy_1_1is_zafl_2_1op_addafm_2_1q2afu_1_1t2afz_1_1Lcall_f''''''''''''_f''''''''''''_Int2_d ;
  \CTf''''''''''''_f''''''''''''_Int_t  \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int3_1sc_0_7_1q1aft_1_1t1afy_1_1is_zafl_2_1op_addafm_2_1q2afu_1_1t2afz_1_1Lcall_f''''''''''''_f''''''''''''_Int2_bufchan_buf ;
  assign \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int3_1sc_0_7_1q1aft_1_1t1afy_1_1is_zafl_2_1op_addafm_2_1q2afu_1_1t2afz_1_1Lcall_f''''''''''''_f''''''''''''_Int2_bufchan_r  = (! \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int3_1sc_0_7_1q1aft_1_1t1afy_1_1is_zafl_2_1op_addafm_2_1q2afu_1_1t2afz_1_1Lcall_f''''''''''''_f''''''''''''_Int2_bufchan_buf [0]);
  assign lizzieLet63_1_argbuf_d = (\lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int3_1sc_0_7_1q1aft_1_1t1afy_1_1is_zafl_2_1op_addafm_2_1q2afu_1_1t2afz_1_1Lcall_f''''''''''''_f''''''''''''_Int2_bufchan_buf [0] ? \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int3_1sc_0_7_1q1aft_1_1t1afy_1_1is_zafl_2_1op_addafm_2_1q2afu_1_1t2afz_1_1Lcall_f''''''''''''_f''''''''''''_Int2_bufchan_buf  :
                                   \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int3_1sc_0_7_1q1aft_1_1t1afy_1_1is_zafl_2_1op_addafm_2_1q2afu_1_1t2afz_1_1Lcall_f''''''''''''_f''''''''''''_Int2_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int3_1sc_0_7_1q1aft_1_1t1afy_1_1is_zafl_2_1op_addafm_2_1q2afu_1_1t2afz_1_1Lcall_f''''''''''''_f''''''''''''_Int2_bufchan_buf  <= {115'd0,
                                                                                                                                                                                        1'd0};
    else
      if ((lizzieLet63_1_argbuf_r && \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int3_1sc_0_7_1q1aft_1_1t1afy_1_1is_zafl_2_1op_addafm_2_1q2afu_1_1t2afz_1_1Lcall_f''''''''''''_f''''''''''''_Int2_bufchan_buf [0]))
        \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int3_1sc_0_7_1q1aft_1_1t1afy_1_1is_zafl_2_1op_addafm_2_1q2afu_1_1t2afz_1_1Lcall_f''''''''''''_f''''''''''''_Int2_bufchan_buf  <= {115'd0,
                                                                                                                                                                                          1'd0};
      else if (((! lizzieLet63_1_argbuf_r) && (! \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int3_1sc_0_7_1q1aft_1_1t1afy_1_1is_zafl_2_1op_addafm_2_1q2afu_1_1t2afz_1_1Lcall_f''''''''''''_f''''''''''''_Int2_bufchan_buf [0])))
        \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int3_1sc_0_7_1q1aft_1_1t1afy_1_1is_zafl_2_1op_addafm_2_1q2afu_1_1t2afz_1_1Lcall_f''''''''''''_f''''''''''''_Int2_bufchan_buf  <= \lizzieLet62_4Lcall_f''''''''''''_f''''''''''''_Int3_1sc_0_7_1q1aft_1_1t1afy_1_1is_zafl_2_1op_addafm_2_1q2afu_1_1t2afz_1_1Lcall_f''''''''''''_f''''''''''''_Int2_bufchan_d ;
  
  /* fork (Ty Pointer_QTree_Int) : (lizzieLet62_4Lf''''''''''''_f''''''''''''_Intsbos,Pointer_QTree_Int) > [(lizzieLet62_4Lf''''''''''''_f''''''''''''_Intsbos_1_merge_merge_fork_1,Pointer_QTree_Int),
                                                                                                       (lizzieLet62_4Lf''''''''''''_f''''''''''''_Intsbos_1_merge_merge_fork_2,Pointer_QTree_Int)] */
  logic [1:0] \lizzieLet62_4Lf''''''''''''_f''''''''''''_Intsbos_emitted ;
  logic [1:0] \lizzieLet62_4Lf''''''''''''_f''''''''''''_Intsbos_done ;
  assign \lizzieLet62_4Lf''''''''''''_f''''''''''''_Intsbos_1_merge_merge_fork_1_d  = {\lizzieLet62_4Lf''''''''''''_f''''''''''''_Intsbos_d [16:1],
                                                                                       (\lizzieLet62_4Lf''''''''''''_f''''''''''''_Intsbos_d [0] && (! \lizzieLet62_4Lf''''''''''''_f''''''''''''_Intsbos_emitted [0]))};
  assign \lizzieLet62_4Lf''''''''''''_f''''''''''''_Intsbos_1_merge_merge_fork_2_d  = {\lizzieLet62_4Lf''''''''''''_f''''''''''''_Intsbos_d [16:1],
                                                                                       (\lizzieLet62_4Lf''''''''''''_f''''''''''''_Intsbos_d [0] && (! \lizzieLet62_4Lf''''''''''''_f''''''''''''_Intsbos_emitted [1]))};
  assign \lizzieLet62_4Lf''''''''''''_f''''''''''''_Intsbos_done  = (\lizzieLet62_4Lf''''''''''''_f''''''''''''_Intsbos_emitted  | ({\lizzieLet62_4Lf''''''''''''_f''''''''''''_Intsbos_1_merge_merge_fork_2_d [0],
                                                                                                                                     \lizzieLet62_4Lf''''''''''''_f''''''''''''_Intsbos_1_merge_merge_fork_1_d [0]} & {\lizzieLet62_4Lf''''''''''''_f''''''''''''_Intsbos_1_merge_merge_fork_2_r ,
                                                                                                                                                                                                                       \lizzieLet62_4Lf''''''''''''_f''''''''''''_Intsbos_1_merge_merge_fork_1_r }));
  assign \lizzieLet62_4Lf''''''''''''_f''''''''''''_Intsbos_r  = (& \lizzieLet62_4Lf''''''''''''_f''''''''''''_Intsbos_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet62_4Lf''''''''''''_f''''''''''''_Intsbos_emitted  <= 2'd0;
    else
      \lizzieLet62_4Lf''''''''''''_f''''''''''''_Intsbos_emitted  <= (\lizzieLet62_4Lf''''''''''''_f''''''''''''_Intsbos_r  ? 2'd0 :
                                                                      \lizzieLet62_4Lf''''''''''''_f''''''''''''_Intsbos_done );
  
  /* togo (Ty Pointer_QTree_Int) : (lizzieLet62_4Lf''''''''''''_f''''''''''''_Intsbos_1_merge_merge_fork_1,Pointer_QTree_Int) > (call_f''''''''''''_f''''''''''''_Int_goConst,Go) */
  assign \call_f''''''''''''_f''''''''''''_Int_goConst_d  = \lizzieLet62_4Lf''''''''''''_f''''''''''''_Intsbos_1_merge_merge_fork_1_d [0];
  assign \lizzieLet62_4Lf''''''''''''_f''''''''''''_Intsbos_1_merge_merge_fork_1_r  = \call_f''''''''''''_f''''''''''''_Int_goConst_r ;
  
  /* destruct (Ty CTf_f_Int,
          Dcon Lcall_f_f_Int0) : (lizzieLet67_1Lcall_f_f_Int0,CTf_f_Int) > [(es_35_destruct,Pointer_QTree_Int),
                                                                            (es_36_1_destruct,Pointer_QTree_Int),
                                                                            (es_37_2_destruct,Pointer_QTree_Int),
                                                                            (sc_0_14_destruct,Pointer_CTf_f_Int)] */
  logic [3:0] lizzieLet67_1Lcall_f_f_Int0_emitted;
  logic [3:0] lizzieLet67_1Lcall_f_f_Int0_done;
  assign es_35_destruct_d = {lizzieLet67_1Lcall_f_f_Int0_d[19:4],
                             (lizzieLet67_1Lcall_f_f_Int0_d[0] && (! lizzieLet67_1Lcall_f_f_Int0_emitted[0]))};
  assign es_36_1_destruct_d = {lizzieLet67_1Lcall_f_f_Int0_d[35:20],
                               (lizzieLet67_1Lcall_f_f_Int0_d[0] && (! lizzieLet67_1Lcall_f_f_Int0_emitted[1]))};
  assign es_37_2_destruct_d = {lizzieLet67_1Lcall_f_f_Int0_d[51:36],
                               (lizzieLet67_1Lcall_f_f_Int0_d[0] && (! lizzieLet67_1Lcall_f_f_Int0_emitted[2]))};
  assign sc_0_14_destruct_d = {lizzieLet67_1Lcall_f_f_Int0_d[67:52],
                               (lizzieLet67_1Lcall_f_f_Int0_d[0] && (! lizzieLet67_1Lcall_f_f_Int0_emitted[3]))};
  assign lizzieLet67_1Lcall_f_f_Int0_done = (lizzieLet67_1Lcall_f_f_Int0_emitted | ({sc_0_14_destruct_d[0],
                                                                                     es_37_2_destruct_d[0],
                                                                                     es_36_1_destruct_d[0],
                                                                                     es_35_destruct_d[0]} & {sc_0_14_destruct_r,
                                                                                                             es_37_2_destruct_r,
                                                                                                             es_36_1_destruct_r,
                                                                                                             es_35_destruct_r}));
  assign lizzieLet67_1Lcall_f_f_Int0_r = (& lizzieLet67_1Lcall_f_f_Int0_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet67_1Lcall_f_f_Int0_emitted <= 4'd0;
    else
      lizzieLet67_1Lcall_f_f_Int0_emitted <= (lizzieLet67_1Lcall_f_f_Int0_r ? 4'd0 :
                                              lizzieLet67_1Lcall_f_f_Int0_done);
  
  /* destruct (Ty CTf_f_Int,
          Dcon Lcall_f_f_Int1) : (lizzieLet67_1Lcall_f_f_Int1,CTf_f_Int) > [(es_36_destruct,Pointer_QTree_Int),
                                                                            (es_37_1_destruct,Pointer_QTree_Int),
                                                                            (sc_0_13_destruct,Pointer_CTf_f_Int),
                                                                            (q1af0_3_destruct,Pointer_QTree_Int),
                                                                            (t1afa_3_destruct,Pointer_QTree_Int),
                                                                            (t1'aff_3_destruct,Pointer_QTree_Int),
                                                                            (is_zaet_4_destruct,MyDTInt_Bool),
                                                                            (op_addaeu_4_destruct,MyDTInt_Int_Int)] */
  logic [7:0] lizzieLet67_1Lcall_f_f_Int1_emitted;
  logic [7:0] lizzieLet67_1Lcall_f_f_Int1_done;
  assign es_36_destruct_d = {lizzieLet67_1Lcall_f_f_Int1_d[19:4],
                             (lizzieLet67_1Lcall_f_f_Int1_d[0] && (! lizzieLet67_1Lcall_f_f_Int1_emitted[0]))};
  assign es_37_1_destruct_d = {lizzieLet67_1Lcall_f_f_Int1_d[35:20],
                               (lizzieLet67_1Lcall_f_f_Int1_d[0] && (! lizzieLet67_1Lcall_f_f_Int1_emitted[1]))};
  assign sc_0_13_destruct_d = {lizzieLet67_1Lcall_f_f_Int1_d[51:36],
                               (lizzieLet67_1Lcall_f_f_Int1_d[0] && (! lizzieLet67_1Lcall_f_f_Int1_emitted[2]))};
  assign q1af0_3_destruct_d = {lizzieLet67_1Lcall_f_f_Int1_d[67:52],
                               (lizzieLet67_1Lcall_f_f_Int1_d[0] && (! lizzieLet67_1Lcall_f_f_Int1_emitted[3]))};
  assign t1afa_3_destruct_d = {lizzieLet67_1Lcall_f_f_Int1_d[83:68],
                               (lizzieLet67_1Lcall_f_f_Int1_d[0] && (! lizzieLet67_1Lcall_f_f_Int1_emitted[4]))};
  assign \t1'aff_3_destruct_d  = {lizzieLet67_1Lcall_f_f_Int1_d[99:84],
                                  (lizzieLet67_1Lcall_f_f_Int1_d[0] && (! lizzieLet67_1Lcall_f_f_Int1_emitted[5]))};
  assign is_zaet_4_destruct_d = (lizzieLet67_1Lcall_f_f_Int1_d[0] && (! lizzieLet67_1Lcall_f_f_Int1_emitted[6]));
  assign op_addaeu_4_destruct_d = (lizzieLet67_1Lcall_f_f_Int1_d[0] && (! lizzieLet67_1Lcall_f_f_Int1_emitted[7]));
  assign lizzieLet67_1Lcall_f_f_Int1_done = (lizzieLet67_1Lcall_f_f_Int1_emitted | ({op_addaeu_4_destruct_d[0],
                                                                                     is_zaet_4_destruct_d[0],
                                                                                     \t1'aff_3_destruct_d [0],
                                                                                     t1afa_3_destruct_d[0],
                                                                                     q1af0_3_destruct_d[0],
                                                                                     sc_0_13_destruct_d[0],
                                                                                     es_37_1_destruct_d[0],
                                                                                     es_36_destruct_d[0]} & {op_addaeu_4_destruct_r,
                                                                                                             is_zaet_4_destruct_r,
                                                                                                             \t1'aff_3_destruct_r ,
                                                                                                             t1afa_3_destruct_r,
                                                                                                             q1af0_3_destruct_r,
                                                                                                             sc_0_13_destruct_r,
                                                                                                             es_37_1_destruct_r,
                                                                                                             es_36_destruct_r}));
  assign lizzieLet67_1Lcall_f_f_Int1_r = (& lizzieLet67_1Lcall_f_f_Int1_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet67_1Lcall_f_f_Int1_emitted <= 8'd0;
    else
      lizzieLet67_1Lcall_f_f_Int1_emitted <= (lizzieLet67_1Lcall_f_f_Int1_r ? 8'd0 :
                                              lizzieLet67_1Lcall_f_f_Int1_done);
  
  /* destruct (Ty CTf_f_Int,
          Dcon Lcall_f_f_Int2) : (lizzieLet67_1Lcall_f_f_Int2,CTf_f_Int) > [(es_37_destruct,Pointer_QTree_Int),
                                                                            (sc_0_12_destruct,Pointer_CTf_f_Int),
                                                                            (q1af0_2_destruct,Pointer_QTree_Int),
                                                                            (t1afa_2_destruct,Pointer_QTree_Int),
                                                                            (t1'aff_2_destruct,Pointer_QTree_Int),
                                                                            (is_zaet_3_destruct,MyDTInt_Bool),
                                                                            (op_addaeu_3_destruct,MyDTInt_Int_Int),
                                                                            (q2af1_2_destruct,Pointer_QTree_Int),
                                                                            (t2afb_2_destruct,Pointer_QTree_Int),
                                                                            (t2'afg_2_destruct,Pointer_QTree_Int)] */
  logic [9:0] lizzieLet67_1Lcall_f_f_Int2_emitted;
  logic [9:0] lizzieLet67_1Lcall_f_f_Int2_done;
  assign es_37_destruct_d = {lizzieLet67_1Lcall_f_f_Int2_d[19:4],
                             (lizzieLet67_1Lcall_f_f_Int2_d[0] && (! lizzieLet67_1Lcall_f_f_Int2_emitted[0]))};
  assign sc_0_12_destruct_d = {lizzieLet67_1Lcall_f_f_Int2_d[35:20],
                               (lizzieLet67_1Lcall_f_f_Int2_d[0] && (! lizzieLet67_1Lcall_f_f_Int2_emitted[1]))};
  assign q1af0_2_destruct_d = {lizzieLet67_1Lcall_f_f_Int2_d[51:36],
                               (lizzieLet67_1Lcall_f_f_Int2_d[0] && (! lizzieLet67_1Lcall_f_f_Int2_emitted[2]))};
  assign t1afa_2_destruct_d = {lizzieLet67_1Lcall_f_f_Int2_d[67:52],
                               (lizzieLet67_1Lcall_f_f_Int2_d[0] && (! lizzieLet67_1Lcall_f_f_Int2_emitted[3]))};
  assign \t1'aff_2_destruct_d  = {lizzieLet67_1Lcall_f_f_Int2_d[83:68],
                                  (lizzieLet67_1Lcall_f_f_Int2_d[0] && (! lizzieLet67_1Lcall_f_f_Int2_emitted[4]))};
  assign is_zaet_3_destruct_d = (lizzieLet67_1Lcall_f_f_Int2_d[0] && (! lizzieLet67_1Lcall_f_f_Int2_emitted[5]));
  assign op_addaeu_3_destruct_d = (lizzieLet67_1Lcall_f_f_Int2_d[0] && (! lizzieLet67_1Lcall_f_f_Int2_emitted[6]));
  assign q2af1_2_destruct_d = {lizzieLet67_1Lcall_f_f_Int2_d[99:84],
                               (lizzieLet67_1Lcall_f_f_Int2_d[0] && (! lizzieLet67_1Lcall_f_f_Int2_emitted[7]))};
  assign t2afb_2_destruct_d = {lizzieLet67_1Lcall_f_f_Int2_d[115:100],
                               (lizzieLet67_1Lcall_f_f_Int2_d[0] && (! lizzieLet67_1Lcall_f_f_Int2_emitted[8]))};
  assign \t2'afg_2_destruct_d  = {lizzieLet67_1Lcall_f_f_Int2_d[131:116],
                                  (lizzieLet67_1Lcall_f_f_Int2_d[0] && (! lizzieLet67_1Lcall_f_f_Int2_emitted[9]))};
  assign lizzieLet67_1Lcall_f_f_Int2_done = (lizzieLet67_1Lcall_f_f_Int2_emitted | ({\t2'afg_2_destruct_d [0],
                                                                                     t2afb_2_destruct_d[0],
                                                                                     q2af1_2_destruct_d[0],
                                                                                     op_addaeu_3_destruct_d[0],
                                                                                     is_zaet_3_destruct_d[0],
                                                                                     \t1'aff_2_destruct_d [0],
                                                                                     t1afa_2_destruct_d[0],
                                                                                     q1af0_2_destruct_d[0],
                                                                                     sc_0_12_destruct_d[0],
                                                                                     es_37_destruct_d[0]} & {\t2'afg_2_destruct_r ,
                                                                                                             t2afb_2_destruct_r,
                                                                                                             q2af1_2_destruct_r,
                                                                                                             op_addaeu_3_destruct_r,
                                                                                                             is_zaet_3_destruct_r,
                                                                                                             \t1'aff_2_destruct_r ,
                                                                                                             t1afa_2_destruct_r,
                                                                                                             q1af0_2_destruct_r,
                                                                                                             sc_0_12_destruct_r,
                                                                                                             es_37_destruct_r}));
  assign lizzieLet67_1Lcall_f_f_Int2_r = (& lizzieLet67_1Lcall_f_f_Int2_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet67_1Lcall_f_f_Int2_emitted <= 10'd0;
    else
      lizzieLet67_1Lcall_f_f_Int2_emitted <= (lizzieLet67_1Lcall_f_f_Int2_r ? 10'd0 :
                                              lizzieLet67_1Lcall_f_f_Int2_done);
  
  /* destruct (Ty CTf_f_Int,
          Dcon Lcall_f_f_Int3) : (lizzieLet67_1Lcall_f_f_Int3,CTf_f_Int) > [(sc_0_11_destruct,Pointer_CTf_f_Int),
                                                                            (q1af0_1_destruct,Pointer_QTree_Int),
                                                                            (t1afa_1_destruct,Pointer_QTree_Int),
                                                                            (t1'aff_1_destruct,Pointer_QTree_Int),
                                                                            (is_zaet_2_destruct,MyDTInt_Bool),
                                                                            (op_addaeu_2_destruct,MyDTInt_Int_Int),
                                                                            (q2af1_1_destruct,Pointer_QTree_Int),
                                                                            (t2afb_1_destruct,Pointer_QTree_Int),
                                                                            (t2'afg_1_destruct,Pointer_QTree_Int),
                                                                            (q3af2_1_destruct,Pointer_QTree_Int),
                                                                            (t3afc_1_destruct,Pointer_QTree_Int),
                                                                            (t3'afh_1_destruct,Pointer_QTree_Int)] */
  logic [11:0] lizzieLet67_1Lcall_f_f_Int3_emitted;
  logic [11:0] lizzieLet67_1Lcall_f_f_Int3_done;
  assign sc_0_11_destruct_d = {lizzieLet67_1Lcall_f_f_Int3_d[19:4],
                               (lizzieLet67_1Lcall_f_f_Int3_d[0] && (! lizzieLet67_1Lcall_f_f_Int3_emitted[0]))};
  assign q1af0_1_destruct_d = {lizzieLet67_1Lcall_f_f_Int3_d[35:20],
                               (lizzieLet67_1Lcall_f_f_Int3_d[0] && (! lizzieLet67_1Lcall_f_f_Int3_emitted[1]))};
  assign t1afa_1_destruct_d = {lizzieLet67_1Lcall_f_f_Int3_d[51:36],
                               (lizzieLet67_1Lcall_f_f_Int3_d[0] && (! lizzieLet67_1Lcall_f_f_Int3_emitted[2]))};
  assign \t1'aff_1_destruct_d  = {lizzieLet67_1Lcall_f_f_Int3_d[67:52],
                                  (lizzieLet67_1Lcall_f_f_Int3_d[0] && (! lizzieLet67_1Lcall_f_f_Int3_emitted[3]))};
  assign is_zaet_2_destruct_d = (lizzieLet67_1Lcall_f_f_Int3_d[0] && (! lizzieLet67_1Lcall_f_f_Int3_emitted[4]));
  assign op_addaeu_2_destruct_d = (lizzieLet67_1Lcall_f_f_Int3_d[0] && (! lizzieLet67_1Lcall_f_f_Int3_emitted[5]));
  assign q2af1_1_destruct_d = {lizzieLet67_1Lcall_f_f_Int3_d[83:68],
                               (lizzieLet67_1Lcall_f_f_Int3_d[0] && (! lizzieLet67_1Lcall_f_f_Int3_emitted[6]))};
  assign t2afb_1_destruct_d = {lizzieLet67_1Lcall_f_f_Int3_d[99:84],
                               (lizzieLet67_1Lcall_f_f_Int3_d[0] && (! lizzieLet67_1Lcall_f_f_Int3_emitted[7]))};
  assign \t2'afg_1_destruct_d  = {lizzieLet67_1Lcall_f_f_Int3_d[115:100],
                                  (lizzieLet67_1Lcall_f_f_Int3_d[0] && (! lizzieLet67_1Lcall_f_f_Int3_emitted[8]))};
  assign q3af2_1_destruct_d = {lizzieLet67_1Lcall_f_f_Int3_d[131:116],
                               (lizzieLet67_1Lcall_f_f_Int3_d[0] && (! lizzieLet67_1Lcall_f_f_Int3_emitted[9]))};
  assign t3afc_1_destruct_d = {lizzieLet67_1Lcall_f_f_Int3_d[147:132],
                               (lizzieLet67_1Lcall_f_f_Int3_d[0] && (! lizzieLet67_1Lcall_f_f_Int3_emitted[10]))};
  assign \t3'afh_1_destruct_d  = {lizzieLet67_1Lcall_f_f_Int3_d[163:148],
                                  (lizzieLet67_1Lcall_f_f_Int3_d[0] && (! lizzieLet67_1Lcall_f_f_Int3_emitted[11]))};
  assign lizzieLet67_1Lcall_f_f_Int3_done = (lizzieLet67_1Lcall_f_f_Int3_emitted | ({\t3'afh_1_destruct_d [0],
                                                                                     t3afc_1_destruct_d[0],
                                                                                     q3af2_1_destruct_d[0],
                                                                                     \t2'afg_1_destruct_d [0],
                                                                                     t2afb_1_destruct_d[0],
                                                                                     q2af1_1_destruct_d[0],
                                                                                     op_addaeu_2_destruct_d[0],
                                                                                     is_zaet_2_destruct_d[0],
                                                                                     \t1'aff_1_destruct_d [0],
                                                                                     t1afa_1_destruct_d[0],
                                                                                     q1af0_1_destruct_d[0],
                                                                                     sc_0_11_destruct_d[0]} & {\t3'afh_1_destruct_r ,
                                                                                                               t3afc_1_destruct_r,
                                                                                                               q3af2_1_destruct_r,
                                                                                                               \t2'afg_1_destruct_r ,
                                                                                                               t2afb_1_destruct_r,
                                                                                                               q2af1_1_destruct_r,
                                                                                                               op_addaeu_2_destruct_r,
                                                                                                               is_zaet_2_destruct_r,
                                                                                                               \t1'aff_1_destruct_r ,
                                                                                                               t1afa_1_destruct_r,
                                                                                                               q1af0_1_destruct_r,
                                                                                                               sc_0_11_destruct_r}));
  assign lizzieLet67_1Lcall_f_f_Int3_r = (& lizzieLet67_1Lcall_f_f_Int3_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet67_1Lcall_f_f_Int3_emitted <= 12'd0;
    else
      lizzieLet67_1Lcall_f_f_Int3_emitted <= (lizzieLet67_1Lcall_f_f_Int3_r ? 12'd0 :
                                              lizzieLet67_1Lcall_f_f_Int3_done);
  
  /* demux (Ty CTf_f_Int,
       Ty CTf_f_Int) : (lizzieLet67_2,CTf_f_Int) (lizzieLet67_1,CTf_f_Int) > [(_53,CTf_f_Int),
                                                                              (lizzieLet67_1Lcall_f_f_Int3,CTf_f_Int),
                                                                              (lizzieLet67_1Lcall_f_f_Int2,CTf_f_Int),
                                                                              (lizzieLet67_1Lcall_f_f_Int1,CTf_f_Int),
                                                                              (lizzieLet67_1Lcall_f_f_Int0,CTf_f_Int)] */
  logic [4:0] lizzieLet67_1_onehotd;
  always_comb
    if ((lizzieLet67_2_d[0] && lizzieLet67_1_d[0]))
      unique case (lizzieLet67_2_d[3:1])
        3'd0: lizzieLet67_1_onehotd = 5'd1;
        3'd1: lizzieLet67_1_onehotd = 5'd2;
        3'd2: lizzieLet67_1_onehotd = 5'd4;
        3'd3: lizzieLet67_1_onehotd = 5'd8;
        3'd4: lizzieLet67_1_onehotd = 5'd16;
        default: lizzieLet67_1_onehotd = 5'd0;
      endcase
    else lizzieLet67_1_onehotd = 5'd0;
  assign _53_d = {lizzieLet67_1_d[163:1], lizzieLet67_1_onehotd[0]};
  assign lizzieLet67_1Lcall_f_f_Int3_d = {lizzieLet67_1_d[163:1],
                                          lizzieLet67_1_onehotd[1]};
  assign lizzieLet67_1Lcall_f_f_Int2_d = {lizzieLet67_1_d[163:1],
                                          lizzieLet67_1_onehotd[2]};
  assign lizzieLet67_1Lcall_f_f_Int1_d = {lizzieLet67_1_d[163:1],
                                          lizzieLet67_1_onehotd[3]};
  assign lizzieLet67_1Lcall_f_f_Int0_d = {lizzieLet67_1_d[163:1],
                                          lizzieLet67_1_onehotd[4]};
  assign lizzieLet67_1_r = (| (lizzieLet67_1_onehotd & {lizzieLet67_1Lcall_f_f_Int0_r,
                                                        lizzieLet67_1Lcall_f_f_Int1_r,
                                                        lizzieLet67_1Lcall_f_f_Int2_r,
                                                        lizzieLet67_1Lcall_f_f_Int3_r,
                                                        _53_r}));
  assign lizzieLet67_2_r = lizzieLet67_1_r;
  
  /* demux (Ty CTf_f_Int,
       Ty Go) : (lizzieLet67_3,CTf_f_Int) (go_15_goMux_data,Go) > [(_52,Go),
                                                                   (lizzieLet67_3Lcall_f_f_Int3,Go),
                                                                   (lizzieLet67_3Lcall_f_f_Int2,Go),
                                                                   (lizzieLet67_3Lcall_f_f_Int1,Go),
                                                                   (lizzieLet67_3Lcall_f_f_Int0,Go)] */
  logic [4:0] go_15_goMux_data_onehotd;
  always_comb
    if ((lizzieLet67_3_d[0] && go_15_goMux_data_d[0]))
      unique case (lizzieLet67_3_d[3:1])
        3'd0: go_15_goMux_data_onehotd = 5'd1;
        3'd1: go_15_goMux_data_onehotd = 5'd2;
        3'd2: go_15_goMux_data_onehotd = 5'd4;
        3'd3: go_15_goMux_data_onehotd = 5'd8;
        3'd4: go_15_goMux_data_onehotd = 5'd16;
        default: go_15_goMux_data_onehotd = 5'd0;
      endcase
    else go_15_goMux_data_onehotd = 5'd0;
  assign _52_d = go_15_goMux_data_onehotd[0];
  assign lizzieLet67_3Lcall_f_f_Int3_d = go_15_goMux_data_onehotd[1];
  assign lizzieLet67_3Lcall_f_f_Int2_d = go_15_goMux_data_onehotd[2];
  assign lizzieLet67_3Lcall_f_f_Int1_d = go_15_goMux_data_onehotd[3];
  assign lizzieLet67_3Lcall_f_f_Int0_d = go_15_goMux_data_onehotd[4];
  assign go_15_goMux_data_r = (| (go_15_goMux_data_onehotd & {lizzieLet67_3Lcall_f_f_Int0_r,
                                                              lizzieLet67_3Lcall_f_f_Int1_r,
                                                              lizzieLet67_3Lcall_f_f_Int2_r,
                                                              lizzieLet67_3Lcall_f_f_Int3_r,
                                                              _52_r}));
  assign lizzieLet67_3_r = go_15_goMux_data_r;
  
  /* buf (Ty Go) : (lizzieLet67_3Lcall_f_f_Int0,Go) > (lizzieLet67_3Lcall_f_f_Int0_1_argbuf,Go) */
  Go_t lizzieLet67_3Lcall_f_f_Int0_bufchan_d;
  logic lizzieLet67_3Lcall_f_f_Int0_bufchan_r;
  assign lizzieLet67_3Lcall_f_f_Int0_r = ((! lizzieLet67_3Lcall_f_f_Int0_bufchan_d[0]) || lizzieLet67_3Lcall_f_f_Int0_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet67_3Lcall_f_f_Int0_bufchan_d <= 1'd0;
    else
      if (lizzieLet67_3Lcall_f_f_Int0_r)
        lizzieLet67_3Lcall_f_f_Int0_bufchan_d <= lizzieLet67_3Lcall_f_f_Int0_d;
  Go_t lizzieLet67_3Lcall_f_f_Int0_bufchan_buf;
  assign lizzieLet67_3Lcall_f_f_Int0_bufchan_r = (! lizzieLet67_3Lcall_f_f_Int0_bufchan_buf[0]);
  assign lizzieLet67_3Lcall_f_f_Int0_1_argbuf_d = (lizzieLet67_3Lcall_f_f_Int0_bufchan_buf[0] ? lizzieLet67_3Lcall_f_f_Int0_bufchan_buf :
                                                   lizzieLet67_3Lcall_f_f_Int0_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet67_3Lcall_f_f_Int0_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet67_3Lcall_f_f_Int0_1_argbuf_r && lizzieLet67_3Lcall_f_f_Int0_bufchan_buf[0]))
        lizzieLet67_3Lcall_f_f_Int0_bufchan_buf <= 1'd0;
      else if (((! lizzieLet67_3Lcall_f_f_Int0_1_argbuf_r) && (! lizzieLet67_3Lcall_f_f_Int0_bufchan_buf[0])))
        lizzieLet67_3Lcall_f_f_Int0_bufchan_buf <= lizzieLet67_3Lcall_f_f_Int0_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet67_3Lcall_f_f_Int1,Go) > (lizzieLet67_3Lcall_f_f_Int1_1_argbuf,Go) */
  Go_t lizzieLet67_3Lcall_f_f_Int1_bufchan_d;
  logic lizzieLet67_3Lcall_f_f_Int1_bufchan_r;
  assign lizzieLet67_3Lcall_f_f_Int1_r = ((! lizzieLet67_3Lcall_f_f_Int1_bufchan_d[0]) || lizzieLet67_3Lcall_f_f_Int1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet67_3Lcall_f_f_Int1_bufchan_d <= 1'd0;
    else
      if (lizzieLet67_3Lcall_f_f_Int1_r)
        lizzieLet67_3Lcall_f_f_Int1_bufchan_d <= lizzieLet67_3Lcall_f_f_Int1_d;
  Go_t lizzieLet67_3Lcall_f_f_Int1_bufchan_buf;
  assign lizzieLet67_3Lcall_f_f_Int1_bufchan_r = (! lizzieLet67_3Lcall_f_f_Int1_bufchan_buf[0]);
  assign lizzieLet67_3Lcall_f_f_Int1_1_argbuf_d = (lizzieLet67_3Lcall_f_f_Int1_bufchan_buf[0] ? lizzieLet67_3Lcall_f_f_Int1_bufchan_buf :
                                                   lizzieLet67_3Lcall_f_f_Int1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet67_3Lcall_f_f_Int1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet67_3Lcall_f_f_Int1_1_argbuf_r && lizzieLet67_3Lcall_f_f_Int1_bufchan_buf[0]))
        lizzieLet67_3Lcall_f_f_Int1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet67_3Lcall_f_f_Int1_1_argbuf_r) && (! lizzieLet67_3Lcall_f_f_Int1_bufchan_buf[0])))
        lizzieLet67_3Lcall_f_f_Int1_bufchan_buf <= lizzieLet67_3Lcall_f_f_Int1_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet67_3Lcall_f_f_Int2,Go) > (lizzieLet67_3Lcall_f_f_Int2_1_argbuf,Go) */
  Go_t lizzieLet67_3Lcall_f_f_Int2_bufchan_d;
  logic lizzieLet67_3Lcall_f_f_Int2_bufchan_r;
  assign lizzieLet67_3Lcall_f_f_Int2_r = ((! lizzieLet67_3Lcall_f_f_Int2_bufchan_d[0]) || lizzieLet67_3Lcall_f_f_Int2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet67_3Lcall_f_f_Int2_bufchan_d <= 1'd0;
    else
      if (lizzieLet67_3Lcall_f_f_Int2_r)
        lizzieLet67_3Lcall_f_f_Int2_bufchan_d <= lizzieLet67_3Lcall_f_f_Int2_d;
  Go_t lizzieLet67_3Lcall_f_f_Int2_bufchan_buf;
  assign lizzieLet67_3Lcall_f_f_Int2_bufchan_r = (! lizzieLet67_3Lcall_f_f_Int2_bufchan_buf[0]);
  assign lizzieLet67_3Lcall_f_f_Int2_1_argbuf_d = (lizzieLet67_3Lcall_f_f_Int2_bufchan_buf[0] ? lizzieLet67_3Lcall_f_f_Int2_bufchan_buf :
                                                   lizzieLet67_3Lcall_f_f_Int2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet67_3Lcall_f_f_Int2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet67_3Lcall_f_f_Int2_1_argbuf_r && lizzieLet67_3Lcall_f_f_Int2_bufchan_buf[0]))
        lizzieLet67_3Lcall_f_f_Int2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet67_3Lcall_f_f_Int2_1_argbuf_r) && (! lizzieLet67_3Lcall_f_f_Int2_bufchan_buf[0])))
        lizzieLet67_3Lcall_f_f_Int2_bufchan_buf <= lizzieLet67_3Lcall_f_f_Int2_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet67_3Lcall_f_f_Int3,Go) > (lizzieLet67_3Lcall_f_f_Int3_1_argbuf,Go) */
  Go_t lizzieLet67_3Lcall_f_f_Int3_bufchan_d;
  logic lizzieLet67_3Lcall_f_f_Int3_bufchan_r;
  assign lizzieLet67_3Lcall_f_f_Int3_r = ((! lizzieLet67_3Lcall_f_f_Int3_bufchan_d[0]) || lizzieLet67_3Lcall_f_f_Int3_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet67_3Lcall_f_f_Int3_bufchan_d <= 1'd0;
    else
      if (lizzieLet67_3Lcall_f_f_Int3_r)
        lizzieLet67_3Lcall_f_f_Int3_bufchan_d <= lizzieLet67_3Lcall_f_f_Int3_d;
  Go_t lizzieLet67_3Lcall_f_f_Int3_bufchan_buf;
  assign lizzieLet67_3Lcall_f_f_Int3_bufchan_r = (! lizzieLet67_3Lcall_f_f_Int3_bufchan_buf[0]);
  assign lizzieLet67_3Lcall_f_f_Int3_1_argbuf_d = (lizzieLet67_3Lcall_f_f_Int3_bufchan_buf[0] ? lizzieLet67_3Lcall_f_f_Int3_bufchan_buf :
                                                   lizzieLet67_3Lcall_f_f_Int3_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet67_3Lcall_f_f_Int3_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet67_3Lcall_f_f_Int3_1_argbuf_r && lizzieLet67_3Lcall_f_f_Int3_bufchan_buf[0]))
        lizzieLet67_3Lcall_f_f_Int3_bufchan_buf <= 1'd0;
      else if (((! lizzieLet67_3Lcall_f_f_Int3_1_argbuf_r) && (! lizzieLet67_3Lcall_f_f_Int3_bufchan_buf[0])))
        lizzieLet67_3Lcall_f_f_Int3_bufchan_buf <= lizzieLet67_3Lcall_f_f_Int3_bufchan_d;
  
  /* demux (Ty CTf_f_Int,
       Ty Pointer_QTree_Int) : (lizzieLet67_4,CTf_f_Int) (srtarg_0_2_goMux_mux,Pointer_QTree_Int) > [(lizzieLet67_4Lf_f_Intsbos,Pointer_QTree_Int),
                                                                                                     (lizzieLet67_4Lcall_f_f_Int3,Pointer_QTree_Int),
                                                                                                     (lizzieLet67_4Lcall_f_f_Int2,Pointer_QTree_Int),
                                                                                                     (lizzieLet67_4Lcall_f_f_Int1,Pointer_QTree_Int),
                                                                                                     (lizzieLet67_4Lcall_f_f_Int0,Pointer_QTree_Int)] */
  logic [4:0] srtarg_0_2_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet67_4_d[0] && srtarg_0_2_goMux_mux_d[0]))
      unique case (lizzieLet67_4_d[3:1])
        3'd0: srtarg_0_2_goMux_mux_onehotd = 5'd1;
        3'd1: srtarg_0_2_goMux_mux_onehotd = 5'd2;
        3'd2: srtarg_0_2_goMux_mux_onehotd = 5'd4;
        3'd3: srtarg_0_2_goMux_mux_onehotd = 5'd8;
        3'd4: srtarg_0_2_goMux_mux_onehotd = 5'd16;
        default: srtarg_0_2_goMux_mux_onehotd = 5'd0;
      endcase
    else srtarg_0_2_goMux_mux_onehotd = 5'd0;
  assign lizzieLet67_4Lf_f_Intsbos_d = {srtarg_0_2_goMux_mux_d[16:1],
                                        srtarg_0_2_goMux_mux_onehotd[0]};
  assign lizzieLet67_4Lcall_f_f_Int3_d = {srtarg_0_2_goMux_mux_d[16:1],
                                          srtarg_0_2_goMux_mux_onehotd[1]};
  assign lizzieLet67_4Lcall_f_f_Int2_d = {srtarg_0_2_goMux_mux_d[16:1],
                                          srtarg_0_2_goMux_mux_onehotd[2]};
  assign lizzieLet67_4Lcall_f_f_Int1_d = {srtarg_0_2_goMux_mux_d[16:1],
                                          srtarg_0_2_goMux_mux_onehotd[3]};
  assign lizzieLet67_4Lcall_f_f_Int0_d = {srtarg_0_2_goMux_mux_d[16:1],
                                          srtarg_0_2_goMux_mux_onehotd[4]};
  assign srtarg_0_2_goMux_mux_r = (| (srtarg_0_2_goMux_mux_onehotd & {lizzieLet67_4Lcall_f_f_Int0_r,
                                                                      lizzieLet67_4Lcall_f_f_Int1_r,
                                                                      lizzieLet67_4Lcall_f_f_Int2_r,
                                                                      lizzieLet67_4Lcall_f_f_Int3_r,
                                                                      lizzieLet67_4Lf_f_Intsbos_r}));
  assign lizzieLet67_4_r = srtarg_0_2_goMux_mux_r;
  
  /* dcon (Ty QTree_Int,
      Dcon QNode_Int) : [(lizzieLet67_4Lcall_f_f_Int0,Pointer_QTree_Int),
                         (es_35_destruct,Pointer_QTree_Int),
                         (es_36_1_destruct,Pointer_QTree_Int),
                         (es_37_2_destruct,Pointer_QTree_Int)] > (lizzieLet67_4Lcall_f_f_Int0_1es_35_1es_36_1_1es_37_2_1QNode_Int,QTree_Int) */
  assign lizzieLet67_4Lcall_f_f_Int0_1es_35_1es_36_1_1es_37_2_1QNode_Int_d = QNode_Int_dc((& {lizzieLet67_4Lcall_f_f_Int0_d[0],
                                                                                              es_35_destruct_d[0],
                                                                                              es_36_1_destruct_d[0],
                                                                                              es_37_2_destruct_d[0]}), lizzieLet67_4Lcall_f_f_Int0_d, es_35_destruct_d, es_36_1_destruct_d, es_37_2_destruct_d);
  assign {lizzieLet67_4Lcall_f_f_Int0_r,
          es_35_destruct_r,
          es_36_1_destruct_r,
          es_37_2_destruct_r} = {4 {(lizzieLet67_4Lcall_f_f_Int0_1es_35_1es_36_1_1es_37_2_1QNode_Int_r && lizzieLet67_4Lcall_f_f_Int0_1es_35_1es_36_1_1es_37_2_1QNode_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (lizzieLet67_4Lcall_f_f_Int0_1es_35_1es_36_1_1es_37_2_1QNode_Int,QTree_Int) > (lizzieLet71_1_argbuf,QTree_Int) */
  QTree_Int_t lizzieLet67_4Lcall_f_f_Int0_1es_35_1es_36_1_1es_37_2_1QNode_Int_bufchan_d;
  logic lizzieLet67_4Lcall_f_f_Int0_1es_35_1es_36_1_1es_37_2_1QNode_Int_bufchan_r;
  assign lizzieLet67_4Lcall_f_f_Int0_1es_35_1es_36_1_1es_37_2_1QNode_Int_r = ((! lizzieLet67_4Lcall_f_f_Int0_1es_35_1es_36_1_1es_37_2_1QNode_Int_bufchan_d[0]) || lizzieLet67_4Lcall_f_f_Int0_1es_35_1es_36_1_1es_37_2_1QNode_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet67_4Lcall_f_f_Int0_1es_35_1es_36_1_1es_37_2_1QNode_Int_bufchan_d <= {66'd0,
                                                                                    1'd0};
    else
      if (lizzieLet67_4Lcall_f_f_Int0_1es_35_1es_36_1_1es_37_2_1QNode_Int_r)
        lizzieLet67_4Lcall_f_f_Int0_1es_35_1es_36_1_1es_37_2_1QNode_Int_bufchan_d <= lizzieLet67_4Lcall_f_f_Int0_1es_35_1es_36_1_1es_37_2_1QNode_Int_d;
  QTree_Int_t lizzieLet67_4Lcall_f_f_Int0_1es_35_1es_36_1_1es_37_2_1QNode_Int_bufchan_buf;
  assign lizzieLet67_4Lcall_f_f_Int0_1es_35_1es_36_1_1es_37_2_1QNode_Int_bufchan_r = (! lizzieLet67_4Lcall_f_f_Int0_1es_35_1es_36_1_1es_37_2_1QNode_Int_bufchan_buf[0]);
  assign lizzieLet71_1_argbuf_d = (lizzieLet67_4Lcall_f_f_Int0_1es_35_1es_36_1_1es_37_2_1QNode_Int_bufchan_buf[0] ? lizzieLet67_4Lcall_f_f_Int0_1es_35_1es_36_1_1es_37_2_1QNode_Int_bufchan_buf :
                                   lizzieLet67_4Lcall_f_f_Int0_1es_35_1es_36_1_1es_37_2_1QNode_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet67_4Lcall_f_f_Int0_1es_35_1es_36_1_1es_37_2_1QNode_Int_bufchan_buf <= {66'd0,
                                                                                      1'd0};
    else
      if ((lizzieLet71_1_argbuf_r && lizzieLet67_4Lcall_f_f_Int0_1es_35_1es_36_1_1es_37_2_1QNode_Int_bufchan_buf[0]))
        lizzieLet67_4Lcall_f_f_Int0_1es_35_1es_36_1_1es_37_2_1QNode_Int_bufchan_buf <= {66'd0,
                                                                                        1'd0};
      else if (((! lizzieLet71_1_argbuf_r) && (! lizzieLet67_4Lcall_f_f_Int0_1es_35_1es_36_1_1es_37_2_1QNode_Int_bufchan_buf[0])))
        lizzieLet67_4Lcall_f_f_Int0_1es_35_1es_36_1_1es_37_2_1QNode_Int_bufchan_buf <= lizzieLet67_4Lcall_f_f_Int0_1es_35_1es_36_1_1es_37_2_1QNode_Int_bufchan_d;
  
  /* dcon (Ty CTf_f_Int,
      Dcon Lcall_f_f_Int0) : [(lizzieLet67_4Lcall_f_f_Int1,Pointer_QTree_Int),
                              (es_36_destruct,Pointer_QTree_Int),
                              (es_37_1_destruct,Pointer_QTree_Int),
                              (sc_0_13_destruct,Pointer_CTf_f_Int)] > (lizzieLet67_4Lcall_f_f_Int1_1es_36_1es_37_1_1sc_0_13_1Lcall_f_f_Int0,CTf_f_Int) */
  assign lizzieLet67_4Lcall_f_f_Int1_1es_36_1es_37_1_1sc_0_13_1Lcall_f_f_Int0_d = Lcall_f_f_Int0_dc((& {lizzieLet67_4Lcall_f_f_Int1_d[0],
                                                                                                        es_36_destruct_d[0],
                                                                                                        es_37_1_destruct_d[0],
                                                                                                        sc_0_13_destruct_d[0]}), lizzieLet67_4Lcall_f_f_Int1_d, es_36_destruct_d, es_37_1_destruct_d, sc_0_13_destruct_d);
  assign {lizzieLet67_4Lcall_f_f_Int1_r,
          es_36_destruct_r,
          es_37_1_destruct_r,
          sc_0_13_destruct_r} = {4 {(lizzieLet67_4Lcall_f_f_Int1_1es_36_1es_37_1_1sc_0_13_1Lcall_f_f_Int0_r && lizzieLet67_4Lcall_f_f_Int1_1es_36_1es_37_1_1sc_0_13_1Lcall_f_f_Int0_d[0])}};
  
  /* buf (Ty CTf_f_Int) : (lizzieLet67_4Lcall_f_f_Int1_1es_36_1es_37_1_1sc_0_13_1Lcall_f_f_Int0,CTf_f_Int) > (lizzieLet70_1_argbuf,CTf_f_Int) */
  CTf_f_Int_t lizzieLet67_4Lcall_f_f_Int1_1es_36_1es_37_1_1sc_0_13_1Lcall_f_f_Int0_bufchan_d;
  logic lizzieLet67_4Lcall_f_f_Int1_1es_36_1es_37_1_1sc_0_13_1Lcall_f_f_Int0_bufchan_r;
  assign lizzieLet67_4Lcall_f_f_Int1_1es_36_1es_37_1_1sc_0_13_1Lcall_f_f_Int0_r = ((! lizzieLet67_4Lcall_f_f_Int1_1es_36_1es_37_1_1sc_0_13_1Lcall_f_f_Int0_bufchan_d[0]) || lizzieLet67_4Lcall_f_f_Int1_1es_36_1es_37_1_1sc_0_13_1Lcall_f_f_Int0_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet67_4Lcall_f_f_Int1_1es_36_1es_37_1_1sc_0_13_1Lcall_f_f_Int0_bufchan_d <= {163'd0,
                                                                                         1'd0};
    else
      if (lizzieLet67_4Lcall_f_f_Int1_1es_36_1es_37_1_1sc_0_13_1Lcall_f_f_Int0_r)
        lizzieLet67_4Lcall_f_f_Int1_1es_36_1es_37_1_1sc_0_13_1Lcall_f_f_Int0_bufchan_d <= lizzieLet67_4Lcall_f_f_Int1_1es_36_1es_37_1_1sc_0_13_1Lcall_f_f_Int0_d;
  CTf_f_Int_t lizzieLet67_4Lcall_f_f_Int1_1es_36_1es_37_1_1sc_0_13_1Lcall_f_f_Int0_bufchan_buf;
  assign lizzieLet67_4Lcall_f_f_Int1_1es_36_1es_37_1_1sc_0_13_1Lcall_f_f_Int0_bufchan_r = (! lizzieLet67_4Lcall_f_f_Int1_1es_36_1es_37_1_1sc_0_13_1Lcall_f_f_Int0_bufchan_buf[0]);
  assign lizzieLet70_1_argbuf_d = (lizzieLet67_4Lcall_f_f_Int1_1es_36_1es_37_1_1sc_0_13_1Lcall_f_f_Int0_bufchan_buf[0] ? lizzieLet67_4Lcall_f_f_Int1_1es_36_1es_37_1_1sc_0_13_1Lcall_f_f_Int0_bufchan_buf :
                                   lizzieLet67_4Lcall_f_f_Int1_1es_36_1es_37_1_1sc_0_13_1Lcall_f_f_Int0_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet67_4Lcall_f_f_Int1_1es_36_1es_37_1_1sc_0_13_1Lcall_f_f_Int0_bufchan_buf <= {163'd0,
                                                                                           1'd0};
    else
      if ((lizzieLet70_1_argbuf_r && lizzieLet67_4Lcall_f_f_Int1_1es_36_1es_37_1_1sc_0_13_1Lcall_f_f_Int0_bufchan_buf[0]))
        lizzieLet67_4Lcall_f_f_Int1_1es_36_1es_37_1_1sc_0_13_1Lcall_f_f_Int0_bufchan_buf <= {163'd0,
                                                                                             1'd0};
      else if (((! lizzieLet70_1_argbuf_r) && (! lizzieLet67_4Lcall_f_f_Int1_1es_36_1es_37_1_1sc_0_13_1Lcall_f_f_Int0_bufchan_buf[0])))
        lizzieLet67_4Lcall_f_f_Int1_1es_36_1es_37_1_1sc_0_13_1Lcall_f_f_Int0_bufchan_buf <= lizzieLet67_4Lcall_f_f_Int1_1es_36_1es_37_1_1sc_0_13_1Lcall_f_f_Int0_bufchan_d;
  
  /* dcon (Ty CTf_f_Int,
      Dcon Lcall_f_f_Int1) : [(lizzieLet67_4Lcall_f_f_Int2,Pointer_QTree_Int),
                              (es_37_destruct,Pointer_QTree_Int),
                              (sc_0_12_destruct,Pointer_CTf_f_Int),
                              (q1af0_2_destruct,Pointer_QTree_Int),
                              (t1afa_2_destruct,Pointer_QTree_Int),
                              (t1'aff_2_destruct,Pointer_QTree_Int),
                              (is_zaet_3_1,MyDTInt_Bool),
                              (op_addaeu_3_1,MyDTInt_Int_Int)] > (lizzieLet67_4Lcall_f_f_Int2_1es_37_1sc_0_12_1q1af0_2_1t1afa_2_1t1'aff_2_1is_zaet_3_1op_addaeu_3_1Lcall_f_f_Int1,CTf_f_Int) */
  assign \lizzieLet67_4Lcall_f_f_Int2_1es_37_1sc_0_12_1q1af0_2_1t1afa_2_1t1'aff_2_1is_zaet_3_1op_addaeu_3_1Lcall_f_f_Int1_d  = Lcall_f_f_Int1_dc((& {lizzieLet67_4Lcall_f_f_Int2_d[0],
                                                                                                                                                     es_37_destruct_d[0],
                                                                                                                                                     sc_0_12_destruct_d[0],
                                                                                                                                                     q1af0_2_destruct_d[0],
                                                                                                                                                     t1afa_2_destruct_d[0],
                                                                                                                                                     \t1'aff_2_destruct_d [0],
                                                                                                                                                     is_zaet_3_1_d[0],
                                                                                                                                                     op_addaeu_3_1_d[0]}), lizzieLet67_4Lcall_f_f_Int2_d, es_37_destruct_d, sc_0_12_destruct_d, q1af0_2_destruct_d, t1afa_2_destruct_d, \t1'aff_2_destruct_d , is_zaet_3_1_d, op_addaeu_3_1_d);
  assign {lizzieLet67_4Lcall_f_f_Int2_r,
          es_37_destruct_r,
          sc_0_12_destruct_r,
          q1af0_2_destruct_r,
          t1afa_2_destruct_r,
          \t1'aff_2_destruct_r ,
          is_zaet_3_1_r,
          op_addaeu_3_1_r} = {8 {(\lizzieLet67_4Lcall_f_f_Int2_1es_37_1sc_0_12_1q1af0_2_1t1afa_2_1t1'aff_2_1is_zaet_3_1op_addaeu_3_1Lcall_f_f_Int1_r  && \lizzieLet67_4Lcall_f_f_Int2_1es_37_1sc_0_12_1q1af0_2_1t1afa_2_1t1'aff_2_1is_zaet_3_1op_addaeu_3_1Lcall_f_f_Int1_d [0])}};
  
  /* buf (Ty CTf_f_Int) : (lizzieLet67_4Lcall_f_f_Int2_1es_37_1sc_0_12_1q1af0_2_1t1afa_2_1t1'aff_2_1is_zaet_3_1op_addaeu_3_1Lcall_f_f_Int1,CTf_f_Int) > (lizzieLet69_1_argbuf,CTf_f_Int) */
  CTf_f_Int_t \lizzieLet67_4Lcall_f_f_Int2_1es_37_1sc_0_12_1q1af0_2_1t1afa_2_1t1'aff_2_1is_zaet_3_1op_addaeu_3_1Lcall_f_f_Int1_bufchan_d ;
  logic \lizzieLet67_4Lcall_f_f_Int2_1es_37_1sc_0_12_1q1af0_2_1t1afa_2_1t1'aff_2_1is_zaet_3_1op_addaeu_3_1Lcall_f_f_Int1_bufchan_r ;
  assign \lizzieLet67_4Lcall_f_f_Int2_1es_37_1sc_0_12_1q1af0_2_1t1afa_2_1t1'aff_2_1is_zaet_3_1op_addaeu_3_1Lcall_f_f_Int1_r  = ((! \lizzieLet67_4Lcall_f_f_Int2_1es_37_1sc_0_12_1q1af0_2_1t1afa_2_1t1'aff_2_1is_zaet_3_1op_addaeu_3_1Lcall_f_f_Int1_bufchan_d [0]) || \lizzieLet67_4Lcall_f_f_Int2_1es_37_1sc_0_12_1q1af0_2_1t1afa_2_1t1'aff_2_1is_zaet_3_1op_addaeu_3_1Lcall_f_f_Int1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet67_4Lcall_f_f_Int2_1es_37_1sc_0_12_1q1af0_2_1t1afa_2_1t1'aff_2_1is_zaet_3_1op_addaeu_3_1Lcall_f_f_Int1_bufchan_d  <= {163'd0,
                                                                                                                                      1'd0};
    else
      if (\lizzieLet67_4Lcall_f_f_Int2_1es_37_1sc_0_12_1q1af0_2_1t1afa_2_1t1'aff_2_1is_zaet_3_1op_addaeu_3_1Lcall_f_f_Int1_r )
        \lizzieLet67_4Lcall_f_f_Int2_1es_37_1sc_0_12_1q1af0_2_1t1afa_2_1t1'aff_2_1is_zaet_3_1op_addaeu_3_1Lcall_f_f_Int1_bufchan_d  <= \lizzieLet67_4Lcall_f_f_Int2_1es_37_1sc_0_12_1q1af0_2_1t1afa_2_1t1'aff_2_1is_zaet_3_1op_addaeu_3_1Lcall_f_f_Int1_d ;
  CTf_f_Int_t \lizzieLet67_4Lcall_f_f_Int2_1es_37_1sc_0_12_1q1af0_2_1t1afa_2_1t1'aff_2_1is_zaet_3_1op_addaeu_3_1Lcall_f_f_Int1_bufchan_buf ;
  assign \lizzieLet67_4Lcall_f_f_Int2_1es_37_1sc_0_12_1q1af0_2_1t1afa_2_1t1'aff_2_1is_zaet_3_1op_addaeu_3_1Lcall_f_f_Int1_bufchan_r  = (! \lizzieLet67_4Lcall_f_f_Int2_1es_37_1sc_0_12_1q1af0_2_1t1afa_2_1t1'aff_2_1is_zaet_3_1op_addaeu_3_1Lcall_f_f_Int1_bufchan_buf [0]);
  assign lizzieLet69_1_argbuf_d = (\lizzieLet67_4Lcall_f_f_Int2_1es_37_1sc_0_12_1q1af0_2_1t1afa_2_1t1'aff_2_1is_zaet_3_1op_addaeu_3_1Lcall_f_f_Int1_bufchan_buf [0] ? \lizzieLet67_4Lcall_f_f_Int2_1es_37_1sc_0_12_1q1af0_2_1t1afa_2_1t1'aff_2_1is_zaet_3_1op_addaeu_3_1Lcall_f_f_Int1_bufchan_buf  :
                                   \lizzieLet67_4Lcall_f_f_Int2_1es_37_1sc_0_12_1q1af0_2_1t1afa_2_1t1'aff_2_1is_zaet_3_1op_addaeu_3_1Lcall_f_f_Int1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet67_4Lcall_f_f_Int2_1es_37_1sc_0_12_1q1af0_2_1t1afa_2_1t1'aff_2_1is_zaet_3_1op_addaeu_3_1Lcall_f_f_Int1_bufchan_buf  <= {163'd0,
                                                                                                                                        1'd0};
    else
      if ((lizzieLet69_1_argbuf_r && \lizzieLet67_4Lcall_f_f_Int2_1es_37_1sc_0_12_1q1af0_2_1t1afa_2_1t1'aff_2_1is_zaet_3_1op_addaeu_3_1Lcall_f_f_Int1_bufchan_buf [0]))
        \lizzieLet67_4Lcall_f_f_Int2_1es_37_1sc_0_12_1q1af0_2_1t1afa_2_1t1'aff_2_1is_zaet_3_1op_addaeu_3_1Lcall_f_f_Int1_bufchan_buf  <= {163'd0,
                                                                                                                                          1'd0};
      else if (((! lizzieLet69_1_argbuf_r) && (! \lizzieLet67_4Lcall_f_f_Int2_1es_37_1sc_0_12_1q1af0_2_1t1afa_2_1t1'aff_2_1is_zaet_3_1op_addaeu_3_1Lcall_f_f_Int1_bufchan_buf [0])))
        \lizzieLet67_4Lcall_f_f_Int2_1es_37_1sc_0_12_1q1af0_2_1t1afa_2_1t1'aff_2_1is_zaet_3_1op_addaeu_3_1Lcall_f_f_Int1_bufchan_buf  <= \lizzieLet67_4Lcall_f_f_Int2_1es_37_1sc_0_12_1q1af0_2_1t1afa_2_1t1'aff_2_1is_zaet_3_1op_addaeu_3_1Lcall_f_f_Int1_bufchan_d ;
  
  /* dcon (Ty CTf_f_Int,
      Dcon Lcall_f_f_Int2) : [(lizzieLet67_4Lcall_f_f_Int3,Pointer_QTree_Int),
                              (sc_0_11_destruct,Pointer_CTf_f_Int),
                              (q1af0_1_destruct,Pointer_QTree_Int),
                              (t1afa_1_destruct,Pointer_QTree_Int),
                              (t1'aff_1_destruct,Pointer_QTree_Int),
                              (is_zaet_2_1,MyDTInt_Bool),
                              (op_addaeu_2_1,MyDTInt_Int_Int),
                              (q2af1_1_destruct,Pointer_QTree_Int),
                              (t2afb_1_destruct,Pointer_QTree_Int),
                              (t2'afg_1_destruct,Pointer_QTree_Int)] > (lizzieLet67_4Lcall_f_f_Int3_1sc_0_11_1q1af0_1_1t1afa_1_1t1'aff_1_1is_zaet_2_1op_addaeu_2_1q2af1_1_1t2afb_1_1t2'afg_1_1Lcall_f_f_Int2,CTf_f_Int) */
  assign \lizzieLet67_4Lcall_f_f_Int3_1sc_0_11_1q1af0_1_1t1afa_1_1t1'aff_1_1is_zaet_2_1op_addaeu_2_1q2af1_1_1t2afb_1_1t2'afg_1_1Lcall_f_f_Int2_d  = Lcall_f_f_Int2_dc((& {lizzieLet67_4Lcall_f_f_Int3_d[0],
                                                                                                                                                                          sc_0_11_destruct_d[0],
                                                                                                                                                                          q1af0_1_destruct_d[0],
                                                                                                                                                                          t1afa_1_destruct_d[0],
                                                                                                                                                                          \t1'aff_1_destruct_d [0],
                                                                                                                                                                          is_zaet_2_1_d[0],
                                                                                                                                                                          op_addaeu_2_1_d[0],
                                                                                                                                                                          q2af1_1_destruct_d[0],
                                                                                                                                                                          t2afb_1_destruct_d[0],
                                                                                                                                                                          \t2'afg_1_destruct_d [0]}), lizzieLet67_4Lcall_f_f_Int3_d, sc_0_11_destruct_d, q1af0_1_destruct_d, t1afa_1_destruct_d, \t1'aff_1_destruct_d , is_zaet_2_1_d, op_addaeu_2_1_d, q2af1_1_destruct_d, t2afb_1_destruct_d, \t2'afg_1_destruct_d );
  assign {lizzieLet67_4Lcall_f_f_Int3_r,
          sc_0_11_destruct_r,
          q1af0_1_destruct_r,
          t1afa_1_destruct_r,
          \t1'aff_1_destruct_r ,
          is_zaet_2_1_r,
          op_addaeu_2_1_r,
          q2af1_1_destruct_r,
          t2afb_1_destruct_r,
          \t2'afg_1_destruct_r } = {10 {(\lizzieLet67_4Lcall_f_f_Int3_1sc_0_11_1q1af0_1_1t1afa_1_1t1'aff_1_1is_zaet_2_1op_addaeu_2_1q2af1_1_1t2afb_1_1t2'afg_1_1Lcall_f_f_Int2_r  && \lizzieLet67_4Lcall_f_f_Int3_1sc_0_11_1q1af0_1_1t1afa_1_1t1'aff_1_1is_zaet_2_1op_addaeu_2_1q2af1_1_1t2afb_1_1t2'afg_1_1Lcall_f_f_Int2_d [0])}};
  
  /* buf (Ty CTf_f_Int) : (lizzieLet67_4Lcall_f_f_Int3_1sc_0_11_1q1af0_1_1t1afa_1_1t1'aff_1_1is_zaet_2_1op_addaeu_2_1q2af1_1_1t2afb_1_1t2'afg_1_1Lcall_f_f_Int2,CTf_f_Int) > (lizzieLet68_1_argbuf,CTf_f_Int) */
  CTf_f_Int_t \lizzieLet67_4Lcall_f_f_Int3_1sc_0_11_1q1af0_1_1t1afa_1_1t1'aff_1_1is_zaet_2_1op_addaeu_2_1q2af1_1_1t2afb_1_1t2'afg_1_1Lcall_f_f_Int2_bufchan_d ;
  logic \lizzieLet67_4Lcall_f_f_Int3_1sc_0_11_1q1af0_1_1t1afa_1_1t1'aff_1_1is_zaet_2_1op_addaeu_2_1q2af1_1_1t2afb_1_1t2'afg_1_1Lcall_f_f_Int2_bufchan_r ;
  assign \lizzieLet67_4Lcall_f_f_Int3_1sc_0_11_1q1af0_1_1t1afa_1_1t1'aff_1_1is_zaet_2_1op_addaeu_2_1q2af1_1_1t2afb_1_1t2'afg_1_1Lcall_f_f_Int2_r  = ((! \lizzieLet67_4Lcall_f_f_Int3_1sc_0_11_1q1af0_1_1t1afa_1_1t1'aff_1_1is_zaet_2_1op_addaeu_2_1q2af1_1_1t2afb_1_1t2'afg_1_1Lcall_f_f_Int2_bufchan_d [0]) || \lizzieLet67_4Lcall_f_f_Int3_1sc_0_11_1q1af0_1_1t1afa_1_1t1'aff_1_1is_zaet_2_1op_addaeu_2_1q2af1_1_1t2afb_1_1t2'afg_1_1Lcall_f_f_Int2_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet67_4Lcall_f_f_Int3_1sc_0_11_1q1af0_1_1t1afa_1_1t1'aff_1_1is_zaet_2_1op_addaeu_2_1q2af1_1_1t2afb_1_1t2'afg_1_1Lcall_f_f_Int2_bufchan_d  <= {163'd0,
                                                                                                                                                           1'd0};
    else
      if (\lizzieLet67_4Lcall_f_f_Int3_1sc_0_11_1q1af0_1_1t1afa_1_1t1'aff_1_1is_zaet_2_1op_addaeu_2_1q2af1_1_1t2afb_1_1t2'afg_1_1Lcall_f_f_Int2_r )
        \lizzieLet67_4Lcall_f_f_Int3_1sc_0_11_1q1af0_1_1t1afa_1_1t1'aff_1_1is_zaet_2_1op_addaeu_2_1q2af1_1_1t2afb_1_1t2'afg_1_1Lcall_f_f_Int2_bufchan_d  <= \lizzieLet67_4Lcall_f_f_Int3_1sc_0_11_1q1af0_1_1t1afa_1_1t1'aff_1_1is_zaet_2_1op_addaeu_2_1q2af1_1_1t2afb_1_1t2'afg_1_1Lcall_f_f_Int2_d ;
  CTf_f_Int_t \lizzieLet67_4Lcall_f_f_Int3_1sc_0_11_1q1af0_1_1t1afa_1_1t1'aff_1_1is_zaet_2_1op_addaeu_2_1q2af1_1_1t2afb_1_1t2'afg_1_1Lcall_f_f_Int2_bufchan_buf ;
  assign \lizzieLet67_4Lcall_f_f_Int3_1sc_0_11_1q1af0_1_1t1afa_1_1t1'aff_1_1is_zaet_2_1op_addaeu_2_1q2af1_1_1t2afb_1_1t2'afg_1_1Lcall_f_f_Int2_bufchan_r  = (! \lizzieLet67_4Lcall_f_f_Int3_1sc_0_11_1q1af0_1_1t1afa_1_1t1'aff_1_1is_zaet_2_1op_addaeu_2_1q2af1_1_1t2afb_1_1t2'afg_1_1Lcall_f_f_Int2_bufchan_buf [0]);
  assign lizzieLet68_1_argbuf_d = (\lizzieLet67_4Lcall_f_f_Int3_1sc_0_11_1q1af0_1_1t1afa_1_1t1'aff_1_1is_zaet_2_1op_addaeu_2_1q2af1_1_1t2afb_1_1t2'afg_1_1Lcall_f_f_Int2_bufchan_buf [0] ? \lizzieLet67_4Lcall_f_f_Int3_1sc_0_11_1q1af0_1_1t1afa_1_1t1'aff_1_1is_zaet_2_1op_addaeu_2_1q2af1_1_1t2afb_1_1t2'afg_1_1Lcall_f_f_Int2_bufchan_buf  :
                                   \lizzieLet67_4Lcall_f_f_Int3_1sc_0_11_1q1af0_1_1t1afa_1_1t1'aff_1_1is_zaet_2_1op_addaeu_2_1q2af1_1_1t2afb_1_1t2'afg_1_1Lcall_f_f_Int2_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet67_4Lcall_f_f_Int3_1sc_0_11_1q1af0_1_1t1afa_1_1t1'aff_1_1is_zaet_2_1op_addaeu_2_1q2af1_1_1t2afb_1_1t2'afg_1_1Lcall_f_f_Int2_bufchan_buf  <= {163'd0,
                                                                                                                                                             1'd0};
    else
      if ((lizzieLet68_1_argbuf_r && \lizzieLet67_4Lcall_f_f_Int3_1sc_0_11_1q1af0_1_1t1afa_1_1t1'aff_1_1is_zaet_2_1op_addaeu_2_1q2af1_1_1t2afb_1_1t2'afg_1_1Lcall_f_f_Int2_bufchan_buf [0]))
        \lizzieLet67_4Lcall_f_f_Int3_1sc_0_11_1q1af0_1_1t1afa_1_1t1'aff_1_1is_zaet_2_1op_addaeu_2_1q2af1_1_1t2afb_1_1t2'afg_1_1Lcall_f_f_Int2_bufchan_buf  <= {163'd0,
                                                                                                                                                               1'd0};
      else if (((! lizzieLet68_1_argbuf_r) && (! \lizzieLet67_4Lcall_f_f_Int3_1sc_0_11_1q1af0_1_1t1afa_1_1t1'aff_1_1is_zaet_2_1op_addaeu_2_1q2af1_1_1t2afb_1_1t2'afg_1_1Lcall_f_f_Int2_bufchan_buf [0])))
        \lizzieLet67_4Lcall_f_f_Int3_1sc_0_11_1q1af0_1_1t1afa_1_1t1'aff_1_1is_zaet_2_1op_addaeu_2_1q2af1_1_1t2afb_1_1t2'afg_1_1Lcall_f_f_Int2_bufchan_buf  <= \lizzieLet67_4Lcall_f_f_Int3_1sc_0_11_1q1af0_1_1t1afa_1_1t1'aff_1_1is_zaet_2_1op_addaeu_2_1q2af1_1_1t2afb_1_1t2'afg_1_1Lcall_f_f_Int2_bufchan_d ;
  
  /* fork (Ty Pointer_QTree_Int) : (lizzieLet67_4Lf_f_Intsbos,Pointer_QTree_Int) > [(lizzieLet67_4Lf_f_Intsbos_1_merge_merge_merge_fork_1,Pointer_QTree_Int),
                                                                               (lizzieLet67_4Lf_f_Intsbos_1_merge_merge_merge_fork_2,Pointer_QTree_Int)] */
  logic [1:0] lizzieLet67_4Lf_f_Intsbos_emitted;
  logic [1:0] lizzieLet67_4Lf_f_Intsbos_done;
  assign lizzieLet67_4Lf_f_Intsbos_1_merge_merge_merge_fork_1_d = {lizzieLet67_4Lf_f_Intsbos_d[16:1],
                                                                   (lizzieLet67_4Lf_f_Intsbos_d[0] && (! lizzieLet67_4Lf_f_Intsbos_emitted[0]))};
  assign lizzieLet67_4Lf_f_Intsbos_1_merge_merge_merge_fork_2_d = {lizzieLet67_4Lf_f_Intsbos_d[16:1],
                                                                   (lizzieLet67_4Lf_f_Intsbos_d[0] && (! lizzieLet67_4Lf_f_Intsbos_emitted[1]))};
  assign lizzieLet67_4Lf_f_Intsbos_done = (lizzieLet67_4Lf_f_Intsbos_emitted | ({lizzieLet67_4Lf_f_Intsbos_1_merge_merge_merge_fork_2_d[0],
                                                                                 lizzieLet67_4Lf_f_Intsbos_1_merge_merge_merge_fork_1_d[0]} & {lizzieLet67_4Lf_f_Intsbos_1_merge_merge_merge_fork_2_r,
                                                                                                                                               lizzieLet67_4Lf_f_Intsbos_1_merge_merge_merge_fork_1_r}));
  assign lizzieLet67_4Lf_f_Intsbos_r = (& lizzieLet67_4Lf_f_Intsbos_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet67_4Lf_f_Intsbos_emitted <= 2'd0;
    else
      lizzieLet67_4Lf_f_Intsbos_emitted <= (lizzieLet67_4Lf_f_Intsbos_r ? 2'd0 :
                                            lizzieLet67_4Lf_f_Intsbos_done);
  
  /* togo (Ty Pointer_QTree_Int) : (lizzieLet67_4Lf_f_Intsbos_1_merge_merge_merge_fork_1,Pointer_QTree_Int) > (call_f_f_Int_goConst,Go) */
  assign call_f_f_Int_goConst_d = lizzieLet67_4Lf_f_Intsbos_1_merge_merge_merge_fork_1_d[0];
  assign lizzieLet67_4Lf_f_Intsbos_1_merge_merge_merge_fork_1_r = call_f_f_Int_goConst_r;
  
  /* buf (Ty Pointer_QTree_Int) : (lizzieLet67_4Lf_f_Intsbos_1_merge_merge_merge_fork_2,Pointer_QTree_Int) > (f_f_Int_resbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t lizzieLet67_4Lf_f_Intsbos_1_merge_merge_merge_fork_2_bufchan_d;
  logic lizzieLet67_4Lf_f_Intsbos_1_merge_merge_merge_fork_2_bufchan_r;
  assign lizzieLet67_4Lf_f_Intsbos_1_merge_merge_merge_fork_2_r = ((! lizzieLet67_4Lf_f_Intsbos_1_merge_merge_merge_fork_2_bufchan_d[0]) || lizzieLet67_4Lf_f_Intsbos_1_merge_merge_merge_fork_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet67_4Lf_f_Intsbos_1_merge_merge_merge_fork_2_bufchan_d <= {16'd0,
                                                                         1'd0};
    else
      if (lizzieLet67_4Lf_f_Intsbos_1_merge_merge_merge_fork_2_r)
        lizzieLet67_4Lf_f_Intsbos_1_merge_merge_merge_fork_2_bufchan_d <= lizzieLet67_4Lf_f_Intsbos_1_merge_merge_merge_fork_2_d;
  Pointer_QTree_Int_t lizzieLet67_4Lf_f_Intsbos_1_merge_merge_merge_fork_2_bufchan_buf;
  assign lizzieLet67_4Lf_f_Intsbos_1_merge_merge_merge_fork_2_bufchan_r = (! lizzieLet67_4Lf_f_Intsbos_1_merge_merge_merge_fork_2_bufchan_buf[0]);
  assign f_f_Int_resbuf_d = (lizzieLet67_4Lf_f_Intsbos_1_merge_merge_merge_fork_2_bufchan_buf[0] ? lizzieLet67_4Lf_f_Intsbos_1_merge_merge_merge_fork_2_bufchan_buf :
                             lizzieLet67_4Lf_f_Intsbos_1_merge_merge_merge_fork_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet67_4Lf_f_Intsbos_1_merge_merge_merge_fork_2_bufchan_buf <= {16'd0,
                                                                           1'd0};
    else
      if ((f_f_Int_resbuf_r && lizzieLet67_4Lf_f_Intsbos_1_merge_merge_merge_fork_2_bufchan_buf[0]))
        lizzieLet67_4Lf_f_Intsbos_1_merge_merge_merge_fork_2_bufchan_buf <= {16'd0,
                                                                             1'd0};
      else if (((! f_f_Int_resbuf_r) && (! lizzieLet67_4Lf_f_Intsbos_1_merge_merge_merge_fork_2_bufchan_buf[0])))
        lizzieLet67_4Lf_f_Intsbos_1_merge_merge_merge_fork_2_bufchan_buf <= lizzieLet67_4Lf_f_Intsbos_1_merge_merge_merge_fork_2_bufchan_d;
  
  /* destruct (Ty QTree_Int,
          Dcon QNode_Int) : (lizzieLet6_1QNode_Int,QTree_Int) > [(q1aft_destruct,Pointer_QTree_Int),
                                                                 (q2afu_destruct,Pointer_QTree_Int),
                                                                 (q3afv_destruct,Pointer_QTree_Int),
                                                                 (q5afw_destruct,Pointer_QTree_Int)] */
  logic [3:0] lizzieLet6_1QNode_Int_emitted;
  logic [3:0] lizzieLet6_1QNode_Int_done;
  assign q1aft_destruct_d = {lizzieLet6_1QNode_Int_d[18:3],
                             (lizzieLet6_1QNode_Int_d[0] && (! lizzieLet6_1QNode_Int_emitted[0]))};
  assign q2afu_destruct_d = {lizzieLet6_1QNode_Int_d[34:19],
                             (lizzieLet6_1QNode_Int_d[0] && (! lizzieLet6_1QNode_Int_emitted[1]))};
  assign q3afv_destruct_d = {lizzieLet6_1QNode_Int_d[50:35],
                             (lizzieLet6_1QNode_Int_d[0] && (! lizzieLet6_1QNode_Int_emitted[2]))};
  assign q5afw_destruct_d = {lizzieLet6_1QNode_Int_d[66:51],
                             (lizzieLet6_1QNode_Int_d[0] && (! lizzieLet6_1QNode_Int_emitted[3]))};
  assign lizzieLet6_1QNode_Int_done = (lizzieLet6_1QNode_Int_emitted | ({q5afw_destruct_d[0],
                                                                         q3afv_destruct_d[0],
                                                                         q2afu_destruct_d[0],
                                                                         q1aft_destruct_d[0]} & {q5afw_destruct_r,
                                                                                                 q3afv_destruct_r,
                                                                                                 q2afu_destruct_r,
                                                                                                 q1aft_destruct_r}));
  assign lizzieLet6_1QNode_Int_r = (& lizzieLet6_1QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_1QNode_Int_emitted <= 4'd0;
    else
      lizzieLet6_1QNode_Int_emitted <= (lizzieLet6_1QNode_Int_r ? 4'd0 :
                                        lizzieLet6_1QNode_Int_done);
  
  /* destruct (Ty QTree_Int,
          Dcon QVal_Int) : (lizzieLet6_1QVal_Int,QTree_Int) > [(v1afn_destruct,Int)] */
  assign v1afn_destruct_d = {lizzieLet6_1QVal_Int_d[34:3],
                             lizzieLet6_1QVal_Int_d[0]};
  assign lizzieLet6_1QVal_Int_r = v1afn_destruct_r;
  
  /* demux (Ty QTree_Int,
       Ty QTree_Int) : (lizzieLet6_2,QTree_Int) (lizzieLet6_1,QTree_Int) > [(_51,QTree_Int),
                                                                            (lizzieLet6_1QVal_Int,QTree_Int),
                                                                            (lizzieLet6_1QNode_Int,QTree_Int),
                                                                            (_50,QTree_Int)] */
  logic [3:0] lizzieLet6_1_onehotd;
  always_comb
    if ((lizzieLet6_2_d[0] && lizzieLet6_1_d[0]))
      unique case (lizzieLet6_2_d[2:1])
        2'd0: lizzieLet6_1_onehotd = 4'd1;
        2'd1: lizzieLet6_1_onehotd = 4'd2;
        2'd2: lizzieLet6_1_onehotd = 4'd4;
        2'd3: lizzieLet6_1_onehotd = 4'd8;
        default: lizzieLet6_1_onehotd = 4'd0;
      endcase
    else lizzieLet6_1_onehotd = 4'd0;
  assign _51_d = {lizzieLet6_1_d[66:1], lizzieLet6_1_onehotd[0]};
  assign lizzieLet6_1QVal_Int_d = {lizzieLet6_1_d[66:1],
                                   lizzieLet6_1_onehotd[1]};
  assign lizzieLet6_1QNode_Int_d = {lizzieLet6_1_d[66:1],
                                    lizzieLet6_1_onehotd[2]};
  assign _50_d = {lizzieLet6_1_d[66:1], lizzieLet6_1_onehotd[3]};
  assign lizzieLet6_1_r = (| (lizzieLet6_1_onehotd & {_50_r,
                                                      lizzieLet6_1QNode_Int_r,
                                                      lizzieLet6_1QVal_Int_r,
                                                      _51_r}));
  assign lizzieLet6_2_r = lizzieLet6_1_r;
  
  /* demux (Ty QTree_Int,
       Ty Go) : (lizzieLet6_3,QTree_Int) (go_9_goMux_data,Go) > [(lizzieLet6_3QNone_Int,Go),
                                                                 (lizzieLet6_3QVal_Int,Go),
                                                                 (lizzieLet6_3QNode_Int,Go),
                                                                 (lizzieLet6_3QError_Int,Go)] */
  logic [3:0] go_9_goMux_data_onehotd;
  always_comb
    if ((lizzieLet6_3_d[0] && go_9_goMux_data_d[0]))
      unique case (lizzieLet6_3_d[2:1])
        2'd0: go_9_goMux_data_onehotd = 4'd1;
        2'd1: go_9_goMux_data_onehotd = 4'd2;
        2'd2: go_9_goMux_data_onehotd = 4'd4;
        2'd3: go_9_goMux_data_onehotd = 4'd8;
        default: go_9_goMux_data_onehotd = 4'd0;
      endcase
    else go_9_goMux_data_onehotd = 4'd0;
  assign lizzieLet6_3QNone_Int_d = go_9_goMux_data_onehotd[0];
  assign lizzieLet6_3QVal_Int_d = go_9_goMux_data_onehotd[1];
  assign lizzieLet6_3QNode_Int_d = go_9_goMux_data_onehotd[2];
  assign lizzieLet6_3QError_Int_d = go_9_goMux_data_onehotd[3];
  assign go_9_goMux_data_r = (| (go_9_goMux_data_onehotd & {lizzieLet6_3QError_Int_r,
                                                            lizzieLet6_3QNode_Int_r,
                                                            lizzieLet6_3QVal_Int_r,
                                                            lizzieLet6_3QNone_Int_r}));
  assign lizzieLet6_3_r = go_9_goMux_data_r;
  
  /* fork (Ty Go) : (lizzieLet6_3QError_Int,Go) > [(lizzieLet6_3QError_Int_1,Go),
                                              (lizzieLet6_3QError_Int_2,Go)] */
  logic [1:0] lizzieLet6_3QError_Int_emitted;
  logic [1:0] lizzieLet6_3QError_Int_done;
  assign lizzieLet6_3QError_Int_1_d = (lizzieLet6_3QError_Int_d[0] && (! lizzieLet6_3QError_Int_emitted[0]));
  assign lizzieLet6_3QError_Int_2_d = (lizzieLet6_3QError_Int_d[0] && (! lizzieLet6_3QError_Int_emitted[1]));
  assign lizzieLet6_3QError_Int_done = (lizzieLet6_3QError_Int_emitted | ({lizzieLet6_3QError_Int_2_d[0],
                                                                           lizzieLet6_3QError_Int_1_d[0]} & {lizzieLet6_3QError_Int_2_r,
                                                                                                             lizzieLet6_3QError_Int_1_r}));
  assign lizzieLet6_3QError_Int_r = (& lizzieLet6_3QError_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_3QError_Int_emitted <= 2'd0;
    else
      lizzieLet6_3QError_Int_emitted <= (lizzieLet6_3QError_Int_r ? 2'd0 :
                                         lizzieLet6_3QError_Int_done);
  
  /* dcon (Ty QTree_Int,
      Dcon QError_Int) : [(lizzieLet6_3QError_Int_1,Go)] > (lizzieLet6_3QError_Int_1QError_Int,QTree_Int) */
  assign lizzieLet6_3QError_Int_1QError_Int_d = QError_Int_dc((& {lizzieLet6_3QError_Int_1_d[0]}), lizzieLet6_3QError_Int_1_d);
  assign {lizzieLet6_3QError_Int_1_r} = {1 {(lizzieLet6_3QError_Int_1QError_Int_r && lizzieLet6_3QError_Int_1QError_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (lizzieLet6_3QError_Int_1QError_Int,QTree_Int) > (lizzieLet16_1_argbuf,QTree_Int) */
  QTree_Int_t lizzieLet6_3QError_Int_1QError_Int_bufchan_d;
  logic lizzieLet6_3QError_Int_1QError_Int_bufchan_r;
  assign lizzieLet6_3QError_Int_1QError_Int_r = ((! lizzieLet6_3QError_Int_1QError_Int_bufchan_d[0]) || lizzieLet6_3QError_Int_1QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_3QError_Int_1QError_Int_bufchan_d <= {66'd0, 1'd0};
    else
      if (lizzieLet6_3QError_Int_1QError_Int_r)
        lizzieLet6_3QError_Int_1QError_Int_bufchan_d <= lizzieLet6_3QError_Int_1QError_Int_d;
  QTree_Int_t lizzieLet6_3QError_Int_1QError_Int_bufchan_buf;
  assign lizzieLet6_3QError_Int_1QError_Int_bufchan_r = (! lizzieLet6_3QError_Int_1QError_Int_bufchan_buf[0]);
  assign lizzieLet16_1_argbuf_d = (lizzieLet6_3QError_Int_1QError_Int_bufchan_buf[0] ? lizzieLet6_3QError_Int_1QError_Int_bufchan_buf :
                                   lizzieLet6_3QError_Int_1QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_3QError_Int_1QError_Int_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((lizzieLet16_1_argbuf_r && lizzieLet6_3QError_Int_1QError_Int_bufchan_buf[0]))
        lizzieLet6_3QError_Int_1QError_Int_bufchan_buf <= {66'd0, 1'd0};
      else if (((! lizzieLet16_1_argbuf_r) && (! lizzieLet6_3QError_Int_1QError_Int_bufchan_buf[0])))
        lizzieLet6_3QError_Int_1QError_Int_bufchan_buf <= lizzieLet6_3QError_Int_1QError_Int_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet6_3QError_Int_2,Go) > (lizzieLet6_3QError_Int_2_argbuf,Go) */
  Go_t lizzieLet6_3QError_Int_2_bufchan_d;
  logic lizzieLet6_3QError_Int_2_bufchan_r;
  assign lizzieLet6_3QError_Int_2_r = ((! lizzieLet6_3QError_Int_2_bufchan_d[0]) || lizzieLet6_3QError_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_3QError_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet6_3QError_Int_2_r)
        lizzieLet6_3QError_Int_2_bufchan_d <= lizzieLet6_3QError_Int_2_d;
  Go_t lizzieLet6_3QError_Int_2_bufchan_buf;
  assign lizzieLet6_3QError_Int_2_bufchan_r = (! lizzieLet6_3QError_Int_2_bufchan_buf[0]);
  assign lizzieLet6_3QError_Int_2_argbuf_d = (lizzieLet6_3QError_Int_2_bufchan_buf[0] ? lizzieLet6_3QError_Int_2_bufchan_buf :
                                              lizzieLet6_3QError_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_3QError_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet6_3QError_Int_2_argbuf_r && lizzieLet6_3QError_Int_2_bufchan_buf[0]))
        lizzieLet6_3QError_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet6_3QError_Int_2_argbuf_r) && (! lizzieLet6_3QError_Int_2_bufchan_buf[0])))
        lizzieLet6_3QError_Int_2_bufchan_buf <= lizzieLet6_3QError_Int_2_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet6_3QNone_Int,Go) > (lizzieLet6_3QNone_Int_1_argbuf,Go) */
  Go_t lizzieLet6_3QNone_Int_bufchan_d;
  logic lizzieLet6_3QNone_Int_bufchan_r;
  assign lizzieLet6_3QNone_Int_r = ((! lizzieLet6_3QNone_Int_bufchan_d[0]) || lizzieLet6_3QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_3QNone_Int_bufchan_d <= 1'd0;
    else
      if (lizzieLet6_3QNone_Int_r)
        lizzieLet6_3QNone_Int_bufchan_d <= lizzieLet6_3QNone_Int_d;
  Go_t lizzieLet6_3QNone_Int_bufchan_buf;
  assign lizzieLet6_3QNone_Int_bufchan_r = (! lizzieLet6_3QNone_Int_bufchan_buf[0]);
  assign lizzieLet6_3QNone_Int_1_argbuf_d = (lizzieLet6_3QNone_Int_bufchan_buf[0] ? lizzieLet6_3QNone_Int_bufchan_buf :
                                             lizzieLet6_3QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_3QNone_Int_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet6_3QNone_Int_1_argbuf_r && lizzieLet6_3QNone_Int_bufchan_buf[0]))
        lizzieLet6_3QNone_Int_bufchan_buf <= 1'd0;
      else if (((! lizzieLet6_3QNone_Int_1_argbuf_r) && (! lizzieLet6_3QNone_Int_bufchan_buf[0])))
        lizzieLet6_3QNone_Int_bufchan_buf <= lizzieLet6_3QNone_Int_bufchan_d;
  
  /* mergectrl (Ty C11,Ty Go) : [(lizzieLet6_3QNone_Int_1_argbuf,Go),
                            (lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int0_1_argbuf,Go),
                            (lizzieLet6_5QVal_Int_3QNone_Int_1_argbuf,Go),
                            (es_2_1MyFalse_1_argbuf,Go),
                            (es_2_1MyTrue_2_argbuf,Go),
                            (lizzieLet6_5QVal_Int_3QNode_Int_2_argbuf,Go),
                            (lizzieLet6_5QVal_Int_3QError_Int_2_argbuf,Go),
                            (lizzieLet6_5QNode_Int_3QNone_Int_1_argbuf,Go),
                            (lizzieLet6_5QNode_Int_3QVal_Int_2_argbuf,Go),
                            (lizzieLet6_5QNode_Int_3QError_Int_2_argbuf,Go),
                            (lizzieLet6_3QError_Int_2_argbuf,Go)] > (go_14_goMux_choice,C11) (go_14_goMux_data,Go) */
  logic [10:0] lizzieLet6_3QNone_Int_1_argbuf_select_d;
  assign lizzieLet6_3QNone_Int_1_argbuf_select_d = ((| lizzieLet6_3QNone_Int_1_argbuf_select_q) ? lizzieLet6_3QNone_Int_1_argbuf_select_q :
                                                    (lizzieLet6_3QNone_Int_1_argbuf_d[0] ? 11'd1 :
                                                     (\lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int0_1_argbuf_d [0] ? 11'd2 :
                                                      (lizzieLet6_5QVal_Int_3QNone_Int_1_argbuf_d[0] ? 11'd4 :
                                                       (es_2_1MyFalse_1_argbuf_d[0] ? 11'd8 :
                                                        (es_2_1MyTrue_2_argbuf_d[0] ? 11'd16 :
                                                         (lizzieLet6_5QVal_Int_3QNode_Int_2_argbuf_d[0] ? 11'd32 :
                                                          (lizzieLet6_5QVal_Int_3QError_Int_2_argbuf_d[0] ? 11'd64 :
                                                           (lizzieLet6_5QNode_Int_3QNone_Int_1_argbuf_d[0] ? 11'd128 :
                                                            (lizzieLet6_5QNode_Int_3QVal_Int_2_argbuf_d[0] ? 11'd256 :
                                                             (lizzieLet6_5QNode_Int_3QError_Int_2_argbuf_d[0] ? 11'd512 :
                                                              (lizzieLet6_3QError_Int_2_argbuf_d[0] ? 11'd1024 :
                                                               11'd0))))))))))));
  logic [10:0] lizzieLet6_3QNone_Int_1_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_3QNone_Int_1_argbuf_select_q <= 11'd0;
    else
      lizzieLet6_3QNone_Int_1_argbuf_select_q <= (lizzieLet6_3QNone_Int_1_argbuf_done ? 11'd0 :
                                                  lizzieLet6_3QNone_Int_1_argbuf_select_d);
  logic [1:0] lizzieLet6_3QNone_Int_1_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_3QNone_Int_1_argbuf_emit_q <= 2'd0;
    else
      lizzieLet6_3QNone_Int_1_argbuf_emit_q <= (lizzieLet6_3QNone_Int_1_argbuf_done ? 2'd0 :
                                                lizzieLet6_3QNone_Int_1_argbuf_emit_d);
  logic [1:0] lizzieLet6_3QNone_Int_1_argbuf_emit_d;
  assign lizzieLet6_3QNone_Int_1_argbuf_emit_d = (lizzieLet6_3QNone_Int_1_argbuf_emit_q | ({go_14_goMux_choice_d[0],
                                                                                            go_14_goMux_data_d[0]} & {go_14_goMux_choice_r,
                                                                                                                      go_14_goMux_data_r}));
  logic lizzieLet6_3QNone_Int_1_argbuf_done;
  assign lizzieLet6_3QNone_Int_1_argbuf_done = (& lizzieLet6_3QNone_Int_1_argbuf_emit_d);
  assign {lizzieLet6_3QError_Int_2_argbuf_r,
          lizzieLet6_5QNode_Int_3QError_Int_2_argbuf_r,
          lizzieLet6_5QNode_Int_3QVal_Int_2_argbuf_r,
          lizzieLet6_5QNode_Int_3QNone_Int_1_argbuf_r,
          lizzieLet6_5QVal_Int_3QError_Int_2_argbuf_r,
          lizzieLet6_5QVal_Int_3QNode_Int_2_argbuf_r,
          es_2_1MyTrue_2_argbuf_r,
          es_2_1MyFalse_1_argbuf_r,
          lizzieLet6_5QVal_Int_3QNone_Int_1_argbuf_r,
          \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int0_1_argbuf_r ,
          lizzieLet6_3QNone_Int_1_argbuf_r} = (lizzieLet6_3QNone_Int_1_argbuf_done ? lizzieLet6_3QNone_Int_1_argbuf_select_d :
                                               11'd0);
  assign go_14_goMux_data_d = ((lizzieLet6_3QNone_Int_1_argbuf_select_d[0] && (! lizzieLet6_3QNone_Int_1_argbuf_emit_q[0])) ? lizzieLet6_3QNone_Int_1_argbuf_d :
                               ((lizzieLet6_3QNone_Int_1_argbuf_select_d[1] && (! lizzieLet6_3QNone_Int_1_argbuf_emit_q[0])) ? \lizzieLet62_3Lcall_f''''''''''''_f''''''''''''_Int0_1_argbuf_d  :
                                ((lizzieLet6_3QNone_Int_1_argbuf_select_d[2] && (! lizzieLet6_3QNone_Int_1_argbuf_emit_q[0])) ? lizzieLet6_5QVal_Int_3QNone_Int_1_argbuf_d :
                                 ((lizzieLet6_3QNone_Int_1_argbuf_select_d[3] && (! lizzieLet6_3QNone_Int_1_argbuf_emit_q[0])) ? es_2_1MyFalse_1_argbuf_d :
                                  ((lizzieLet6_3QNone_Int_1_argbuf_select_d[4] && (! lizzieLet6_3QNone_Int_1_argbuf_emit_q[0])) ? es_2_1MyTrue_2_argbuf_d :
                                   ((lizzieLet6_3QNone_Int_1_argbuf_select_d[5] && (! lizzieLet6_3QNone_Int_1_argbuf_emit_q[0])) ? lizzieLet6_5QVal_Int_3QNode_Int_2_argbuf_d :
                                    ((lizzieLet6_3QNone_Int_1_argbuf_select_d[6] && (! lizzieLet6_3QNone_Int_1_argbuf_emit_q[0])) ? lizzieLet6_5QVal_Int_3QError_Int_2_argbuf_d :
                                     ((lizzieLet6_3QNone_Int_1_argbuf_select_d[7] && (! lizzieLet6_3QNone_Int_1_argbuf_emit_q[0])) ? lizzieLet6_5QNode_Int_3QNone_Int_1_argbuf_d :
                                      ((lizzieLet6_3QNone_Int_1_argbuf_select_d[8] && (! lizzieLet6_3QNone_Int_1_argbuf_emit_q[0])) ? lizzieLet6_5QNode_Int_3QVal_Int_2_argbuf_d :
                                       ((lizzieLet6_3QNone_Int_1_argbuf_select_d[9] && (! lizzieLet6_3QNone_Int_1_argbuf_emit_q[0])) ? lizzieLet6_5QNode_Int_3QError_Int_2_argbuf_d :
                                        ((lizzieLet6_3QNone_Int_1_argbuf_select_d[10] && (! lizzieLet6_3QNone_Int_1_argbuf_emit_q[0])) ? lizzieLet6_3QError_Int_2_argbuf_d :
                                         1'd0)))))))))));
  assign go_14_goMux_choice_d = ((lizzieLet6_3QNone_Int_1_argbuf_select_d[0] && (! lizzieLet6_3QNone_Int_1_argbuf_emit_q[1])) ? C1_11_dc(1'd1) :
                                 ((lizzieLet6_3QNone_Int_1_argbuf_select_d[1] && (! lizzieLet6_3QNone_Int_1_argbuf_emit_q[1])) ? C2_11_dc(1'd1) :
                                  ((lizzieLet6_3QNone_Int_1_argbuf_select_d[2] && (! lizzieLet6_3QNone_Int_1_argbuf_emit_q[1])) ? C3_11_dc(1'd1) :
                                   ((lizzieLet6_3QNone_Int_1_argbuf_select_d[3] && (! lizzieLet6_3QNone_Int_1_argbuf_emit_q[1])) ? C4_11_dc(1'd1) :
                                    ((lizzieLet6_3QNone_Int_1_argbuf_select_d[4] && (! lizzieLet6_3QNone_Int_1_argbuf_emit_q[1])) ? C5_11_dc(1'd1) :
                                     ((lizzieLet6_3QNone_Int_1_argbuf_select_d[5] && (! lizzieLet6_3QNone_Int_1_argbuf_emit_q[1])) ? C6_11_dc(1'd1) :
                                      ((lizzieLet6_3QNone_Int_1_argbuf_select_d[6] && (! lizzieLet6_3QNone_Int_1_argbuf_emit_q[1])) ? C7_11_dc(1'd1) :
                                       ((lizzieLet6_3QNone_Int_1_argbuf_select_d[7] && (! lizzieLet6_3QNone_Int_1_argbuf_emit_q[1])) ? C8_11_dc(1'd1) :
                                        ((lizzieLet6_3QNone_Int_1_argbuf_select_d[8] && (! lizzieLet6_3QNone_Int_1_argbuf_emit_q[1])) ? C9_11_dc(1'd1) :
                                         ((lizzieLet6_3QNone_Int_1_argbuf_select_d[9] && (! lizzieLet6_3QNone_Int_1_argbuf_emit_q[1])) ? C10_11_dc(1'd1) :
                                          ((lizzieLet6_3QNone_Int_1_argbuf_select_d[10] && (! lizzieLet6_3QNone_Int_1_argbuf_emit_q[1])) ? C11_11_dc(1'd1) :
                                           {4'd0, 1'd0})))))))))));
  
  /* demux (Ty QTree_Int,
       Ty MyDTInt_Bool) : (lizzieLet6_4,QTree_Int) (is_zafl_goMux_mux,MyDTInt_Bool) > [(_49,MyDTInt_Bool),
                                                                                       (lizzieLet6_4QVal_Int,MyDTInt_Bool),
                                                                                       (lizzieLet6_4QNode_Int,MyDTInt_Bool),
                                                                                       (_48,MyDTInt_Bool)] */
  logic [3:0] is_zafl_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet6_4_d[0] && is_zafl_goMux_mux_d[0]))
      unique case (lizzieLet6_4_d[2:1])
        2'd0: is_zafl_goMux_mux_onehotd = 4'd1;
        2'd1: is_zafl_goMux_mux_onehotd = 4'd2;
        2'd2: is_zafl_goMux_mux_onehotd = 4'd4;
        2'd3: is_zafl_goMux_mux_onehotd = 4'd8;
        default: is_zafl_goMux_mux_onehotd = 4'd0;
      endcase
    else is_zafl_goMux_mux_onehotd = 4'd0;
  assign _49_d = is_zafl_goMux_mux_onehotd[0];
  assign lizzieLet6_4QVal_Int_d = is_zafl_goMux_mux_onehotd[1];
  assign lizzieLet6_4QNode_Int_d = is_zafl_goMux_mux_onehotd[2];
  assign _48_d = is_zafl_goMux_mux_onehotd[3];
  assign is_zafl_goMux_mux_r = (| (is_zafl_goMux_mux_onehotd & {_48_r,
                                                                lizzieLet6_4QNode_Int_r,
                                                                lizzieLet6_4QVal_Int_r,
                                                                _49_r}));
  assign lizzieLet6_4_r = is_zafl_goMux_mux_r;
  
  /* demux (Ty QTree_Int,
       Ty QTree_Int) : (lizzieLet6_5,QTree_Int) (readPointer_QTree_Intt4afk_1_argbuf_rwb,QTree_Int) > [(_47,QTree_Int),
                                                                                                       (lizzieLet6_5QVal_Int,QTree_Int),
                                                                                                       (lizzieLet6_5QNode_Int,QTree_Int),
                                                                                                       (_46,QTree_Int)] */
  logic [3:0] readPointer_QTree_Intt4afk_1_argbuf_rwb_onehotd;
  always_comb
    if ((lizzieLet6_5_d[0] && readPointer_QTree_Intt4afk_1_argbuf_rwb_d[0]))
      unique case (lizzieLet6_5_d[2:1])
        2'd0: readPointer_QTree_Intt4afk_1_argbuf_rwb_onehotd = 4'd1;
        2'd1: readPointer_QTree_Intt4afk_1_argbuf_rwb_onehotd = 4'd2;
        2'd2: readPointer_QTree_Intt4afk_1_argbuf_rwb_onehotd = 4'd4;
        2'd3: readPointer_QTree_Intt4afk_1_argbuf_rwb_onehotd = 4'd8;
        default: readPointer_QTree_Intt4afk_1_argbuf_rwb_onehotd = 4'd0;
      endcase
    else readPointer_QTree_Intt4afk_1_argbuf_rwb_onehotd = 4'd0;
  assign _47_d = {readPointer_QTree_Intt4afk_1_argbuf_rwb_d[66:1],
                  readPointer_QTree_Intt4afk_1_argbuf_rwb_onehotd[0]};
  assign lizzieLet6_5QVal_Int_d = {readPointer_QTree_Intt4afk_1_argbuf_rwb_d[66:1],
                                   readPointer_QTree_Intt4afk_1_argbuf_rwb_onehotd[1]};
  assign lizzieLet6_5QNode_Int_d = {readPointer_QTree_Intt4afk_1_argbuf_rwb_d[66:1],
                                    readPointer_QTree_Intt4afk_1_argbuf_rwb_onehotd[2]};
  assign _46_d = {readPointer_QTree_Intt4afk_1_argbuf_rwb_d[66:1],
                  readPointer_QTree_Intt4afk_1_argbuf_rwb_onehotd[3]};
  assign readPointer_QTree_Intt4afk_1_argbuf_rwb_r = (| (readPointer_QTree_Intt4afk_1_argbuf_rwb_onehotd & {_46_r,
                                                                                                            lizzieLet6_5QNode_Int_r,
                                                                                                            lizzieLet6_5QVal_Int_r,
                                                                                                            _47_r}));
  assign lizzieLet6_5_r = readPointer_QTree_Intt4afk_1_argbuf_rwb_r;
  
  /* fork (Ty QTree_Int) : (lizzieLet6_5QNode_Int,QTree_Int) > [(lizzieLet6_5QNode_Int_1,QTree_Int),
                                                           (lizzieLet6_5QNode_Int_2,QTree_Int),
                                                           (lizzieLet6_5QNode_Int_3,QTree_Int),
                                                           (lizzieLet6_5QNode_Int_4,QTree_Int),
                                                           (lizzieLet6_5QNode_Int_5,QTree_Int),
                                                           (lizzieLet6_5QNode_Int_6,QTree_Int),
                                                           (lizzieLet6_5QNode_Int_7,QTree_Int),
                                                           (lizzieLet6_5QNode_Int_8,QTree_Int),
                                                           (lizzieLet6_5QNode_Int_9,QTree_Int),
                                                           (lizzieLet6_5QNode_Int_10,QTree_Int),
                                                           (lizzieLet6_5QNode_Int_11,QTree_Int)] */
  logic [10:0] lizzieLet6_5QNode_Int_emitted;
  logic [10:0] lizzieLet6_5QNode_Int_done;
  assign lizzieLet6_5QNode_Int_1_d = {lizzieLet6_5QNode_Int_d[66:1],
                                      (lizzieLet6_5QNode_Int_d[0] && (! lizzieLet6_5QNode_Int_emitted[0]))};
  assign lizzieLet6_5QNode_Int_2_d = {lizzieLet6_5QNode_Int_d[66:1],
                                      (lizzieLet6_5QNode_Int_d[0] && (! lizzieLet6_5QNode_Int_emitted[1]))};
  assign lizzieLet6_5QNode_Int_3_d = {lizzieLet6_5QNode_Int_d[66:1],
                                      (lizzieLet6_5QNode_Int_d[0] && (! lizzieLet6_5QNode_Int_emitted[2]))};
  assign lizzieLet6_5QNode_Int_4_d = {lizzieLet6_5QNode_Int_d[66:1],
                                      (lizzieLet6_5QNode_Int_d[0] && (! lizzieLet6_5QNode_Int_emitted[3]))};
  assign lizzieLet6_5QNode_Int_5_d = {lizzieLet6_5QNode_Int_d[66:1],
                                      (lizzieLet6_5QNode_Int_d[0] && (! lizzieLet6_5QNode_Int_emitted[4]))};
  assign lizzieLet6_5QNode_Int_6_d = {lizzieLet6_5QNode_Int_d[66:1],
                                      (lizzieLet6_5QNode_Int_d[0] && (! lizzieLet6_5QNode_Int_emitted[5]))};
  assign lizzieLet6_5QNode_Int_7_d = {lizzieLet6_5QNode_Int_d[66:1],
                                      (lizzieLet6_5QNode_Int_d[0] && (! lizzieLet6_5QNode_Int_emitted[6]))};
  assign lizzieLet6_5QNode_Int_8_d = {lizzieLet6_5QNode_Int_d[66:1],
                                      (lizzieLet6_5QNode_Int_d[0] && (! lizzieLet6_5QNode_Int_emitted[7]))};
  assign lizzieLet6_5QNode_Int_9_d = {lizzieLet6_5QNode_Int_d[66:1],
                                      (lizzieLet6_5QNode_Int_d[0] && (! lizzieLet6_5QNode_Int_emitted[8]))};
  assign lizzieLet6_5QNode_Int_10_d = {lizzieLet6_5QNode_Int_d[66:1],
                                       (lizzieLet6_5QNode_Int_d[0] && (! lizzieLet6_5QNode_Int_emitted[9]))};
  assign lizzieLet6_5QNode_Int_11_d = {lizzieLet6_5QNode_Int_d[66:1],
                                       (lizzieLet6_5QNode_Int_d[0] && (! lizzieLet6_5QNode_Int_emitted[10]))};
  assign lizzieLet6_5QNode_Int_done = (lizzieLet6_5QNode_Int_emitted | ({lizzieLet6_5QNode_Int_11_d[0],
                                                                         lizzieLet6_5QNode_Int_10_d[0],
                                                                         lizzieLet6_5QNode_Int_9_d[0],
                                                                         lizzieLet6_5QNode_Int_8_d[0],
                                                                         lizzieLet6_5QNode_Int_7_d[0],
                                                                         lizzieLet6_5QNode_Int_6_d[0],
                                                                         lizzieLet6_5QNode_Int_5_d[0],
                                                                         lizzieLet6_5QNode_Int_4_d[0],
                                                                         lizzieLet6_5QNode_Int_3_d[0],
                                                                         lizzieLet6_5QNode_Int_2_d[0],
                                                                         lizzieLet6_5QNode_Int_1_d[0]} & {lizzieLet6_5QNode_Int_11_r,
                                                                                                          lizzieLet6_5QNode_Int_10_r,
                                                                                                          lizzieLet6_5QNode_Int_9_r,
                                                                                                          lizzieLet6_5QNode_Int_8_r,
                                                                                                          lizzieLet6_5QNode_Int_7_r,
                                                                                                          lizzieLet6_5QNode_Int_6_r,
                                                                                                          lizzieLet6_5QNode_Int_5_r,
                                                                                                          lizzieLet6_5QNode_Int_4_r,
                                                                                                          lizzieLet6_5QNode_Int_3_r,
                                                                                                          lizzieLet6_5QNode_Int_2_r,
                                                                                                          lizzieLet6_5QNode_Int_1_r}));
  assign lizzieLet6_5QNode_Int_r = (& lizzieLet6_5QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_5QNode_Int_emitted <= 11'd0;
    else
      lizzieLet6_5QNode_Int_emitted <= (lizzieLet6_5QNode_Int_r ? 11'd0 :
                                        lizzieLet6_5QNode_Int_done);
  
  /* demux (Ty QTree_Int,
       Ty Pointer_QTree_Int) : (lizzieLet6_5QNode_Int_10,QTree_Int) (q3afv_destruct,Pointer_QTree_Int) > [(_45,Pointer_QTree_Int),
                                                                                                          (_44,Pointer_QTree_Int),
                                                                                                          (lizzieLet6_5QNode_Int_10QNode_Int,Pointer_QTree_Int),
                                                                                                          (_43,Pointer_QTree_Int)] */
  logic [3:0] q3afv_destruct_onehotd;
  always_comb
    if ((lizzieLet6_5QNode_Int_10_d[0] && q3afv_destruct_d[0]))
      unique case (lizzieLet6_5QNode_Int_10_d[2:1])
        2'd0: q3afv_destruct_onehotd = 4'd1;
        2'd1: q3afv_destruct_onehotd = 4'd2;
        2'd2: q3afv_destruct_onehotd = 4'd4;
        2'd3: q3afv_destruct_onehotd = 4'd8;
        default: q3afv_destruct_onehotd = 4'd0;
      endcase
    else q3afv_destruct_onehotd = 4'd0;
  assign _45_d = {q3afv_destruct_d[16:1], q3afv_destruct_onehotd[0]};
  assign _44_d = {q3afv_destruct_d[16:1], q3afv_destruct_onehotd[1]};
  assign lizzieLet6_5QNode_Int_10QNode_Int_d = {q3afv_destruct_d[16:1],
                                                q3afv_destruct_onehotd[2]};
  assign _43_d = {q3afv_destruct_d[16:1], q3afv_destruct_onehotd[3]};
  assign q3afv_destruct_r = (| (q3afv_destruct_onehotd & {_43_r,
                                                          lizzieLet6_5QNode_Int_10QNode_Int_r,
                                                          _44_r,
                                                          _45_r}));
  assign lizzieLet6_5QNode_Int_10_r = q3afv_destruct_r;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_QTree_Int) : (lizzieLet6_5QNode_Int_11,QTree_Int) (q5afw_destruct,Pointer_QTree_Int) > [(_42,Pointer_QTree_Int),
                                                                                                          (_41,Pointer_QTree_Int),
                                                                                                          (lizzieLet6_5QNode_Int_11QNode_Int,Pointer_QTree_Int),
                                                                                                          (_40,Pointer_QTree_Int)] */
  logic [3:0] q5afw_destruct_onehotd;
  always_comb
    if ((lizzieLet6_5QNode_Int_11_d[0] && q5afw_destruct_d[0]))
      unique case (lizzieLet6_5QNode_Int_11_d[2:1])
        2'd0: q5afw_destruct_onehotd = 4'd1;
        2'd1: q5afw_destruct_onehotd = 4'd2;
        2'd2: q5afw_destruct_onehotd = 4'd4;
        2'd3: q5afw_destruct_onehotd = 4'd8;
        default: q5afw_destruct_onehotd = 4'd0;
      endcase
    else q5afw_destruct_onehotd = 4'd0;
  assign _42_d = {q5afw_destruct_d[16:1], q5afw_destruct_onehotd[0]};
  assign _41_d = {q5afw_destruct_d[16:1], q5afw_destruct_onehotd[1]};
  assign lizzieLet6_5QNode_Int_11QNode_Int_d = {q5afw_destruct_d[16:1],
                                                q5afw_destruct_onehotd[2]};
  assign _40_d = {q5afw_destruct_d[16:1], q5afw_destruct_onehotd[3]};
  assign q5afw_destruct_r = (| (q5afw_destruct_onehotd & {_40_r,
                                                          lizzieLet6_5QNode_Int_11QNode_Int_r,
                                                          _41_r,
                                                          _42_r}));
  assign lizzieLet6_5QNode_Int_11_r = q5afw_destruct_r;
  
  /* buf (Ty Pointer_QTree_Int) : (lizzieLet6_5QNode_Int_11QNode_Int,Pointer_QTree_Int) > (lizzieLet6_5QNode_Int_11QNode_Int_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t lizzieLet6_5QNode_Int_11QNode_Int_bufchan_d;
  logic lizzieLet6_5QNode_Int_11QNode_Int_bufchan_r;
  assign lizzieLet6_5QNode_Int_11QNode_Int_r = ((! lizzieLet6_5QNode_Int_11QNode_Int_bufchan_d[0]) || lizzieLet6_5QNode_Int_11QNode_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_5QNode_Int_11QNode_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet6_5QNode_Int_11QNode_Int_r)
        lizzieLet6_5QNode_Int_11QNode_Int_bufchan_d <= lizzieLet6_5QNode_Int_11QNode_Int_d;
  Pointer_QTree_Int_t lizzieLet6_5QNode_Int_11QNode_Int_bufchan_buf;
  assign lizzieLet6_5QNode_Int_11QNode_Int_bufchan_r = (! lizzieLet6_5QNode_Int_11QNode_Int_bufchan_buf[0]);
  assign lizzieLet6_5QNode_Int_11QNode_Int_1_argbuf_d = (lizzieLet6_5QNode_Int_11QNode_Int_bufchan_buf[0] ? lizzieLet6_5QNode_Int_11QNode_Int_bufchan_buf :
                                                         lizzieLet6_5QNode_Int_11QNode_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_5QNode_Int_11QNode_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet6_5QNode_Int_11QNode_Int_1_argbuf_r && lizzieLet6_5QNode_Int_11QNode_Int_bufchan_buf[0]))
        lizzieLet6_5QNode_Int_11QNode_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet6_5QNode_Int_11QNode_Int_1_argbuf_r) && (! lizzieLet6_5QNode_Int_11QNode_Int_bufchan_buf[0])))
        lizzieLet6_5QNode_Int_11QNode_Int_bufchan_buf <= lizzieLet6_5QNode_Int_11QNode_Int_bufchan_d;
  
  /* destruct (Ty QTree_Int,
          Dcon QNode_Int) : (lizzieLet6_5QNode_Int_1QNode_Int,QTree_Int) > [(t1afy_destruct,Pointer_QTree_Int),
                                                                            (t2afz_destruct,Pointer_QTree_Int),
                                                                            (t3afA_destruct,Pointer_QTree_Int),
                                                                            (t5afB_destruct,Pointer_QTree_Int)] */
  logic [3:0] lizzieLet6_5QNode_Int_1QNode_Int_emitted;
  logic [3:0] lizzieLet6_5QNode_Int_1QNode_Int_done;
  assign t1afy_destruct_d = {lizzieLet6_5QNode_Int_1QNode_Int_d[18:3],
                             (lizzieLet6_5QNode_Int_1QNode_Int_d[0] && (! lizzieLet6_5QNode_Int_1QNode_Int_emitted[0]))};
  assign t2afz_destruct_d = {lizzieLet6_5QNode_Int_1QNode_Int_d[34:19],
                             (lizzieLet6_5QNode_Int_1QNode_Int_d[0] && (! lizzieLet6_5QNode_Int_1QNode_Int_emitted[1]))};
  assign t3afA_destruct_d = {lizzieLet6_5QNode_Int_1QNode_Int_d[50:35],
                             (lizzieLet6_5QNode_Int_1QNode_Int_d[0] && (! lizzieLet6_5QNode_Int_1QNode_Int_emitted[2]))};
  assign t5afB_destruct_d = {lizzieLet6_5QNode_Int_1QNode_Int_d[66:51],
                             (lizzieLet6_5QNode_Int_1QNode_Int_d[0] && (! lizzieLet6_5QNode_Int_1QNode_Int_emitted[3]))};
  assign lizzieLet6_5QNode_Int_1QNode_Int_done = (lizzieLet6_5QNode_Int_1QNode_Int_emitted | ({t5afB_destruct_d[0],
                                                                                               t3afA_destruct_d[0],
                                                                                               t2afz_destruct_d[0],
                                                                                               t1afy_destruct_d[0]} & {t5afB_destruct_r,
                                                                                                                       t3afA_destruct_r,
                                                                                                                       t2afz_destruct_r,
                                                                                                                       t1afy_destruct_r}));
  assign lizzieLet6_5QNode_Int_1QNode_Int_r = (& lizzieLet6_5QNode_Int_1QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_5QNode_Int_1QNode_Int_emitted <= 4'd0;
    else
      lizzieLet6_5QNode_Int_1QNode_Int_emitted <= (lizzieLet6_5QNode_Int_1QNode_Int_r ? 4'd0 :
                                                   lizzieLet6_5QNode_Int_1QNode_Int_done);
  
  /* demux (Ty QTree_Int,
       Ty QTree_Int) : (lizzieLet6_5QNode_Int_2,QTree_Int) (lizzieLet6_5QNode_Int_1,QTree_Int) > [(_39,QTree_Int),
                                                                                                  (_38,QTree_Int),
                                                                                                  (lizzieLet6_5QNode_Int_1QNode_Int,QTree_Int),
                                                                                                  (_37,QTree_Int)] */
  logic [3:0] lizzieLet6_5QNode_Int_1_onehotd;
  always_comb
    if ((lizzieLet6_5QNode_Int_2_d[0] && lizzieLet6_5QNode_Int_1_d[0]))
      unique case (lizzieLet6_5QNode_Int_2_d[2:1])
        2'd0: lizzieLet6_5QNode_Int_1_onehotd = 4'd1;
        2'd1: lizzieLet6_5QNode_Int_1_onehotd = 4'd2;
        2'd2: lizzieLet6_5QNode_Int_1_onehotd = 4'd4;
        2'd3: lizzieLet6_5QNode_Int_1_onehotd = 4'd8;
        default: lizzieLet6_5QNode_Int_1_onehotd = 4'd0;
      endcase
    else lizzieLet6_5QNode_Int_1_onehotd = 4'd0;
  assign _39_d = {lizzieLet6_5QNode_Int_1_d[66:1],
                  lizzieLet6_5QNode_Int_1_onehotd[0]};
  assign _38_d = {lizzieLet6_5QNode_Int_1_d[66:1],
                  lizzieLet6_5QNode_Int_1_onehotd[1]};
  assign lizzieLet6_5QNode_Int_1QNode_Int_d = {lizzieLet6_5QNode_Int_1_d[66:1],
                                               lizzieLet6_5QNode_Int_1_onehotd[2]};
  assign _37_d = {lizzieLet6_5QNode_Int_1_d[66:1],
                  lizzieLet6_5QNode_Int_1_onehotd[3]};
  assign lizzieLet6_5QNode_Int_1_r = (| (lizzieLet6_5QNode_Int_1_onehotd & {_37_r,
                                                                            lizzieLet6_5QNode_Int_1QNode_Int_r,
                                                                            _38_r,
                                                                            _39_r}));
  assign lizzieLet6_5QNode_Int_2_r = lizzieLet6_5QNode_Int_1_r;
  
  /* demux (Ty QTree_Int,
       Ty Go) : (lizzieLet6_5QNode_Int_3,QTree_Int) (lizzieLet6_3QNode_Int,Go) > [(lizzieLet6_5QNode_Int_3QNone_Int,Go),
                                                                                  (lizzieLet6_5QNode_Int_3QVal_Int,Go),
                                                                                  (lizzieLet6_5QNode_Int_3QNode_Int,Go),
                                                                                  (lizzieLet6_5QNode_Int_3QError_Int,Go)] */
  logic [3:0] lizzieLet6_3QNode_Int_onehotd;
  always_comb
    if ((lizzieLet6_5QNode_Int_3_d[0] && lizzieLet6_3QNode_Int_d[0]))
      unique case (lizzieLet6_5QNode_Int_3_d[2:1])
        2'd0: lizzieLet6_3QNode_Int_onehotd = 4'd1;
        2'd1: lizzieLet6_3QNode_Int_onehotd = 4'd2;
        2'd2: lizzieLet6_3QNode_Int_onehotd = 4'd4;
        2'd3: lizzieLet6_3QNode_Int_onehotd = 4'd8;
        default: lizzieLet6_3QNode_Int_onehotd = 4'd0;
      endcase
    else lizzieLet6_3QNode_Int_onehotd = 4'd0;
  assign lizzieLet6_5QNode_Int_3QNone_Int_d = lizzieLet6_3QNode_Int_onehotd[0];
  assign lizzieLet6_5QNode_Int_3QVal_Int_d = lizzieLet6_3QNode_Int_onehotd[1];
  assign lizzieLet6_5QNode_Int_3QNode_Int_d = lizzieLet6_3QNode_Int_onehotd[2];
  assign lizzieLet6_5QNode_Int_3QError_Int_d = lizzieLet6_3QNode_Int_onehotd[3];
  assign lizzieLet6_3QNode_Int_r = (| (lizzieLet6_3QNode_Int_onehotd & {lizzieLet6_5QNode_Int_3QError_Int_r,
                                                                        lizzieLet6_5QNode_Int_3QNode_Int_r,
                                                                        lizzieLet6_5QNode_Int_3QVal_Int_r,
                                                                        lizzieLet6_5QNode_Int_3QNone_Int_r}));
  assign lizzieLet6_5QNode_Int_3_r = lizzieLet6_3QNode_Int_r;
  
  /* fork (Ty Go) : (lizzieLet6_5QNode_Int_3QError_Int,Go) > [(lizzieLet6_5QNode_Int_3QError_Int_1,Go),
                                                         (lizzieLet6_5QNode_Int_3QError_Int_2,Go)] */
  logic [1:0] lizzieLet6_5QNode_Int_3QError_Int_emitted;
  logic [1:0] lizzieLet6_5QNode_Int_3QError_Int_done;
  assign lizzieLet6_5QNode_Int_3QError_Int_1_d = (lizzieLet6_5QNode_Int_3QError_Int_d[0] && (! lizzieLet6_5QNode_Int_3QError_Int_emitted[0]));
  assign lizzieLet6_5QNode_Int_3QError_Int_2_d = (lizzieLet6_5QNode_Int_3QError_Int_d[0] && (! lizzieLet6_5QNode_Int_3QError_Int_emitted[1]));
  assign lizzieLet6_5QNode_Int_3QError_Int_done = (lizzieLet6_5QNode_Int_3QError_Int_emitted | ({lizzieLet6_5QNode_Int_3QError_Int_2_d[0],
                                                                                                 lizzieLet6_5QNode_Int_3QError_Int_1_d[0]} & {lizzieLet6_5QNode_Int_3QError_Int_2_r,
                                                                                                                                              lizzieLet6_5QNode_Int_3QError_Int_1_r}));
  assign lizzieLet6_5QNode_Int_3QError_Int_r = (& lizzieLet6_5QNode_Int_3QError_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_5QNode_Int_3QError_Int_emitted <= 2'd0;
    else
      lizzieLet6_5QNode_Int_3QError_Int_emitted <= (lizzieLet6_5QNode_Int_3QError_Int_r ? 2'd0 :
                                                    lizzieLet6_5QNode_Int_3QError_Int_done);
  
  /* dcon (Ty QTree_Int,
      Dcon QError_Int) : [(lizzieLet6_5QNode_Int_3QError_Int_1,Go)] > (lizzieLet6_5QNode_Int_3QError_Int_1QError_Int,QTree_Int) */
  assign lizzieLet6_5QNode_Int_3QError_Int_1QError_Int_d = QError_Int_dc((& {lizzieLet6_5QNode_Int_3QError_Int_1_d[0]}), lizzieLet6_5QNode_Int_3QError_Int_1_d);
  assign {lizzieLet6_5QNode_Int_3QError_Int_1_r} = {1 {(lizzieLet6_5QNode_Int_3QError_Int_1QError_Int_r && lizzieLet6_5QNode_Int_3QError_Int_1QError_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (lizzieLet6_5QNode_Int_3QError_Int_1QError_Int,QTree_Int) > (lizzieLet15_1_argbuf,QTree_Int) */
  QTree_Int_t lizzieLet6_5QNode_Int_3QError_Int_1QError_Int_bufchan_d;
  logic lizzieLet6_5QNode_Int_3QError_Int_1QError_Int_bufchan_r;
  assign lizzieLet6_5QNode_Int_3QError_Int_1QError_Int_r = ((! lizzieLet6_5QNode_Int_3QError_Int_1QError_Int_bufchan_d[0]) || lizzieLet6_5QNode_Int_3QError_Int_1QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_5QNode_Int_3QError_Int_1QError_Int_bufchan_d <= {66'd0,
                                                                  1'd0};
    else
      if (lizzieLet6_5QNode_Int_3QError_Int_1QError_Int_r)
        lizzieLet6_5QNode_Int_3QError_Int_1QError_Int_bufchan_d <= lizzieLet6_5QNode_Int_3QError_Int_1QError_Int_d;
  QTree_Int_t lizzieLet6_5QNode_Int_3QError_Int_1QError_Int_bufchan_buf;
  assign lizzieLet6_5QNode_Int_3QError_Int_1QError_Int_bufchan_r = (! lizzieLet6_5QNode_Int_3QError_Int_1QError_Int_bufchan_buf[0]);
  assign lizzieLet15_1_argbuf_d = (lizzieLet6_5QNode_Int_3QError_Int_1QError_Int_bufchan_buf[0] ? lizzieLet6_5QNode_Int_3QError_Int_1QError_Int_bufchan_buf :
                                   lizzieLet6_5QNode_Int_3QError_Int_1QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_5QNode_Int_3QError_Int_1QError_Int_bufchan_buf <= {66'd0,
                                                                    1'd0};
    else
      if ((lizzieLet15_1_argbuf_r && lizzieLet6_5QNode_Int_3QError_Int_1QError_Int_bufchan_buf[0]))
        lizzieLet6_5QNode_Int_3QError_Int_1QError_Int_bufchan_buf <= {66'd0,
                                                                      1'd0};
      else if (((! lizzieLet15_1_argbuf_r) && (! lizzieLet6_5QNode_Int_3QError_Int_1QError_Int_bufchan_buf[0])))
        lizzieLet6_5QNode_Int_3QError_Int_1QError_Int_bufchan_buf <= lizzieLet6_5QNode_Int_3QError_Int_1QError_Int_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet6_5QNode_Int_3QError_Int_2,Go) > (lizzieLet6_5QNode_Int_3QError_Int_2_argbuf,Go) */
  Go_t lizzieLet6_5QNode_Int_3QError_Int_2_bufchan_d;
  logic lizzieLet6_5QNode_Int_3QError_Int_2_bufchan_r;
  assign lizzieLet6_5QNode_Int_3QError_Int_2_r = ((! lizzieLet6_5QNode_Int_3QError_Int_2_bufchan_d[0]) || lizzieLet6_5QNode_Int_3QError_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_5QNode_Int_3QError_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet6_5QNode_Int_3QError_Int_2_r)
        lizzieLet6_5QNode_Int_3QError_Int_2_bufchan_d <= lizzieLet6_5QNode_Int_3QError_Int_2_d;
  Go_t lizzieLet6_5QNode_Int_3QError_Int_2_bufchan_buf;
  assign lizzieLet6_5QNode_Int_3QError_Int_2_bufchan_r = (! lizzieLet6_5QNode_Int_3QError_Int_2_bufchan_buf[0]);
  assign lizzieLet6_5QNode_Int_3QError_Int_2_argbuf_d = (lizzieLet6_5QNode_Int_3QError_Int_2_bufchan_buf[0] ? lizzieLet6_5QNode_Int_3QError_Int_2_bufchan_buf :
                                                         lizzieLet6_5QNode_Int_3QError_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_5QNode_Int_3QError_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet6_5QNode_Int_3QError_Int_2_argbuf_r && lizzieLet6_5QNode_Int_3QError_Int_2_bufchan_buf[0]))
        lizzieLet6_5QNode_Int_3QError_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet6_5QNode_Int_3QError_Int_2_argbuf_r) && (! lizzieLet6_5QNode_Int_3QError_Int_2_bufchan_buf[0])))
        lizzieLet6_5QNode_Int_3QError_Int_2_bufchan_buf <= lizzieLet6_5QNode_Int_3QError_Int_2_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet6_5QNode_Int_3QNode_Int,Go) > (lizzieLet6_5QNode_Int_3QNode_Int_1_argbuf,Go) */
  Go_t lizzieLet6_5QNode_Int_3QNode_Int_bufchan_d;
  logic lizzieLet6_5QNode_Int_3QNode_Int_bufchan_r;
  assign lizzieLet6_5QNode_Int_3QNode_Int_r = ((! lizzieLet6_5QNode_Int_3QNode_Int_bufchan_d[0]) || lizzieLet6_5QNode_Int_3QNode_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_5QNode_Int_3QNode_Int_bufchan_d <= 1'd0;
    else
      if (lizzieLet6_5QNode_Int_3QNode_Int_r)
        lizzieLet6_5QNode_Int_3QNode_Int_bufchan_d <= lizzieLet6_5QNode_Int_3QNode_Int_d;
  Go_t lizzieLet6_5QNode_Int_3QNode_Int_bufchan_buf;
  assign lizzieLet6_5QNode_Int_3QNode_Int_bufchan_r = (! lizzieLet6_5QNode_Int_3QNode_Int_bufchan_buf[0]);
  assign lizzieLet6_5QNode_Int_3QNode_Int_1_argbuf_d = (lizzieLet6_5QNode_Int_3QNode_Int_bufchan_buf[0] ? lizzieLet6_5QNode_Int_3QNode_Int_bufchan_buf :
                                                        lizzieLet6_5QNode_Int_3QNode_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_5QNode_Int_3QNode_Int_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet6_5QNode_Int_3QNode_Int_1_argbuf_r && lizzieLet6_5QNode_Int_3QNode_Int_bufchan_buf[0]))
        lizzieLet6_5QNode_Int_3QNode_Int_bufchan_buf <= 1'd0;
      else if (((! lizzieLet6_5QNode_Int_3QNode_Int_1_argbuf_r) && (! lizzieLet6_5QNode_Int_3QNode_Int_bufchan_buf[0])))
        lizzieLet6_5QNode_Int_3QNode_Int_bufchan_buf <= lizzieLet6_5QNode_Int_3QNode_Int_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet6_5QNode_Int_3QNone_Int,Go) > (lizzieLet6_5QNode_Int_3QNone_Int_1_argbuf,Go) */
  Go_t lizzieLet6_5QNode_Int_3QNone_Int_bufchan_d;
  logic lizzieLet6_5QNode_Int_3QNone_Int_bufchan_r;
  assign lizzieLet6_5QNode_Int_3QNone_Int_r = ((! lizzieLet6_5QNode_Int_3QNone_Int_bufchan_d[0]) || lizzieLet6_5QNode_Int_3QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_5QNode_Int_3QNone_Int_bufchan_d <= 1'd0;
    else
      if (lizzieLet6_5QNode_Int_3QNone_Int_r)
        lizzieLet6_5QNode_Int_3QNone_Int_bufchan_d <= lizzieLet6_5QNode_Int_3QNone_Int_d;
  Go_t lizzieLet6_5QNode_Int_3QNone_Int_bufchan_buf;
  assign lizzieLet6_5QNode_Int_3QNone_Int_bufchan_r = (! lizzieLet6_5QNode_Int_3QNone_Int_bufchan_buf[0]);
  assign lizzieLet6_5QNode_Int_3QNone_Int_1_argbuf_d = (lizzieLet6_5QNode_Int_3QNone_Int_bufchan_buf[0] ? lizzieLet6_5QNode_Int_3QNone_Int_bufchan_buf :
                                                        lizzieLet6_5QNode_Int_3QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_5QNode_Int_3QNone_Int_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet6_5QNode_Int_3QNone_Int_1_argbuf_r && lizzieLet6_5QNode_Int_3QNone_Int_bufchan_buf[0]))
        lizzieLet6_5QNode_Int_3QNone_Int_bufchan_buf <= 1'd0;
      else if (((! lizzieLet6_5QNode_Int_3QNone_Int_1_argbuf_r) && (! lizzieLet6_5QNode_Int_3QNone_Int_bufchan_buf[0])))
        lizzieLet6_5QNode_Int_3QNone_Int_bufchan_buf <= lizzieLet6_5QNode_Int_3QNone_Int_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet6_5QNode_Int_3QVal_Int,Go) > [(lizzieLet6_5QNode_Int_3QVal_Int_1,Go),
                                                       (lizzieLet6_5QNode_Int_3QVal_Int_2,Go)] */
  logic [1:0] lizzieLet6_5QNode_Int_3QVal_Int_emitted;
  logic [1:0] lizzieLet6_5QNode_Int_3QVal_Int_done;
  assign lizzieLet6_5QNode_Int_3QVal_Int_1_d = (lizzieLet6_5QNode_Int_3QVal_Int_d[0] && (! lizzieLet6_5QNode_Int_3QVal_Int_emitted[0]));
  assign lizzieLet6_5QNode_Int_3QVal_Int_2_d = (lizzieLet6_5QNode_Int_3QVal_Int_d[0] && (! lizzieLet6_5QNode_Int_3QVal_Int_emitted[1]));
  assign lizzieLet6_5QNode_Int_3QVal_Int_done = (lizzieLet6_5QNode_Int_3QVal_Int_emitted | ({lizzieLet6_5QNode_Int_3QVal_Int_2_d[0],
                                                                                             lizzieLet6_5QNode_Int_3QVal_Int_1_d[0]} & {lizzieLet6_5QNode_Int_3QVal_Int_2_r,
                                                                                                                                        lizzieLet6_5QNode_Int_3QVal_Int_1_r}));
  assign lizzieLet6_5QNode_Int_3QVal_Int_r = (& lizzieLet6_5QNode_Int_3QVal_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_5QNode_Int_3QVal_Int_emitted <= 2'd0;
    else
      lizzieLet6_5QNode_Int_3QVal_Int_emitted <= (lizzieLet6_5QNode_Int_3QVal_Int_r ? 2'd0 :
                                                  lizzieLet6_5QNode_Int_3QVal_Int_done);
  
  /* dcon (Ty QTree_Int,
      Dcon QError_Int) : [(lizzieLet6_5QNode_Int_3QVal_Int_1,Go)] > (lizzieLet6_5QNode_Int_3QVal_Int_1QError_Int,QTree_Int) */
  assign lizzieLet6_5QNode_Int_3QVal_Int_1QError_Int_d = QError_Int_dc((& {lizzieLet6_5QNode_Int_3QVal_Int_1_d[0]}), lizzieLet6_5QNode_Int_3QVal_Int_1_d);
  assign {lizzieLet6_5QNode_Int_3QVal_Int_1_r} = {1 {(lizzieLet6_5QNode_Int_3QVal_Int_1QError_Int_r && lizzieLet6_5QNode_Int_3QVal_Int_1QError_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (lizzieLet6_5QNode_Int_3QVal_Int_1QError_Int,QTree_Int) > (lizzieLet13_1_argbuf,QTree_Int) */
  QTree_Int_t lizzieLet6_5QNode_Int_3QVal_Int_1QError_Int_bufchan_d;
  logic lizzieLet6_5QNode_Int_3QVal_Int_1QError_Int_bufchan_r;
  assign lizzieLet6_5QNode_Int_3QVal_Int_1QError_Int_r = ((! lizzieLet6_5QNode_Int_3QVal_Int_1QError_Int_bufchan_d[0]) || lizzieLet6_5QNode_Int_3QVal_Int_1QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_5QNode_Int_3QVal_Int_1QError_Int_bufchan_d <= {66'd0,
                                                                1'd0};
    else
      if (lizzieLet6_5QNode_Int_3QVal_Int_1QError_Int_r)
        lizzieLet6_5QNode_Int_3QVal_Int_1QError_Int_bufchan_d <= lizzieLet6_5QNode_Int_3QVal_Int_1QError_Int_d;
  QTree_Int_t lizzieLet6_5QNode_Int_3QVal_Int_1QError_Int_bufchan_buf;
  assign lizzieLet6_5QNode_Int_3QVal_Int_1QError_Int_bufchan_r = (! lizzieLet6_5QNode_Int_3QVal_Int_1QError_Int_bufchan_buf[0]);
  assign lizzieLet13_1_argbuf_d = (lizzieLet6_5QNode_Int_3QVal_Int_1QError_Int_bufchan_buf[0] ? lizzieLet6_5QNode_Int_3QVal_Int_1QError_Int_bufchan_buf :
                                   lizzieLet6_5QNode_Int_3QVal_Int_1QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_5QNode_Int_3QVal_Int_1QError_Int_bufchan_buf <= {66'd0,
                                                                  1'd0};
    else
      if ((lizzieLet13_1_argbuf_r && lizzieLet6_5QNode_Int_3QVal_Int_1QError_Int_bufchan_buf[0]))
        lizzieLet6_5QNode_Int_3QVal_Int_1QError_Int_bufchan_buf <= {66'd0,
                                                                    1'd0};
      else if (((! lizzieLet13_1_argbuf_r) && (! lizzieLet6_5QNode_Int_3QVal_Int_1QError_Int_bufchan_buf[0])))
        lizzieLet6_5QNode_Int_3QVal_Int_1QError_Int_bufchan_buf <= lizzieLet6_5QNode_Int_3QVal_Int_1QError_Int_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet6_5QNode_Int_3QVal_Int_2,Go) > (lizzieLet6_5QNode_Int_3QVal_Int_2_argbuf,Go) */
  Go_t lizzieLet6_5QNode_Int_3QVal_Int_2_bufchan_d;
  logic lizzieLet6_5QNode_Int_3QVal_Int_2_bufchan_r;
  assign lizzieLet6_5QNode_Int_3QVal_Int_2_r = ((! lizzieLet6_5QNode_Int_3QVal_Int_2_bufchan_d[0]) || lizzieLet6_5QNode_Int_3QVal_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_5QNode_Int_3QVal_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet6_5QNode_Int_3QVal_Int_2_r)
        lizzieLet6_5QNode_Int_3QVal_Int_2_bufchan_d <= lizzieLet6_5QNode_Int_3QVal_Int_2_d;
  Go_t lizzieLet6_5QNode_Int_3QVal_Int_2_bufchan_buf;
  assign lizzieLet6_5QNode_Int_3QVal_Int_2_bufchan_r = (! lizzieLet6_5QNode_Int_3QVal_Int_2_bufchan_buf[0]);
  assign lizzieLet6_5QNode_Int_3QVal_Int_2_argbuf_d = (lizzieLet6_5QNode_Int_3QVal_Int_2_bufchan_buf[0] ? lizzieLet6_5QNode_Int_3QVal_Int_2_bufchan_buf :
                                                       lizzieLet6_5QNode_Int_3QVal_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_5QNode_Int_3QVal_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet6_5QNode_Int_3QVal_Int_2_argbuf_r && lizzieLet6_5QNode_Int_3QVal_Int_2_bufchan_buf[0]))
        lizzieLet6_5QNode_Int_3QVal_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet6_5QNode_Int_3QVal_Int_2_argbuf_r) && (! lizzieLet6_5QNode_Int_3QVal_Int_2_bufchan_buf[0])))
        lizzieLet6_5QNode_Int_3QVal_Int_2_bufchan_buf <= lizzieLet6_5QNode_Int_3QVal_Int_2_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty MyDTInt_Bool) : (lizzieLet6_5QNode_Int_4,QTree_Int) (lizzieLet6_4QNode_Int,MyDTInt_Bool) > [(_36,MyDTInt_Bool),
                                                                                                      (_35,MyDTInt_Bool),
                                                                                                      (lizzieLet6_5QNode_Int_4QNode_Int,MyDTInt_Bool),
                                                                                                      (_34,MyDTInt_Bool)] */
  logic [3:0] lizzieLet6_4QNode_Int_onehotd;
  always_comb
    if ((lizzieLet6_5QNode_Int_4_d[0] && lizzieLet6_4QNode_Int_d[0]))
      unique case (lizzieLet6_5QNode_Int_4_d[2:1])
        2'd0: lizzieLet6_4QNode_Int_onehotd = 4'd1;
        2'd1: lizzieLet6_4QNode_Int_onehotd = 4'd2;
        2'd2: lizzieLet6_4QNode_Int_onehotd = 4'd4;
        2'd3: lizzieLet6_4QNode_Int_onehotd = 4'd8;
        default: lizzieLet6_4QNode_Int_onehotd = 4'd0;
      endcase
    else lizzieLet6_4QNode_Int_onehotd = 4'd0;
  assign _36_d = lizzieLet6_4QNode_Int_onehotd[0];
  assign _35_d = lizzieLet6_4QNode_Int_onehotd[1];
  assign lizzieLet6_5QNode_Int_4QNode_Int_d = lizzieLet6_4QNode_Int_onehotd[2];
  assign _34_d = lizzieLet6_4QNode_Int_onehotd[3];
  assign lizzieLet6_4QNode_Int_r = (| (lizzieLet6_4QNode_Int_onehotd & {_34_r,
                                                                        lizzieLet6_5QNode_Int_4QNode_Int_r,
                                                                        _35_r,
                                                                        _36_r}));
  assign lizzieLet6_5QNode_Int_4_r = lizzieLet6_4QNode_Int_r;
  
  /* fork (Ty MyDTInt_Bool) : (lizzieLet6_5QNode_Int_4QNode_Int,MyDTInt_Bool) > [(lizzieLet6_5QNode_Int_4QNode_Int_1,MyDTInt_Bool),
                                                                            (lizzieLet6_5QNode_Int_4QNode_Int_2,MyDTInt_Bool)] */
  logic [1:0] lizzieLet6_5QNode_Int_4QNode_Int_emitted;
  logic [1:0] lizzieLet6_5QNode_Int_4QNode_Int_done;
  assign lizzieLet6_5QNode_Int_4QNode_Int_1_d = (lizzieLet6_5QNode_Int_4QNode_Int_d[0] && (! lizzieLet6_5QNode_Int_4QNode_Int_emitted[0]));
  assign lizzieLet6_5QNode_Int_4QNode_Int_2_d = (lizzieLet6_5QNode_Int_4QNode_Int_d[0] && (! lizzieLet6_5QNode_Int_4QNode_Int_emitted[1]));
  assign lizzieLet6_5QNode_Int_4QNode_Int_done = (lizzieLet6_5QNode_Int_4QNode_Int_emitted | ({lizzieLet6_5QNode_Int_4QNode_Int_2_d[0],
                                                                                               lizzieLet6_5QNode_Int_4QNode_Int_1_d[0]} & {lizzieLet6_5QNode_Int_4QNode_Int_2_r,
                                                                                                                                           lizzieLet6_5QNode_Int_4QNode_Int_1_r}));
  assign lizzieLet6_5QNode_Int_4QNode_Int_r = (& lizzieLet6_5QNode_Int_4QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_5QNode_Int_4QNode_Int_emitted <= 2'd0;
    else
      lizzieLet6_5QNode_Int_4QNode_Int_emitted <= (lizzieLet6_5QNode_Int_4QNode_Int_r ? 2'd0 :
                                                   lizzieLet6_5QNode_Int_4QNode_Int_done);
  
  /* buf (Ty MyDTInt_Bool) : (lizzieLet6_5QNode_Int_4QNode_Int_2,MyDTInt_Bool) > (lizzieLet6_5QNode_Int_4QNode_Int_2_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t lizzieLet6_5QNode_Int_4QNode_Int_2_bufchan_d;
  logic lizzieLet6_5QNode_Int_4QNode_Int_2_bufchan_r;
  assign lizzieLet6_5QNode_Int_4QNode_Int_2_r = ((! lizzieLet6_5QNode_Int_4QNode_Int_2_bufchan_d[0]) || lizzieLet6_5QNode_Int_4QNode_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_5QNode_Int_4QNode_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet6_5QNode_Int_4QNode_Int_2_r)
        lizzieLet6_5QNode_Int_4QNode_Int_2_bufchan_d <= lizzieLet6_5QNode_Int_4QNode_Int_2_d;
  MyDTInt_Bool_t lizzieLet6_5QNode_Int_4QNode_Int_2_bufchan_buf;
  assign lizzieLet6_5QNode_Int_4QNode_Int_2_bufchan_r = (! lizzieLet6_5QNode_Int_4QNode_Int_2_bufchan_buf[0]);
  assign lizzieLet6_5QNode_Int_4QNode_Int_2_argbuf_d = (lizzieLet6_5QNode_Int_4QNode_Int_2_bufchan_buf[0] ? lizzieLet6_5QNode_Int_4QNode_Int_2_bufchan_buf :
                                                        lizzieLet6_5QNode_Int_4QNode_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_5QNode_Int_4QNode_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet6_5QNode_Int_4QNode_Int_2_argbuf_r && lizzieLet6_5QNode_Int_4QNode_Int_2_bufchan_buf[0]))
        lizzieLet6_5QNode_Int_4QNode_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet6_5QNode_Int_4QNode_Int_2_argbuf_r) && (! lizzieLet6_5QNode_Int_4QNode_Int_2_bufchan_buf[0])))
        lizzieLet6_5QNode_Int_4QNode_Int_2_bufchan_buf <= lizzieLet6_5QNode_Int_4QNode_Int_2_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty MyDTInt_Int_Int) : (lizzieLet6_5QNode_Int_5,QTree_Int) (lizzieLet6_6QNode_Int,MyDTInt_Int_Int) > [(_33,MyDTInt_Int_Int),
                                                                                                            (_32,MyDTInt_Int_Int),
                                                                                                            (lizzieLet6_5QNode_Int_5QNode_Int,MyDTInt_Int_Int),
                                                                                                            (_31,MyDTInt_Int_Int)] */
  logic [3:0] lizzieLet6_6QNode_Int_onehotd;
  always_comb
    if ((lizzieLet6_5QNode_Int_5_d[0] && lizzieLet6_6QNode_Int_d[0]))
      unique case (lizzieLet6_5QNode_Int_5_d[2:1])
        2'd0: lizzieLet6_6QNode_Int_onehotd = 4'd1;
        2'd1: lizzieLet6_6QNode_Int_onehotd = 4'd2;
        2'd2: lizzieLet6_6QNode_Int_onehotd = 4'd4;
        2'd3: lizzieLet6_6QNode_Int_onehotd = 4'd8;
        default: lizzieLet6_6QNode_Int_onehotd = 4'd0;
      endcase
    else lizzieLet6_6QNode_Int_onehotd = 4'd0;
  assign _33_d = lizzieLet6_6QNode_Int_onehotd[0];
  assign _32_d = lizzieLet6_6QNode_Int_onehotd[1];
  assign lizzieLet6_5QNode_Int_5QNode_Int_d = lizzieLet6_6QNode_Int_onehotd[2];
  assign _31_d = lizzieLet6_6QNode_Int_onehotd[3];
  assign lizzieLet6_6QNode_Int_r = (| (lizzieLet6_6QNode_Int_onehotd & {_31_r,
                                                                        lizzieLet6_5QNode_Int_5QNode_Int_r,
                                                                        _32_r,
                                                                        _33_r}));
  assign lizzieLet6_5QNode_Int_5_r = lizzieLet6_6QNode_Int_r;
  
  /* fork (Ty MyDTInt_Int_Int) : (lizzieLet6_5QNode_Int_5QNode_Int,MyDTInt_Int_Int) > [(lizzieLet6_5QNode_Int_5QNode_Int_1,MyDTInt_Int_Int),
                                                                                  (lizzieLet6_5QNode_Int_5QNode_Int_2,MyDTInt_Int_Int)] */
  logic [1:0] lizzieLet6_5QNode_Int_5QNode_Int_emitted;
  logic [1:0] lizzieLet6_5QNode_Int_5QNode_Int_done;
  assign lizzieLet6_5QNode_Int_5QNode_Int_1_d = (lizzieLet6_5QNode_Int_5QNode_Int_d[0] && (! lizzieLet6_5QNode_Int_5QNode_Int_emitted[0]));
  assign lizzieLet6_5QNode_Int_5QNode_Int_2_d = (lizzieLet6_5QNode_Int_5QNode_Int_d[0] && (! lizzieLet6_5QNode_Int_5QNode_Int_emitted[1]));
  assign lizzieLet6_5QNode_Int_5QNode_Int_done = (lizzieLet6_5QNode_Int_5QNode_Int_emitted | ({lizzieLet6_5QNode_Int_5QNode_Int_2_d[0],
                                                                                               lizzieLet6_5QNode_Int_5QNode_Int_1_d[0]} & {lizzieLet6_5QNode_Int_5QNode_Int_2_r,
                                                                                                                                           lizzieLet6_5QNode_Int_5QNode_Int_1_r}));
  assign lizzieLet6_5QNode_Int_5QNode_Int_r = (& lizzieLet6_5QNode_Int_5QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_5QNode_Int_5QNode_Int_emitted <= 2'd0;
    else
      lizzieLet6_5QNode_Int_5QNode_Int_emitted <= (lizzieLet6_5QNode_Int_5QNode_Int_r ? 2'd0 :
                                                   lizzieLet6_5QNode_Int_5QNode_Int_done);
  
  /* buf (Ty MyDTInt_Int_Int) : (lizzieLet6_5QNode_Int_5QNode_Int_2,MyDTInt_Int_Int) > (lizzieLet6_5QNode_Int_5QNode_Int_2_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t lizzieLet6_5QNode_Int_5QNode_Int_2_bufchan_d;
  logic lizzieLet6_5QNode_Int_5QNode_Int_2_bufchan_r;
  assign lizzieLet6_5QNode_Int_5QNode_Int_2_r = ((! lizzieLet6_5QNode_Int_5QNode_Int_2_bufchan_d[0]) || lizzieLet6_5QNode_Int_5QNode_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_5QNode_Int_5QNode_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet6_5QNode_Int_5QNode_Int_2_r)
        lizzieLet6_5QNode_Int_5QNode_Int_2_bufchan_d <= lizzieLet6_5QNode_Int_5QNode_Int_2_d;
  MyDTInt_Int_Int_t lizzieLet6_5QNode_Int_5QNode_Int_2_bufchan_buf;
  assign lizzieLet6_5QNode_Int_5QNode_Int_2_bufchan_r = (! lizzieLet6_5QNode_Int_5QNode_Int_2_bufchan_buf[0]);
  assign lizzieLet6_5QNode_Int_5QNode_Int_2_argbuf_d = (lizzieLet6_5QNode_Int_5QNode_Int_2_bufchan_buf[0] ? lizzieLet6_5QNode_Int_5QNode_Int_2_bufchan_buf :
                                                        lizzieLet6_5QNode_Int_5QNode_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_5QNode_Int_5QNode_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet6_5QNode_Int_5QNode_Int_2_argbuf_r && lizzieLet6_5QNode_Int_5QNode_Int_2_bufchan_buf[0]))
        lizzieLet6_5QNode_Int_5QNode_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet6_5QNode_Int_5QNode_Int_2_argbuf_r) && (! lizzieLet6_5QNode_Int_5QNode_Int_2_bufchan_buf[0])))
        lizzieLet6_5QNode_Int_5QNode_Int_2_bufchan_buf <= lizzieLet6_5QNode_Int_5QNode_Int_2_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_QTree_Int) : (lizzieLet6_5QNode_Int_6,QTree_Int) (lizzieLet6_7QNode_Int,Pointer_QTree_Int) > [(lizzieLet6_5QNode_Int_6QNone_Int,Pointer_QTree_Int),
                                                                                                                (_30,Pointer_QTree_Int),
                                                                                                                (_29,Pointer_QTree_Int),
                                                                                                                (_28,Pointer_QTree_Int)] */
  logic [3:0] lizzieLet6_7QNode_Int_onehotd;
  always_comb
    if ((lizzieLet6_5QNode_Int_6_d[0] && lizzieLet6_7QNode_Int_d[0]))
      unique case (lizzieLet6_5QNode_Int_6_d[2:1])
        2'd0: lizzieLet6_7QNode_Int_onehotd = 4'd1;
        2'd1: lizzieLet6_7QNode_Int_onehotd = 4'd2;
        2'd2: lizzieLet6_7QNode_Int_onehotd = 4'd4;
        2'd3: lizzieLet6_7QNode_Int_onehotd = 4'd8;
        default: lizzieLet6_7QNode_Int_onehotd = 4'd0;
      endcase
    else lizzieLet6_7QNode_Int_onehotd = 4'd0;
  assign lizzieLet6_5QNode_Int_6QNone_Int_d = {lizzieLet6_7QNode_Int_d[16:1],
                                               lizzieLet6_7QNode_Int_onehotd[0]};
  assign _30_d = {lizzieLet6_7QNode_Int_d[16:1],
                  lizzieLet6_7QNode_Int_onehotd[1]};
  assign _29_d = {lizzieLet6_7QNode_Int_d[16:1],
                  lizzieLet6_7QNode_Int_onehotd[2]};
  assign _28_d = {lizzieLet6_7QNode_Int_d[16:1],
                  lizzieLet6_7QNode_Int_onehotd[3]};
  assign lizzieLet6_7QNode_Int_r = (| (lizzieLet6_7QNode_Int_onehotd & {_28_r,
                                                                        _29_r,
                                                                        _30_r,
                                                                        lizzieLet6_5QNode_Int_6QNone_Int_r}));
  assign lizzieLet6_5QNode_Int_6_r = lizzieLet6_7QNode_Int_r;
  
  /* buf (Ty Pointer_QTree_Int) : (lizzieLet6_5QNode_Int_6QNone_Int,Pointer_QTree_Int) > (lizzieLet6_5QNode_Int_6QNone_Int_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t lizzieLet6_5QNode_Int_6QNone_Int_bufchan_d;
  logic lizzieLet6_5QNode_Int_6QNone_Int_bufchan_r;
  assign lizzieLet6_5QNode_Int_6QNone_Int_r = ((! lizzieLet6_5QNode_Int_6QNone_Int_bufchan_d[0]) || lizzieLet6_5QNode_Int_6QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_5QNode_Int_6QNone_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet6_5QNode_Int_6QNone_Int_r)
        lizzieLet6_5QNode_Int_6QNone_Int_bufchan_d <= lizzieLet6_5QNode_Int_6QNone_Int_d;
  Pointer_QTree_Int_t lizzieLet6_5QNode_Int_6QNone_Int_bufchan_buf;
  assign lizzieLet6_5QNode_Int_6QNone_Int_bufchan_r = (! lizzieLet6_5QNode_Int_6QNone_Int_bufchan_buf[0]);
  assign lizzieLet6_5QNode_Int_6QNone_Int_1_argbuf_d = (lizzieLet6_5QNode_Int_6QNone_Int_bufchan_buf[0] ? lizzieLet6_5QNode_Int_6QNone_Int_bufchan_buf :
                                                        lizzieLet6_5QNode_Int_6QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_5QNode_Int_6QNone_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet6_5QNode_Int_6QNone_Int_1_argbuf_r && lizzieLet6_5QNode_Int_6QNone_Int_bufchan_buf[0]))
        lizzieLet6_5QNode_Int_6QNone_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet6_5QNode_Int_6QNone_Int_1_argbuf_r) && (! lizzieLet6_5QNode_Int_6QNone_Int_bufchan_buf[0])))
        lizzieLet6_5QNode_Int_6QNone_Int_bufchan_buf <= lizzieLet6_5QNode_Int_6QNone_Int_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_CTf''''''''''''_f''''''''''''_Int) : (lizzieLet6_5QNode_Int_7,QTree_Int) (lizzieLet6_8QNode_Int,Pointer_CTf''''''''''''_f''''''''''''_Int) > [(lizzieLet6_5QNode_Int_7QNone_Int,Pointer_CTf''''''''''''_f''''''''''''_Int),
                                                                                                                                                                (lizzieLet6_5QNode_Int_7QVal_Int,Pointer_CTf''''''''''''_f''''''''''''_Int),
                                                                                                                                                                (lizzieLet6_5QNode_Int_7QNode_Int,Pointer_CTf''''''''''''_f''''''''''''_Int),
                                                                                                                                                                (lizzieLet6_5QNode_Int_7QError_Int,Pointer_CTf''''''''''''_f''''''''''''_Int)] */
  logic [3:0] lizzieLet6_8QNode_Int_onehotd;
  always_comb
    if ((lizzieLet6_5QNode_Int_7_d[0] && lizzieLet6_8QNode_Int_d[0]))
      unique case (lizzieLet6_5QNode_Int_7_d[2:1])
        2'd0: lizzieLet6_8QNode_Int_onehotd = 4'd1;
        2'd1: lizzieLet6_8QNode_Int_onehotd = 4'd2;
        2'd2: lizzieLet6_8QNode_Int_onehotd = 4'd4;
        2'd3: lizzieLet6_8QNode_Int_onehotd = 4'd8;
        default: lizzieLet6_8QNode_Int_onehotd = 4'd0;
      endcase
    else lizzieLet6_8QNode_Int_onehotd = 4'd0;
  assign lizzieLet6_5QNode_Int_7QNone_Int_d = {lizzieLet6_8QNode_Int_d[16:1],
                                               lizzieLet6_8QNode_Int_onehotd[0]};
  assign lizzieLet6_5QNode_Int_7QVal_Int_d = {lizzieLet6_8QNode_Int_d[16:1],
                                              lizzieLet6_8QNode_Int_onehotd[1]};
  assign lizzieLet6_5QNode_Int_7QNode_Int_d = {lizzieLet6_8QNode_Int_d[16:1],
                                               lizzieLet6_8QNode_Int_onehotd[2]};
  assign lizzieLet6_5QNode_Int_7QError_Int_d = {lizzieLet6_8QNode_Int_d[16:1],
                                                lizzieLet6_8QNode_Int_onehotd[3]};
  assign lizzieLet6_8QNode_Int_r = (| (lizzieLet6_8QNode_Int_onehotd & {lizzieLet6_5QNode_Int_7QError_Int_r,
                                                                        lizzieLet6_5QNode_Int_7QNode_Int_r,
                                                                        lizzieLet6_5QNode_Int_7QVal_Int_r,
                                                                        lizzieLet6_5QNode_Int_7QNone_Int_r}));
  assign lizzieLet6_5QNode_Int_7_r = lizzieLet6_8QNode_Int_r;
  
  /* buf (Ty Pointer_CTf''''''''''''_f''''''''''''_Int) : (lizzieLet6_5QNode_Int_7QError_Int,Pointer_CTf''''''''''''_f''''''''''''_Int) > (lizzieLet6_5QNode_Int_7QError_Int_1_argbuf,Pointer_CTf''''''''''''_f''''''''''''_Int) */
  \Pointer_CTf''''''''''''_f''''''''''''_Int_t  lizzieLet6_5QNode_Int_7QError_Int_bufchan_d;
  logic lizzieLet6_5QNode_Int_7QError_Int_bufchan_r;
  assign lizzieLet6_5QNode_Int_7QError_Int_r = ((! lizzieLet6_5QNode_Int_7QError_Int_bufchan_d[0]) || lizzieLet6_5QNode_Int_7QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_5QNode_Int_7QError_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet6_5QNode_Int_7QError_Int_r)
        lizzieLet6_5QNode_Int_7QError_Int_bufchan_d <= lizzieLet6_5QNode_Int_7QError_Int_d;
  \Pointer_CTf''''''''''''_f''''''''''''_Int_t  lizzieLet6_5QNode_Int_7QError_Int_bufchan_buf;
  assign lizzieLet6_5QNode_Int_7QError_Int_bufchan_r = (! lizzieLet6_5QNode_Int_7QError_Int_bufchan_buf[0]);
  assign lizzieLet6_5QNode_Int_7QError_Int_1_argbuf_d = (lizzieLet6_5QNode_Int_7QError_Int_bufchan_buf[0] ? lizzieLet6_5QNode_Int_7QError_Int_bufchan_buf :
                                                         lizzieLet6_5QNode_Int_7QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_5QNode_Int_7QError_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet6_5QNode_Int_7QError_Int_1_argbuf_r && lizzieLet6_5QNode_Int_7QError_Int_bufchan_buf[0]))
        lizzieLet6_5QNode_Int_7QError_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet6_5QNode_Int_7QError_Int_1_argbuf_r) && (! lizzieLet6_5QNode_Int_7QError_Int_bufchan_buf[0])))
        lizzieLet6_5QNode_Int_7QError_Int_bufchan_buf <= lizzieLet6_5QNode_Int_7QError_Int_bufchan_d;
  
  /* dcon (Ty CTf''''''''''''_f''''''''''''_Int,
      Dcon Lcall_f''''''''''''_f''''''''''''_Int3) : [(lizzieLet6_5QNode_Int_7QNode_Int,Pointer_CTf''''''''''''_f''''''''''''_Int),
                                                      (lizzieLet6_5QNode_Int_8QNode_Int,Pointer_QTree_Int),
                                                      (t1afy_destruct,Pointer_QTree_Int),
                                                      (lizzieLet6_5QNode_Int_4QNode_Int_1,MyDTInt_Bool),
                                                      (lizzieLet6_5QNode_Int_5QNode_Int_1,MyDTInt_Int_Int),
                                                      (lizzieLet6_5QNode_Int_9QNode_Int,Pointer_QTree_Int),
                                                      (t2afz_destruct,Pointer_QTree_Int),
                                                      (lizzieLet6_5QNode_Int_10QNode_Int,Pointer_QTree_Int),
                                                      (t3afA_destruct,Pointer_QTree_Int)] > (lizzieLet6_5QNode_Int_7QNode_Int_1lizzieLet6_5QNode_Int_8QNode_Int_1t1afy_1lizzieLet6_5QNode_Int_4QNode_Int_1lizzieLet6_5QNode_Int_5QNode_Int_1lizzieLet6_5QNode_Int_9QNode_Int_1t2afz_1lizzieLet6_5QNode_Int_10QNode_Int_1t3afA_1Lcall_f''''''''''''_f''''''''''''_Int3,CTf''''''''''''_f''''''''''''_Int) */
  assign \lizzieLet6_5QNode_Int_7QNode_Int_1lizzieLet6_5QNode_Int_8QNode_Int_1t1afy_1lizzieLet6_5QNode_Int_4QNode_Int_1lizzieLet6_5QNode_Int_5QNode_Int_1lizzieLet6_5QNode_Int_9QNode_Int_1t2afz_1lizzieLet6_5QNode_Int_10QNode_Int_1t3afA_1Lcall_f''''''''''''_f''''''''''''_Int3_d  = \Lcall_f''''''''''''_f''''''''''''_Int3_dc ((& {lizzieLet6_5QNode_Int_7QNode_Int_d[0],
                                                                                                                                                                                                                                                                                                                                        lizzieLet6_5QNode_Int_8QNode_Int_d[0],
                                                                                                                                                                                                                                                                                                                                        t1afy_destruct_d[0],
                                                                                                                                                                                                                                                                                                                                        lizzieLet6_5QNode_Int_4QNode_Int_1_d[0],
                                                                                                                                                                                                                                                                                                                                        lizzieLet6_5QNode_Int_5QNode_Int_1_d[0],
                                                                                                                                                                                                                                                                                                                                        lizzieLet6_5QNode_Int_9QNode_Int_d[0],
                                                                                                                                                                                                                                                                                                                                        t2afz_destruct_d[0],
                                                                                                                                                                                                                                                                                                                                        lizzieLet6_5QNode_Int_10QNode_Int_d[0],
                                                                                                                                                                                                                                                                                                                                        t3afA_destruct_d[0]}), lizzieLet6_5QNode_Int_7QNode_Int_d, lizzieLet6_5QNode_Int_8QNode_Int_d, t1afy_destruct_d, lizzieLet6_5QNode_Int_4QNode_Int_1_d, lizzieLet6_5QNode_Int_5QNode_Int_1_d, lizzieLet6_5QNode_Int_9QNode_Int_d, t2afz_destruct_d, lizzieLet6_5QNode_Int_10QNode_Int_d, t3afA_destruct_d);
  assign {lizzieLet6_5QNode_Int_7QNode_Int_r,
          lizzieLet6_5QNode_Int_8QNode_Int_r,
          t1afy_destruct_r,
          lizzieLet6_5QNode_Int_4QNode_Int_1_r,
          lizzieLet6_5QNode_Int_5QNode_Int_1_r,
          lizzieLet6_5QNode_Int_9QNode_Int_r,
          t2afz_destruct_r,
          lizzieLet6_5QNode_Int_10QNode_Int_r,
          t3afA_destruct_r} = {9 {(\lizzieLet6_5QNode_Int_7QNode_Int_1lizzieLet6_5QNode_Int_8QNode_Int_1t1afy_1lizzieLet6_5QNode_Int_4QNode_Int_1lizzieLet6_5QNode_Int_5QNode_Int_1lizzieLet6_5QNode_Int_9QNode_Int_1t2afz_1lizzieLet6_5QNode_Int_10QNode_Int_1t3afA_1Lcall_f''''''''''''_f''''''''''''_Int3_r  && \lizzieLet6_5QNode_Int_7QNode_Int_1lizzieLet6_5QNode_Int_8QNode_Int_1t1afy_1lizzieLet6_5QNode_Int_4QNode_Int_1lizzieLet6_5QNode_Int_5QNode_Int_1lizzieLet6_5QNode_Int_9QNode_Int_1t2afz_1lizzieLet6_5QNode_Int_10QNode_Int_1t3afA_1Lcall_f''''''''''''_f''''''''''''_Int3_d [0])}};
  
  /* buf (Ty CTf''''''''''''_f''''''''''''_Int) : (lizzieLet6_5QNode_Int_7QNode_Int_1lizzieLet6_5QNode_Int_8QNode_Int_1t1afy_1lizzieLet6_5QNode_Int_4QNode_Int_1lizzieLet6_5QNode_Int_5QNode_Int_1lizzieLet6_5QNode_Int_9QNode_Int_1t2afz_1lizzieLet6_5QNode_Int_10QNode_Int_1t3afA_1Lcall_f''''''''''''_f''''''''''''_Int3,CTf''''''''''''_f''''''''''''_Int) > (lizzieLet14_1_argbuf,CTf''''''''''''_f''''''''''''_Int) */
  \CTf''''''''''''_f''''''''''''_Int_t  \lizzieLet6_5QNode_Int_7QNode_Int_1lizzieLet6_5QNode_Int_8QNode_Int_1t1afy_1lizzieLet6_5QNode_Int_4QNode_Int_1lizzieLet6_5QNode_Int_5QNode_Int_1lizzieLet6_5QNode_Int_9QNode_Int_1t2afz_1lizzieLet6_5QNode_Int_10QNode_Int_1t3afA_1Lcall_f''''''''''''_f''''''''''''_Int3_bufchan_d ;
  logic \lizzieLet6_5QNode_Int_7QNode_Int_1lizzieLet6_5QNode_Int_8QNode_Int_1t1afy_1lizzieLet6_5QNode_Int_4QNode_Int_1lizzieLet6_5QNode_Int_5QNode_Int_1lizzieLet6_5QNode_Int_9QNode_Int_1t2afz_1lizzieLet6_5QNode_Int_10QNode_Int_1t3afA_1Lcall_f''''''''''''_f''''''''''''_Int3_bufchan_r ;
  assign \lizzieLet6_5QNode_Int_7QNode_Int_1lizzieLet6_5QNode_Int_8QNode_Int_1t1afy_1lizzieLet6_5QNode_Int_4QNode_Int_1lizzieLet6_5QNode_Int_5QNode_Int_1lizzieLet6_5QNode_Int_9QNode_Int_1t2afz_1lizzieLet6_5QNode_Int_10QNode_Int_1t3afA_1Lcall_f''''''''''''_f''''''''''''_Int3_r  = ((! \lizzieLet6_5QNode_Int_7QNode_Int_1lizzieLet6_5QNode_Int_8QNode_Int_1t1afy_1lizzieLet6_5QNode_Int_4QNode_Int_1lizzieLet6_5QNode_Int_5QNode_Int_1lizzieLet6_5QNode_Int_9QNode_Int_1t2afz_1lizzieLet6_5QNode_Int_10QNode_Int_1t3afA_1Lcall_f''''''''''''_f''''''''''''_Int3_bufchan_d [0]) || \lizzieLet6_5QNode_Int_7QNode_Int_1lizzieLet6_5QNode_Int_8QNode_Int_1t1afy_1lizzieLet6_5QNode_Int_4QNode_Int_1lizzieLet6_5QNode_Int_5QNode_Int_1lizzieLet6_5QNode_Int_9QNode_Int_1t2afz_1lizzieLet6_5QNode_Int_10QNode_Int_1t3afA_1Lcall_f''''''''''''_f''''''''''''_Int3_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet6_5QNode_Int_7QNode_Int_1lizzieLet6_5QNode_Int_8QNode_Int_1t1afy_1lizzieLet6_5QNode_Int_4QNode_Int_1lizzieLet6_5QNode_Int_5QNode_Int_1lizzieLet6_5QNode_Int_9QNode_Int_1t2afz_1lizzieLet6_5QNode_Int_10QNode_Int_1t3afA_1Lcall_f''''''''''''_f''''''''''''_Int3_bufchan_d  <= {115'd0,
                                                                                                                                                                                                                                                                                               1'd0};
    else
      if (\lizzieLet6_5QNode_Int_7QNode_Int_1lizzieLet6_5QNode_Int_8QNode_Int_1t1afy_1lizzieLet6_5QNode_Int_4QNode_Int_1lizzieLet6_5QNode_Int_5QNode_Int_1lizzieLet6_5QNode_Int_9QNode_Int_1t2afz_1lizzieLet6_5QNode_Int_10QNode_Int_1t3afA_1Lcall_f''''''''''''_f''''''''''''_Int3_r )
        \lizzieLet6_5QNode_Int_7QNode_Int_1lizzieLet6_5QNode_Int_8QNode_Int_1t1afy_1lizzieLet6_5QNode_Int_4QNode_Int_1lizzieLet6_5QNode_Int_5QNode_Int_1lizzieLet6_5QNode_Int_9QNode_Int_1t2afz_1lizzieLet6_5QNode_Int_10QNode_Int_1t3afA_1Lcall_f''''''''''''_f''''''''''''_Int3_bufchan_d  <= \lizzieLet6_5QNode_Int_7QNode_Int_1lizzieLet6_5QNode_Int_8QNode_Int_1t1afy_1lizzieLet6_5QNode_Int_4QNode_Int_1lizzieLet6_5QNode_Int_5QNode_Int_1lizzieLet6_5QNode_Int_9QNode_Int_1t2afz_1lizzieLet6_5QNode_Int_10QNode_Int_1t3afA_1Lcall_f''''''''''''_f''''''''''''_Int3_d ;
  \CTf''''''''''''_f''''''''''''_Int_t  \lizzieLet6_5QNode_Int_7QNode_Int_1lizzieLet6_5QNode_Int_8QNode_Int_1t1afy_1lizzieLet6_5QNode_Int_4QNode_Int_1lizzieLet6_5QNode_Int_5QNode_Int_1lizzieLet6_5QNode_Int_9QNode_Int_1t2afz_1lizzieLet6_5QNode_Int_10QNode_Int_1t3afA_1Lcall_f''''''''''''_f''''''''''''_Int3_bufchan_buf ;
  assign \lizzieLet6_5QNode_Int_7QNode_Int_1lizzieLet6_5QNode_Int_8QNode_Int_1t1afy_1lizzieLet6_5QNode_Int_4QNode_Int_1lizzieLet6_5QNode_Int_5QNode_Int_1lizzieLet6_5QNode_Int_9QNode_Int_1t2afz_1lizzieLet6_5QNode_Int_10QNode_Int_1t3afA_1Lcall_f''''''''''''_f''''''''''''_Int3_bufchan_r  = (! \lizzieLet6_5QNode_Int_7QNode_Int_1lizzieLet6_5QNode_Int_8QNode_Int_1t1afy_1lizzieLet6_5QNode_Int_4QNode_Int_1lizzieLet6_5QNode_Int_5QNode_Int_1lizzieLet6_5QNode_Int_9QNode_Int_1t2afz_1lizzieLet6_5QNode_Int_10QNode_Int_1t3afA_1Lcall_f''''''''''''_f''''''''''''_Int3_bufchan_buf [0]);
  assign lizzieLet14_1_argbuf_d = (\lizzieLet6_5QNode_Int_7QNode_Int_1lizzieLet6_5QNode_Int_8QNode_Int_1t1afy_1lizzieLet6_5QNode_Int_4QNode_Int_1lizzieLet6_5QNode_Int_5QNode_Int_1lizzieLet6_5QNode_Int_9QNode_Int_1t2afz_1lizzieLet6_5QNode_Int_10QNode_Int_1t3afA_1Lcall_f''''''''''''_f''''''''''''_Int3_bufchan_buf [0] ? \lizzieLet6_5QNode_Int_7QNode_Int_1lizzieLet6_5QNode_Int_8QNode_Int_1t1afy_1lizzieLet6_5QNode_Int_4QNode_Int_1lizzieLet6_5QNode_Int_5QNode_Int_1lizzieLet6_5QNode_Int_9QNode_Int_1t2afz_1lizzieLet6_5QNode_Int_10QNode_Int_1t3afA_1Lcall_f''''''''''''_f''''''''''''_Int3_bufchan_buf  :
                                   \lizzieLet6_5QNode_Int_7QNode_Int_1lizzieLet6_5QNode_Int_8QNode_Int_1t1afy_1lizzieLet6_5QNode_Int_4QNode_Int_1lizzieLet6_5QNode_Int_5QNode_Int_1lizzieLet6_5QNode_Int_9QNode_Int_1t2afz_1lizzieLet6_5QNode_Int_10QNode_Int_1t3afA_1Lcall_f''''''''''''_f''''''''''''_Int3_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet6_5QNode_Int_7QNode_Int_1lizzieLet6_5QNode_Int_8QNode_Int_1t1afy_1lizzieLet6_5QNode_Int_4QNode_Int_1lizzieLet6_5QNode_Int_5QNode_Int_1lizzieLet6_5QNode_Int_9QNode_Int_1t2afz_1lizzieLet6_5QNode_Int_10QNode_Int_1t3afA_1Lcall_f''''''''''''_f''''''''''''_Int3_bufchan_buf  <= {115'd0,
                                                                                                                                                                                                                                                                                                 1'd0};
    else
      if ((lizzieLet14_1_argbuf_r && \lizzieLet6_5QNode_Int_7QNode_Int_1lizzieLet6_5QNode_Int_8QNode_Int_1t1afy_1lizzieLet6_5QNode_Int_4QNode_Int_1lizzieLet6_5QNode_Int_5QNode_Int_1lizzieLet6_5QNode_Int_9QNode_Int_1t2afz_1lizzieLet6_5QNode_Int_10QNode_Int_1t3afA_1Lcall_f''''''''''''_f''''''''''''_Int3_bufchan_buf [0]))
        \lizzieLet6_5QNode_Int_7QNode_Int_1lizzieLet6_5QNode_Int_8QNode_Int_1t1afy_1lizzieLet6_5QNode_Int_4QNode_Int_1lizzieLet6_5QNode_Int_5QNode_Int_1lizzieLet6_5QNode_Int_9QNode_Int_1t2afz_1lizzieLet6_5QNode_Int_10QNode_Int_1t3afA_1Lcall_f''''''''''''_f''''''''''''_Int3_bufchan_buf  <= {115'd0,
                                                                                                                                                                                                                                                                                                   1'd0};
      else if (((! lizzieLet14_1_argbuf_r) && (! \lizzieLet6_5QNode_Int_7QNode_Int_1lizzieLet6_5QNode_Int_8QNode_Int_1t1afy_1lizzieLet6_5QNode_Int_4QNode_Int_1lizzieLet6_5QNode_Int_5QNode_Int_1lizzieLet6_5QNode_Int_9QNode_Int_1t2afz_1lizzieLet6_5QNode_Int_10QNode_Int_1t3afA_1Lcall_f''''''''''''_f''''''''''''_Int3_bufchan_buf [0])))
        \lizzieLet6_5QNode_Int_7QNode_Int_1lizzieLet6_5QNode_Int_8QNode_Int_1t1afy_1lizzieLet6_5QNode_Int_4QNode_Int_1lizzieLet6_5QNode_Int_5QNode_Int_1lizzieLet6_5QNode_Int_9QNode_Int_1t2afz_1lizzieLet6_5QNode_Int_10QNode_Int_1t3afA_1Lcall_f''''''''''''_f''''''''''''_Int3_bufchan_buf  <= \lizzieLet6_5QNode_Int_7QNode_Int_1lizzieLet6_5QNode_Int_8QNode_Int_1t1afy_1lizzieLet6_5QNode_Int_4QNode_Int_1lizzieLet6_5QNode_Int_5QNode_Int_1lizzieLet6_5QNode_Int_9QNode_Int_1t2afz_1lizzieLet6_5QNode_Int_10QNode_Int_1t3afA_1Lcall_f''''''''''''_f''''''''''''_Int3_bufchan_d ;
  
  /* buf (Ty Pointer_CTf''''''''''''_f''''''''''''_Int) : (lizzieLet6_5QNode_Int_7QNone_Int,Pointer_CTf''''''''''''_f''''''''''''_Int) > (lizzieLet6_5QNode_Int_7QNone_Int_1_argbuf,Pointer_CTf''''''''''''_f''''''''''''_Int) */
  \Pointer_CTf''''''''''''_f''''''''''''_Int_t  lizzieLet6_5QNode_Int_7QNone_Int_bufchan_d;
  logic lizzieLet6_5QNode_Int_7QNone_Int_bufchan_r;
  assign lizzieLet6_5QNode_Int_7QNone_Int_r = ((! lizzieLet6_5QNode_Int_7QNone_Int_bufchan_d[0]) || lizzieLet6_5QNode_Int_7QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_5QNode_Int_7QNone_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet6_5QNode_Int_7QNone_Int_r)
        lizzieLet6_5QNode_Int_7QNone_Int_bufchan_d <= lizzieLet6_5QNode_Int_7QNone_Int_d;
  \Pointer_CTf''''''''''''_f''''''''''''_Int_t  lizzieLet6_5QNode_Int_7QNone_Int_bufchan_buf;
  assign lizzieLet6_5QNode_Int_7QNone_Int_bufchan_r = (! lizzieLet6_5QNode_Int_7QNone_Int_bufchan_buf[0]);
  assign lizzieLet6_5QNode_Int_7QNone_Int_1_argbuf_d = (lizzieLet6_5QNode_Int_7QNone_Int_bufchan_buf[0] ? lizzieLet6_5QNode_Int_7QNone_Int_bufchan_buf :
                                                        lizzieLet6_5QNode_Int_7QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_5QNode_Int_7QNone_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet6_5QNode_Int_7QNone_Int_1_argbuf_r && lizzieLet6_5QNode_Int_7QNone_Int_bufchan_buf[0]))
        lizzieLet6_5QNode_Int_7QNone_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet6_5QNode_Int_7QNone_Int_1_argbuf_r) && (! lizzieLet6_5QNode_Int_7QNone_Int_bufchan_buf[0])))
        lizzieLet6_5QNode_Int_7QNone_Int_bufchan_buf <= lizzieLet6_5QNode_Int_7QNone_Int_bufchan_d;
  
  /* buf (Ty Pointer_CTf''''''''''''_f''''''''''''_Int) : (lizzieLet6_5QNode_Int_7QVal_Int,Pointer_CTf''''''''''''_f''''''''''''_Int) > (lizzieLet6_5QNode_Int_7QVal_Int_1_argbuf,Pointer_CTf''''''''''''_f''''''''''''_Int) */
  \Pointer_CTf''''''''''''_f''''''''''''_Int_t  lizzieLet6_5QNode_Int_7QVal_Int_bufchan_d;
  logic lizzieLet6_5QNode_Int_7QVal_Int_bufchan_r;
  assign lizzieLet6_5QNode_Int_7QVal_Int_r = ((! lizzieLet6_5QNode_Int_7QVal_Int_bufchan_d[0]) || lizzieLet6_5QNode_Int_7QVal_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_5QNode_Int_7QVal_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet6_5QNode_Int_7QVal_Int_r)
        lizzieLet6_5QNode_Int_7QVal_Int_bufchan_d <= lizzieLet6_5QNode_Int_7QVal_Int_d;
  \Pointer_CTf''''''''''''_f''''''''''''_Int_t  lizzieLet6_5QNode_Int_7QVal_Int_bufchan_buf;
  assign lizzieLet6_5QNode_Int_7QVal_Int_bufchan_r = (! lizzieLet6_5QNode_Int_7QVal_Int_bufchan_buf[0]);
  assign lizzieLet6_5QNode_Int_7QVal_Int_1_argbuf_d = (lizzieLet6_5QNode_Int_7QVal_Int_bufchan_buf[0] ? lizzieLet6_5QNode_Int_7QVal_Int_bufchan_buf :
                                                       lizzieLet6_5QNode_Int_7QVal_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_5QNode_Int_7QVal_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet6_5QNode_Int_7QVal_Int_1_argbuf_r && lizzieLet6_5QNode_Int_7QVal_Int_bufchan_buf[0]))
        lizzieLet6_5QNode_Int_7QVal_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet6_5QNode_Int_7QVal_Int_1_argbuf_r) && (! lizzieLet6_5QNode_Int_7QVal_Int_bufchan_buf[0])))
        lizzieLet6_5QNode_Int_7QVal_Int_bufchan_buf <= lizzieLet6_5QNode_Int_7QVal_Int_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_QTree_Int) : (lizzieLet6_5QNode_Int_8,QTree_Int) (q1aft_destruct,Pointer_QTree_Int) > [(_27,Pointer_QTree_Int),
                                                                                                         (_26,Pointer_QTree_Int),
                                                                                                         (lizzieLet6_5QNode_Int_8QNode_Int,Pointer_QTree_Int),
                                                                                                         (_25,Pointer_QTree_Int)] */
  logic [3:0] q1aft_destruct_onehotd;
  always_comb
    if ((lizzieLet6_5QNode_Int_8_d[0] && q1aft_destruct_d[0]))
      unique case (lizzieLet6_5QNode_Int_8_d[2:1])
        2'd0: q1aft_destruct_onehotd = 4'd1;
        2'd1: q1aft_destruct_onehotd = 4'd2;
        2'd2: q1aft_destruct_onehotd = 4'd4;
        2'd3: q1aft_destruct_onehotd = 4'd8;
        default: q1aft_destruct_onehotd = 4'd0;
      endcase
    else q1aft_destruct_onehotd = 4'd0;
  assign _27_d = {q1aft_destruct_d[16:1], q1aft_destruct_onehotd[0]};
  assign _26_d = {q1aft_destruct_d[16:1], q1aft_destruct_onehotd[1]};
  assign lizzieLet6_5QNode_Int_8QNode_Int_d = {q1aft_destruct_d[16:1],
                                               q1aft_destruct_onehotd[2]};
  assign _25_d = {q1aft_destruct_d[16:1], q1aft_destruct_onehotd[3]};
  assign q1aft_destruct_r = (| (q1aft_destruct_onehotd & {_25_r,
                                                          lizzieLet6_5QNode_Int_8QNode_Int_r,
                                                          _26_r,
                                                          _27_r}));
  assign lizzieLet6_5QNode_Int_8_r = q1aft_destruct_r;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_QTree_Int) : (lizzieLet6_5QNode_Int_9,QTree_Int) (q2afu_destruct,Pointer_QTree_Int) > [(_24,Pointer_QTree_Int),
                                                                                                         (_23,Pointer_QTree_Int),
                                                                                                         (lizzieLet6_5QNode_Int_9QNode_Int,Pointer_QTree_Int),
                                                                                                         (_22,Pointer_QTree_Int)] */
  logic [3:0] q2afu_destruct_onehotd;
  always_comb
    if ((lizzieLet6_5QNode_Int_9_d[0] && q2afu_destruct_d[0]))
      unique case (lizzieLet6_5QNode_Int_9_d[2:1])
        2'd0: q2afu_destruct_onehotd = 4'd1;
        2'd1: q2afu_destruct_onehotd = 4'd2;
        2'd2: q2afu_destruct_onehotd = 4'd4;
        2'd3: q2afu_destruct_onehotd = 4'd8;
        default: q2afu_destruct_onehotd = 4'd0;
      endcase
    else q2afu_destruct_onehotd = 4'd0;
  assign _24_d = {q2afu_destruct_d[16:1], q2afu_destruct_onehotd[0]};
  assign _23_d = {q2afu_destruct_d[16:1], q2afu_destruct_onehotd[1]};
  assign lizzieLet6_5QNode_Int_9QNode_Int_d = {q2afu_destruct_d[16:1],
                                               q2afu_destruct_onehotd[2]};
  assign _22_d = {q2afu_destruct_d[16:1], q2afu_destruct_onehotd[3]};
  assign q2afu_destruct_r = (| (q2afu_destruct_onehotd & {_22_r,
                                                          lizzieLet6_5QNode_Int_9QNode_Int_r,
                                                          _23_r,
                                                          _24_r}));
  assign lizzieLet6_5QNode_Int_9_r = q2afu_destruct_r;
  
  /* fork (Ty QTree_Int) : (lizzieLet6_5QVal_Int,QTree_Int) > [(lizzieLet6_5QVal_Int_1,QTree_Int),
                                                          (lizzieLet6_5QVal_Int_2,QTree_Int),
                                                          (lizzieLet6_5QVal_Int_3,QTree_Int),
                                                          (lizzieLet6_5QVal_Int_4,QTree_Int),
                                                          (lizzieLet6_5QVal_Int_5,QTree_Int),
                                                          (lizzieLet6_5QVal_Int_6,QTree_Int),
                                                          (lizzieLet6_5QVal_Int_7,QTree_Int),
                                                          (lizzieLet6_5QVal_Int_8,QTree_Int)] */
  logic [7:0] lizzieLet6_5QVal_Int_emitted;
  logic [7:0] lizzieLet6_5QVal_Int_done;
  assign lizzieLet6_5QVal_Int_1_d = {lizzieLet6_5QVal_Int_d[66:1],
                                     (lizzieLet6_5QVal_Int_d[0] && (! lizzieLet6_5QVal_Int_emitted[0]))};
  assign lizzieLet6_5QVal_Int_2_d = {lizzieLet6_5QVal_Int_d[66:1],
                                     (lizzieLet6_5QVal_Int_d[0] && (! lizzieLet6_5QVal_Int_emitted[1]))};
  assign lizzieLet6_5QVal_Int_3_d = {lizzieLet6_5QVal_Int_d[66:1],
                                     (lizzieLet6_5QVal_Int_d[0] && (! lizzieLet6_5QVal_Int_emitted[2]))};
  assign lizzieLet6_5QVal_Int_4_d = {lizzieLet6_5QVal_Int_d[66:1],
                                     (lizzieLet6_5QVal_Int_d[0] && (! lizzieLet6_5QVal_Int_emitted[3]))};
  assign lizzieLet6_5QVal_Int_5_d = {lizzieLet6_5QVal_Int_d[66:1],
                                     (lizzieLet6_5QVal_Int_d[0] && (! lizzieLet6_5QVal_Int_emitted[4]))};
  assign lizzieLet6_5QVal_Int_6_d = {lizzieLet6_5QVal_Int_d[66:1],
                                     (lizzieLet6_5QVal_Int_d[0] && (! lizzieLet6_5QVal_Int_emitted[5]))};
  assign lizzieLet6_5QVal_Int_7_d = {lizzieLet6_5QVal_Int_d[66:1],
                                     (lizzieLet6_5QVal_Int_d[0] && (! lizzieLet6_5QVal_Int_emitted[6]))};
  assign lizzieLet6_5QVal_Int_8_d = {lizzieLet6_5QVal_Int_d[66:1],
                                     (lizzieLet6_5QVal_Int_d[0] && (! lizzieLet6_5QVal_Int_emitted[7]))};
  assign lizzieLet6_5QVal_Int_done = (lizzieLet6_5QVal_Int_emitted | ({lizzieLet6_5QVal_Int_8_d[0],
                                                                       lizzieLet6_5QVal_Int_7_d[0],
                                                                       lizzieLet6_5QVal_Int_6_d[0],
                                                                       lizzieLet6_5QVal_Int_5_d[0],
                                                                       lizzieLet6_5QVal_Int_4_d[0],
                                                                       lizzieLet6_5QVal_Int_3_d[0],
                                                                       lizzieLet6_5QVal_Int_2_d[0],
                                                                       lizzieLet6_5QVal_Int_1_d[0]} & {lizzieLet6_5QVal_Int_8_r,
                                                                                                       lizzieLet6_5QVal_Int_7_r,
                                                                                                       lizzieLet6_5QVal_Int_6_r,
                                                                                                       lizzieLet6_5QVal_Int_5_r,
                                                                                                       lizzieLet6_5QVal_Int_4_r,
                                                                                                       lizzieLet6_5QVal_Int_3_r,
                                                                                                       lizzieLet6_5QVal_Int_2_r,
                                                                                                       lizzieLet6_5QVal_Int_1_r}));
  assign lizzieLet6_5QVal_Int_r = (& lizzieLet6_5QVal_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_5QVal_Int_emitted <= 8'd0;
    else
      lizzieLet6_5QVal_Int_emitted <= (lizzieLet6_5QVal_Int_r ? 8'd0 :
                                       lizzieLet6_5QVal_Int_done);
  
  /* destruct (Ty QTree_Int,
          Dcon QVal_Int) : (lizzieLet6_5QVal_Int_1QVal_Int,QTree_Int) > [(vafo_destruct,Int)] */
  assign vafo_destruct_d = {lizzieLet6_5QVal_Int_1QVal_Int_d[34:3],
                            lizzieLet6_5QVal_Int_1QVal_Int_d[0]};
  assign lizzieLet6_5QVal_Int_1QVal_Int_r = vafo_destruct_r;
  
  /* demux (Ty QTree_Int,
       Ty QTree_Int) : (lizzieLet6_5QVal_Int_2,QTree_Int) (lizzieLet6_5QVal_Int_1,QTree_Int) > [(_21,QTree_Int),
                                                                                                (lizzieLet6_5QVal_Int_1QVal_Int,QTree_Int),
                                                                                                (_20,QTree_Int),
                                                                                                (_19,QTree_Int)] */
  logic [3:0] lizzieLet6_5QVal_Int_1_onehotd;
  always_comb
    if ((lizzieLet6_5QVal_Int_2_d[0] && lizzieLet6_5QVal_Int_1_d[0]))
      unique case (lizzieLet6_5QVal_Int_2_d[2:1])
        2'd0: lizzieLet6_5QVal_Int_1_onehotd = 4'd1;
        2'd1: lizzieLet6_5QVal_Int_1_onehotd = 4'd2;
        2'd2: lizzieLet6_5QVal_Int_1_onehotd = 4'd4;
        2'd3: lizzieLet6_5QVal_Int_1_onehotd = 4'd8;
        default: lizzieLet6_5QVal_Int_1_onehotd = 4'd0;
      endcase
    else lizzieLet6_5QVal_Int_1_onehotd = 4'd0;
  assign _21_d = {lizzieLet6_5QVal_Int_1_d[66:1],
                  lizzieLet6_5QVal_Int_1_onehotd[0]};
  assign lizzieLet6_5QVal_Int_1QVal_Int_d = {lizzieLet6_5QVal_Int_1_d[66:1],
                                             lizzieLet6_5QVal_Int_1_onehotd[1]};
  assign _20_d = {lizzieLet6_5QVal_Int_1_d[66:1],
                  lizzieLet6_5QVal_Int_1_onehotd[2]};
  assign _19_d = {lizzieLet6_5QVal_Int_1_d[66:1],
                  lizzieLet6_5QVal_Int_1_onehotd[3]};
  assign lizzieLet6_5QVal_Int_1_r = (| (lizzieLet6_5QVal_Int_1_onehotd & {_19_r,
                                                                          _20_r,
                                                                          lizzieLet6_5QVal_Int_1QVal_Int_r,
                                                                          _21_r}));
  assign lizzieLet6_5QVal_Int_2_r = lizzieLet6_5QVal_Int_1_r;
  
  /* demux (Ty QTree_Int,
       Ty Go) : (lizzieLet6_5QVal_Int_3,QTree_Int) (lizzieLet6_3QVal_Int,Go) > [(lizzieLet6_5QVal_Int_3QNone_Int,Go),
                                                                                (lizzieLet6_5QVal_Int_3QVal_Int,Go),
                                                                                (lizzieLet6_5QVal_Int_3QNode_Int,Go),
                                                                                (lizzieLet6_5QVal_Int_3QError_Int,Go)] */
  logic [3:0] lizzieLet6_3QVal_Int_onehotd;
  always_comb
    if ((lizzieLet6_5QVal_Int_3_d[0] && lizzieLet6_3QVal_Int_d[0]))
      unique case (lizzieLet6_5QVal_Int_3_d[2:1])
        2'd0: lizzieLet6_3QVal_Int_onehotd = 4'd1;
        2'd1: lizzieLet6_3QVal_Int_onehotd = 4'd2;
        2'd2: lizzieLet6_3QVal_Int_onehotd = 4'd4;
        2'd3: lizzieLet6_3QVal_Int_onehotd = 4'd8;
        default: lizzieLet6_3QVal_Int_onehotd = 4'd0;
      endcase
    else lizzieLet6_3QVal_Int_onehotd = 4'd0;
  assign lizzieLet6_5QVal_Int_3QNone_Int_d = lizzieLet6_3QVal_Int_onehotd[0];
  assign lizzieLet6_5QVal_Int_3QVal_Int_d = lizzieLet6_3QVal_Int_onehotd[1];
  assign lizzieLet6_5QVal_Int_3QNode_Int_d = lizzieLet6_3QVal_Int_onehotd[2];
  assign lizzieLet6_5QVal_Int_3QError_Int_d = lizzieLet6_3QVal_Int_onehotd[3];
  assign lizzieLet6_3QVal_Int_r = (| (lizzieLet6_3QVal_Int_onehotd & {lizzieLet6_5QVal_Int_3QError_Int_r,
                                                                      lizzieLet6_5QVal_Int_3QNode_Int_r,
                                                                      lizzieLet6_5QVal_Int_3QVal_Int_r,
                                                                      lizzieLet6_5QVal_Int_3QNone_Int_r}));
  assign lizzieLet6_5QVal_Int_3_r = lizzieLet6_3QVal_Int_r;
  
  /* fork (Ty Go) : (lizzieLet6_5QVal_Int_3QError_Int,Go) > [(lizzieLet6_5QVal_Int_3QError_Int_1,Go),
                                                        (lizzieLet6_5QVal_Int_3QError_Int_2,Go)] */
  logic [1:0] lizzieLet6_5QVal_Int_3QError_Int_emitted;
  logic [1:0] lizzieLet6_5QVal_Int_3QError_Int_done;
  assign lizzieLet6_5QVal_Int_3QError_Int_1_d = (lizzieLet6_5QVal_Int_3QError_Int_d[0] && (! lizzieLet6_5QVal_Int_3QError_Int_emitted[0]));
  assign lizzieLet6_5QVal_Int_3QError_Int_2_d = (lizzieLet6_5QVal_Int_3QError_Int_d[0] && (! lizzieLet6_5QVal_Int_3QError_Int_emitted[1]));
  assign lizzieLet6_5QVal_Int_3QError_Int_done = (lizzieLet6_5QVal_Int_3QError_Int_emitted | ({lizzieLet6_5QVal_Int_3QError_Int_2_d[0],
                                                                                               lizzieLet6_5QVal_Int_3QError_Int_1_d[0]} & {lizzieLet6_5QVal_Int_3QError_Int_2_r,
                                                                                                                                           lizzieLet6_5QVal_Int_3QError_Int_1_r}));
  assign lizzieLet6_5QVal_Int_3QError_Int_r = (& lizzieLet6_5QVal_Int_3QError_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_5QVal_Int_3QError_Int_emitted <= 2'd0;
    else
      lizzieLet6_5QVal_Int_3QError_Int_emitted <= (lizzieLet6_5QVal_Int_3QError_Int_r ? 2'd0 :
                                                   lizzieLet6_5QVal_Int_3QError_Int_done);
  
  /* dcon (Ty QTree_Int,
      Dcon QError_Int) : [(lizzieLet6_5QVal_Int_3QError_Int_1,Go)] > (lizzieLet6_5QVal_Int_3QError_Int_1QError_Int,QTree_Int) */
  assign lizzieLet6_5QVal_Int_3QError_Int_1QError_Int_d = QError_Int_dc((& {lizzieLet6_5QVal_Int_3QError_Int_1_d[0]}), lizzieLet6_5QVal_Int_3QError_Int_1_d);
  assign {lizzieLet6_5QVal_Int_3QError_Int_1_r} = {1 {(lizzieLet6_5QVal_Int_3QError_Int_1QError_Int_r && lizzieLet6_5QVal_Int_3QError_Int_1QError_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (lizzieLet6_5QVal_Int_3QError_Int_1QError_Int,QTree_Int) > (lizzieLet11_1_argbuf,QTree_Int) */
  QTree_Int_t lizzieLet6_5QVal_Int_3QError_Int_1QError_Int_bufchan_d;
  logic lizzieLet6_5QVal_Int_3QError_Int_1QError_Int_bufchan_r;
  assign lizzieLet6_5QVal_Int_3QError_Int_1QError_Int_r = ((! lizzieLet6_5QVal_Int_3QError_Int_1QError_Int_bufchan_d[0]) || lizzieLet6_5QVal_Int_3QError_Int_1QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_5QVal_Int_3QError_Int_1QError_Int_bufchan_d <= {66'd0,
                                                                 1'd0};
    else
      if (lizzieLet6_5QVal_Int_3QError_Int_1QError_Int_r)
        lizzieLet6_5QVal_Int_3QError_Int_1QError_Int_bufchan_d <= lizzieLet6_5QVal_Int_3QError_Int_1QError_Int_d;
  QTree_Int_t lizzieLet6_5QVal_Int_3QError_Int_1QError_Int_bufchan_buf;
  assign lizzieLet6_5QVal_Int_3QError_Int_1QError_Int_bufchan_r = (! lizzieLet6_5QVal_Int_3QError_Int_1QError_Int_bufchan_buf[0]);
  assign lizzieLet11_1_argbuf_d = (lizzieLet6_5QVal_Int_3QError_Int_1QError_Int_bufchan_buf[0] ? lizzieLet6_5QVal_Int_3QError_Int_1QError_Int_bufchan_buf :
                                   lizzieLet6_5QVal_Int_3QError_Int_1QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_5QVal_Int_3QError_Int_1QError_Int_bufchan_buf <= {66'd0,
                                                                   1'd0};
    else
      if ((lizzieLet11_1_argbuf_r && lizzieLet6_5QVal_Int_3QError_Int_1QError_Int_bufchan_buf[0]))
        lizzieLet6_5QVal_Int_3QError_Int_1QError_Int_bufchan_buf <= {66'd0,
                                                                     1'd0};
      else if (((! lizzieLet11_1_argbuf_r) && (! lizzieLet6_5QVal_Int_3QError_Int_1QError_Int_bufchan_buf[0])))
        lizzieLet6_5QVal_Int_3QError_Int_1QError_Int_bufchan_buf <= lizzieLet6_5QVal_Int_3QError_Int_1QError_Int_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet6_5QVal_Int_3QError_Int_2,Go) > (lizzieLet6_5QVal_Int_3QError_Int_2_argbuf,Go) */
  Go_t lizzieLet6_5QVal_Int_3QError_Int_2_bufchan_d;
  logic lizzieLet6_5QVal_Int_3QError_Int_2_bufchan_r;
  assign lizzieLet6_5QVal_Int_3QError_Int_2_r = ((! lizzieLet6_5QVal_Int_3QError_Int_2_bufchan_d[0]) || lizzieLet6_5QVal_Int_3QError_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_5QVal_Int_3QError_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet6_5QVal_Int_3QError_Int_2_r)
        lizzieLet6_5QVal_Int_3QError_Int_2_bufchan_d <= lizzieLet6_5QVal_Int_3QError_Int_2_d;
  Go_t lizzieLet6_5QVal_Int_3QError_Int_2_bufchan_buf;
  assign lizzieLet6_5QVal_Int_3QError_Int_2_bufchan_r = (! lizzieLet6_5QVal_Int_3QError_Int_2_bufchan_buf[0]);
  assign lizzieLet6_5QVal_Int_3QError_Int_2_argbuf_d = (lizzieLet6_5QVal_Int_3QError_Int_2_bufchan_buf[0] ? lizzieLet6_5QVal_Int_3QError_Int_2_bufchan_buf :
                                                        lizzieLet6_5QVal_Int_3QError_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_5QVal_Int_3QError_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet6_5QVal_Int_3QError_Int_2_argbuf_r && lizzieLet6_5QVal_Int_3QError_Int_2_bufchan_buf[0]))
        lizzieLet6_5QVal_Int_3QError_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet6_5QVal_Int_3QError_Int_2_argbuf_r) && (! lizzieLet6_5QVal_Int_3QError_Int_2_bufchan_buf[0])))
        lizzieLet6_5QVal_Int_3QError_Int_2_bufchan_buf <= lizzieLet6_5QVal_Int_3QError_Int_2_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet6_5QVal_Int_3QNode_Int,Go) > [(lizzieLet6_5QVal_Int_3QNode_Int_1,Go),
                                                       (lizzieLet6_5QVal_Int_3QNode_Int_2,Go)] */
  logic [1:0] lizzieLet6_5QVal_Int_3QNode_Int_emitted;
  logic [1:0] lizzieLet6_5QVal_Int_3QNode_Int_done;
  assign lizzieLet6_5QVal_Int_3QNode_Int_1_d = (lizzieLet6_5QVal_Int_3QNode_Int_d[0] && (! lizzieLet6_5QVal_Int_3QNode_Int_emitted[0]));
  assign lizzieLet6_5QVal_Int_3QNode_Int_2_d = (lizzieLet6_5QVal_Int_3QNode_Int_d[0] && (! lizzieLet6_5QVal_Int_3QNode_Int_emitted[1]));
  assign lizzieLet6_5QVal_Int_3QNode_Int_done = (lizzieLet6_5QVal_Int_3QNode_Int_emitted | ({lizzieLet6_5QVal_Int_3QNode_Int_2_d[0],
                                                                                             lizzieLet6_5QVal_Int_3QNode_Int_1_d[0]} & {lizzieLet6_5QVal_Int_3QNode_Int_2_r,
                                                                                                                                        lizzieLet6_5QVal_Int_3QNode_Int_1_r}));
  assign lizzieLet6_5QVal_Int_3QNode_Int_r = (& lizzieLet6_5QVal_Int_3QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_5QVal_Int_3QNode_Int_emitted <= 2'd0;
    else
      lizzieLet6_5QVal_Int_3QNode_Int_emitted <= (lizzieLet6_5QVal_Int_3QNode_Int_r ? 2'd0 :
                                                  lizzieLet6_5QVal_Int_3QNode_Int_done);
  
  /* dcon (Ty QTree_Int,
      Dcon QError_Int) : [(lizzieLet6_5QVal_Int_3QNode_Int_1,Go)] > (lizzieLet6_5QVal_Int_3QNode_Int_1QError_Int,QTree_Int) */
  assign lizzieLet6_5QVal_Int_3QNode_Int_1QError_Int_d = QError_Int_dc((& {lizzieLet6_5QVal_Int_3QNode_Int_1_d[0]}), lizzieLet6_5QVal_Int_3QNode_Int_1_d);
  assign {lizzieLet6_5QVal_Int_3QNode_Int_1_r} = {1 {(lizzieLet6_5QVal_Int_3QNode_Int_1QError_Int_r && lizzieLet6_5QVal_Int_3QNode_Int_1QError_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (lizzieLet6_5QVal_Int_3QNode_Int_1QError_Int,QTree_Int) > (lizzieLet10_1_argbuf,QTree_Int) */
  QTree_Int_t lizzieLet6_5QVal_Int_3QNode_Int_1QError_Int_bufchan_d;
  logic lizzieLet6_5QVal_Int_3QNode_Int_1QError_Int_bufchan_r;
  assign lizzieLet6_5QVal_Int_3QNode_Int_1QError_Int_r = ((! lizzieLet6_5QVal_Int_3QNode_Int_1QError_Int_bufchan_d[0]) || lizzieLet6_5QVal_Int_3QNode_Int_1QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_5QVal_Int_3QNode_Int_1QError_Int_bufchan_d <= {66'd0,
                                                                1'd0};
    else
      if (lizzieLet6_5QVal_Int_3QNode_Int_1QError_Int_r)
        lizzieLet6_5QVal_Int_3QNode_Int_1QError_Int_bufchan_d <= lizzieLet6_5QVal_Int_3QNode_Int_1QError_Int_d;
  QTree_Int_t lizzieLet6_5QVal_Int_3QNode_Int_1QError_Int_bufchan_buf;
  assign lizzieLet6_5QVal_Int_3QNode_Int_1QError_Int_bufchan_r = (! lizzieLet6_5QVal_Int_3QNode_Int_1QError_Int_bufchan_buf[0]);
  assign lizzieLet10_1_argbuf_d = (lizzieLet6_5QVal_Int_3QNode_Int_1QError_Int_bufchan_buf[0] ? lizzieLet6_5QVal_Int_3QNode_Int_1QError_Int_bufchan_buf :
                                   lizzieLet6_5QVal_Int_3QNode_Int_1QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_5QVal_Int_3QNode_Int_1QError_Int_bufchan_buf <= {66'd0,
                                                                  1'd0};
    else
      if ((lizzieLet10_1_argbuf_r && lizzieLet6_5QVal_Int_3QNode_Int_1QError_Int_bufchan_buf[0]))
        lizzieLet6_5QVal_Int_3QNode_Int_1QError_Int_bufchan_buf <= {66'd0,
                                                                    1'd0};
      else if (((! lizzieLet10_1_argbuf_r) && (! lizzieLet6_5QVal_Int_3QNode_Int_1QError_Int_bufchan_buf[0])))
        lizzieLet6_5QVal_Int_3QNode_Int_1QError_Int_bufchan_buf <= lizzieLet6_5QVal_Int_3QNode_Int_1QError_Int_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet6_5QVal_Int_3QNode_Int_2,Go) > (lizzieLet6_5QVal_Int_3QNode_Int_2_argbuf,Go) */
  Go_t lizzieLet6_5QVal_Int_3QNode_Int_2_bufchan_d;
  logic lizzieLet6_5QVal_Int_3QNode_Int_2_bufchan_r;
  assign lizzieLet6_5QVal_Int_3QNode_Int_2_r = ((! lizzieLet6_5QVal_Int_3QNode_Int_2_bufchan_d[0]) || lizzieLet6_5QVal_Int_3QNode_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_5QVal_Int_3QNode_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet6_5QVal_Int_3QNode_Int_2_r)
        lizzieLet6_5QVal_Int_3QNode_Int_2_bufchan_d <= lizzieLet6_5QVal_Int_3QNode_Int_2_d;
  Go_t lizzieLet6_5QVal_Int_3QNode_Int_2_bufchan_buf;
  assign lizzieLet6_5QVal_Int_3QNode_Int_2_bufchan_r = (! lizzieLet6_5QVal_Int_3QNode_Int_2_bufchan_buf[0]);
  assign lizzieLet6_5QVal_Int_3QNode_Int_2_argbuf_d = (lizzieLet6_5QVal_Int_3QNode_Int_2_bufchan_buf[0] ? lizzieLet6_5QVal_Int_3QNode_Int_2_bufchan_buf :
                                                       lizzieLet6_5QVal_Int_3QNode_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_5QVal_Int_3QNode_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet6_5QVal_Int_3QNode_Int_2_argbuf_r && lizzieLet6_5QVal_Int_3QNode_Int_2_bufchan_buf[0]))
        lizzieLet6_5QVal_Int_3QNode_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet6_5QVal_Int_3QNode_Int_2_argbuf_r) && (! lizzieLet6_5QVal_Int_3QNode_Int_2_bufchan_buf[0])))
        lizzieLet6_5QVal_Int_3QNode_Int_2_bufchan_buf <= lizzieLet6_5QVal_Int_3QNode_Int_2_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet6_5QVal_Int_3QNone_Int,Go) > (lizzieLet6_5QVal_Int_3QNone_Int_1_argbuf,Go) */
  Go_t lizzieLet6_5QVal_Int_3QNone_Int_bufchan_d;
  logic lizzieLet6_5QVal_Int_3QNone_Int_bufchan_r;
  assign lizzieLet6_5QVal_Int_3QNone_Int_r = ((! lizzieLet6_5QVal_Int_3QNone_Int_bufchan_d[0]) || lizzieLet6_5QVal_Int_3QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_5QVal_Int_3QNone_Int_bufchan_d <= 1'd0;
    else
      if (lizzieLet6_5QVal_Int_3QNone_Int_r)
        lizzieLet6_5QVal_Int_3QNone_Int_bufchan_d <= lizzieLet6_5QVal_Int_3QNone_Int_d;
  Go_t lizzieLet6_5QVal_Int_3QNone_Int_bufchan_buf;
  assign lizzieLet6_5QVal_Int_3QNone_Int_bufchan_r = (! lizzieLet6_5QVal_Int_3QNone_Int_bufchan_buf[0]);
  assign lizzieLet6_5QVal_Int_3QNone_Int_1_argbuf_d = (lizzieLet6_5QVal_Int_3QNone_Int_bufchan_buf[0] ? lizzieLet6_5QVal_Int_3QNone_Int_bufchan_buf :
                                                       lizzieLet6_5QVal_Int_3QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_5QVal_Int_3QNone_Int_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet6_5QVal_Int_3QNone_Int_1_argbuf_r && lizzieLet6_5QVal_Int_3QNone_Int_bufchan_buf[0]))
        lizzieLet6_5QVal_Int_3QNone_Int_bufchan_buf <= 1'd0;
      else if (((! lizzieLet6_5QVal_Int_3QNone_Int_1_argbuf_r) && (! lizzieLet6_5QVal_Int_3QNone_Int_bufchan_buf[0])))
        lizzieLet6_5QVal_Int_3QNone_Int_bufchan_buf <= lizzieLet6_5QVal_Int_3QNone_Int_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet6_5QVal_Int_3QVal_Int,Go) > [(lizzieLet6_5QVal_Int_3QVal_Int_1,Go),
                                                      (lizzieLet6_5QVal_Int_3QVal_Int_2,Go)] */
  logic [1:0] lizzieLet6_5QVal_Int_3QVal_Int_emitted;
  logic [1:0] lizzieLet6_5QVal_Int_3QVal_Int_done;
  assign lizzieLet6_5QVal_Int_3QVal_Int_1_d = (lizzieLet6_5QVal_Int_3QVal_Int_d[0] && (! lizzieLet6_5QVal_Int_3QVal_Int_emitted[0]));
  assign lizzieLet6_5QVal_Int_3QVal_Int_2_d = (lizzieLet6_5QVal_Int_3QVal_Int_d[0] && (! lizzieLet6_5QVal_Int_3QVal_Int_emitted[1]));
  assign lizzieLet6_5QVal_Int_3QVal_Int_done = (lizzieLet6_5QVal_Int_3QVal_Int_emitted | ({lizzieLet6_5QVal_Int_3QVal_Int_2_d[0],
                                                                                           lizzieLet6_5QVal_Int_3QVal_Int_1_d[0]} & {lizzieLet6_5QVal_Int_3QVal_Int_2_r,
                                                                                                                                     lizzieLet6_5QVal_Int_3QVal_Int_1_r}));
  assign lizzieLet6_5QVal_Int_3QVal_Int_r = (& lizzieLet6_5QVal_Int_3QVal_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_5QVal_Int_3QVal_Int_emitted <= 2'd0;
    else
      lizzieLet6_5QVal_Int_3QVal_Int_emitted <= (lizzieLet6_5QVal_Int_3QVal_Int_r ? 2'd0 :
                                                 lizzieLet6_5QVal_Int_3QVal_Int_done);
  
  /* buf (Ty Go) : (lizzieLet6_5QVal_Int_3QVal_Int_1,Go) > (lizzieLet6_5QVal_Int_3QVal_Int_1_argbuf,Go) */
  Go_t lizzieLet6_5QVal_Int_3QVal_Int_1_bufchan_d;
  logic lizzieLet6_5QVal_Int_3QVal_Int_1_bufchan_r;
  assign lizzieLet6_5QVal_Int_3QVal_Int_1_r = ((! lizzieLet6_5QVal_Int_3QVal_Int_1_bufchan_d[0]) || lizzieLet6_5QVal_Int_3QVal_Int_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_5QVal_Int_3QVal_Int_1_bufchan_d <= 1'd0;
    else
      if (lizzieLet6_5QVal_Int_3QVal_Int_1_r)
        lizzieLet6_5QVal_Int_3QVal_Int_1_bufchan_d <= lizzieLet6_5QVal_Int_3QVal_Int_1_d;
  Go_t lizzieLet6_5QVal_Int_3QVal_Int_1_bufchan_buf;
  assign lizzieLet6_5QVal_Int_3QVal_Int_1_bufchan_r = (! lizzieLet6_5QVal_Int_3QVal_Int_1_bufchan_buf[0]);
  assign lizzieLet6_5QVal_Int_3QVal_Int_1_argbuf_d = (lizzieLet6_5QVal_Int_3QVal_Int_1_bufchan_buf[0] ? lizzieLet6_5QVal_Int_3QVal_Int_1_bufchan_buf :
                                                      lizzieLet6_5QVal_Int_3QVal_Int_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_5QVal_Int_3QVal_Int_1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet6_5QVal_Int_3QVal_Int_1_argbuf_r && lizzieLet6_5QVal_Int_3QVal_Int_1_bufchan_buf[0]))
        lizzieLet6_5QVal_Int_3QVal_Int_1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet6_5QVal_Int_3QVal_Int_1_argbuf_r) && (! lizzieLet6_5QVal_Int_3QVal_Int_1_bufchan_buf[0])))
        lizzieLet6_5QVal_Int_3QVal_Int_1_bufchan_buf <= lizzieLet6_5QVal_Int_3QVal_Int_1_bufchan_d;
  
  /* dcon (Ty TupGo___MyDTInt_Bool___Int,
      Dcon TupGo___MyDTInt_Bool___Int) : [(lizzieLet6_5QVal_Int_3QVal_Int_1_argbuf,Go),
                                          (lizzieLet6_5QVal_Int_4QVal_Int_1_argbuf,MyDTInt_Bool),
                                          (es_1_1_argbuf,Int)] > (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int2,TupGo___MyDTInt_Bool___Int) */
  assign applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int2_d = TupGo___MyDTInt_Bool___Int_dc((& {lizzieLet6_5QVal_Int_3QVal_Int_1_argbuf_d[0],
                                                                                            lizzieLet6_5QVal_Int_4QVal_Int_1_argbuf_d[0],
                                                                                            es_1_1_argbuf_d[0]}), lizzieLet6_5QVal_Int_3QVal_Int_1_argbuf_d, lizzieLet6_5QVal_Int_4QVal_Int_1_argbuf_d, es_1_1_argbuf_d);
  assign {lizzieLet6_5QVal_Int_3QVal_Int_1_argbuf_r,
          lizzieLet6_5QVal_Int_4QVal_Int_1_argbuf_r,
          es_1_1_argbuf_r} = {3 {(applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int2_r && applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int2_d[0])}};
  
  /* demux (Ty QTree_Int,
       Ty MyDTInt_Bool) : (lizzieLet6_5QVal_Int_4,QTree_Int) (lizzieLet6_4QVal_Int,MyDTInt_Bool) > [(_18,MyDTInt_Bool),
                                                                                                    (lizzieLet6_5QVal_Int_4QVal_Int,MyDTInt_Bool),
                                                                                                    (_17,MyDTInt_Bool),
                                                                                                    (_16,MyDTInt_Bool)] */
  logic [3:0] lizzieLet6_4QVal_Int_onehotd;
  always_comb
    if ((lizzieLet6_5QVal_Int_4_d[0] && lizzieLet6_4QVal_Int_d[0]))
      unique case (lizzieLet6_5QVal_Int_4_d[2:1])
        2'd0: lizzieLet6_4QVal_Int_onehotd = 4'd1;
        2'd1: lizzieLet6_4QVal_Int_onehotd = 4'd2;
        2'd2: lizzieLet6_4QVal_Int_onehotd = 4'd4;
        2'd3: lizzieLet6_4QVal_Int_onehotd = 4'd8;
        default: lizzieLet6_4QVal_Int_onehotd = 4'd0;
      endcase
    else lizzieLet6_4QVal_Int_onehotd = 4'd0;
  assign _18_d = lizzieLet6_4QVal_Int_onehotd[0];
  assign lizzieLet6_5QVal_Int_4QVal_Int_d = lizzieLet6_4QVal_Int_onehotd[1];
  assign _17_d = lizzieLet6_4QVal_Int_onehotd[2];
  assign _16_d = lizzieLet6_4QVal_Int_onehotd[3];
  assign lizzieLet6_4QVal_Int_r = (| (lizzieLet6_4QVal_Int_onehotd & {_16_r,
                                                                      _17_r,
                                                                      lizzieLet6_5QVal_Int_4QVal_Int_r,
                                                                      _18_r}));
  assign lizzieLet6_5QVal_Int_4_r = lizzieLet6_4QVal_Int_r;
  
  /* buf (Ty MyDTInt_Bool) : (lizzieLet6_5QVal_Int_4QVal_Int,MyDTInt_Bool) > (lizzieLet6_5QVal_Int_4QVal_Int_1_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t lizzieLet6_5QVal_Int_4QVal_Int_bufchan_d;
  logic lizzieLet6_5QVal_Int_4QVal_Int_bufchan_r;
  assign lizzieLet6_5QVal_Int_4QVal_Int_r = ((! lizzieLet6_5QVal_Int_4QVal_Int_bufchan_d[0]) || lizzieLet6_5QVal_Int_4QVal_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_5QVal_Int_4QVal_Int_bufchan_d <= 1'd0;
    else
      if (lizzieLet6_5QVal_Int_4QVal_Int_r)
        lizzieLet6_5QVal_Int_4QVal_Int_bufchan_d <= lizzieLet6_5QVal_Int_4QVal_Int_d;
  MyDTInt_Bool_t lizzieLet6_5QVal_Int_4QVal_Int_bufchan_buf;
  assign lizzieLet6_5QVal_Int_4QVal_Int_bufchan_r = (! lizzieLet6_5QVal_Int_4QVal_Int_bufchan_buf[0]);
  assign lizzieLet6_5QVal_Int_4QVal_Int_1_argbuf_d = (lizzieLet6_5QVal_Int_4QVal_Int_bufchan_buf[0] ? lizzieLet6_5QVal_Int_4QVal_Int_bufchan_buf :
                                                      lizzieLet6_5QVal_Int_4QVal_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_5QVal_Int_4QVal_Int_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet6_5QVal_Int_4QVal_Int_1_argbuf_r && lizzieLet6_5QVal_Int_4QVal_Int_bufchan_buf[0]))
        lizzieLet6_5QVal_Int_4QVal_Int_bufchan_buf <= 1'd0;
      else if (((! lizzieLet6_5QVal_Int_4QVal_Int_1_argbuf_r) && (! lizzieLet6_5QVal_Int_4QVal_Int_bufchan_buf[0])))
        lizzieLet6_5QVal_Int_4QVal_Int_bufchan_buf <= lizzieLet6_5QVal_Int_4QVal_Int_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty MyDTInt_Int_Int) : (lizzieLet6_5QVal_Int_5,QTree_Int) (lizzieLet6_6QVal_Int,MyDTInt_Int_Int) > [(_15,MyDTInt_Int_Int),
                                                                                                          (lizzieLet6_5QVal_Int_5QVal_Int,MyDTInt_Int_Int),
                                                                                                          (_14,MyDTInt_Int_Int),
                                                                                                          (_13,MyDTInt_Int_Int)] */
  logic [3:0] lizzieLet6_6QVal_Int_onehotd;
  always_comb
    if ((lizzieLet6_5QVal_Int_5_d[0] && lizzieLet6_6QVal_Int_d[0]))
      unique case (lizzieLet6_5QVal_Int_5_d[2:1])
        2'd0: lizzieLet6_6QVal_Int_onehotd = 4'd1;
        2'd1: lizzieLet6_6QVal_Int_onehotd = 4'd2;
        2'd2: lizzieLet6_6QVal_Int_onehotd = 4'd4;
        2'd3: lizzieLet6_6QVal_Int_onehotd = 4'd8;
        default: lizzieLet6_6QVal_Int_onehotd = 4'd0;
      endcase
    else lizzieLet6_6QVal_Int_onehotd = 4'd0;
  assign _15_d = lizzieLet6_6QVal_Int_onehotd[0];
  assign lizzieLet6_5QVal_Int_5QVal_Int_d = lizzieLet6_6QVal_Int_onehotd[1];
  assign _14_d = lizzieLet6_6QVal_Int_onehotd[2];
  assign _13_d = lizzieLet6_6QVal_Int_onehotd[3];
  assign lizzieLet6_6QVal_Int_r = (| (lizzieLet6_6QVal_Int_onehotd & {_13_r,
                                                                      _14_r,
                                                                      lizzieLet6_5QVal_Int_5QVal_Int_r,
                                                                      _15_r}));
  assign lizzieLet6_5QVal_Int_5_r = lizzieLet6_6QVal_Int_r;
  
  /* fork (Ty MyDTInt_Int_Int) : (lizzieLet6_5QVal_Int_5QVal_Int,MyDTInt_Int_Int) > [(lizzieLet6_5QVal_Int_5QVal_Int_1,MyDTInt_Int_Int),
                                                                                (lizzieLet6_5QVal_Int_5QVal_Int_2,MyDTInt_Int_Int)] */
  logic [1:0] lizzieLet6_5QVal_Int_5QVal_Int_emitted;
  logic [1:0] lizzieLet6_5QVal_Int_5QVal_Int_done;
  assign lizzieLet6_5QVal_Int_5QVal_Int_1_d = (lizzieLet6_5QVal_Int_5QVal_Int_d[0] && (! lizzieLet6_5QVal_Int_5QVal_Int_emitted[0]));
  assign lizzieLet6_5QVal_Int_5QVal_Int_2_d = (lizzieLet6_5QVal_Int_5QVal_Int_d[0] && (! lizzieLet6_5QVal_Int_5QVal_Int_emitted[1]));
  assign lizzieLet6_5QVal_Int_5QVal_Int_done = (lizzieLet6_5QVal_Int_5QVal_Int_emitted | ({lizzieLet6_5QVal_Int_5QVal_Int_2_d[0],
                                                                                           lizzieLet6_5QVal_Int_5QVal_Int_1_d[0]} & {lizzieLet6_5QVal_Int_5QVal_Int_2_r,
                                                                                                                                     lizzieLet6_5QVal_Int_5QVal_Int_1_r}));
  assign lizzieLet6_5QVal_Int_5QVal_Int_r = (& lizzieLet6_5QVal_Int_5QVal_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_5QVal_Int_5QVal_Int_emitted <= 2'd0;
    else
      lizzieLet6_5QVal_Int_5QVal_Int_emitted <= (lizzieLet6_5QVal_Int_5QVal_Int_r ? 2'd0 :
                                                 lizzieLet6_5QVal_Int_5QVal_Int_done);
  
  /* buf (Ty MyDTInt_Int_Int) : (lizzieLet6_5QVal_Int_5QVal_Int_1,MyDTInt_Int_Int) > (lizzieLet6_5QVal_Int_5QVal_Int_1_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t lizzieLet6_5QVal_Int_5QVal_Int_1_bufchan_d;
  logic lizzieLet6_5QVal_Int_5QVal_Int_1_bufchan_r;
  assign lizzieLet6_5QVal_Int_5QVal_Int_1_r = ((! lizzieLet6_5QVal_Int_5QVal_Int_1_bufchan_d[0]) || lizzieLet6_5QVal_Int_5QVal_Int_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_5QVal_Int_5QVal_Int_1_bufchan_d <= 1'd0;
    else
      if (lizzieLet6_5QVal_Int_5QVal_Int_1_r)
        lizzieLet6_5QVal_Int_5QVal_Int_1_bufchan_d <= lizzieLet6_5QVal_Int_5QVal_Int_1_d;
  MyDTInt_Int_Int_t lizzieLet6_5QVal_Int_5QVal_Int_1_bufchan_buf;
  assign lizzieLet6_5QVal_Int_5QVal_Int_1_bufchan_r = (! lizzieLet6_5QVal_Int_5QVal_Int_1_bufchan_buf[0]);
  assign lizzieLet6_5QVal_Int_5QVal_Int_1_argbuf_d = (lizzieLet6_5QVal_Int_5QVal_Int_1_bufchan_buf[0] ? lizzieLet6_5QVal_Int_5QVal_Int_1_bufchan_buf :
                                                      lizzieLet6_5QVal_Int_5QVal_Int_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_5QVal_Int_5QVal_Int_1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet6_5QVal_Int_5QVal_Int_1_argbuf_r && lizzieLet6_5QVal_Int_5QVal_Int_1_bufchan_buf[0]))
        lizzieLet6_5QVal_Int_5QVal_Int_1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet6_5QVal_Int_5QVal_Int_1_argbuf_r) && (! lizzieLet6_5QVal_Int_5QVal_Int_1_bufchan_buf[0])))
        lizzieLet6_5QVal_Int_5QVal_Int_1_bufchan_buf <= lizzieLet6_5QVal_Int_5QVal_Int_1_bufchan_d;
  
  /* dcon (Ty TupMyDTInt_Int_Int___Int___Int,
      Dcon TupMyDTInt_Int_Int___Int___Int) : [(lizzieLet6_5QVal_Int_5QVal_Int_1_argbuf,MyDTInt_Int_Int),
                                              (lizzieLet6_5QVal_Int_8QVal_Int_1_argbuf,Int),
                                              (vafo_1_argbuf,Int)] > (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int3,TupMyDTInt_Int_Int___Int___Int) */
  assign applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int3_d = TupMyDTInt_Int_Int___Int___Int_dc((& {lizzieLet6_5QVal_Int_5QVal_Int_1_argbuf_d[0],
                                                                                                       lizzieLet6_5QVal_Int_8QVal_Int_1_argbuf_d[0],
                                                                                                       vafo_1_argbuf_d[0]}), lizzieLet6_5QVal_Int_5QVal_Int_1_argbuf_d, lizzieLet6_5QVal_Int_8QVal_Int_1_argbuf_d, vafo_1_argbuf_d);
  assign {lizzieLet6_5QVal_Int_5QVal_Int_1_argbuf_r,
          lizzieLet6_5QVal_Int_8QVal_Int_1_argbuf_r,
          vafo_1_argbuf_r} = {3 {(applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int3_r && applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int3_d[0])}};
  
  /* demux (Ty QTree_Int,
       Ty Pointer_QTree_Int) : (lizzieLet6_5QVal_Int_6,QTree_Int) (lizzieLet6_7QVal_Int,Pointer_QTree_Int) > [(lizzieLet6_5QVal_Int_6QNone_Int,Pointer_QTree_Int),
                                                                                                              (_12,Pointer_QTree_Int),
                                                                                                              (_11,Pointer_QTree_Int),
                                                                                                              (_10,Pointer_QTree_Int)] */
  logic [3:0] lizzieLet6_7QVal_Int_onehotd;
  always_comb
    if ((lizzieLet6_5QVal_Int_6_d[0] && lizzieLet6_7QVal_Int_d[0]))
      unique case (lizzieLet6_5QVal_Int_6_d[2:1])
        2'd0: lizzieLet6_7QVal_Int_onehotd = 4'd1;
        2'd1: lizzieLet6_7QVal_Int_onehotd = 4'd2;
        2'd2: lizzieLet6_7QVal_Int_onehotd = 4'd4;
        2'd3: lizzieLet6_7QVal_Int_onehotd = 4'd8;
        default: lizzieLet6_7QVal_Int_onehotd = 4'd0;
      endcase
    else lizzieLet6_7QVal_Int_onehotd = 4'd0;
  assign lizzieLet6_5QVal_Int_6QNone_Int_d = {lizzieLet6_7QVal_Int_d[16:1],
                                              lizzieLet6_7QVal_Int_onehotd[0]};
  assign _12_d = {lizzieLet6_7QVal_Int_d[16:1],
                  lizzieLet6_7QVal_Int_onehotd[1]};
  assign _11_d = {lizzieLet6_7QVal_Int_d[16:1],
                  lizzieLet6_7QVal_Int_onehotd[2]};
  assign _10_d = {lizzieLet6_7QVal_Int_d[16:1],
                  lizzieLet6_7QVal_Int_onehotd[3]};
  assign lizzieLet6_7QVal_Int_r = (| (lizzieLet6_7QVal_Int_onehotd & {_10_r,
                                                                      _11_r,
                                                                      _12_r,
                                                                      lizzieLet6_5QVal_Int_6QNone_Int_r}));
  assign lizzieLet6_5QVal_Int_6_r = lizzieLet6_7QVal_Int_r;
  
  /* buf (Ty Pointer_QTree_Int) : (lizzieLet6_5QVal_Int_6QNone_Int,Pointer_QTree_Int) > (lizzieLet6_5QVal_Int_6QNone_Int_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t lizzieLet6_5QVal_Int_6QNone_Int_bufchan_d;
  logic lizzieLet6_5QVal_Int_6QNone_Int_bufchan_r;
  assign lizzieLet6_5QVal_Int_6QNone_Int_r = ((! lizzieLet6_5QVal_Int_6QNone_Int_bufchan_d[0]) || lizzieLet6_5QVal_Int_6QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_5QVal_Int_6QNone_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet6_5QVal_Int_6QNone_Int_r)
        lizzieLet6_5QVal_Int_6QNone_Int_bufchan_d <= lizzieLet6_5QVal_Int_6QNone_Int_d;
  Pointer_QTree_Int_t lizzieLet6_5QVal_Int_6QNone_Int_bufchan_buf;
  assign lizzieLet6_5QVal_Int_6QNone_Int_bufchan_r = (! lizzieLet6_5QVal_Int_6QNone_Int_bufchan_buf[0]);
  assign lizzieLet6_5QVal_Int_6QNone_Int_1_argbuf_d = (lizzieLet6_5QVal_Int_6QNone_Int_bufchan_buf[0] ? lizzieLet6_5QVal_Int_6QNone_Int_bufchan_buf :
                                                       lizzieLet6_5QVal_Int_6QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_5QVal_Int_6QNone_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet6_5QVal_Int_6QNone_Int_1_argbuf_r && lizzieLet6_5QVal_Int_6QNone_Int_bufchan_buf[0]))
        lizzieLet6_5QVal_Int_6QNone_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet6_5QVal_Int_6QNone_Int_1_argbuf_r) && (! lizzieLet6_5QVal_Int_6QNone_Int_bufchan_buf[0])))
        lizzieLet6_5QVal_Int_6QNone_Int_bufchan_buf <= lizzieLet6_5QVal_Int_6QNone_Int_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_CTf''''''''''''_f''''''''''''_Int) : (lizzieLet6_5QVal_Int_7,QTree_Int) (lizzieLet6_8QVal_Int,Pointer_CTf''''''''''''_f''''''''''''_Int) > [(lizzieLet6_5QVal_Int_7QNone_Int,Pointer_CTf''''''''''''_f''''''''''''_Int),
                                                                                                                                                              (lizzieLet6_5QVal_Int_7QVal_Int,Pointer_CTf''''''''''''_f''''''''''''_Int),
                                                                                                                                                              (lizzieLet6_5QVal_Int_7QNode_Int,Pointer_CTf''''''''''''_f''''''''''''_Int),
                                                                                                                                                              (lizzieLet6_5QVal_Int_7QError_Int,Pointer_CTf''''''''''''_f''''''''''''_Int)] */
  logic [3:0] lizzieLet6_8QVal_Int_onehotd;
  always_comb
    if ((lizzieLet6_5QVal_Int_7_d[0] && lizzieLet6_8QVal_Int_d[0]))
      unique case (lizzieLet6_5QVal_Int_7_d[2:1])
        2'd0: lizzieLet6_8QVal_Int_onehotd = 4'd1;
        2'd1: lizzieLet6_8QVal_Int_onehotd = 4'd2;
        2'd2: lizzieLet6_8QVal_Int_onehotd = 4'd4;
        2'd3: lizzieLet6_8QVal_Int_onehotd = 4'd8;
        default: lizzieLet6_8QVal_Int_onehotd = 4'd0;
      endcase
    else lizzieLet6_8QVal_Int_onehotd = 4'd0;
  assign lizzieLet6_5QVal_Int_7QNone_Int_d = {lizzieLet6_8QVal_Int_d[16:1],
                                              lizzieLet6_8QVal_Int_onehotd[0]};
  assign lizzieLet6_5QVal_Int_7QVal_Int_d = {lizzieLet6_8QVal_Int_d[16:1],
                                             lizzieLet6_8QVal_Int_onehotd[1]};
  assign lizzieLet6_5QVal_Int_7QNode_Int_d = {lizzieLet6_8QVal_Int_d[16:1],
                                              lizzieLet6_8QVal_Int_onehotd[2]};
  assign lizzieLet6_5QVal_Int_7QError_Int_d = {lizzieLet6_8QVal_Int_d[16:1],
                                               lizzieLet6_8QVal_Int_onehotd[3]};
  assign lizzieLet6_8QVal_Int_r = (| (lizzieLet6_8QVal_Int_onehotd & {lizzieLet6_5QVal_Int_7QError_Int_r,
                                                                      lizzieLet6_5QVal_Int_7QNode_Int_r,
                                                                      lizzieLet6_5QVal_Int_7QVal_Int_r,
                                                                      lizzieLet6_5QVal_Int_7QNone_Int_r}));
  assign lizzieLet6_5QVal_Int_7_r = lizzieLet6_8QVal_Int_r;
  
  /* buf (Ty Pointer_CTf''''''''''''_f''''''''''''_Int) : (lizzieLet6_5QVal_Int_7QError_Int,Pointer_CTf''''''''''''_f''''''''''''_Int) > (lizzieLet6_5QVal_Int_7QError_Int_1_argbuf,Pointer_CTf''''''''''''_f''''''''''''_Int) */
  \Pointer_CTf''''''''''''_f''''''''''''_Int_t  lizzieLet6_5QVal_Int_7QError_Int_bufchan_d;
  logic lizzieLet6_5QVal_Int_7QError_Int_bufchan_r;
  assign lizzieLet6_5QVal_Int_7QError_Int_r = ((! lizzieLet6_5QVal_Int_7QError_Int_bufchan_d[0]) || lizzieLet6_5QVal_Int_7QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_5QVal_Int_7QError_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet6_5QVal_Int_7QError_Int_r)
        lizzieLet6_5QVal_Int_7QError_Int_bufchan_d <= lizzieLet6_5QVal_Int_7QError_Int_d;
  \Pointer_CTf''''''''''''_f''''''''''''_Int_t  lizzieLet6_5QVal_Int_7QError_Int_bufchan_buf;
  assign lizzieLet6_5QVal_Int_7QError_Int_bufchan_r = (! lizzieLet6_5QVal_Int_7QError_Int_bufchan_buf[0]);
  assign lizzieLet6_5QVal_Int_7QError_Int_1_argbuf_d = (lizzieLet6_5QVal_Int_7QError_Int_bufchan_buf[0] ? lizzieLet6_5QVal_Int_7QError_Int_bufchan_buf :
                                                        lizzieLet6_5QVal_Int_7QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_5QVal_Int_7QError_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet6_5QVal_Int_7QError_Int_1_argbuf_r && lizzieLet6_5QVal_Int_7QError_Int_bufchan_buf[0]))
        lizzieLet6_5QVal_Int_7QError_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet6_5QVal_Int_7QError_Int_1_argbuf_r) && (! lizzieLet6_5QVal_Int_7QError_Int_bufchan_buf[0])))
        lizzieLet6_5QVal_Int_7QError_Int_bufchan_buf <= lizzieLet6_5QVal_Int_7QError_Int_bufchan_d;
  
  /* buf (Ty Pointer_CTf''''''''''''_f''''''''''''_Int) : (lizzieLet6_5QVal_Int_7QNode_Int,Pointer_CTf''''''''''''_f''''''''''''_Int) > (lizzieLet6_5QVal_Int_7QNode_Int_1_argbuf,Pointer_CTf''''''''''''_f''''''''''''_Int) */
  \Pointer_CTf''''''''''''_f''''''''''''_Int_t  lizzieLet6_5QVal_Int_7QNode_Int_bufchan_d;
  logic lizzieLet6_5QVal_Int_7QNode_Int_bufchan_r;
  assign lizzieLet6_5QVal_Int_7QNode_Int_r = ((! lizzieLet6_5QVal_Int_7QNode_Int_bufchan_d[0]) || lizzieLet6_5QVal_Int_7QNode_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_5QVal_Int_7QNode_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet6_5QVal_Int_7QNode_Int_r)
        lizzieLet6_5QVal_Int_7QNode_Int_bufchan_d <= lizzieLet6_5QVal_Int_7QNode_Int_d;
  \Pointer_CTf''''''''''''_f''''''''''''_Int_t  lizzieLet6_5QVal_Int_7QNode_Int_bufchan_buf;
  assign lizzieLet6_5QVal_Int_7QNode_Int_bufchan_r = (! lizzieLet6_5QVal_Int_7QNode_Int_bufchan_buf[0]);
  assign lizzieLet6_5QVal_Int_7QNode_Int_1_argbuf_d = (lizzieLet6_5QVal_Int_7QNode_Int_bufchan_buf[0] ? lizzieLet6_5QVal_Int_7QNode_Int_bufchan_buf :
                                                       lizzieLet6_5QVal_Int_7QNode_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_5QVal_Int_7QNode_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet6_5QVal_Int_7QNode_Int_1_argbuf_r && lizzieLet6_5QVal_Int_7QNode_Int_bufchan_buf[0]))
        lizzieLet6_5QVal_Int_7QNode_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet6_5QVal_Int_7QNode_Int_1_argbuf_r) && (! lizzieLet6_5QVal_Int_7QNode_Int_bufchan_buf[0])))
        lizzieLet6_5QVal_Int_7QNode_Int_bufchan_buf <= lizzieLet6_5QVal_Int_7QNode_Int_bufchan_d;
  
  /* buf (Ty Pointer_CTf''''''''''''_f''''''''''''_Int) : (lizzieLet6_5QVal_Int_7QNone_Int,Pointer_CTf''''''''''''_f''''''''''''_Int) > (lizzieLet6_5QVal_Int_7QNone_Int_1_argbuf,Pointer_CTf''''''''''''_f''''''''''''_Int) */
  \Pointer_CTf''''''''''''_f''''''''''''_Int_t  lizzieLet6_5QVal_Int_7QNone_Int_bufchan_d;
  logic lizzieLet6_5QVal_Int_7QNone_Int_bufchan_r;
  assign lizzieLet6_5QVal_Int_7QNone_Int_r = ((! lizzieLet6_5QVal_Int_7QNone_Int_bufchan_d[0]) || lizzieLet6_5QVal_Int_7QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_5QVal_Int_7QNone_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet6_5QVal_Int_7QNone_Int_r)
        lizzieLet6_5QVal_Int_7QNone_Int_bufchan_d <= lizzieLet6_5QVal_Int_7QNone_Int_d;
  \Pointer_CTf''''''''''''_f''''''''''''_Int_t  lizzieLet6_5QVal_Int_7QNone_Int_bufchan_buf;
  assign lizzieLet6_5QVal_Int_7QNone_Int_bufchan_r = (! lizzieLet6_5QVal_Int_7QNone_Int_bufchan_buf[0]);
  assign lizzieLet6_5QVal_Int_7QNone_Int_1_argbuf_d = (lizzieLet6_5QVal_Int_7QNone_Int_bufchan_buf[0] ? lizzieLet6_5QVal_Int_7QNone_Int_bufchan_buf :
                                                       lizzieLet6_5QVal_Int_7QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_5QVal_Int_7QNone_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet6_5QVal_Int_7QNone_Int_1_argbuf_r && lizzieLet6_5QVal_Int_7QNone_Int_bufchan_buf[0]))
        lizzieLet6_5QVal_Int_7QNone_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet6_5QVal_Int_7QNone_Int_1_argbuf_r) && (! lizzieLet6_5QVal_Int_7QNone_Int_bufchan_buf[0])))
        lizzieLet6_5QVal_Int_7QNone_Int_bufchan_buf <= lizzieLet6_5QVal_Int_7QNone_Int_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Int) : (lizzieLet6_5QVal_Int_8,QTree_Int) (v1afn_destruct,Int) > [(_9,Int),
                                                                            (lizzieLet6_5QVal_Int_8QVal_Int,Int),
                                                                            (_8,Int),
                                                                            (_7,Int)] */
  logic [3:0] v1afn_destruct_onehotd;
  always_comb
    if ((lizzieLet6_5QVal_Int_8_d[0] && v1afn_destruct_d[0]))
      unique case (lizzieLet6_5QVal_Int_8_d[2:1])
        2'd0: v1afn_destruct_onehotd = 4'd1;
        2'd1: v1afn_destruct_onehotd = 4'd2;
        2'd2: v1afn_destruct_onehotd = 4'd4;
        2'd3: v1afn_destruct_onehotd = 4'd8;
        default: v1afn_destruct_onehotd = 4'd0;
      endcase
    else v1afn_destruct_onehotd = 4'd0;
  assign _9_d = {v1afn_destruct_d[32:1], v1afn_destruct_onehotd[0]};
  assign lizzieLet6_5QVal_Int_8QVal_Int_d = {v1afn_destruct_d[32:1],
                                             v1afn_destruct_onehotd[1]};
  assign _8_d = {v1afn_destruct_d[32:1], v1afn_destruct_onehotd[2]};
  assign _7_d = {v1afn_destruct_d[32:1], v1afn_destruct_onehotd[3]};
  assign v1afn_destruct_r = (| (v1afn_destruct_onehotd & {_7_r,
                                                          _8_r,
                                                          lizzieLet6_5QVal_Int_8QVal_Int_r,
                                                          _9_r}));
  assign lizzieLet6_5QVal_Int_8_r = v1afn_destruct_r;
  
  /* fork (Ty Int) : (lizzieLet6_5QVal_Int_8QVal_Int,Int) > [(lizzieLet6_5QVal_Int_8QVal_Int_1,Int),
                                                        (lizzieLet6_5QVal_Int_8QVal_Int_2,Int)] */
  logic [1:0] lizzieLet6_5QVal_Int_8QVal_Int_emitted;
  logic [1:0] lizzieLet6_5QVal_Int_8QVal_Int_done;
  assign lizzieLet6_5QVal_Int_8QVal_Int_1_d = {lizzieLet6_5QVal_Int_8QVal_Int_d[32:1],
                                               (lizzieLet6_5QVal_Int_8QVal_Int_d[0] && (! lizzieLet6_5QVal_Int_8QVal_Int_emitted[0]))};
  assign lizzieLet6_5QVal_Int_8QVal_Int_2_d = {lizzieLet6_5QVal_Int_8QVal_Int_d[32:1],
                                               (lizzieLet6_5QVal_Int_8QVal_Int_d[0] && (! lizzieLet6_5QVal_Int_8QVal_Int_emitted[1]))};
  assign lizzieLet6_5QVal_Int_8QVal_Int_done = (lizzieLet6_5QVal_Int_8QVal_Int_emitted | ({lizzieLet6_5QVal_Int_8QVal_Int_2_d[0],
                                                                                           lizzieLet6_5QVal_Int_8QVal_Int_1_d[0]} & {lizzieLet6_5QVal_Int_8QVal_Int_2_r,
                                                                                                                                     lizzieLet6_5QVal_Int_8QVal_Int_1_r}));
  assign lizzieLet6_5QVal_Int_8QVal_Int_r = (& lizzieLet6_5QVal_Int_8QVal_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_5QVal_Int_8QVal_Int_emitted <= 2'd0;
    else
      lizzieLet6_5QVal_Int_8QVal_Int_emitted <= (lizzieLet6_5QVal_Int_8QVal_Int_r ? 2'd0 :
                                                 lizzieLet6_5QVal_Int_8QVal_Int_done);
  
  /* buf (Ty Int) : (lizzieLet6_5QVal_Int_8QVal_Int_1,Int) > (lizzieLet6_5QVal_Int_8QVal_Int_1_argbuf,Int) */
  Int_t lizzieLet6_5QVal_Int_8QVal_Int_1_bufchan_d;
  logic lizzieLet6_5QVal_Int_8QVal_Int_1_bufchan_r;
  assign lizzieLet6_5QVal_Int_8QVal_Int_1_r = ((! lizzieLet6_5QVal_Int_8QVal_Int_1_bufchan_d[0]) || lizzieLet6_5QVal_Int_8QVal_Int_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_5QVal_Int_8QVal_Int_1_bufchan_d <= {32'd0, 1'd0};
    else
      if (lizzieLet6_5QVal_Int_8QVal_Int_1_r)
        lizzieLet6_5QVal_Int_8QVal_Int_1_bufchan_d <= lizzieLet6_5QVal_Int_8QVal_Int_1_d;
  Int_t lizzieLet6_5QVal_Int_8QVal_Int_1_bufchan_buf;
  assign lizzieLet6_5QVal_Int_8QVal_Int_1_bufchan_r = (! lizzieLet6_5QVal_Int_8QVal_Int_1_bufchan_buf[0]);
  assign lizzieLet6_5QVal_Int_8QVal_Int_1_argbuf_d = (lizzieLet6_5QVal_Int_8QVal_Int_1_bufchan_buf[0] ? lizzieLet6_5QVal_Int_8QVal_Int_1_bufchan_buf :
                                                      lizzieLet6_5QVal_Int_8QVal_Int_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_5QVal_Int_8QVal_Int_1_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((lizzieLet6_5QVal_Int_8QVal_Int_1_argbuf_r && lizzieLet6_5QVal_Int_8QVal_Int_1_bufchan_buf[0]))
        lizzieLet6_5QVal_Int_8QVal_Int_1_bufchan_buf <= {32'd0, 1'd0};
      else if (((! lizzieLet6_5QVal_Int_8QVal_Int_1_argbuf_r) && (! lizzieLet6_5QVal_Int_8QVal_Int_1_bufchan_buf[0])))
        lizzieLet6_5QVal_Int_8QVal_Int_1_bufchan_buf <= lizzieLet6_5QVal_Int_8QVal_Int_1_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty MyDTInt_Int_Int) : (lizzieLet6_6,QTree_Int) (op_addafm_goMux_mux,MyDTInt_Int_Int) > [(_6,MyDTInt_Int_Int),
                                                                                               (lizzieLet6_6QVal_Int,MyDTInt_Int_Int),
                                                                                               (lizzieLet6_6QNode_Int,MyDTInt_Int_Int),
                                                                                               (_5,MyDTInt_Int_Int)] */
  logic [3:0] op_addafm_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet6_6_d[0] && op_addafm_goMux_mux_d[0]))
      unique case (lizzieLet6_6_d[2:1])
        2'd0: op_addafm_goMux_mux_onehotd = 4'd1;
        2'd1: op_addafm_goMux_mux_onehotd = 4'd2;
        2'd2: op_addafm_goMux_mux_onehotd = 4'd4;
        2'd3: op_addafm_goMux_mux_onehotd = 4'd8;
        default: op_addafm_goMux_mux_onehotd = 4'd0;
      endcase
    else op_addafm_goMux_mux_onehotd = 4'd0;
  assign _6_d = op_addafm_goMux_mux_onehotd[0];
  assign lizzieLet6_6QVal_Int_d = op_addafm_goMux_mux_onehotd[1];
  assign lizzieLet6_6QNode_Int_d = op_addafm_goMux_mux_onehotd[2];
  assign _5_d = op_addafm_goMux_mux_onehotd[3];
  assign op_addafm_goMux_mux_r = (| (op_addafm_goMux_mux_onehotd & {_5_r,
                                                                    lizzieLet6_6QNode_Int_r,
                                                                    lizzieLet6_6QVal_Int_r,
                                                                    _6_r}));
  assign lizzieLet6_6_r = op_addafm_goMux_mux_r;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_QTree_Int) : (lizzieLet6_7,QTree_Int) (q4afj_2,Pointer_QTree_Int) > [(_4,Pointer_QTree_Int),
                                                                                       (lizzieLet6_7QVal_Int,Pointer_QTree_Int),
                                                                                       (lizzieLet6_7QNode_Int,Pointer_QTree_Int),
                                                                                       (_3,Pointer_QTree_Int)] */
  logic [3:0] q4afj_2_onehotd;
  always_comb
    if ((lizzieLet6_7_d[0] && q4afj_2_d[0]))
      unique case (lizzieLet6_7_d[2:1])
        2'd0: q4afj_2_onehotd = 4'd1;
        2'd1: q4afj_2_onehotd = 4'd2;
        2'd2: q4afj_2_onehotd = 4'd4;
        2'd3: q4afj_2_onehotd = 4'd8;
        default: q4afj_2_onehotd = 4'd0;
      endcase
    else q4afj_2_onehotd = 4'd0;
  assign _4_d = {q4afj_2_d[16:1], q4afj_2_onehotd[0]};
  assign lizzieLet6_7QVal_Int_d = {q4afj_2_d[16:1],
                                   q4afj_2_onehotd[1]};
  assign lizzieLet6_7QNode_Int_d = {q4afj_2_d[16:1],
                                    q4afj_2_onehotd[2]};
  assign _3_d = {q4afj_2_d[16:1], q4afj_2_onehotd[3]};
  assign q4afj_2_r = (| (q4afj_2_onehotd & {_3_r,
                                            lizzieLet6_7QNode_Int_r,
                                            lizzieLet6_7QVal_Int_r,
                                            _4_r}));
  assign lizzieLet6_7_r = q4afj_2_r;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_CTf''''''''''''_f''''''''''''_Int) : (lizzieLet6_8,QTree_Int) (sc_0_1_goMux_mux,Pointer_CTf''''''''''''_f''''''''''''_Int) > [(lizzieLet6_8QNone_Int,Pointer_CTf''''''''''''_f''''''''''''_Int),
                                                                                                                                                (lizzieLet6_8QVal_Int,Pointer_CTf''''''''''''_f''''''''''''_Int),
                                                                                                                                                (lizzieLet6_8QNode_Int,Pointer_CTf''''''''''''_f''''''''''''_Int),
                                                                                                                                                (lizzieLet6_8QError_Int,Pointer_CTf''''''''''''_f''''''''''''_Int)] */
  logic [3:0] sc_0_1_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet6_8_d[0] && sc_0_1_goMux_mux_d[0]))
      unique case (lizzieLet6_8_d[2:1])
        2'd0: sc_0_1_goMux_mux_onehotd = 4'd1;
        2'd1: sc_0_1_goMux_mux_onehotd = 4'd2;
        2'd2: sc_0_1_goMux_mux_onehotd = 4'd4;
        2'd3: sc_0_1_goMux_mux_onehotd = 4'd8;
        default: sc_0_1_goMux_mux_onehotd = 4'd0;
      endcase
    else sc_0_1_goMux_mux_onehotd = 4'd0;
  assign lizzieLet6_8QNone_Int_d = {sc_0_1_goMux_mux_d[16:1],
                                    sc_0_1_goMux_mux_onehotd[0]};
  assign lizzieLet6_8QVal_Int_d = {sc_0_1_goMux_mux_d[16:1],
                                   sc_0_1_goMux_mux_onehotd[1]};
  assign lizzieLet6_8QNode_Int_d = {sc_0_1_goMux_mux_d[16:1],
                                    sc_0_1_goMux_mux_onehotd[2]};
  assign lizzieLet6_8QError_Int_d = {sc_0_1_goMux_mux_d[16:1],
                                     sc_0_1_goMux_mux_onehotd[3]};
  assign sc_0_1_goMux_mux_r = (| (sc_0_1_goMux_mux_onehotd & {lizzieLet6_8QError_Int_r,
                                                              lizzieLet6_8QNode_Int_r,
                                                              lizzieLet6_8QVal_Int_r,
                                                              lizzieLet6_8QNone_Int_r}));
  assign lizzieLet6_8_r = sc_0_1_goMux_mux_r;
  
  /* buf (Ty Pointer_CTf''''''''''''_f''''''''''''_Int) : (lizzieLet6_8QError_Int,Pointer_CTf''''''''''''_f''''''''''''_Int) > (lizzieLet6_8QError_Int_1_argbuf,Pointer_CTf''''''''''''_f''''''''''''_Int) */
  \Pointer_CTf''''''''''''_f''''''''''''_Int_t  lizzieLet6_8QError_Int_bufchan_d;
  logic lizzieLet6_8QError_Int_bufchan_r;
  assign lizzieLet6_8QError_Int_r = ((! lizzieLet6_8QError_Int_bufchan_d[0]) || lizzieLet6_8QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_8QError_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet6_8QError_Int_r)
        lizzieLet6_8QError_Int_bufchan_d <= lizzieLet6_8QError_Int_d;
  \Pointer_CTf''''''''''''_f''''''''''''_Int_t  lizzieLet6_8QError_Int_bufchan_buf;
  assign lizzieLet6_8QError_Int_bufchan_r = (! lizzieLet6_8QError_Int_bufchan_buf[0]);
  assign lizzieLet6_8QError_Int_1_argbuf_d = (lizzieLet6_8QError_Int_bufchan_buf[0] ? lizzieLet6_8QError_Int_bufchan_buf :
                                              lizzieLet6_8QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_8QError_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet6_8QError_Int_1_argbuf_r && lizzieLet6_8QError_Int_bufchan_buf[0]))
        lizzieLet6_8QError_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet6_8QError_Int_1_argbuf_r) && (! lizzieLet6_8QError_Int_bufchan_buf[0])))
        lizzieLet6_8QError_Int_bufchan_buf <= lizzieLet6_8QError_Int_bufchan_d;
  
  /* buf (Ty Pointer_CTf''''''''''''_f''''''''''''_Int) : (lizzieLet6_8QNone_Int,Pointer_CTf''''''''''''_f''''''''''''_Int) > (lizzieLet6_8QNone_Int_1_argbuf,Pointer_CTf''''''''''''_f''''''''''''_Int) */
  \Pointer_CTf''''''''''''_f''''''''''''_Int_t  lizzieLet6_8QNone_Int_bufchan_d;
  logic lizzieLet6_8QNone_Int_bufchan_r;
  assign lizzieLet6_8QNone_Int_r = ((! lizzieLet6_8QNone_Int_bufchan_d[0]) || lizzieLet6_8QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_8QNone_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet6_8QNone_Int_r)
        lizzieLet6_8QNone_Int_bufchan_d <= lizzieLet6_8QNone_Int_d;
  \Pointer_CTf''''''''''''_f''''''''''''_Int_t  lizzieLet6_8QNone_Int_bufchan_buf;
  assign lizzieLet6_8QNone_Int_bufchan_r = (! lizzieLet6_8QNone_Int_bufchan_buf[0]);
  assign lizzieLet6_8QNone_Int_1_argbuf_d = (lizzieLet6_8QNone_Int_bufchan_buf[0] ? lizzieLet6_8QNone_Int_bufchan_buf :
                                             lizzieLet6_8QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_8QNone_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet6_8QNone_Int_1_argbuf_r && lizzieLet6_8QNone_Int_bufchan_buf[0]))
        lizzieLet6_8QNone_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet6_8QNone_Int_1_argbuf_r) && (! lizzieLet6_8QNone_Int_bufchan_buf[0])))
        lizzieLet6_8QNone_Int_bufchan_buf <= lizzieLet6_8QNone_Int_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_QTree_Int) : (lizzieLet6_9,QTree_Int) (t4afk_2,Pointer_QTree_Int) > [(lizzieLet6_9QNone_Int,Pointer_QTree_Int),
                                                                                       (_2,Pointer_QTree_Int),
                                                                                       (_1,Pointer_QTree_Int),
                                                                                       (_0,Pointer_QTree_Int)] */
  logic [3:0] t4afk_2_onehotd;
  always_comb
    if ((lizzieLet6_9_d[0] && t4afk_2_d[0]))
      unique case (lizzieLet6_9_d[2:1])
        2'd0: t4afk_2_onehotd = 4'd1;
        2'd1: t4afk_2_onehotd = 4'd2;
        2'd2: t4afk_2_onehotd = 4'd4;
        2'd3: t4afk_2_onehotd = 4'd8;
        default: t4afk_2_onehotd = 4'd0;
      endcase
    else t4afk_2_onehotd = 4'd0;
  assign lizzieLet6_9QNone_Int_d = {t4afk_2_d[16:1],
                                    t4afk_2_onehotd[0]};
  assign _2_d = {t4afk_2_d[16:1], t4afk_2_onehotd[1]};
  assign _1_d = {t4afk_2_d[16:1], t4afk_2_onehotd[2]};
  assign _0_d = {t4afk_2_d[16:1], t4afk_2_onehotd[3]};
  assign t4afk_2_r = (| (t4afk_2_onehotd & {_0_r,
                                            _1_r,
                                            _2_r,
                                            lizzieLet6_9QNone_Int_r}));
  assign lizzieLet6_9_r = t4afk_2_r;
  
  /* buf (Ty Pointer_QTree_Int) : (lizzieLet6_9QNone_Int,Pointer_QTree_Int) > (lizzieLet6_9QNone_Int_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t lizzieLet6_9QNone_Int_bufchan_d;
  logic lizzieLet6_9QNone_Int_bufchan_r;
  assign lizzieLet6_9QNone_Int_r = ((! lizzieLet6_9QNone_Int_bufchan_d[0]) || lizzieLet6_9QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_9QNone_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet6_9QNone_Int_r)
        lizzieLet6_9QNone_Int_bufchan_d <= lizzieLet6_9QNone_Int_d;
  Pointer_QTree_Int_t lizzieLet6_9QNone_Int_bufchan_buf;
  assign lizzieLet6_9QNone_Int_bufchan_r = (! lizzieLet6_9QNone_Int_bufchan_buf[0]);
  assign lizzieLet6_9QNone_Int_1_argbuf_d = (lizzieLet6_9QNone_Int_bufchan_buf[0] ? lizzieLet6_9QNone_Int_bufchan_buf :
                                             lizzieLet6_9QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_9QNone_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet6_9QNone_Int_1_argbuf_r && lizzieLet6_9QNone_Int_bufchan_buf[0]))
        lizzieLet6_9QNone_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet6_9QNone_Int_1_argbuf_r) && (! lizzieLet6_9QNone_Int_bufchan_buf[0])))
        lizzieLet6_9QNone_Int_bufchan_buf <= lizzieLet6_9QNone_Int_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (m1aeq_1,Pointer_QTree_Int) > (m1aeq_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t m1aeq_1_bufchan_d;
  logic m1aeq_1_bufchan_r;
  assign m1aeq_1_r = ((! m1aeq_1_bufchan_d[0]) || m1aeq_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m1aeq_1_bufchan_d <= {16'd0, 1'd0};
    else if (m1aeq_1_r) m1aeq_1_bufchan_d <= m1aeq_1_d;
  Pointer_QTree_Int_t m1aeq_1_bufchan_buf;
  assign m1aeq_1_bufchan_r = (! m1aeq_1_bufchan_buf[0]);
  assign m1aeq_1_argbuf_d = (m1aeq_1_bufchan_buf[0] ? m1aeq_1_bufchan_buf :
                             m1aeq_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m1aeq_1_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((m1aeq_1_argbuf_r && m1aeq_1_bufchan_buf[0]))
        m1aeq_1_bufchan_buf <= {16'd0, 1'd0};
      else if (((! m1aeq_1_argbuf_r) && (! m1aeq_1_bufchan_buf[0])))
        m1aeq_1_bufchan_buf <= m1aeq_1_bufchan_d;
  
  /* fork (Ty Pointer_QTree_Int) : (m1aeq_goMux_mux,Pointer_QTree_Int) > [(m1aeq_1,Pointer_QTree_Int),
                                                                     (m1aeq_2,Pointer_QTree_Int)] */
  logic [1:0] m1aeq_goMux_mux_emitted;
  logic [1:0] m1aeq_goMux_mux_done;
  assign m1aeq_1_d = {m1aeq_goMux_mux_d[16:1],
                      (m1aeq_goMux_mux_d[0] && (! m1aeq_goMux_mux_emitted[0]))};
  assign m1aeq_2_d = {m1aeq_goMux_mux_d[16:1],
                      (m1aeq_goMux_mux_d[0] && (! m1aeq_goMux_mux_emitted[1]))};
  assign m1aeq_goMux_mux_done = (m1aeq_goMux_mux_emitted | ({m1aeq_2_d[0],
                                                             m1aeq_1_d[0]} & {m1aeq_2_r,
                                                                              m1aeq_1_r}));
  assign m1aeq_goMux_mux_r = (& m1aeq_goMux_mux_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m1aeq_goMux_mux_emitted <= 2'd0;
    else
      m1aeq_goMux_mux_emitted <= (m1aeq_goMux_mux_r ? 2'd0 :
                                  m1aeq_goMux_mux_done);
  
  /* buf (Ty Pointer_QTree_Int) : (m2aer_1,Pointer_QTree_Int) > (m2aer_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t m2aer_1_bufchan_d;
  logic m2aer_1_bufchan_r;
  assign m2aer_1_r = ((! m2aer_1_bufchan_d[0]) || m2aer_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m2aer_1_bufchan_d <= {16'd0, 1'd0};
    else if (m2aer_1_r) m2aer_1_bufchan_d <= m2aer_1_d;
  Pointer_QTree_Int_t m2aer_1_bufchan_buf;
  assign m2aer_1_bufchan_r = (! m2aer_1_bufchan_buf[0]);
  assign m2aer_1_argbuf_d = (m2aer_1_bufchan_buf[0] ? m2aer_1_bufchan_buf :
                             m2aer_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m2aer_1_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((m2aer_1_argbuf_r && m2aer_1_bufchan_buf[0]))
        m2aer_1_bufchan_buf <= {16'd0, 1'd0};
      else if (((! m2aer_1_argbuf_r) && (! m2aer_1_bufchan_buf[0])))
        m2aer_1_bufchan_buf <= m2aer_1_bufchan_d;
  
  /* fork (Ty Pointer_QTree_Int) : (m2aer_goMux_mux,Pointer_QTree_Int) > [(m2aer_1,Pointer_QTree_Int),
                                                                     (m2aer_2,Pointer_QTree_Int)] */
  logic [1:0] m2aer_goMux_mux_emitted;
  logic [1:0] m2aer_goMux_mux_done;
  assign m2aer_1_d = {m2aer_goMux_mux_d[16:1],
                      (m2aer_goMux_mux_d[0] && (! m2aer_goMux_mux_emitted[0]))};
  assign m2aer_2_d = {m2aer_goMux_mux_d[16:1],
                      (m2aer_goMux_mux_d[0] && (! m2aer_goMux_mux_emitted[1]))};
  assign m2aer_goMux_mux_done = (m2aer_goMux_mux_emitted | ({m2aer_2_d[0],
                                                             m2aer_1_d[0]} & {m2aer_2_r,
                                                                              m2aer_1_r}));
  assign m2aer_goMux_mux_r = (& m2aer_goMux_mux_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m2aer_goMux_mux_emitted <= 2'd0;
    else
      m2aer_goMux_mux_emitted <= (m2aer_goMux_mux_r ? 2'd0 :
                                  m2aer_goMux_mux_done);
  
  /* buf (Ty Pointer_QTree_Int) : (m3aes_1,Pointer_QTree_Int) > (m3aes_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t m3aes_1_bufchan_d;
  logic m3aes_1_bufchan_r;
  assign m3aes_1_r = ((! m3aes_1_bufchan_d[0]) || m3aes_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m3aes_1_bufchan_d <= {16'd0, 1'd0};
    else if (m3aes_1_r) m3aes_1_bufchan_d <= m3aes_1_d;
  Pointer_QTree_Int_t m3aes_1_bufchan_buf;
  assign m3aes_1_bufchan_r = (! m3aes_1_bufchan_buf[0]);
  assign m3aes_1_argbuf_d = (m3aes_1_bufchan_buf[0] ? m3aes_1_bufchan_buf :
                             m3aes_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m3aes_1_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((m3aes_1_argbuf_r && m3aes_1_bufchan_buf[0]))
        m3aes_1_bufchan_buf <= {16'd0, 1'd0};
      else if (((! m3aes_1_argbuf_r) && (! m3aes_1_bufchan_buf[0])))
        m3aes_1_bufchan_buf <= m3aes_1_bufchan_d;
  
  /* fork (Ty Pointer_QTree_Int) : (m3aes_goMux_mux,Pointer_QTree_Int) > [(m3aes_1,Pointer_QTree_Int),
                                                                     (m3aes_2,Pointer_QTree_Int)] */
  logic [1:0] m3aes_goMux_mux_emitted;
  logic [1:0] m3aes_goMux_mux_done;
  assign m3aes_1_d = {m3aes_goMux_mux_d[16:1],
                      (m3aes_goMux_mux_d[0] && (! m3aes_goMux_mux_emitted[0]))};
  assign m3aes_2_d = {m3aes_goMux_mux_d[16:1],
                      (m3aes_goMux_mux_d[0] && (! m3aes_goMux_mux_emitted[1]))};
  assign m3aes_goMux_mux_done = (m3aes_goMux_mux_emitted | ({m3aes_2_d[0],
                                                             m3aes_1_d[0]} & {m3aes_2_r,
                                                                              m3aes_1_r}));
  assign m3aes_goMux_mux_r = (& m3aes_goMux_mux_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m3aes_goMux_mux_emitted <= 2'd0;
    else
      m3aes_goMux_mux_emitted <= (m3aes_goMux_mux_r ? 2'd0 :
                                  m3aes_goMux_mux_done);
  
  /* buf (Ty MyDTInt_Int_Int) : (op_addaeu_2_2,MyDTInt_Int_Int) > (op_addaeu_2_2_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t op_addaeu_2_2_bufchan_d;
  logic op_addaeu_2_2_bufchan_r;
  assign op_addaeu_2_2_r = ((! op_addaeu_2_2_bufchan_d[0]) || op_addaeu_2_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) op_addaeu_2_2_bufchan_d <= 1'd0;
    else
      if (op_addaeu_2_2_r) op_addaeu_2_2_bufchan_d <= op_addaeu_2_2_d;
  MyDTInt_Int_Int_t op_addaeu_2_2_bufchan_buf;
  assign op_addaeu_2_2_bufchan_r = (! op_addaeu_2_2_bufchan_buf[0]);
  assign op_addaeu_2_2_argbuf_d = (op_addaeu_2_2_bufchan_buf[0] ? op_addaeu_2_2_bufchan_buf :
                                   op_addaeu_2_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) op_addaeu_2_2_bufchan_buf <= 1'd0;
    else
      if ((op_addaeu_2_2_argbuf_r && op_addaeu_2_2_bufchan_buf[0]))
        op_addaeu_2_2_bufchan_buf <= 1'd0;
      else if (((! op_addaeu_2_2_argbuf_r) && (! op_addaeu_2_2_bufchan_buf[0])))
        op_addaeu_2_2_bufchan_buf <= op_addaeu_2_2_bufchan_d;
  
  /* fork (Ty MyDTInt_Int_Int) : (op_addaeu_2_destruct,MyDTInt_Int_Int) > [(op_addaeu_2_1,MyDTInt_Int_Int),
                                                                      (op_addaeu_2_2,MyDTInt_Int_Int)] */
  logic [1:0] op_addaeu_2_destruct_emitted;
  logic [1:0] op_addaeu_2_destruct_done;
  assign op_addaeu_2_1_d = (op_addaeu_2_destruct_d[0] && (! op_addaeu_2_destruct_emitted[0]));
  assign op_addaeu_2_2_d = (op_addaeu_2_destruct_d[0] && (! op_addaeu_2_destruct_emitted[1]));
  assign op_addaeu_2_destruct_done = (op_addaeu_2_destruct_emitted | ({op_addaeu_2_2_d[0],
                                                                       op_addaeu_2_1_d[0]} & {op_addaeu_2_2_r,
                                                                                              op_addaeu_2_1_r}));
  assign op_addaeu_2_destruct_r = (& op_addaeu_2_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) op_addaeu_2_destruct_emitted <= 2'd0;
    else
      op_addaeu_2_destruct_emitted <= (op_addaeu_2_destruct_r ? 2'd0 :
                                       op_addaeu_2_destruct_done);
  
  /* buf (Ty MyDTInt_Int_Int) : (op_addaeu_3_2,MyDTInt_Int_Int) > (op_addaeu_3_2_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t op_addaeu_3_2_bufchan_d;
  logic op_addaeu_3_2_bufchan_r;
  assign op_addaeu_3_2_r = ((! op_addaeu_3_2_bufchan_d[0]) || op_addaeu_3_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) op_addaeu_3_2_bufchan_d <= 1'd0;
    else
      if (op_addaeu_3_2_r) op_addaeu_3_2_bufchan_d <= op_addaeu_3_2_d;
  MyDTInt_Int_Int_t op_addaeu_3_2_bufchan_buf;
  assign op_addaeu_3_2_bufchan_r = (! op_addaeu_3_2_bufchan_buf[0]);
  assign op_addaeu_3_2_argbuf_d = (op_addaeu_3_2_bufchan_buf[0] ? op_addaeu_3_2_bufchan_buf :
                                   op_addaeu_3_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) op_addaeu_3_2_bufchan_buf <= 1'd0;
    else
      if ((op_addaeu_3_2_argbuf_r && op_addaeu_3_2_bufchan_buf[0]))
        op_addaeu_3_2_bufchan_buf <= 1'd0;
      else if (((! op_addaeu_3_2_argbuf_r) && (! op_addaeu_3_2_bufchan_buf[0])))
        op_addaeu_3_2_bufchan_buf <= op_addaeu_3_2_bufchan_d;
  
  /* fork (Ty MyDTInt_Int_Int) : (op_addaeu_3_destruct,MyDTInt_Int_Int) > [(op_addaeu_3_1,MyDTInt_Int_Int),
                                                                      (op_addaeu_3_2,MyDTInt_Int_Int)] */
  logic [1:0] op_addaeu_3_destruct_emitted;
  logic [1:0] op_addaeu_3_destruct_done;
  assign op_addaeu_3_1_d = (op_addaeu_3_destruct_d[0] && (! op_addaeu_3_destruct_emitted[0]));
  assign op_addaeu_3_2_d = (op_addaeu_3_destruct_d[0] && (! op_addaeu_3_destruct_emitted[1]));
  assign op_addaeu_3_destruct_done = (op_addaeu_3_destruct_emitted | ({op_addaeu_3_2_d[0],
                                                                       op_addaeu_3_1_d[0]} & {op_addaeu_3_2_r,
                                                                                              op_addaeu_3_1_r}));
  assign op_addaeu_3_destruct_r = (& op_addaeu_3_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) op_addaeu_3_destruct_emitted <= 2'd0;
    else
      op_addaeu_3_destruct_emitted <= (op_addaeu_3_destruct_r ? 2'd0 :
                                       op_addaeu_3_destruct_done);
  
  /* buf (Ty MyDTInt_Int_Int) : (op_addaeu_4_destruct,MyDTInt_Int_Int) > (op_addaeu_4_1_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t op_addaeu_4_destruct_bufchan_d;
  logic op_addaeu_4_destruct_bufchan_r;
  assign op_addaeu_4_destruct_r = ((! op_addaeu_4_destruct_bufchan_d[0]) || op_addaeu_4_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) op_addaeu_4_destruct_bufchan_d <= 1'd0;
    else
      if (op_addaeu_4_destruct_r)
        op_addaeu_4_destruct_bufchan_d <= op_addaeu_4_destruct_d;
  MyDTInt_Int_Int_t op_addaeu_4_destruct_bufchan_buf;
  assign op_addaeu_4_destruct_bufchan_r = (! op_addaeu_4_destruct_bufchan_buf[0]);
  assign op_addaeu_4_1_argbuf_d = (op_addaeu_4_destruct_bufchan_buf[0] ? op_addaeu_4_destruct_bufchan_buf :
                                   op_addaeu_4_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) op_addaeu_4_destruct_bufchan_buf <= 1'd0;
    else
      if ((op_addaeu_4_1_argbuf_r && op_addaeu_4_destruct_bufchan_buf[0]))
        op_addaeu_4_destruct_bufchan_buf <= 1'd0;
      else if (((! op_addaeu_4_1_argbuf_r) && (! op_addaeu_4_destruct_bufchan_buf[0])))
        op_addaeu_4_destruct_bufchan_buf <= op_addaeu_4_destruct_bufchan_d;
  
  /* buf (Ty MyDTInt_Int_Int) : (op_addafm_2_2,MyDTInt_Int_Int) > (op_addafm_2_2_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t op_addafm_2_2_bufchan_d;
  logic op_addafm_2_2_bufchan_r;
  assign op_addafm_2_2_r = ((! op_addafm_2_2_bufchan_d[0]) || op_addafm_2_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) op_addafm_2_2_bufchan_d <= 1'd0;
    else
      if (op_addafm_2_2_r) op_addafm_2_2_bufchan_d <= op_addafm_2_2_d;
  MyDTInt_Int_Int_t op_addafm_2_2_bufchan_buf;
  assign op_addafm_2_2_bufchan_r = (! op_addafm_2_2_bufchan_buf[0]);
  assign op_addafm_2_2_argbuf_d = (op_addafm_2_2_bufchan_buf[0] ? op_addafm_2_2_bufchan_buf :
                                   op_addafm_2_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) op_addafm_2_2_bufchan_buf <= 1'd0;
    else
      if ((op_addafm_2_2_argbuf_r && op_addafm_2_2_bufchan_buf[0]))
        op_addafm_2_2_bufchan_buf <= 1'd0;
      else if (((! op_addafm_2_2_argbuf_r) && (! op_addafm_2_2_bufchan_buf[0])))
        op_addafm_2_2_bufchan_buf <= op_addafm_2_2_bufchan_d;
  
  /* fork (Ty MyDTInt_Int_Int) : (op_addafm_2_destruct,MyDTInt_Int_Int) > [(op_addafm_2_1,MyDTInt_Int_Int),
                                                                      (op_addafm_2_2,MyDTInt_Int_Int)] */
  logic [1:0] op_addafm_2_destruct_emitted;
  logic [1:0] op_addafm_2_destruct_done;
  assign op_addafm_2_1_d = (op_addafm_2_destruct_d[0] && (! op_addafm_2_destruct_emitted[0]));
  assign op_addafm_2_2_d = (op_addafm_2_destruct_d[0] && (! op_addafm_2_destruct_emitted[1]));
  assign op_addafm_2_destruct_done = (op_addafm_2_destruct_emitted | ({op_addafm_2_2_d[0],
                                                                       op_addafm_2_1_d[0]} & {op_addafm_2_2_r,
                                                                                              op_addafm_2_1_r}));
  assign op_addafm_2_destruct_r = (& op_addafm_2_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) op_addafm_2_destruct_emitted <= 2'd0;
    else
      op_addafm_2_destruct_emitted <= (op_addafm_2_destruct_r ? 2'd0 :
                                       op_addafm_2_destruct_done);
  
  /* buf (Ty MyDTInt_Int_Int) : (op_addafm_3_2,MyDTInt_Int_Int) > (op_addafm_3_2_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t op_addafm_3_2_bufchan_d;
  logic op_addafm_3_2_bufchan_r;
  assign op_addafm_3_2_r = ((! op_addafm_3_2_bufchan_d[0]) || op_addafm_3_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) op_addafm_3_2_bufchan_d <= 1'd0;
    else
      if (op_addafm_3_2_r) op_addafm_3_2_bufchan_d <= op_addafm_3_2_d;
  MyDTInt_Int_Int_t op_addafm_3_2_bufchan_buf;
  assign op_addafm_3_2_bufchan_r = (! op_addafm_3_2_bufchan_buf[0]);
  assign op_addafm_3_2_argbuf_d = (op_addafm_3_2_bufchan_buf[0] ? op_addafm_3_2_bufchan_buf :
                                   op_addafm_3_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) op_addafm_3_2_bufchan_buf <= 1'd0;
    else
      if ((op_addafm_3_2_argbuf_r && op_addafm_3_2_bufchan_buf[0]))
        op_addafm_3_2_bufchan_buf <= 1'd0;
      else if (((! op_addafm_3_2_argbuf_r) && (! op_addafm_3_2_bufchan_buf[0])))
        op_addafm_3_2_bufchan_buf <= op_addafm_3_2_bufchan_d;
  
  /* fork (Ty MyDTInt_Int_Int) : (op_addafm_3_destruct,MyDTInt_Int_Int) > [(op_addafm_3_1,MyDTInt_Int_Int),
                                                                      (op_addafm_3_2,MyDTInt_Int_Int)] */
  logic [1:0] op_addafm_3_destruct_emitted;
  logic [1:0] op_addafm_3_destruct_done;
  assign op_addafm_3_1_d = (op_addafm_3_destruct_d[0] && (! op_addafm_3_destruct_emitted[0]));
  assign op_addafm_3_2_d = (op_addafm_3_destruct_d[0] && (! op_addafm_3_destruct_emitted[1]));
  assign op_addafm_3_destruct_done = (op_addafm_3_destruct_emitted | ({op_addafm_3_2_d[0],
                                                                       op_addafm_3_1_d[0]} & {op_addafm_3_2_r,
                                                                                              op_addafm_3_1_r}));
  assign op_addafm_3_destruct_r = (& op_addafm_3_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) op_addafm_3_destruct_emitted <= 2'd0;
    else
      op_addafm_3_destruct_emitted <= (op_addafm_3_destruct_r ? 2'd0 :
                                       op_addafm_3_destruct_done);
  
  /* buf (Ty MyDTInt_Int_Int) : (op_addafm_4_destruct,MyDTInt_Int_Int) > (op_addafm_4_1_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t op_addafm_4_destruct_bufchan_d;
  logic op_addafm_4_destruct_bufchan_r;
  assign op_addafm_4_destruct_r = ((! op_addafm_4_destruct_bufchan_d[0]) || op_addafm_4_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) op_addafm_4_destruct_bufchan_d <= 1'd0;
    else
      if (op_addafm_4_destruct_r)
        op_addafm_4_destruct_bufchan_d <= op_addafm_4_destruct_d;
  MyDTInt_Int_Int_t op_addafm_4_destruct_bufchan_buf;
  assign op_addafm_4_destruct_bufchan_r = (! op_addafm_4_destruct_bufchan_buf[0]);
  assign op_addafm_4_1_argbuf_d = (op_addafm_4_destruct_bufchan_buf[0] ? op_addafm_4_destruct_bufchan_buf :
                                   op_addafm_4_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) op_addafm_4_destruct_bufchan_buf <= 1'd0;
    else
      if ((op_addafm_4_1_argbuf_r && op_addafm_4_destruct_bufchan_buf[0]))
        op_addafm_4_destruct_bufchan_buf <= 1'd0;
      else if (((! op_addafm_4_1_argbuf_r) && (! op_addafm_4_destruct_bufchan_buf[0])))
        op_addafm_4_destruct_bufchan_buf <= op_addafm_4_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (q1a8r_destruct,Pointer_QTree_Int) > (q1a8r_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t q1a8r_destruct_bufchan_d;
  logic q1a8r_destruct_bufchan_r;
  assign q1a8r_destruct_r = ((! q1a8r_destruct_bufchan_d[0]) || q1a8r_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q1a8r_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q1a8r_destruct_r) q1a8r_destruct_bufchan_d <= q1a8r_destruct_d;
  Pointer_QTree_Int_t q1a8r_destruct_bufchan_buf;
  assign q1a8r_destruct_bufchan_r = (! q1a8r_destruct_bufchan_buf[0]);
  assign q1a8r_1_argbuf_d = (q1a8r_destruct_bufchan_buf[0] ? q1a8r_destruct_bufchan_buf :
                             q1a8r_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q1a8r_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q1a8r_1_argbuf_r && q1a8r_destruct_bufchan_buf[0]))
        q1a8r_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q1a8r_1_argbuf_r) && (! q1a8r_destruct_bufchan_buf[0])))
        q1a8r_destruct_bufchan_buf <= q1a8r_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (q1af0_3_destruct,Pointer_QTree_Int) > (q1af0_3_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t q1af0_3_destruct_bufchan_d;
  logic q1af0_3_destruct_bufchan_r;
  assign q1af0_3_destruct_r = ((! q1af0_3_destruct_bufchan_d[0]) || q1af0_3_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q1af0_3_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q1af0_3_destruct_r)
        q1af0_3_destruct_bufchan_d <= q1af0_3_destruct_d;
  Pointer_QTree_Int_t q1af0_3_destruct_bufchan_buf;
  assign q1af0_3_destruct_bufchan_r = (! q1af0_3_destruct_bufchan_buf[0]);
  assign q1af0_3_1_argbuf_d = (q1af0_3_destruct_bufchan_buf[0] ? q1af0_3_destruct_bufchan_buf :
                               q1af0_3_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q1af0_3_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q1af0_3_1_argbuf_r && q1af0_3_destruct_bufchan_buf[0]))
        q1af0_3_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q1af0_3_1_argbuf_r) && (! q1af0_3_destruct_bufchan_buf[0])))
        q1af0_3_destruct_bufchan_buf <= q1af0_3_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (q1aft_3_destruct,Pointer_QTree_Int) > (q1aft_3_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t q1aft_3_destruct_bufchan_d;
  logic q1aft_3_destruct_bufchan_r;
  assign q1aft_3_destruct_r = ((! q1aft_3_destruct_bufchan_d[0]) || q1aft_3_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q1aft_3_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q1aft_3_destruct_r)
        q1aft_3_destruct_bufchan_d <= q1aft_3_destruct_d;
  Pointer_QTree_Int_t q1aft_3_destruct_bufchan_buf;
  assign q1aft_3_destruct_bufchan_r = (! q1aft_3_destruct_bufchan_buf[0]);
  assign q1aft_3_1_argbuf_d = (q1aft_3_destruct_bufchan_buf[0] ? q1aft_3_destruct_bufchan_buf :
                               q1aft_3_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q1aft_3_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q1aft_3_1_argbuf_r && q1aft_3_destruct_bufchan_buf[0]))
        q1aft_3_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q1aft_3_1_argbuf_r) && (! q1aft_3_destruct_bufchan_buf[0])))
        q1aft_3_destruct_bufchan_buf <= q1aft_3_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (q2a8s_1_destruct,Pointer_QTree_Int) > (q2a8s_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t q2a8s_1_destruct_bufchan_d;
  logic q2a8s_1_destruct_bufchan_r;
  assign q2a8s_1_destruct_r = ((! q2a8s_1_destruct_bufchan_d[0]) || q2a8s_1_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q2a8s_1_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q2a8s_1_destruct_r)
        q2a8s_1_destruct_bufchan_d <= q2a8s_1_destruct_d;
  Pointer_QTree_Int_t q2a8s_1_destruct_bufchan_buf;
  assign q2a8s_1_destruct_bufchan_r = (! q2a8s_1_destruct_bufchan_buf[0]);
  assign q2a8s_1_1_argbuf_d = (q2a8s_1_destruct_bufchan_buf[0] ? q2a8s_1_destruct_bufchan_buf :
                               q2a8s_1_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q2a8s_1_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q2a8s_1_1_argbuf_r && q2a8s_1_destruct_bufchan_buf[0]))
        q2a8s_1_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q2a8s_1_1_argbuf_r) && (! q2a8s_1_destruct_bufchan_buf[0])))
        q2a8s_1_destruct_bufchan_buf <= q2a8s_1_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (q2af1_2_destruct,Pointer_QTree_Int) > (q2af1_2_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t q2af1_2_destruct_bufchan_d;
  logic q2af1_2_destruct_bufchan_r;
  assign q2af1_2_destruct_r = ((! q2af1_2_destruct_bufchan_d[0]) || q2af1_2_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q2af1_2_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q2af1_2_destruct_r)
        q2af1_2_destruct_bufchan_d <= q2af1_2_destruct_d;
  Pointer_QTree_Int_t q2af1_2_destruct_bufchan_buf;
  assign q2af1_2_destruct_bufchan_r = (! q2af1_2_destruct_bufchan_buf[0]);
  assign q2af1_2_1_argbuf_d = (q2af1_2_destruct_bufchan_buf[0] ? q2af1_2_destruct_bufchan_buf :
                               q2af1_2_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q2af1_2_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q2af1_2_1_argbuf_r && q2af1_2_destruct_bufchan_buf[0]))
        q2af1_2_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q2af1_2_1_argbuf_r) && (! q2af1_2_destruct_bufchan_buf[0])))
        q2af1_2_destruct_bufchan_buf <= q2af1_2_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (q2afu_2_destruct,Pointer_QTree_Int) > (q2afu_2_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t q2afu_2_destruct_bufchan_d;
  logic q2afu_2_destruct_bufchan_r;
  assign q2afu_2_destruct_r = ((! q2afu_2_destruct_bufchan_d[0]) || q2afu_2_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q2afu_2_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q2afu_2_destruct_r)
        q2afu_2_destruct_bufchan_d <= q2afu_2_destruct_d;
  Pointer_QTree_Int_t q2afu_2_destruct_bufchan_buf;
  assign q2afu_2_destruct_bufchan_r = (! q2afu_2_destruct_bufchan_buf[0]);
  assign q2afu_2_1_argbuf_d = (q2afu_2_destruct_bufchan_buf[0] ? q2afu_2_destruct_bufchan_buf :
                               q2afu_2_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q2afu_2_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q2afu_2_1_argbuf_r && q2afu_2_destruct_bufchan_buf[0]))
        q2afu_2_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q2afu_2_1_argbuf_r) && (! q2afu_2_destruct_bufchan_buf[0])))
        q2afu_2_destruct_bufchan_buf <= q2afu_2_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (q3a8t_2_destruct,Pointer_QTree_Int) > (q3a8t_2_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t q3a8t_2_destruct_bufchan_d;
  logic q3a8t_2_destruct_bufchan_r;
  assign q3a8t_2_destruct_r = ((! q3a8t_2_destruct_bufchan_d[0]) || q3a8t_2_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q3a8t_2_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q3a8t_2_destruct_r)
        q3a8t_2_destruct_bufchan_d <= q3a8t_2_destruct_d;
  Pointer_QTree_Int_t q3a8t_2_destruct_bufchan_buf;
  assign q3a8t_2_destruct_bufchan_r = (! q3a8t_2_destruct_bufchan_buf[0]);
  assign q3a8t_2_1_argbuf_d = (q3a8t_2_destruct_bufchan_buf[0] ? q3a8t_2_destruct_bufchan_buf :
                               q3a8t_2_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q3a8t_2_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q3a8t_2_1_argbuf_r && q3a8t_2_destruct_bufchan_buf[0]))
        q3a8t_2_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q3a8t_2_1_argbuf_r) && (! q3a8t_2_destruct_bufchan_buf[0])))
        q3a8t_2_destruct_bufchan_buf <= q3a8t_2_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (q3af2_1_destruct,Pointer_QTree_Int) > (q3af2_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t q3af2_1_destruct_bufchan_d;
  logic q3af2_1_destruct_bufchan_r;
  assign q3af2_1_destruct_r = ((! q3af2_1_destruct_bufchan_d[0]) || q3af2_1_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q3af2_1_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q3af2_1_destruct_r)
        q3af2_1_destruct_bufchan_d <= q3af2_1_destruct_d;
  Pointer_QTree_Int_t q3af2_1_destruct_bufchan_buf;
  assign q3af2_1_destruct_bufchan_r = (! q3af2_1_destruct_bufchan_buf[0]);
  assign q3af2_1_1_argbuf_d = (q3af2_1_destruct_bufchan_buf[0] ? q3af2_1_destruct_bufchan_buf :
                               q3af2_1_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q3af2_1_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q3af2_1_1_argbuf_r && q3af2_1_destruct_bufchan_buf[0]))
        q3af2_1_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q3af2_1_1_argbuf_r) && (! q3af2_1_destruct_bufchan_buf[0])))
        q3af2_1_destruct_bufchan_buf <= q3af2_1_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (q3afv_1_destruct,Pointer_QTree_Int) > (q3afv_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t q3afv_1_destruct_bufchan_d;
  logic q3afv_1_destruct_bufchan_r;
  assign q3afv_1_destruct_r = ((! q3afv_1_destruct_bufchan_d[0]) || q3afv_1_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q3afv_1_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q3afv_1_destruct_r)
        q3afv_1_destruct_bufchan_d <= q3afv_1_destruct_d;
  Pointer_QTree_Int_t q3afv_1_destruct_bufchan_buf;
  assign q3afv_1_destruct_bufchan_r = (! q3afv_1_destruct_bufchan_buf[0]);
  assign q3afv_1_1_argbuf_d = (q3afv_1_destruct_bufchan_buf[0] ? q3afv_1_destruct_bufchan_buf :
                               q3afv_1_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q3afv_1_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q3afv_1_1_argbuf_r && q3afv_1_destruct_bufchan_buf[0]))
        q3afv_1_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q3afv_1_1_argbuf_r) && (! q3afv_1_destruct_bufchan_buf[0])))
        q3afv_1_destruct_bufchan_buf <= q3afv_1_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (q4a8u_3_destruct,Pointer_QTree_Int) > (q4a8u_3_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t q4a8u_3_destruct_bufchan_d;
  logic q4a8u_3_destruct_bufchan_r;
  assign q4a8u_3_destruct_r = ((! q4a8u_3_destruct_bufchan_d[0]) || q4a8u_3_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q4a8u_3_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q4a8u_3_destruct_r)
        q4a8u_3_destruct_bufchan_d <= q4a8u_3_destruct_d;
  Pointer_QTree_Int_t q4a8u_3_destruct_bufchan_buf;
  assign q4a8u_3_destruct_bufchan_r = (! q4a8u_3_destruct_bufchan_buf[0]);
  assign q4a8u_3_1_argbuf_d = (q4a8u_3_destruct_bufchan_buf[0] ? q4a8u_3_destruct_bufchan_buf :
                               q4a8u_3_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q4a8u_3_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q4a8u_3_1_argbuf_r && q4a8u_3_destruct_bufchan_buf[0]))
        q4a8u_3_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q4a8u_3_1_argbuf_r) && (! q4a8u_3_destruct_bufchan_buf[0])))
        q4a8u_3_destruct_bufchan_buf <= q4a8u_3_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (q4afj_1,Pointer_QTree_Int) > (q4afj_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t q4afj_1_bufchan_d;
  logic q4afj_1_bufchan_r;
  assign q4afj_1_r = ((! q4afj_1_bufchan_d[0]) || q4afj_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q4afj_1_bufchan_d <= {16'd0, 1'd0};
    else if (q4afj_1_r) q4afj_1_bufchan_d <= q4afj_1_d;
  Pointer_QTree_Int_t q4afj_1_bufchan_buf;
  assign q4afj_1_bufchan_r = (! q4afj_1_bufchan_buf[0]);
  assign q4afj_1_argbuf_d = (q4afj_1_bufchan_buf[0] ? q4afj_1_bufchan_buf :
                             q4afj_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q4afj_1_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q4afj_1_argbuf_r && q4afj_1_bufchan_buf[0]))
        q4afj_1_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q4afj_1_argbuf_r) && (! q4afj_1_bufchan_buf[0])))
        q4afj_1_bufchan_buf <= q4afj_1_bufchan_d;
  
  /* fork (Ty Pointer_QTree_Int) : (q4afj_goMux_mux,Pointer_QTree_Int) > [(q4afj_1,Pointer_QTree_Int),
                                                                     (q4afj_2,Pointer_QTree_Int)] */
  logic [1:0] q4afj_goMux_mux_emitted;
  logic [1:0] q4afj_goMux_mux_done;
  assign q4afj_1_d = {q4afj_goMux_mux_d[16:1],
                      (q4afj_goMux_mux_d[0] && (! q4afj_goMux_mux_emitted[0]))};
  assign q4afj_2_d = {q4afj_goMux_mux_d[16:1],
                      (q4afj_goMux_mux_d[0] && (! q4afj_goMux_mux_emitted[1]))};
  assign q4afj_goMux_mux_done = (q4afj_goMux_mux_emitted | ({q4afj_2_d[0],
                                                             q4afj_1_d[0]} & {q4afj_2_r,
                                                                              q4afj_1_r}));
  assign q4afj_goMux_mux_r = (& q4afj_goMux_mux_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q4afj_goMux_mux_emitted <= 2'd0;
    else
      q4afj_goMux_mux_emitted <= (q4afj_goMux_mux_r ? 2'd0 :
                                  q4afj_goMux_mux_done);
  
  /* buf (Ty CT$wnnz) : (readPointer_CT$wnnzscfarg_0_1_argbuf,CT$wnnz) > (readPointer_CT$wnnzscfarg_0_1_argbuf_rwb,CT$wnnz) */
  CT$wnnz_t readPointer_CT$wnnzscfarg_0_1_argbuf_bufchan_d;
  logic readPointer_CT$wnnzscfarg_0_1_argbuf_bufchan_r;
  assign readPointer_CT$wnnzscfarg_0_1_argbuf_r = ((! readPointer_CT$wnnzscfarg_0_1_argbuf_bufchan_d[0]) || readPointer_CT$wnnzscfarg_0_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_CT$wnnzscfarg_0_1_argbuf_bufchan_d <= {115'd0, 1'd0};
    else
      if (readPointer_CT$wnnzscfarg_0_1_argbuf_r)
        readPointer_CT$wnnzscfarg_0_1_argbuf_bufchan_d <= readPointer_CT$wnnzscfarg_0_1_argbuf_d;
  CT$wnnz_t readPointer_CT$wnnzscfarg_0_1_argbuf_bufchan_buf;
  assign readPointer_CT$wnnzscfarg_0_1_argbuf_bufchan_r = (! readPointer_CT$wnnzscfarg_0_1_argbuf_bufchan_buf[0]);
  assign readPointer_CT$wnnzscfarg_0_1_argbuf_rwb_d = (readPointer_CT$wnnzscfarg_0_1_argbuf_bufchan_buf[0] ? readPointer_CT$wnnzscfarg_0_1_argbuf_bufchan_buf :
                                                       readPointer_CT$wnnzscfarg_0_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_CT$wnnzscfarg_0_1_argbuf_bufchan_buf <= {115'd0, 1'd0};
    else
      if ((readPointer_CT$wnnzscfarg_0_1_argbuf_rwb_r && readPointer_CT$wnnzscfarg_0_1_argbuf_bufchan_buf[0]))
        readPointer_CT$wnnzscfarg_0_1_argbuf_bufchan_buf <= {115'd0, 1'd0};
      else if (((! readPointer_CT$wnnzscfarg_0_1_argbuf_rwb_r) && (! readPointer_CT$wnnzscfarg_0_1_argbuf_bufchan_buf[0])))
        readPointer_CT$wnnzscfarg_0_1_argbuf_bufchan_buf <= readPointer_CT$wnnzscfarg_0_1_argbuf_bufchan_d;
  
  /* fork (Ty CT$wnnz) : (readPointer_CT$wnnzscfarg_0_1_argbuf_rwb,CT$wnnz) > [(lizzieLet58_1,CT$wnnz),
                                                                          (lizzieLet58_2,CT$wnnz),
                                                                          (lizzieLet58_3,CT$wnnz),
                                                                          (lizzieLet58_4,CT$wnnz)] */
  logic [3:0] readPointer_CT$wnnzscfarg_0_1_argbuf_rwb_emitted;
  logic [3:0] readPointer_CT$wnnzscfarg_0_1_argbuf_rwb_done;
  assign lizzieLet58_1_d = {readPointer_CT$wnnzscfarg_0_1_argbuf_rwb_d[115:1],
                            (readPointer_CT$wnnzscfarg_0_1_argbuf_rwb_d[0] && (! readPointer_CT$wnnzscfarg_0_1_argbuf_rwb_emitted[0]))};
  assign lizzieLet58_2_d = {readPointer_CT$wnnzscfarg_0_1_argbuf_rwb_d[115:1],
                            (readPointer_CT$wnnzscfarg_0_1_argbuf_rwb_d[0] && (! readPointer_CT$wnnzscfarg_0_1_argbuf_rwb_emitted[1]))};
  assign lizzieLet58_3_d = {readPointer_CT$wnnzscfarg_0_1_argbuf_rwb_d[115:1],
                            (readPointer_CT$wnnzscfarg_0_1_argbuf_rwb_d[0] && (! readPointer_CT$wnnzscfarg_0_1_argbuf_rwb_emitted[2]))};
  assign lizzieLet58_4_d = {readPointer_CT$wnnzscfarg_0_1_argbuf_rwb_d[115:1],
                            (readPointer_CT$wnnzscfarg_0_1_argbuf_rwb_d[0] && (! readPointer_CT$wnnzscfarg_0_1_argbuf_rwb_emitted[3]))};
  assign readPointer_CT$wnnzscfarg_0_1_argbuf_rwb_done = (readPointer_CT$wnnzscfarg_0_1_argbuf_rwb_emitted | ({lizzieLet58_4_d[0],
                                                                                                               lizzieLet58_3_d[0],
                                                                                                               lizzieLet58_2_d[0],
                                                                                                               lizzieLet58_1_d[0]} & {lizzieLet58_4_r,
                                                                                                                                      lizzieLet58_3_r,
                                                                                                                                      lizzieLet58_2_r,
                                                                                                                                      lizzieLet58_1_r}));
  assign readPointer_CT$wnnzscfarg_0_1_argbuf_rwb_r = (& readPointer_CT$wnnzscfarg_0_1_argbuf_rwb_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_CT$wnnzscfarg_0_1_argbuf_rwb_emitted <= 4'd0;
    else
      readPointer_CT$wnnzscfarg_0_1_argbuf_rwb_emitted <= (readPointer_CT$wnnzscfarg_0_1_argbuf_rwb_r ? 4'd0 :
                                                           readPointer_CT$wnnzscfarg_0_1_argbuf_rwb_done);
  
  /* buf (Ty CTf''''''''''''_f''''''''''''_Int) : (readPointer_CTf''''''''''''_f''''''''''''_Intscfarg_0_1_1_argbuf,CTf''''''''''''_f''''''''''''_Int) > (readPointer_CTf''''''''''''_f''''''''''''_Intscfarg_0_1_1_argbuf_rwb,CTf''''''''''''_f''''''''''''_Int) */
  \CTf''''''''''''_f''''''''''''_Int_t  \readPointer_CTf''''''''''''_f''''''''''''_Intscfarg_0_1_1_argbuf_bufchan_d ;
  logic \readPointer_CTf''''''''''''_f''''''''''''_Intscfarg_0_1_1_argbuf_bufchan_r ;
  assign \readPointer_CTf''''''''''''_f''''''''''''_Intscfarg_0_1_1_argbuf_r  = ((! \readPointer_CTf''''''''''''_f''''''''''''_Intscfarg_0_1_1_argbuf_bufchan_d [0]) || \readPointer_CTf''''''''''''_f''''''''''''_Intscfarg_0_1_1_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \readPointer_CTf''''''''''''_f''''''''''''_Intscfarg_0_1_1_argbuf_bufchan_d  <= {115'd0,
                                                                                       1'd0};
    else
      if (\readPointer_CTf''''''''''''_f''''''''''''_Intscfarg_0_1_1_argbuf_r )
        \readPointer_CTf''''''''''''_f''''''''''''_Intscfarg_0_1_1_argbuf_bufchan_d  <= \readPointer_CTf''''''''''''_f''''''''''''_Intscfarg_0_1_1_argbuf_d ;
  \CTf''''''''''''_f''''''''''''_Int_t  \readPointer_CTf''''''''''''_f''''''''''''_Intscfarg_0_1_1_argbuf_bufchan_buf ;
  assign \readPointer_CTf''''''''''''_f''''''''''''_Intscfarg_0_1_1_argbuf_bufchan_r  = (! \readPointer_CTf''''''''''''_f''''''''''''_Intscfarg_0_1_1_argbuf_bufchan_buf [0]);
  assign \readPointer_CTf''''''''''''_f''''''''''''_Intscfarg_0_1_1_argbuf_rwb_d  = (\readPointer_CTf''''''''''''_f''''''''''''_Intscfarg_0_1_1_argbuf_bufchan_buf [0] ? \readPointer_CTf''''''''''''_f''''''''''''_Intscfarg_0_1_1_argbuf_bufchan_buf  :
                                                                                     \readPointer_CTf''''''''''''_f''''''''''''_Intscfarg_0_1_1_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \readPointer_CTf''''''''''''_f''''''''''''_Intscfarg_0_1_1_argbuf_bufchan_buf  <= {115'd0,
                                                                                         1'd0};
    else
      if ((\readPointer_CTf''''''''''''_f''''''''''''_Intscfarg_0_1_1_argbuf_rwb_r  && \readPointer_CTf''''''''''''_f''''''''''''_Intscfarg_0_1_1_argbuf_bufchan_buf [0]))
        \readPointer_CTf''''''''''''_f''''''''''''_Intscfarg_0_1_1_argbuf_bufchan_buf  <= {115'd0,
                                                                                           1'd0};
      else if (((! \readPointer_CTf''''''''''''_f''''''''''''_Intscfarg_0_1_1_argbuf_rwb_r ) && (! \readPointer_CTf''''''''''''_f''''''''''''_Intscfarg_0_1_1_argbuf_bufchan_buf [0])))
        \readPointer_CTf''''''''''''_f''''''''''''_Intscfarg_0_1_1_argbuf_bufchan_buf  <= \readPointer_CTf''''''''''''_f''''''''''''_Intscfarg_0_1_1_argbuf_bufchan_d ;
  
  /* fork (Ty CTf''''''''''''_f''''''''''''_Int) : (readPointer_CTf''''''''''''_f''''''''''''_Intscfarg_0_1_1_argbuf_rwb,CTf''''''''''''_f''''''''''''_Int) > [(lizzieLet62_1,CTf''''''''''''_f''''''''''''_Int),
                                                                                                                                                          (lizzieLet62_2,CTf''''''''''''_f''''''''''''_Int),
                                                                                                                                                          (lizzieLet62_3,CTf''''''''''''_f''''''''''''_Int),
                                                                                                                                                          (lizzieLet62_4,CTf''''''''''''_f''''''''''''_Int)] */
  logic [3:0] \readPointer_CTf''''''''''''_f''''''''''''_Intscfarg_0_1_1_argbuf_rwb_emitted ;
  logic [3:0] \readPointer_CTf''''''''''''_f''''''''''''_Intscfarg_0_1_1_argbuf_rwb_done ;
  assign lizzieLet62_1_d = {\readPointer_CTf''''''''''''_f''''''''''''_Intscfarg_0_1_1_argbuf_rwb_d [115:1],
                            (\readPointer_CTf''''''''''''_f''''''''''''_Intscfarg_0_1_1_argbuf_rwb_d [0] && (! \readPointer_CTf''''''''''''_f''''''''''''_Intscfarg_0_1_1_argbuf_rwb_emitted [0]))};
  assign lizzieLet62_2_d = {\readPointer_CTf''''''''''''_f''''''''''''_Intscfarg_0_1_1_argbuf_rwb_d [115:1],
                            (\readPointer_CTf''''''''''''_f''''''''''''_Intscfarg_0_1_1_argbuf_rwb_d [0] && (! \readPointer_CTf''''''''''''_f''''''''''''_Intscfarg_0_1_1_argbuf_rwb_emitted [1]))};
  assign lizzieLet62_3_d = {\readPointer_CTf''''''''''''_f''''''''''''_Intscfarg_0_1_1_argbuf_rwb_d [115:1],
                            (\readPointer_CTf''''''''''''_f''''''''''''_Intscfarg_0_1_1_argbuf_rwb_d [0] && (! \readPointer_CTf''''''''''''_f''''''''''''_Intscfarg_0_1_1_argbuf_rwb_emitted [2]))};
  assign lizzieLet62_4_d = {\readPointer_CTf''''''''''''_f''''''''''''_Intscfarg_0_1_1_argbuf_rwb_d [115:1],
                            (\readPointer_CTf''''''''''''_f''''''''''''_Intscfarg_0_1_1_argbuf_rwb_d [0] && (! \readPointer_CTf''''''''''''_f''''''''''''_Intscfarg_0_1_1_argbuf_rwb_emitted [3]))};
  assign \readPointer_CTf''''''''''''_f''''''''''''_Intscfarg_0_1_1_argbuf_rwb_done  = (\readPointer_CTf''''''''''''_f''''''''''''_Intscfarg_0_1_1_argbuf_rwb_emitted  | ({lizzieLet62_4_d[0],
                                                                                                                                                                           lizzieLet62_3_d[0],
                                                                                                                                                                           lizzieLet62_2_d[0],
                                                                                                                                                                           lizzieLet62_1_d[0]} & {lizzieLet62_4_r,
                                                                                                                                                                                                  lizzieLet62_3_r,
                                                                                                                                                                                                  lizzieLet62_2_r,
                                                                                                                                                                                                  lizzieLet62_1_r}));
  assign \readPointer_CTf''''''''''''_f''''''''''''_Intscfarg_0_1_1_argbuf_rwb_r  = (& \readPointer_CTf''''''''''''_f''''''''''''_Intscfarg_0_1_1_argbuf_rwb_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \readPointer_CTf''''''''''''_f''''''''''''_Intscfarg_0_1_1_argbuf_rwb_emitted  <= 4'd0;
    else
      \readPointer_CTf''''''''''''_f''''''''''''_Intscfarg_0_1_1_argbuf_rwb_emitted  <= (\readPointer_CTf''''''''''''_f''''''''''''_Intscfarg_0_1_1_argbuf_rwb_r  ? 4'd0 :
                                                                                         \readPointer_CTf''''''''''''_f''''''''''''_Intscfarg_0_1_1_argbuf_rwb_done );
  
  /* buf (Ty CTf_f_Int) : (readPointer_CTf_f_Intscfarg_0_2_1_argbuf,CTf_f_Int) > (readPointer_CTf_f_Intscfarg_0_2_1_argbuf_rwb,CTf_f_Int) */
  CTf_f_Int_t readPointer_CTf_f_Intscfarg_0_2_1_argbuf_bufchan_d;
  logic readPointer_CTf_f_Intscfarg_0_2_1_argbuf_bufchan_r;
  assign readPointer_CTf_f_Intscfarg_0_2_1_argbuf_r = ((! readPointer_CTf_f_Intscfarg_0_2_1_argbuf_bufchan_d[0]) || readPointer_CTf_f_Intscfarg_0_2_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_CTf_f_Intscfarg_0_2_1_argbuf_bufchan_d <= {163'd0,
                                                             1'd0};
    else
      if (readPointer_CTf_f_Intscfarg_0_2_1_argbuf_r)
        readPointer_CTf_f_Intscfarg_0_2_1_argbuf_bufchan_d <= readPointer_CTf_f_Intscfarg_0_2_1_argbuf_d;
  CTf_f_Int_t readPointer_CTf_f_Intscfarg_0_2_1_argbuf_bufchan_buf;
  assign readPointer_CTf_f_Intscfarg_0_2_1_argbuf_bufchan_r = (! readPointer_CTf_f_Intscfarg_0_2_1_argbuf_bufchan_buf[0]);
  assign readPointer_CTf_f_Intscfarg_0_2_1_argbuf_rwb_d = (readPointer_CTf_f_Intscfarg_0_2_1_argbuf_bufchan_buf[0] ? readPointer_CTf_f_Intscfarg_0_2_1_argbuf_bufchan_buf :
                                                           readPointer_CTf_f_Intscfarg_0_2_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_CTf_f_Intscfarg_0_2_1_argbuf_bufchan_buf <= {163'd0,
                                                               1'd0};
    else
      if ((readPointer_CTf_f_Intscfarg_0_2_1_argbuf_rwb_r && readPointer_CTf_f_Intscfarg_0_2_1_argbuf_bufchan_buf[0]))
        readPointer_CTf_f_Intscfarg_0_2_1_argbuf_bufchan_buf <= {163'd0,
                                                                 1'd0};
      else if (((! readPointer_CTf_f_Intscfarg_0_2_1_argbuf_rwb_r) && (! readPointer_CTf_f_Intscfarg_0_2_1_argbuf_bufchan_buf[0])))
        readPointer_CTf_f_Intscfarg_0_2_1_argbuf_bufchan_buf <= readPointer_CTf_f_Intscfarg_0_2_1_argbuf_bufchan_d;
  
  /* fork (Ty CTf_f_Int) : (readPointer_CTf_f_Intscfarg_0_2_1_argbuf_rwb,CTf_f_Int) > [(lizzieLet67_1,CTf_f_Int),
                                                                                  (lizzieLet67_2,CTf_f_Int),
                                                                                  (lizzieLet67_3,CTf_f_Int),
                                                                                  (lizzieLet67_4,CTf_f_Int)] */
  logic [3:0] readPointer_CTf_f_Intscfarg_0_2_1_argbuf_rwb_emitted;
  logic [3:0] readPointer_CTf_f_Intscfarg_0_2_1_argbuf_rwb_done;
  assign lizzieLet67_1_d = {readPointer_CTf_f_Intscfarg_0_2_1_argbuf_rwb_d[163:1],
                            (readPointer_CTf_f_Intscfarg_0_2_1_argbuf_rwb_d[0] && (! readPointer_CTf_f_Intscfarg_0_2_1_argbuf_rwb_emitted[0]))};
  assign lizzieLet67_2_d = {readPointer_CTf_f_Intscfarg_0_2_1_argbuf_rwb_d[163:1],
                            (readPointer_CTf_f_Intscfarg_0_2_1_argbuf_rwb_d[0] && (! readPointer_CTf_f_Intscfarg_0_2_1_argbuf_rwb_emitted[1]))};
  assign lizzieLet67_3_d = {readPointer_CTf_f_Intscfarg_0_2_1_argbuf_rwb_d[163:1],
                            (readPointer_CTf_f_Intscfarg_0_2_1_argbuf_rwb_d[0] && (! readPointer_CTf_f_Intscfarg_0_2_1_argbuf_rwb_emitted[2]))};
  assign lizzieLet67_4_d = {readPointer_CTf_f_Intscfarg_0_2_1_argbuf_rwb_d[163:1],
                            (readPointer_CTf_f_Intscfarg_0_2_1_argbuf_rwb_d[0] && (! readPointer_CTf_f_Intscfarg_0_2_1_argbuf_rwb_emitted[3]))};
  assign readPointer_CTf_f_Intscfarg_0_2_1_argbuf_rwb_done = (readPointer_CTf_f_Intscfarg_0_2_1_argbuf_rwb_emitted | ({lizzieLet67_4_d[0],
                                                                                                                       lizzieLet67_3_d[0],
                                                                                                                       lizzieLet67_2_d[0],
                                                                                                                       lizzieLet67_1_d[0]} & {lizzieLet67_4_r,
                                                                                                                                              lizzieLet67_3_r,
                                                                                                                                              lizzieLet67_2_r,
                                                                                                                                              lizzieLet67_1_r}));
  assign readPointer_CTf_f_Intscfarg_0_2_1_argbuf_rwb_r = (& readPointer_CTf_f_Intscfarg_0_2_1_argbuf_rwb_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_CTf_f_Intscfarg_0_2_1_argbuf_rwb_emitted <= 4'd0;
    else
      readPointer_CTf_f_Intscfarg_0_2_1_argbuf_rwb_emitted <= (readPointer_CTf_f_Intscfarg_0_2_1_argbuf_rwb_r ? 4'd0 :
                                                               readPointer_CTf_f_Intscfarg_0_2_1_argbuf_rwb_done);
  
  /* buf (Ty QTree_Int) : (readPointer_QTree_Intm1aeq_1_argbuf,QTree_Int) > (readPointer_QTree_Intm1aeq_1_argbuf_rwb,QTree_Int) */
  QTree_Int_t readPointer_QTree_Intm1aeq_1_argbuf_bufchan_d;
  logic readPointer_QTree_Intm1aeq_1_argbuf_bufchan_r;
  assign readPointer_QTree_Intm1aeq_1_argbuf_r = ((! readPointer_QTree_Intm1aeq_1_argbuf_bufchan_d[0]) || readPointer_QTree_Intm1aeq_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Intm1aeq_1_argbuf_bufchan_d <= {66'd0, 1'd0};
    else
      if (readPointer_QTree_Intm1aeq_1_argbuf_r)
        readPointer_QTree_Intm1aeq_1_argbuf_bufchan_d <= readPointer_QTree_Intm1aeq_1_argbuf_d;
  QTree_Int_t readPointer_QTree_Intm1aeq_1_argbuf_bufchan_buf;
  assign readPointer_QTree_Intm1aeq_1_argbuf_bufchan_r = (! readPointer_QTree_Intm1aeq_1_argbuf_bufchan_buf[0]);
  assign readPointer_QTree_Intm1aeq_1_argbuf_rwb_d = (readPointer_QTree_Intm1aeq_1_argbuf_bufchan_buf[0] ? readPointer_QTree_Intm1aeq_1_argbuf_bufchan_buf :
                                                      readPointer_QTree_Intm1aeq_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Intm1aeq_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((readPointer_QTree_Intm1aeq_1_argbuf_rwb_r && readPointer_QTree_Intm1aeq_1_argbuf_bufchan_buf[0]))
        readPointer_QTree_Intm1aeq_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
      else if (((! readPointer_QTree_Intm1aeq_1_argbuf_rwb_r) && (! readPointer_QTree_Intm1aeq_1_argbuf_bufchan_buf[0])))
        readPointer_QTree_Intm1aeq_1_argbuf_bufchan_buf <= readPointer_QTree_Intm1aeq_1_argbuf_bufchan_d;
  
  /* fork (Ty QTree_Int) : (readPointer_QTree_Intm1aeq_1_argbuf_rwb,QTree_Int) > [(lizzieLet17_1,QTree_Int),
                                                                             (lizzieLet17_2,QTree_Int),
                                                                             (lizzieLet17_3,QTree_Int),
                                                                             (lizzieLet17_4,QTree_Int),
                                                                             (lizzieLet17_5,QTree_Int),
                                                                             (lizzieLet17_6,QTree_Int),
                                                                             (lizzieLet17_7,QTree_Int),
                                                                             (lizzieLet17_8,QTree_Int),
                                                                             (lizzieLet17_9,QTree_Int),
                                                                             (lizzieLet17_10,QTree_Int),
                                                                             (lizzieLet17_11,QTree_Int)] */
  logic [10:0] readPointer_QTree_Intm1aeq_1_argbuf_rwb_emitted;
  logic [10:0] readPointer_QTree_Intm1aeq_1_argbuf_rwb_done;
  assign lizzieLet17_1_d = {readPointer_QTree_Intm1aeq_1_argbuf_rwb_d[66:1],
                            (readPointer_QTree_Intm1aeq_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intm1aeq_1_argbuf_rwb_emitted[0]))};
  assign lizzieLet17_2_d = {readPointer_QTree_Intm1aeq_1_argbuf_rwb_d[66:1],
                            (readPointer_QTree_Intm1aeq_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intm1aeq_1_argbuf_rwb_emitted[1]))};
  assign lizzieLet17_3_d = {readPointer_QTree_Intm1aeq_1_argbuf_rwb_d[66:1],
                            (readPointer_QTree_Intm1aeq_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intm1aeq_1_argbuf_rwb_emitted[2]))};
  assign lizzieLet17_4_d = {readPointer_QTree_Intm1aeq_1_argbuf_rwb_d[66:1],
                            (readPointer_QTree_Intm1aeq_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intm1aeq_1_argbuf_rwb_emitted[3]))};
  assign lizzieLet17_5_d = {readPointer_QTree_Intm1aeq_1_argbuf_rwb_d[66:1],
                            (readPointer_QTree_Intm1aeq_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intm1aeq_1_argbuf_rwb_emitted[4]))};
  assign lizzieLet17_6_d = {readPointer_QTree_Intm1aeq_1_argbuf_rwb_d[66:1],
                            (readPointer_QTree_Intm1aeq_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intm1aeq_1_argbuf_rwb_emitted[5]))};
  assign lizzieLet17_7_d = {readPointer_QTree_Intm1aeq_1_argbuf_rwb_d[66:1],
                            (readPointer_QTree_Intm1aeq_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intm1aeq_1_argbuf_rwb_emitted[6]))};
  assign lizzieLet17_8_d = {readPointer_QTree_Intm1aeq_1_argbuf_rwb_d[66:1],
                            (readPointer_QTree_Intm1aeq_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intm1aeq_1_argbuf_rwb_emitted[7]))};
  assign lizzieLet17_9_d = {readPointer_QTree_Intm1aeq_1_argbuf_rwb_d[66:1],
                            (readPointer_QTree_Intm1aeq_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intm1aeq_1_argbuf_rwb_emitted[8]))};
  assign lizzieLet17_10_d = {readPointer_QTree_Intm1aeq_1_argbuf_rwb_d[66:1],
                             (readPointer_QTree_Intm1aeq_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intm1aeq_1_argbuf_rwb_emitted[9]))};
  assign lizzieLet17_11_d = {readPointer_QTree_Intm1aeq_1_argbuf_rwb_d[66:1],
                             (readPointer_QTree_Intm1aeq_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intm1aeq_1_argbuf_rwb_emitted[10]))};
  assign readPointer_QTree_Intm1aeq_1_argbuf_rwb_done = (readPointer_QTree_Intm1aeq_1_argbuf_rwb_emitted | ({lizzieLet17_11_d[0],
                                                                                                             lizzieLet17_10_d[0],
                                                                                                             lizzieLet17_9_d[0],
                                                                                                             lizzieLet17_8_d[0],
                                                                                                             lizzieLet17_7_d[0],
                                                                                                             lizzieLet17_6_d[0],
                                                                                                             lizzieLet17_5_d[0],
                                                                                                             lizzieLet17_4_d[0],
                                                                                                             lizzieLet17_3_d[0],
                                                                                                             lizzieLet17_2_d[0],
                                                                                                             lizzieLet17_1_d[0]} & {lizzieLet17_11_r,
                                                                                                                                    lizzieLet17_10_r,
                                                                                                                                    lizzieLet17_9_r,
                                                                                                                                    lizzieLet17_8_r,
                                                                                                                                    lizzieLet17_7_r,
                                                                                                                                    lizzieLet17_6_r,
                                                                                                                                    lizzieLet17_5_r,
                                                                                                                                    lizzieLet17_4_r,
                                                                                                                                    lizzieLet17_3_r,
                                                                                                                                    lizzieLet17_2_r,
                                                                                                                                    lizzieLet17_1_r}));
  assign readPointer_QTree_Intm1aeq_1_argbuf_rwb_r = (& readPointer_QTree_Intm1aeq_1_argbuf_rwb_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Intm1aeq_1_argbuf_rwb_emitted <= 11'd0;
    else
      readPointer_QTree_Intm1aeq_1_argbuf_rwb_emitted <= (readPointer_QTree_Intm1aeq_1_argbuf_rwb_r ? 11'd0 :
                                                          readPointer_QTree_Intm1aeq_1_argbuf_rwb_done);
  
  /* buf (Ty QTree_Int) : (readPointer_QTree_Intm2aer_1_argbuf,QTree_Int) > (readPointer_QTree_Intm2aer_1_argbuf_rwb,QTree_Int) */
  QTree_Int_t readPointer_QTree_Intm2aer_1_argbuf_bufchan_d;
  logic readPointer_QTree_Intm2aer_1_argbuf_bufchan_r;
  assign readPointer_QTree_Intm2aer_1_argbuf_r = ((! readPointer_QTree_Intm2aer_1_argbuf_bufchan_d[0]) || readPointer_QTree_Intm2aer_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Intm2aer_1_argbuf_bufchan_d <= {66'd0, 1'd0};
    else
      if (readPointer_QTree_Intm2aer_1_argbuf_r)
        readPointer_QTree_Intm2aer_1_argbuf_bufchan_d <= readPointer_QTree_Intm2aer_1_argbuf_d;
  QTree_Int_t readPointer_QTree_Intm2aer_1_argbuf_bufchan_buf;
  assign readPointer_QTree_Intm2aer_1_argbuf_bufchan_r = (! readPointer_QTree_Intm2aer_1_argbuf_bufchan_buf[0]);
  assign readPointer_QTree_Intm2aer_1_argbuf_rwb_d = (readPointer_QTree_Intm2aer_1_argbuf_bufchan_buf[0] ? readPointer_QTree_Intm2aer_1_argbuf_bufchan_buf :
                                                      readPointer_QTree_Intm2aer_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Intm2aer_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((readPointer_QTree_Intm2aer_1_argbuf_rwb_r && readPointer_QTree_Intm2aer_1_argbuf_bufchan_buf[0]))
        readPointer_QTree_Intm2aer_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
      else if (((! readPointer_QTree_Intm2aer_1_argbuf_rwb_r) && (! readPointer_QTree_Intm2aer_1_argbuf_bufchan_buf[0])))
        readPointer_QTree_Intm2aer_1_argbuf_bufchan_buf <= readPointer_QTree_Intm2aer_1_argbuf_bufchan_d;
  
  /* buf (Ty QTree_Int) : (readPointer_QTree_Intm3aes_1_argbuf,QTree_Int) > (readPointer_QTree_Intm3aes_1_argbuf_rwb,QTree_Int) */
  QTree_Int_t readPointer_QTree_Intm3aes_1_argbuf_bufchan_d;
  logic readPointer_QTree_Intm3aes_1_argbuf_bufchan_r;
  assign readPointer_QTree_Intm3aes_1_argbuf_r = ((! readPointer_QTree_Intm3aes_1_argbuf_bufchan_d[0]) || readPointer_QTree_Intm3aes_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Intm3aes_1_argbuf_bufchan_d <= {66'd0, 1'd0};
    else
      if (readPointer_QTree_Intm3aes_1_argbuf_r)
        readPointer_QTree_Intm3aes_1_argbuf_bufchan_d <= readPointer_QTree_Intm3aes_1_argbuf_d;
  QTree_Int_t readPointer_QTree_Intm3aes_1_argbuf_bufchan_buf;
  assign readPointer_QTree_Intm3aes_1_argbuf_bufchan_r = (! readPointer_QTree_Intm3aes_1_argbuf_bufchan_buf[0]);
  assign readPointer_QTree_Intm3aes_1_argbuf_rwb_d = (readPointer_QTree_Intm3aes_1_argbuf_bufchan_buf[0] ? readPointer_QTree_Intm3aes_1_argbuf_bufchan_buf :
                                                      readPointer_QTree_Intm3aes_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Intm3aes_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((readPointer_QTree_Intm3aes_1_argbuf_rwb_r && readPointer_QTree_Intm3aes_1_argbuf_bufchan_buf[0]))
        readPointer_QTree_Intm3aes_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
      else if (((! readPointer_QTree_Intm3aes_1_argbuf_rwb_r) && (! readPointer_QTree_Intm3aes_1_argbuf_bufchan_buf[0])))
        readPointer_QTree_Intm3aes_1_argbuf_bufchan_buf <= readPointer_QTree_Intm3aes_1_argbuf_bufchan_d;
  
  /* buf (Ty QTree_Int) : (readPointer_QTree_Intq4afj_1_argbuf,QTree_Int) > (readPointer_QTree_Intq4afj_1_argbuf_rwb,QTree_Int) */
  QTree_Int_t readPointer_QTree_Intq4afj_1_argbuf_bufchan_d;
  logic readPointer_QTree_Intq4afj_1_argbuf_bufchan_r;
  assign readPointer_QTree_Intq4afj_1_argbuf_r = ((! readPointer_QTree_Intq4afj_1_argbuf_bufchan_d[0]) || readPointer_QTree_Intq4afj_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Intq4afj_1_argbuf_bufchan_d <= {66'd0, 1'd0};
    else
      if (readPointer_QTree_Intq4afj_1_argbuf_r)
        readPointer_QTree_Intq4afj_1_argbuf_bufchan_d <= readPointer_QTree_Intq4afj_1_argbuf_d;
  QTree_Int_t readPointer_QTree_Intq4afj_1_argbuf_bufchan_buf;
  assign readPointer_QTree_Intq4afj_1_argbuf_bufchan_r = (! readPointer_QTree_Intq4afj_1_argbuf_bufchan_buf[0]);
  assign readPointer_QTree_Intq4afj_1_argbuf_rwb_d = (readPointer_QTree_Intq4afj_1_argbuf_bufchan_buf[0] ? readPointer_QTree_Intq4afj_1_argbuf_bufchan_buf :
                                                      readPointer_QTree_Intq4afj_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Intq4afj_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((readPointer_QTree_Intq4afj_1_argbuf_rwb_r && readPointer_QTree_Intq4afj_1_argbuf_bufchan_buf[0]))
        readPointer_QTree_Intq4afj_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
      else if (((! readPointer_QTree_Intq4afj_1_argbuf_rwb_r) && (! readPointer_QTree_Intq4afj_1_argbuf_bufchan_buf[0])))
        readPointer_QTree_Intq4afj_1_argbuf_bufchan_buf <= readPointer_QTree_Intq4afj_1_argbuf_bufchan_d;
  
  /* fork (Ty QTree_Int) : (readPointer_QTree_Intq4afj_1_argbuf_rwb,QTree_Int) > [(lizzieLet6_1,QTree_Int),
                                                                             (lizzieLet6_2,QTree_Int),
                                                                             (lizzieLet6_3,QTree_Int),
                                                                             (lizzieLet6_4,QTree_Int),
                                                                             (lizzieLet6_5,QTree_Int),
                                                                             (lizzieLet6_6,QTree_Int),
                                                                             (lizzieLet6_7,QTree_Int),
                                                                             (lizzieLet6_8,QTree_Int),
                                                                             (lizzieLet6_9,QTree_Int)] */
  logic [8:0] readPointer_QTree_Intq4afj_1_argbuf_rwb_emitted;
  logic [8:0] readPointer_QTree_Intq4afj_1_argbuf_rwb_done;
  assign lizzieLet6_1_d = {readPointer_QTree_Intq4afj_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_Intq4afj_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intq4afj_1_argbuf_rwb_emitted[0]))};
  assign lizzieLet6_2_d = {readPointer_QTree_Intq4afj_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_Intq4afj_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intq4afj_1_argbuf_rwb_emitted[1]))};
  assign lizzieLet6_3_d = {readPointer_QTree_Intq4afj_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_Intq4afj_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intq4afj_1_argbuf_rwb_emitted[2]))};
  assign lizzieLet6_4_d = {readPointer_QTree_Intq4afj_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_Intq4afj_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intq4afj_1_argbuf_rwb_emitted[3]))};
  assign lizzieLet6_5_d = {readPointer_QTree_Intq4afj_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_Intq4afj_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intq4afj_1_argbuf_rwb_emitted[4]))};
  assign lizzieLet6_6_d = {readPointer_QTree_Intq4afj_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_Intq4afj_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intq4afj_1_argbuf_rwb_emitted[5]))};
  assign lizzieLet6_7_d = {readPointer_QTree_Intq4afj_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_Intq4afj_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intq4afj_1_argbuf_rwb_emitted[6]))};
  assign lizzieLet6_8_d = {readPointer_QTree_Intq4afj_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_Intq4afj_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intq4afj_1_argbuf_rwb_emitted[7]))};
  assign lizzieLet6_9_d = {readPointer_QTree_Intq4afj_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_Intq4afj_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intq4afj_1_argbuf_rwb_emitted[8]))};
  assign readPointer_QTree_Intq4afj_1_argbuf_rwb_done = (readPointer_QTree_Intq4afj_1_argbuf_rwb_emitted | ({lizzieLet6_9_d[0],
                                                                                                             lizzieLet6_8_d[0],
                                                                                                             lizzieLet6_7_d[0],
                                                                                                             lizzieLet6_6_d[0],
                                                                                                             lizzieLet6_5_d[0],
                                                                                                             lizzieLet6_4_d[0],
                                                                                                             lizzieLet6_3_d[0],
                                                                                                             lizzieLet6_2_d[0],
                                                                                                             lizzieLet6_1_d[0]} & {lizzieLet6_9_r,
                                                                                                                                   lizzieLet6_8_r,
                                                                                                                                   lizzieLet6_7_r,
                                                                                                                                   lizzieLet6_6_r,
                                                                                                                                   lizzieLet6_5_r,
                                                                                                                                   lizzieLet6_4_r,
                                                                                                                                   lizzieLet6_3_r,
                                                                                                                                   lizzieLet6_2_r,
                                                                                                                                   lizzieLet6_1_r}));
  assign readPointer_QTree_Intq4afj_1_argbuf_rwb_r = (& readPointer_QTree_Intq4afj_1_argbuf_rwb_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Intq4afj_1_argbuf_rwb_emitted <= 9'd0;
    else
      readPointer_QTree_Intq4afj_1_argbuf_rwb_emitted <= (readPointer_QTree_Intq4afj_1_argbuf_rwb_r ? 9'd0 :
                                                          readPointer_QTree_Intq4afj_1_argbuf_rwb_done);
  
  /* buf (Ty QTree_Int) : (readPointer_QTree_Intt4afk_1_argbuf,QTree_Int) > (readPointer_QTree_Intt4afk_1_argbuf_rwb,QTree_Int) */
  QTree_Int_t readPointer_QTree_Intt4afk_1_argbuf_bufchan_d;
  logic readPointer_QTree_Intt4afk_1_argbuf_bufchan_r;
  assign readPointer_QTree_Intt4afk_1_argbuf_r = ((! readPointer_QTree_Intt4afk_1_argbuf_bufchan_d[0]) || readPointer_QTree_Intt4afk_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Intt4afk_1_argbuf_bufchan_d <= {66'd0, 1'd0};
    else
      if (readPointer_QTree_Intt4afk_1_argbuf_r)
        readPointer_QTree_Intt4afk_1_argbuf_bufchan_d <= readPointer_QTree_Intt4afk_1_argbuf_d;
  QTree_Int_t readPointer_QTree_Intt4afk_1_argbuf_bufchan_buf;
  assign readPointer_QTree_Intt4afk_1_argbuf_bufchan_r = (! readPointer_QTree_Intt4afk_1_argbuf_bufchan_buf[0]);
  assign readPointer_QTree_Intt4afk_1_argbuf_rwb_d = (readPointer_QTree_Intt4afk_1_argbuf_bufchan_buf[0] ? readPointer_QTree_Intt4afk_1_argbuf_bufchan_buf :
                                                      readPointer_QTree_Intt4afk_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Intt4afk_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((readPointer_QTree_Intt4afk_1_argbuf_rwb_r && readPointer_QTree_Intt4afk_1_argbuf_bufchan_buf[0]))
        readPointer_QTree_Intt4afk_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
      else if (((! readPointer_QTree_Intt4afk_1_argbuf_rwb_r) && (! readPointer_QTree_Intt4afk_1_argbuf_bufchan_buf[0])))
        readPointer_QTree_Intt4afk_1_argbuf_bufchan_buf <= readPointer_QTree_Intt4afk_1_argbuf_bufchan_d;
  
  /* buf (Ty QTree_Int) : (readPointer_QTree_Intwsmk_1_1_argbuf,QTree_Int) > (readPointer_QTree_Intwsmk_1_1_argbuf_rwb,QTree_Int) */
  QTree_Int_t readPointer_QTree_Intwsmk_1_1_argbuf_bufchan_d;
  logic readPointer_QTree_Intwsmk_1_1_argbuf_bufchan_r;
  assign readPointer_QTree_Intwsmk_1_1_argbuf_r = ((! readPointer_QTree_Intwsmk_1_1_argbuf_bufchan_d[0]) || readPointer_QTree_Intwsmk_1_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Intwsmk_1_1_argbuf_bufchan_d <= {66'd0, 1'd0};
    else
      if (readPointer_QTree_Intwsmk_1_1_argbuf_r)
        readPointer_QTree_Intwsmk_1_1_argbuf_bufchan_d <= readPointer_QTree_Intwsmk_1_1_argbuf_d;
  QTree_Int_t readPointer_QTree_Intwsmk_1_1_argbuf_bufchan_buf;
  assign readPointer_QTree_Intwsmk_1_1_argbuf_bufchan_r = (! readPointer_QTree_Intwsmk_1_1_argbuf_bufchan_buf[0]);
  assign readPointer_QTree_Intwsmk_1_1_argbuf_rwb_d = (readPointer_QTree_Intwsmk_1_1_argbuf_bufchan_buf[0] ? readPointer_QTree_Intwsmk_1_1_argbuf_bufchan_buf :
                                                       readPointer_QTree_Intwsmk_1_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Intwsmk_1_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((readPointer_QTree_Intwsmk_1_1_argbuf_rwb_r && readPointer_QTree_Intwsmk_1_1_argbuf_bufchan_buf[0]))
        readPointer_QTree_Intwsmk_1_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
      else if (((! readPointer_QTree_Intwsmk_1_1_argbuf_rwb_r) && (! readPointer_QTree_Intwsmk_1_1_argbuf_bufchan_buf[0])))
        readPointer_QTree_Intwsmk_1_1_argbuf_bufchan_buf <= readPointer_QTree_Intwsmk_1_1_argbuf_bufchan_d;
  
  /* fork (Ty QTree_Int) : (readPointer_QTree_Intwsmk_1_1_argbuf_rwb,QTree_Int) > [(lizzieLet4_1,QTree_Int),
                                                                              (lizzieLet4_2,QTree_Int),
                                                                              (lizzieLet4_3,QTree_Int),
                                                                              (lizzieLet4_4,QTree_Int)] */
  logic [3:0] readPointer_QTree_Intwsmk_1_1_argbuf_rwb_emitted;
  logic [3:0] readPointer_QTree_Intwsmk_1_1_argbuf_rwb_done;
  assign lizzieLet4_1_d = {readPointer_QTree_Intwsmk_1_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_Intwsmk_1_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intwsmk_1_1_argbuf_rwb_emitted[0]))};
  assign lizzieLet4_2_d = {readPointer_QTree_Intwsmk_1_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_Intwsmk_1_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intwsmk_1_1_argbuf_rwb_emitted[1]))};
  assign lizzieLet4_3_d = {readPointer_QTree_Intwsmk_1_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_Intwsmk_1_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intwsmk_1_1_argbuf_rwb_emitted[2]))};
  assign lizzieLet4_4_d = {readPointer_QTree_Intwsmk_1_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_Intwsmk_1_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intwsmk_1_1_argbuf_rwb_emitted[3]))};
  assign readPointer_QTree_Intwsmk_1_1_argbuf_rwb_done = (readPointer_QTree_Intwsmk_1_1_argbuf_rwb_emitted | ({lizzieLet4_4_d[0],
                                                                                                               lizzieLet4_3_d[0],
                                                                                                               lizzieLet4_2_d[0],
                                                                                                               lizzieLet4_1_d[0]} & {lizzieLet4_4_r,
                                                                                                                                     lizzieLet4_3_r,
                                                                                                                                     lizzieLet4_2_r,
                                                                                                                                     lizzieLet4_1_r}));
  assign readPointer_QTree_Intwsmk_1_1_argbuf_rwb_r = (& readPointer_QTree_Intwsmk_1_1_argbuf_rwb_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Intwsmk_1_1_argbuf_rwb_emitted <= 4'd0;
    else
      readPointer_QTree_Intwsmk_1_1_argbuf_rwb_emitted <= (readPointer_QTree_Intwsmk_1_1_argbuf_rwb_r ? 4'd0 :
                                                           readPointer_QTree_Intwsmk_1_1_argbuf_rwb_done);
  
  /* buf (Ty Pointer_CTf''''''''''''_f''''''''''''_Int) : (sc_0_10_destruct,Pointer_CTf''''''''''''_f''''''''''''_Int) > (sc_0_10_1_argbuf,Pointer_CTf''''''''''''_f''''''''''''_Int) */
  \Pointer_CTf''''''''''''_f''''''''''''_Int_t  sc_0_10_destruct_bufchan_d;
  logic sc_0_10_destruct_bufchan_r;
  assign sc_0_10_destruct_r = ((! sc_0_10_destruct_bufchan_d[0]) || sc_0_10_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) sc_0_10_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (sc_0_10_destruct_r)
        sc_0_10_destruct_bufchan_d <= sc_0_10_destruct_d;
  \Pointer_CTf''''''''''''_f''''''''''''_Int_t  sc_0_10_destruct_bufchan_buf;
  assign sc_0_10_destruct_bufchan_r = (! sc_0_10_destruct_bufchan_buf[0]);
  assign sc_0_10_1_argbuf_d = (sc_0_10_destruct_bufchan_buf[0] ? sc_0_10_destruct_bufchan_buf :
                               sc_0_10_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) sc_0_10_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((sc_0_10_1_argbuf_r && sc_0_10_destruct_bufchan_buf[0]))
        sc_0_10_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! sc_0_10_1_argbuf_r) && (! sc_0_10_destruct_bufchan_buf[0])))
        sc_0_10_destruct_bufchan_buf <= sc_0_10_destruct_bufchan_d;
  
  /* buf (Ty Pointer_CTf_f_Int) : (sc_0_14_destruct,Pointer_CTf_f_Int) > (sc_0_14_1_argbuf,Pointer_CTf_f_Int) */
  Pointer_CTf_f_Int_t sc_0_14_destruct_bufchan_d;
  logic sc_0_14_destruct_bufchan_r;
  assign sc_0_14_destruct_r = ((! sc_0_14_destruct_bufchan_d[0]) || sc_0_14_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) sc_0_14_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (sc_0_14_destruct_r)
        sc_0_14_destruct_bufchan_d <= sc_0_14_destruct_d;
  Pointer_CTf_f_Int_t sc_0_14_destruct_bufchan_buf;
  assign sc_0_14_destruct_bufchan_r = (! sc_0_14_destruct_bufchan_buf[0]);
  assign sc_0_14_1_argbuf_d = (sc_0_14_destruct_bufchan_buf[0] ? sc_0_14_destruct_bufchan_buf :
                               sc_0_14_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) sc_0_14_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((sc_0_14_1_argbuf_r && sc_0_14_destruct_bufchan_buf[0]))
        sc_0_14_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! sc_0_14_1_argbuf_r) && (! sc_0_14_destruct_bufchan_buf[0])))
        sc_0_14_destruct_bufchan_buf <= sc_0_14_destruct_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz) : (sc_0_6_destruct,Pointer_CT$wnnz) > (sc_0_6_1_argbuf,Pointer_CT$wnnz) */
  Pointer_CT$wnnz_t sc_0_6_destruct_bufchan_d;
  logic sc_0_6_destruct_bufchan_r;
  assign sc_0_6_destruct_r = ((! sc_0_6_destruct_bufchan_d[0]) || sc_0_6_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) sc_0_6_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (sc_0_6_destruct_r)
        sc_0_6_destruct_bufchan_d <= sc_0_6_destruct_d;
  Pointer_CT$wnnz_t sc_0_6_destruct_bufchan_buf;
  assign sc_0_6_destruct_bufchan_r = (! sc_0_6_destruct_bufchan_buf[0]);
  assign sc_0_6_1_argbuf_d = (sc_0_6_destruct_bufchan_buf[0] ? sc_0_6_destruct_bufchan_buf :
                              sc_0_6_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) sc_0_6_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((sc_0_6_1_argbuf_r && sc_0_6_destruct_bufchan_buf[0]))
        sc_0_6_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! sc_0_6_1_argbuf_r) && (! sc_0_6_destruct_bufchan_buf[0])))
        sc_0_6_destruct_bufchan_buf <= sc_0_6_destruct_bufchan_d;
  
  /* buf (Ty Pointer_CTf''''''''''''_f''''''''''''_Int) : (scfarg_0_1_goMux_mux,Pointer_CTf''''''''''''_f''''''''''''_Int) > (scfarg_0_1_1_argbuf,Pointer_CTf''''''''''''_f''''''''''''_Int) */
  \Pointer_CTf''''''''''''_f''''''''''''_Int_t  scfarg_0_1_goMux_mux_bufchan_d;
  logic scfarg_0_1_goMux_mux_bufchan_r;
  assign scfarg_0_1_goMux_mux_r = ((! scfarg_0_1_goMux_mux_bufchan_d[0]) || scfarg_0_1_goMux_mux_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      scfarg_0_1_goMux_mux_bufchan_d <= {16'd0, 1'd0};
    else
      if (scfarg_0_1_goMux_mux_r)
        scfarg_0_1_goMux_mux_bufchan_d <= scfarg_0_1_goMux_mux_d;
  \Pointer_CTf''''''''''''_f''''''''''''_Int_t  scfarg_0_1_goMux_mux_bufchan_buf;
  assign scfarg_0_1_goMux_mux_bufchan_r = (! scfarg_0_1_goMux_mux_bufchan_buf[0]);
  assign scfarg_0_1_1_argbuf_d = (scfarg_0_1_goMux_mux_bufchan_buf[0] ? scfarg_0_1_goMux_mux_bufchan_buf :
                                  scfarg_0_1_goMux_mux_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      scfarg_0_1_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((scfarg_0_1_1_argbuf_r && scfarg_0_1_goMux_mux_bufchan_buf[0]))
        scfarg_0_1_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
      else if (((! scfarg_0_1_1_argbuf_r) && (! scfarg_0_1_goMux_mux_bufchan_buf[0])))
        scfarg_0_1_goMux_mux_bufchan_buf <= scfarg_0_1_goMux_mux_bufchan_d;
  
  /* buf (Ty Pointer_CTf_f_Int) : (scfarg_0_2_goMux_mux,Pointer_CTf_f_Int) > (scfarg_0_2_1_argbuf,Pointer_CTf_f_Int) */
  Pointer_CTf_f_Int_t scfarg_0_2_goMux_mux_bufchan_d;
  logic scfarg_0_2_goMux_mux_bufchan_r;
  assign scfarg_0_2_goMux_mux_r = ((! scfarg_0_2_goMux_mux_bufchan_d[0]) || scfarg_0_2_goMux_mux_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      scfarg_0_2_goMux_mux_bufchan_d <= {16'd0, 1'd0};
    else
      if (scfarg_0_2_goMux_mux_r)
        scfarg_0_2_goMux_mux_bufchan_d <= scfarg_0_2_goMux_mux_d;
  Pointer_CTf_f_Int_t scfarg_0_2_goMux_mux_bufchan_buf;
  assign scfarg_0_2_goMux_mux_bufchan_r = (! scfarg_0_2_goMux_mux_bufchan_buf[0]);
  assign scfarg_0_2_1_argbuf_d = (scfarg_0_2_goMux_mux_bufchan_buf[0] ? scfarg_0_2_goMux_mux_bufchan_buf :
                                  scfarg_0_2_goMux_mux_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      scfarg_0_2_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((scfarg_0_2_1_argbuf_r && scfarg_0_2_goMux_mux_bufchan_buf[0]))
        scfarg_0_2_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
      else if (((! scfarg_0_2_1_argbuf_r) && (! scfarg_0_2_goMux_mux_bufchan_buf[0])))
        scfarg_0_2_goMux_mux_bufchan_buf <= scfarg_0_2_goMux_mux_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz) : (scfarg_0_goMux_mux,Pointer_CT$wnnz) > (scfarg_0_1_argbuf,Pointer_CT$wnnz) */
  Pointer_CT$wnnz_t scfarg_0_goMux_mux_bufchan_d;
  logic scfarg_0_goMux_mux_bufchan_r;
  assign scfarg_0_goMux_mux_r = ((! scfarg_0_goMux_mux_bufchan_d[0]) || scfarg_0_goMux_mux_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) scfarg_0_goMux_mux_bufchan_d <= {16'd0, 1'd0};
    else
      if (scfarg_0_goMux_mux_r)
        scfarg_0_goMux_mux_bufchan_d <= scfarg_0_goMux_mux_d;
  Pointer_CT$wnnz_t scfarg_0_goMux_mux_bufchan_buf;
  assign scfarg_0_goMux_mux_bufchan_r = (! scfarg_0_goMux_mux_bufchan_buf[0]);
  assign scfarg_0_1_argbuf_d = (scfarg_0_goMux_mux_bufchan_buf[0] ? scfarg_0_goMux_mux_bufchan_buf :
                                scfarg_0_goMux_mux_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      scfarg_0_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((scfarg_0_1_argbuf_r && scfarg_0_goMux_mux_bufchan_buf[0]))
        scfarg_0_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
      else if (((! scfarg_0_1_argbuf_r) && (! scfarg_0_goMux_mux_bufchan_buf[0])))
        scfarg_0_goMux_mux_bufchan_buf <= scfarg_0_goMux_mux_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (t1'aff_3_destruct,Pointer_QTree_Int) > (t1'aff_3_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t \t1'aff_3_destruct_bufchan_d ;
  logic \t1'aff_3_destruct_bufchan_r ;
  assign \t1'aff_3_destruct_r  = ((! \t1'aff_3_destruct_bufchan_d [0]) || \t1'aff_3_destruct_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \t1'aff_3_destruct_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\t1'aff_3_destruct_r )
        \t1'aff_3_destruct_bufchan_d  <= \t1'aff_3_destruct_d ;
  Pointer_QTree_Int_t \t1'aff_3_destruct_bufchan_buf ;
  assign \t1'aff_3_destruct_bufchan_r  = (! \t1'aff_3_destruct_bufchan_buf [0]);
  assign \t1'aff_3_1_argbuf_d  = (\t1'aff_3_destruct_bufchan_buf [0] ? \t1'aff_3_destruct_bufchan_buf  :
                                  \t1'aff_3_destruct_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \t1'aff_3_destruct_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((\t1'aff_3_1_argbuf_r  && \t1'aff_3_destruct_bufchan_buf [0]))
        \t1'aff_3_destruct_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! \t1'aff_3_1_argbuf_r ) && (! \t1'aff_3_destruct_bufchan_buf [0])))
        \t1'aff_3_destruct_bufchan_buf  <= \t1'aff_3_destruct_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Int) : (t1aeG_destruct,Pointer_QTree_Int) > (t1aeG_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t t1aeG_destruct_bufchan_d;
  logic t1aeG_destruct_bufchan_r;
  assign t1aeG_destruct_r = ((! t1aeG_destruct_bufchan_d[0]) || t1aeG_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t1aeG_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (t1aeG_destruct_r) t1aeG_destruct_bufchan_d <= t1aeG_destruct_d;
  Pointer_QTree_Int_t t1aeG_destruct_bufchan_buf;
  assign t1aeG_destruct_bufchan_r = (! t1aeG_destruct_bufchan_buf[0]);
  assign t1aeG_1_argbuf_d = (t1aeG_destruct_bufchan_buf[0] ? t1aeG_destruct_bufchan_buf :
                             t1aeG_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t1aeG_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((t1aeG_1_argbuf_r && t1aeG_destruct_bufchan_buf[0]))
        t1aeG_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! t1aeG_1_argbuf_r) && (! t1aeG_destruct_bufchan_buf[0])))
        t1aeG_destruct_bufchan_buf <= t1aeG_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (t1af5_destruct,Pointer_QTree_Int) > (t1af5_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t t1af5_destruct_bufchan_d;
  logic t1af5_destruct_bufchan_r;
  assign t1af5_destruct_r = ((! t1af5_destruct_bufchan_d[0]) || t1af5_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t1af5_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (t1af5_destruct_r) t1af5_destruct_bufchan_d <= t1af5_destruct_d;
  Pointer_QTree_Int_t t1af5_destruct_bufchan_buf;
  assign t1af5_destruct_bufchan_r = (! t1af5_destruct_bufchan_buf[0]);
  assign t1af5_1_argbuf_d = (t1af5_destruct_bufchan_buf[0] ? t1af5_destruct_bufchan_buf :
                             t1af5_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t1af5_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((t1af5_1_argbuf_r && t1af5_destruct_bufchan_buf[0]))
        t1af5_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! t1af5_1_argbuf_r) && (! t1af5_destruct_bufchan_buf[0])))
        t1af5_destruct_bufchan_buf <= t1af5_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (t1afa_3_destruct,Pointer_QTree_Int) > (t1afa_3_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t t1afa_3_destruct_bufchan_d;
  logic t1afa_3_destruct_bufchan_r;
  assign t1afa_3_destruct_r = ((! t1afa_3_destruct_bufchan_d[0]) || t1afa_3_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t1afa_3_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (t1afa_3_destruct_r)
        t1afa_3_destruct_bufchan_d <= t1afa_3_destruct_d;
  Pointer_QTree_Int_t t1afa_3_destruct_bufchan_buf;
  assign t1afa_3_destruct_bufchan_r = (! t1afa_3_destruct_bufchan_buf[0]);
  assign t1afa_3_1_argbuf_d = (t1afa_3_destruct_bufchan_buf[0] ? t1afa_3_destruct_bufchan_buf :
                               t1afa_3_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t1afa_3_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((t1afa_3_1_argbuf_r && t1afa_3_destruct_bufchan_buf[0]))
        t1afa_3_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! t1afa_3_1_argbuf_r) && (! t1afa_3_destruct_bufchan_buf[0])))
        t1afa_3_destruct_bufchan_buf <= t1afa_3_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (t1afy_3_destruct,Pointer_QTree_Int) > (t1afy_3_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t t1afy_3_destruct_bufchan_d;
  logic t1afy_3_destruct_bufchan_r;
  assign t1afy_3_destruct_r = ((! t1afy_3_destruct_bufchan_d[0]) || t1afy_3_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t1afy_3_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (t1afy_3_destruct_r)
        t1afy_3_destruct_bufchan_d <= t1afy_3_destruct_d;
  Pointer_QTree_Int_t t1afy_3_destruct_bufchan_buf;
  assign t1afy_3_destruct_bufchan_r = (! t1afy_3_destruct_bufchan_buf[0]);
  assign t1afy_3_1_argbuf_d = (t1afy_3_destruct_bufchan_buf[0] ? t1afy_3_destruct_bufchan_buf :
                               t1afy_3_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t1afy_3_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((t1afy_3_1_argbuf_r && t1afy_3_destruct_bufchan_buf[0]))
        t1afy_3_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! t1afy_3_1_argbuf_r) && (! t1afy_3_destruct_bufchan_buf[0])))
        t1afy_3_destruct_bufchan_buf <= t1afy_3_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (t2'afg_2_destruct,Pointer_QTree_Int) > (t2'afg_2_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t \t2'afg_2_destruct_bufchan_d ;
  logic \t2'afg_2_destruct_bufchan_r ;
  assign \t2'afg_2_destruct_r  = ((! \t2'afg_2_destruct_bufchan_d [0]) || \t2'afg_2_destruct_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \t2'afg_2_destruct_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\t2'afg_2_destruct_r )
        \t2'afg_2_destruct_bufchan_d  <= \t2'afg_2_destruct_d ;
  Pointer_QTree_Int_t \t2'afg_2_destruct_bufchan_buf ;
  assign \t2'afg_2_destruct_bufchan_r  = (! \t2'afg_2_destruct_bufchan_buf [0]);
  assign \t2'afg_2_1_argbuf_d  = (\t2'afg_2_destruct_bufchan_buf [0] ? \t2'afg_2_destruct_bufchan_buf  :
                                  \t2'afg_2_destruct_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \t2'afg_2_destruct_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((\t2'afg_2_1_argbuf_r  && \t2'afg_2_destruct_bufchan_buf [0]))
        \t2'afg_2_destruct_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! \t2'afg_2_1_argbuf_r ) && (! \t2'afg_2_destruct_bufchan_buf [0])))
        \t2'afg_2_destruct_bufchan_buf  <= \t2'afg_2_destruct_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Int) : (t2aeH_destruct,Pointer_QTree_Int) > (t2aeH_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t t2aeH_destruct_bufchan_d;
  logic t2aeH_destruct_bufchan_r;
  assign t2aeH_destruct_r = ((! t2aeH_destruct_bufchan_d[0]) || t2aeH_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t2aeH_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (t2aeH_destruct_r) t2aeH_destruct_bufchan_d <= t2aeH_destruct_d;
  Pointer_QTree_Int_t t2aeH_destruct_bufchan_buf;
  assign t2aeH_destruct_bufchan_r = (! t2aeH_destruct_bufchan_buf[0]);
  assign t2aeH_1_argbuf_d = (t2aeH_destruct_bufchan_buf[0] ? t2aeH_destruct_bufchan_buf :
                             t2aeH_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t2aeH_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((t2aeH_1_argbuf_r && t2aeH_destruct_bufchan_buf[0]))
        t2aeH_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! t2aeH_1_argbuf_r) && (! t2aeH_destruct_bufchan_buf[0])))
        t2aeH_destruct_bufchan_buf <= t2aeH_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (t2af6_destruct,Pointer_QTree_Int) > (t2af6_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t t2af6_destruct_bufchan_d;
  logic t2af6_destruct_bufchan_r;
  assign t2af6_destruct_r = ((! t2af6_destruct_bufchan_d[0]) || t2af6_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t2af6_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (t2af6_destruct_r) t2af6_destruct_bufchan_d <= t2af6_destruct_d;
  Pointer_QTree_Int_t t2af6_destruct_bufchan_buf;
  assign t2af6_destruct_bufchan_r = (! t2af6_destruct_bufchan_buf[0]);
  assign t2af6_1_argbuf_d = (t2af6_destruct_bufchan_buf[0] ? t2af6_destruct_bufchan_buf :
                             t2af6_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t2af6_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((t2af6_1_argbuf_r && t2af6_destruct_bufchan_buf[0]))
        t2af6_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! t2af6_1_argbuf_r) && (! t2af6_destruct_bufchan_buf[0])))
        t2af6_destruct_bufchan_buf <= t2af6_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (t2afb_2_destruct,Pointer_QTree_Int) > (t2afb_2_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t t2afb_2_destruct_bufchan_d;
  logic t2afb_2_destruct_bufchan_r;
  assign t2afb_2_destruct_r = ((! t2afb_2_destruct_bufchan_d[0]) || t2afb_2_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t2afb_2_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (t2afb_2_destruct_r)
        t2afb_2_destruct_bufchan_d <= t2afb_2_destruct_d;
  Pointer_QTree_Int_t t2afb_2_destruct_bufchan_buf;
  assign t2afb_2_destruct_bufchan_r = (! t2afb_2_destruct_bufchan_buf[0]);
  assign t2afb_2_1_argbuf_d = (t2afb_2_destruct_bufchan_buf[0] ? t2afb_2_destruct_bufchan_buf :
                               t2afb_2_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t2afb_2_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((t2afb_2_1_argbuf_r && t2afb_2_destruct_bufchan_buf[0]))
        t2afb_2_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! t2afb_2_1_argbuf_r) && (! t2afb_2_destruct_bufchan_buf[0])))
        t2afb_2_destruct_bufchan_buf <= t2afb_2_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (t2afz_2_destruct,Pointer_QTree_Int) > (t2afz_2_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t t2afz_2_destruct_bufchan_d;
  logic t2afz_2_destruct_bufchan_r;
  assign t2afz_2_destruct_r = ((! t2afz_2_destruct_bufchan_d[0]) || t2afz_2_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t2afz_2_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (t2afz_2_destruct_r)
        t2afz_2_destruct_bufchan_d <= t2afz_2_destruct_d;
  Pointer_QTree_Int_t t2afz_2_destruct_bufchan_buf;
  assign t2afz_2_destruct_bufchan_r = (! t2afz_2_destruct_bufchan_buf[0]);
  assign t2afz_2_1_argbuf_d = (t2afz_2_destruct_bufchan_buf[0] ? t2afz_2_destruct_bufchan_buf :
                               t2afz_2_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t2afz_2_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((t2afz_2_1_argbuf_r && t2afz_2_destruct_bufchan_buf[0]))
        t2afz_2_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! t2afz_2_1_argbuf_r) && (! t2afz_2_destruct_bufchan_buf[0])))
        t2afz_2_destruct_bufchan_buf <= t2afz_2_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (t3'afh_1_destruct,Pointer_QTree_Int) > (t3'afh_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t \t3'afh_1_destruct_bufchan_d ;
  logic \t3'afh_1_destruct_bufchan_r ;
  assign \t3'afh_1_destruct_r  = ((! \t3'afh_1_destruct_bufchan_d [0]) || \t3'afh_1_destruct_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \t3'afh_1_destruct_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\t3'afh_1_destruct_r )
        \t3'afh_1_destruct_bufchan_d  <= \t3'afh_1_destruct_d ;
  Pointer_QTree_Int_t \t3'afh_1_destruct_bufchan_buf ;
  assign \t3'afh_1_destruct_bufchan_r  = (! \t3'afh_1_destruct_bufchan_buf [0]);
  assign \t3'afh_1_1_argbuf_d  = (\t3'afh_1_destruct_bufchan_buf [0] ? \t3'afh_1_destruct_bufchan_buf  :
                                  \t3'afh_1_destruct_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \t3'afh_1_destruct_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((\t3'afh_1_1_argbuf_r  && \t3'afh_1_destruct_bufchan_buf [0]))
        \t3'afh_1_destruct_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! \t3'afh_1_1_argbuf_r ) && (! \t3'afh_1_destruct_bufchan_buf [0])))
        \t3'afh_1_destruct_bufchan_buf  <= \t3'afh_1_destruct_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Int) : (t3aeI_destruct,Pointer_QTree_Int) > (t3aeI_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t t3aeI_destruct_bufchan_d;
  logic t3aeI_destruct_bufchan_r;
  assign t3aeI_destruct_r = ((! t3aeI_destruct_bufchan_d[0]) || t3aeI_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t3aeI_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (t3aeI_destruct_r) t3aeI_destruct_bufchan_d <= t3aeI_destruct_d;
  Pointer_QTree_Int_t t3aeI_destruct_bufchan_buf;
  assign t3aeI_destruct_bufchan_r = (! t3aeI_destruct_bufchan_buf[0]);
  assign t3aeI_1_argbuf_d = (t3aeI_destruct_bufchan_buf[0] ? t3aeI_destruct_bufchan_buf :
                             t3aeI_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t3aeI_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((t3aeI_1_argbuf_r && t3aeI_destruct_bufchan_buf[0]))
        t3aeI_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! t3aeI_1_argbuf_r) && (! t3aeI_destruct_bufchan_buf[0])))
        t3aeI_destruct_bufchan_buf <= t3aeI_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (t3af7_destruct,Pointer_QTree_Int) > (t3af7_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t t3af7_destruct_bufchan_d;
  logic t3af7_destruct_bufchan_r;
  assign t3af7_destruct_r = ((! t3af7_destruct_bufchan_d[0]) || t3af7_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t3af7_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (t3af7_destruct_r) t3af7_destruct_bufchan_d <= t3af7_destruct_d;
  Pointer_QTree_Int_t t3af7_destruct_bufchan_buf;
  assign t3af7_destruct_bufchan_r = (! t3af7_destruct_bufchan_buf[0]);
  assign t3af7_1_argbuf_d = (t3af7_destruct_bufchan_buf[0] ? t3af7_destruct_bufchan_buf :
                             t3af7_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t3af7_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((t3af7_1_argbuf_r && t3af7_destruct_bufchan_buf[0]))
        t3af7_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! t3af7_1_argbuf_r) && (! t3af7_destruct_bufchan_buf[0])))
        t3af7_destruct_bufchan_buf <= t3af7_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (t3afA_1_destruct,Pointer_QTree_Int) > (t3afA_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t t3afA_1_destruct_bufchan_d;
  logic t3afA_1_destruct_bufchan_r;
  assign t3afA_1_destruct_r = ((! t3afA_1_destruct_bufchan_d[0]) || t3afA_1_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t3afA_1_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (t3afA_1_destruct_r)
        t3afA_1_destruct_bufchan_d <= t3afA_1_destruct_d;
  Pointer_QTree_Int_t t3afA_1_destruct_bufchan_buf;
  assign t3afA_1_destruct_bufchan_r = (! t3afA_1_destruct_bufchan_buf[0]);
  assign t3afA_1_1_argbuf_d = (t3afA_1_destruct_bufchan_buf[0] ? t3afA_1_destruct_bufchan_buf :
                               t3afA_1_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t3afA_1_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((t3afA_1_1_argbuf_r && t3afA_1_destruct_bufchan_buf[0]))
        t3afA_1_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! t3afA_1_1_argbuf_r) && (! t3afA_1_destruct_bufchan_buf[0])))
        t3afA_1_destruct_bufchan_buf <= t3afA_1_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (t3afc_1_destruct,Pointer_QTree_Int) > (t3afc_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t t3afc_1_destruct_bufchan_d;
  logic t3afc_1_destruct_bufchan_r;
  assign t3afc_1_destruct_r = ((! t3afc_1_destruct_bufchan_d[0]) || t3afc_1_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t3afc_1_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (t3afc_1_destruct_r)
        t3afc_1_destruct_bufchan_d <= t3afc_1_destruct_d;
  Pointer_QTree_Int_t t3afc_1_destruct_bufchan_buf;
  assign t3afc_1_destruct_bufchan_r = (! t3afc_1_destruct_bufchan_buf[0]);
  assign t3afc_1_1_argbuf_d = (t3afc_1_destruct_bufchan_buf[0] ? t3afc_1_destruct_bufchan_buf :
                               t3afc_1_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t3afc_1_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((t3afc_1_1_argbuf_r && t3afc_1_destruct_bufchan_buf[0]))
        t3afc_1_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! t3afc_1_1_argbuf_r) && (! t3afc_1_destruct_bufchan_buf[0])))
        t3afc_1_destruct_bufchan_buf <= t3afc_1_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (t4'afi_destruct,Pointer_QTree_Int) > (t4'afi_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t \t4'afi_destruct_bufchan_d ;
  logic \t4'afi_destruct_bufchan_r ;
  assign \t4'afi_destruct_r  = ((! \t4'afi_destruct_bufchan_d [0]) || \t4'afi_destruct_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \t4'afi_destruct_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\t4'afi_destruct_r )
        \t4'afi_destruct_bufchan_d  <= \t4'afi_destruct_d ;
  Pointer_QTree_Int_t \t4'afi_destruct_bufchan_buf ;
  assign \t4'afi_destruct_bufchan_r  = (! \t4'afi_destruct_bufchan_buf [0]);
  assign \t4'afi_1_argbuf_d  = (\t4'afi_destruct_bufchan_buf [0] ? \t4'afi_destruct_bufchan_buf  :
                                \t4'afi_destruct_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \t4'afi_destruct_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((\t4'afi_1_argbuf_r  && \t4'afi_destruct_bufchan_buf [0]))
        \t4'afi_destruct_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! \t4'afi_1_argbuf_r ) && (! \t4'afi_destruct_bufchan_buf [0])))
        \t4'afi_destruct_bufchan_buf  <= \t4'afi_destruct_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Int) : (t4aeJ_destruct,Pointer_QTree_Int) > (t4aeJ_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t t4aeJ_destruct_bufchan_d;
  logic t4aeJ_destruct_bufchan_r;
  assign t4aeJ_destruct_r = ((! t4aeJ_destruct_bufchan_d[0]) || t4aeJ_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t4aeJ_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (t4aeJ_destruct_r) t4aeJ_destruct_bufchan_d <= t4aeJ_destruct_d;
  Pointer_QTree_Int_t t4aeJ_destruct_bufchan_buf;
  assign t4aeJ_destruct_bufchan_r = (! t4aeJ_destruct_bufchan_buf[0]);
  assign t4aeJ_1_argbuf_d = (t4aeJ_destruct_bufchan_buf[0] ? t4aeJ_destruct_bufchan_buf :
                             t4aeJ_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t4aeJ_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((t4aeJ_1_argbuf_r && t4aeJ_destruct_bufchan_buf[0]))
        t4aeJ_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! t4aeJ_1_argbuf_r) && (! t4aeJ_destruct_bufchan_buf[0])))
        t4aeJ_destruct_bufchan_buf <= t4aeJ_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (t4af8_destruct,Pointer_QTree_Int) > (t4af8_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t t4af8_destruct_bufchan_d;
  logic t4af8_destruct_bufchan_r;
  assign t4af8_destruct_r = ((! t4af8_destruct_bufchan_d[0]) || t4af8_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t4af8_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (t4af8_destruct_r) t4af8_destruct_bufchan_d <= t4af8_destruct_d;
  Pointer_QTree_Int_t t4af8_destruct_bufchan_buf;
  assign t4af8_destruct_bufchan_r = (! t4af8_destruct_bufchan_buf[0]);
  assign t4af8_1_argbuf_d = (t4af8_destruct_bufchan_buf[0] ? t4af8_destruct_bufchan_buf :
                             t4af8_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t4af8_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((t4af8_1_argbuf_r && t4af8_destruct_bufchan_buf[0]))
        t4af8_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! t4af8_1_argbuf_r) && (! t4af8_destruct_bufchan_buf[0])))
        t4af8_destruct_bufchan_buf <= t4af8_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (t4afk_1,Pointer_QTree_Int) > (t4afk_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t t4afk_1_bufchan_d;
  logic t4afk_1_bufchan_r;
  assign t4afk_1_r = ((! t4afk_1_bufchan_d[0]) || t4afk_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t4afk_1_bufchan_d <= {16'd0, 1'd0};
    else if (t4afk_1_r) t4afk_1_bufchan_d <= t4afk_1_d;
  Pointer_QTree_Int_t t4afk_1_bufchan_buf;
  assign t4afk_1_bufchan_r = (! t4afk_1_bufchan_buf[0]);
  assign t4afk_1_argbuf_d = (t4afk_1_bufchan_buf[0] ? t4afk_1_bufchan_buf :
                             t4afk_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t4afk_1_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((t4afk_1_argbuf_r && t4afk_1_bufchan_buf[0]))
        t4afk_1_bufchan_buf <= {16'd0, 1'd0};
      else if (((! t4afk_1_argbuf_r) && (! t4afk_1_bufchan_buf[0])))
        t4afk_1_bufchan_buf <= t4afk_1_bufchan_d;
  
  /* fork (Ty Pointer_QTree_Int) : (t4afk_goMux_mux,Pointer_QTree_Int) > [(t4afk_1,Pointer_QTree_Int),
                                                                     (t4afk_2,Pointer_QTree_Int)] */
  logic [1:0] t4afk_goMux_mux_emitted;
  logic [1:0] t4afk_goMux_mux_done;
  assign t4afk_1_d = {t4afk_goMux_mux_d[16:1],
                      (t4afk_goMux_mux_d[0] && (! t4afk_goMux_mux_emitted[0]))};
  assign t4afk_2_d = {t4afk_goMux_mux_d[16:1],
                      (t4afk_goMux_mux_d[0] && (! t4afk_goMux_mux_emitted[1]))};
  assign t4afk_goMux_mux_done = (t4afk_goMux_mux_emitted | ({t4afk_2_d[0],
                                                             t4afk_1_d[0]} & {t4afk_2_r,
                                                                              t4afk_1_r}));
  assign t4afk_goMux_mux_r = (& t4afk_goMux_mux_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t4afk_goMux_mux_emitted <= 2'd0;
    else
      t4afk_goMux_mux_emitted <= (t4afk_goMux_mux_r ? 2'd0 :
                                  t4afk_goMux_mux_done);
  
  /* buf (Ty Pointer_QTree_Int) : (t5afB_destruct,Pointer_QTree_Int) > (t5afB_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t t5afB_destruct_bufchan_d;
  logic t5afB_destruct_bufchan_r;
  assign t5afB_destruct_r = ((! t5afB_destruct_bufchan_d[0]) || t5afB_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t5afB_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (t5afB_destruct_r) t5afB_destruct_bufchan_d <= t5afB_destruct_d;
  Pointer_QTree_Int_t t5afB_destruct_bufchan_buf;
  assign t5afB_destruct_bufchan_r = (! t5afB_destruct_bufchan_buf[0]);
  assign t5afB_1_argbuf_d = (t5afB_destruct_bufchan_buf[0] ? t5afB_destruct_bufchan_buf :
                             t5afB_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t5afB_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((t5afB_1_argbuf_r && t5afB_destruct_bufchan_buf[0]))
        t5afB_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! t5afB_1_argbuf_r) && (! t5afB_destruct_bufchan_buf[0])))
        t5afB_destruct_bufchan_buf <= t5afB_destruct_bufchan_d;
  
  /* buf (Ty Int) : (v'aeR_1,Int) > (v'aeR_1_argbuf,Int) */
  Int_t \v'aeR_1_bufchan_d ;
  logic \v'aeR_1_bufchan_r ;
  assign \v'aeR_1_r  = ((! \v'aeR_1_bufchan_d [0]) || \v'aeR_1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \v'aeR_1_bufchan_d  <= {32'd0, 1'd0};
    else if (\v'aeR_1_r ) \v'aeR_1_bufchan_d  <= \v'aeR_1_d ;
  Int_t \v'aeR_1_bufchan_buf ;
  assign \v'aeR_1_bufchan_r  = (! \v'aeR_1_bufchan_buf [0]);
  assign \v'aeR_1_argbuf_d  = (\v'aeR_1_bufchan_buf [0] ? \v'aeR_1_bufchan_buf  :
                               \v'aeR_1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \v'aeR_1_bufchan_buf  <= {32'd0, 1'd0};
    else
      if ((\v'aeR_1_argbuf_r  && \v'aeR_1_bufchan_buf [0]))
        \v'aeR_1_bufchan_buf  <= {32'd0, 1'd0};
      else if (((! \v'aeR_1_argbuf_r ) && (! \v'aeR_1_bufchan_buf [0])))
        \v'aeR_1_bufchan_buf  <= \v'aeR_1_bufchan_d ;
  
  /* fork (Ty Int) : (v'aeR_destruct,Int) > [(v'aeR_1,Int),
                                        (v'aeR_2,Int)] */
  logic [1:0] \v'aeR_destruct_emitted ;
  logic [1:0] \v'aeR_destruct_done ;
  assign \v'aeR_1_d  = {\v'aeR_destruct_d [32:1],
                        (\v'aeR_destruct_d [0] && (! \v'aeR_destruct_emitted [0]))};
  assign \v'aeR_2_d  = {\v'aeR_destruct_d [32:1],
                        (\v'aeR_destruct_d [0] && (! \v'aeR_destruct_emitted [1]))};
  assign \v'aeR_destruct_done  = (\v'aeR_destruct_emitted  | ({\v'aeR_2_d [0],
                                                               \v'aeR_1_d [0]} & {\v'aeR_2_r ,
                                                                                  \v'aeR_1_r }));
  assign \v'aeR_destruct_r  = (& \v'aeR_destruct_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \v'aeR_destruct_emitted  <= 2'd0;
    else
      \v'aeR_destruct_emitted  <= (\v'aeR_destruct_r  ? 2'd0 :
                                   \v'aeR_destruct_done );
  
  /* buf (Ty Int) : (vaeL_1,Int) > (vaeL_1_argbuf,Int) */
  Int_t vaeL_1_bufchan_d;
  logic vaeL_1_bufchan_r;
  assign vaeL_1_r = ((! vaeL_1_bufchan_d[0]) || vaeL_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) vaeL_1_bufchan_d <= {32'd0, 1'd0};
    else if (vaeL_1_r) vaeL_1_bufchan_d <= vaeL_1_d;
  Int_t vaeL_1_bufchan_buf;
  assign vaeL_1_bufchan_r = (! vaeL_1_bufchan_buf[0]);
  assign vaeL_1_argbuf_d = (vaeL_1_bufchan_buf[0] ? vaeL_1_bufchan_buf :
                            vaeL_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) vaeL_1_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((vaeL_1_argbuf_r && vaeL_1_bufchan_buf[0]))
        vaeL_1_bufchan_buf <= {32'd0, 1'd0};
      else if (((! vaeL_1_argbuf_r) && (! vaeL_1_bufchan_buf[0])))
        vaeL_1_bufchan_buf <= vaeL_1_bufchan_d;
  
  /* fork (Ty Int) : (vaeL_destruct,Int) > [(vaeL_1,Int),(vaeL_2,Int)] */
  logic [1:0] vaeL_destruct_emitted;
  logic [1:0] vaeL_destruct_done;
  assign vaeL_1_d = {vaeL_destruct_d[32:1],
                     (vaeL_destruct_d[0] && (! vaeL_destruct_emitted[0]))};
  assign vaeL_2_d = {vaeL_destruct_d[32:1],
                     (vaeL_destruct_d[0] && (! vaeL_destruct_emitted[1]))};
  assign vaeL_destruct_done = (vaeL_destruct_emitted | ({vaeL_2_d[0],
                                                         vaeL_1_d[0]} & {vaeL_2_r, vaeL_1_r}));
  assign vaeL_destruct_r = (& vaeL_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) vaeL_destruct_emitted <= 2'd0;
    else
      vaeL_destruct_emitted <= (vaeL_destruct_r ? 2'd0 :
                                vaeL_destruct_done);
  
  /* buf (Ty Int) : (vaeQ_1,Int) > (vaeQ_1_argbuf,Int) */
  Int_t vaeQ_1_bufchan_d;
  logic vaeQ_1_bufchan_r;
  assign vaeQ_1_r = ((! vaeQ_1_bufchan_d[0]) || vaeQ_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) vaeQ_1_bufchan_d <= {32'd0, 1'd0};
    else if (vaeQ_1_r) vaeQ_1_bufchan_d <= vaeQ_1_d;
  Int_t vaeQ_1_bufchan_buf;
  assign vaeQ_1_bufchan_r = (! vaeQ_1_bufchan_buf[0]);
  assign vaeQ_1_argbuf_d = (vaeQ_1_bufchan_buf[0] ? vaeQ_1_bufchan_buf :
                            vaeQ_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) vaeQ_1_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((vaeQ_1_argbuf_r && vaeQ_1_bufchan_buf[0]))
        vaeQ_1_bufchan_buf <= {32'd0, 1'd0};
      else if (((! vaeQ_1_argbuf_r) && (! vaeQ_1_bufchan_buf[0])))
        vaeQ_1_bufchan_buf <= vaeQ_1_bufchan_d;
  
  /* fork (Ty Int) : (vaeQ_destruct,Int) > [(vaeQ_1,Int),(vaeQ_2,Int)] */
  logic [1:0] vaeQ_destruct_emitted;
  logic [1:0] vaeQ_destruct_done;
  assign vaeQ_1_d = {vaeQ_destruct_d[32:1],
                     (vaeQ_destruct_d[0] && (! vaeQ_destruct_emitted[0]))};
  assign vaeQ_2_d = {vaeQ_destruct_d[32:1],
                     (vaeQ_destruct_d[0] && (! vaeQ_destruct_emitted[1]))};
  assign vaeQ_destruct_done = (vaeQ_destruct_emitted | ({vaeQ_2_d[0],
                                                         vaeQ_1_d[0]} & {vaeQ_2_r, vaeQ_1_r}));
  assign vaeQ_destruct_r = (& vaeQ_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) vaeQ_destruct_emitted <= 2'd0;
    else
      vaeQ_destruct_emitted <= (vaeQ_destruct_r ? 2'd0 :
                                vaeQ_destruct_done);
  
  /* buf (Ty Int) : (vaew_1,Int) > (vaew_1_argbuf,Int) */
  Int_t vaew_1_bufchan_d;
  logic vaew_1_bufchan_r;
  assign vaew_1_r = ((! vaew_1_bufchan_d[0]) || vaew_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) vaew_1_bufchan_d <= {32'd0, 1'd0};
    else if (vaew_1_r) vaew_1_bufchan_d <= vaew_1_d;
  Int_t vaew_1_bufchan_buf;
  assign vaew_1_bufchan_r = (! vaew_1_bufchan_buf[0]);
  assign vaew_1_argbuf_d = (vaew_1_bufchan_buf[0] ? vaew_1_bufchan_buf :
                            vaew_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) vaew_1_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((vaew_1_argbuf_r && vaew_1_bufchan_buf[0]))
        vaew_1_bufchan_buf <= {32'd0, 1'd0};
      else if (((! vaew_1_argbuf_r) && (! vaew_1_bufchan_buf[0])))
        vaew_1_bufchan_buf <= vaew_1_bufchan_d;
  
  /* fork (Ty Int) : (vaew_destruct,Int) > [(vaew_1,Int),(vaew_2,Int)] */
  logic [1:0] vaew_destruct_emitted;
  logic [1:0] vaew_destruct_done;
  assign vaew_1_d = {vaew_destruct_d[32:1],
                     (vaew_destruct_d[0] && (! vaew_destruct_emitted[0]))};
  assign vaew_2_d = {vaew_destruct_d[32:1],
                     (vaew_destruct_d[0] && (! vaew_destruct_emitted[1]))};
  assign vaew_destruct_done = (vaew_destruct_emitted | ({vaew_2_d[0],
                                                         vaew_1_d[0]} & {vaew_2_r, vaew_1_r}));
  assign vaew_destruct_r = (& vaew_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) vaew_destruct_emitted <= 2'd0;
    else
      vaew_destruct_emitted <= (vaew_destruct_r ? 2'd0 :
                                vaew_destruct_done);
  
  /* buf (Ty Int) : (vafo_1,Int) > (vafo_1_argbuf,Int) */
  Int_t vafo_1_bufchan_d;
  logic vafo_1_bufchan_r;
  assign vafo_1_r = ((! vafo_1_bufchan_d[0]) || vafo_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) vafo_1_bufchan_d <= {32'd0, 1'd0};
    else if (vafo_1_r) vafo_1_bufchan_d <= vafo_1_d;
  Int_t vafo_1_bufchan_buf;
  assign vafo_1_bufchan_r = (! vafo_1_bufchan_buf[0]);
  assign vafo_1_argbuf_d = (vafo_1_bufchan_buf[0] ? vafo_1_bufchan_buf :
                            vafo_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) vafo_1_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((vafo_1_argbuf_r && vafo_1_bufchan_buf[0]))
        vafo_1_bufchan_buf <= {32'd0, 1'd0};
      else if (((! vafo_1_argbuf_r) && (! vafo_1_bufchan_buf[0])))
        vafo_1_bufchan_buf <= vafo_1_bufchan_d;
  
  /* fork (Ty Int) : (vafo_destruct,Int) > [(vafo_1,Int),(vafo_2,Int)] */
  logic [1:0] vafo_destruct_emitted;
  logic [1:0] vafo_destruct_done;
  assign vafo_1_d = {vafo_destruct_d[32:1],
                     (vafo_destruct_d[0] && (! vafo_destruct_emitted[0]))};
  assign vafo_2_d = {vafo_destruct_d[32:1],
                     (vafo_destruct_d[0] && (! vafo_destruct_emitted[1]))};
  assign vafo_destruct_done = (vafo_destruct_emitted | ({vafo_2_d[0],
                                                         vafo_1_d[0]} & {vafo_2_r, vafo_1_r}));
  assign vafo_destruct_r = (& vafo_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) vafo_destruct_emitted <= 2'd0;
    else
      vafo_destruct_emitted <= (vafo_destruct_r ? 2'd0 :
                                vafo_destruct_done);
  
  /* buf (Ty Pointer_CT$wnnz) : (writeCT$wnnzlizzieLet0_1_argbuf,Pointer_CT$wnnz) > (writeCT$wnnzlizzieLet0_1_argbuf_rwb,Pointer_CT$wnnz) */
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet0_1_argbuf_bufchan_d;
  logic writeCT$wnnzlizzieLet0_1_argbuf_bufchan_r;
  assign writeCT$wnnzlizzieLet0_1_argbuf_r = ((! writeCT$wnnzlizzieLet0_1_argbuf_bufchan_d[0]) || writeCT$wnnzlizzieLet0_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnzlizzieLet0_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCT$wnnzlizzieLet0_1_argbuf_r)
        writeCT$wnnzlizzieLet0_1_argbuf_bufchan_d <= writeCT$wnnzlizzieLet0_1_argbuf_d;
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet0_1_argbuf_bufchan_buf;
  assign writeCT$wnnzlizzieLet0_1_argbuf_bufchan_r = (! writeCT$wnnzlizzieLet0_1_argbuf_bufchan_buf[0]);
  assign writeCT$wnnzlizzieLet0_1_argbuf_rwb_d = (writeCT$wnnzlizzieLet0_1_argbuf_bufchan_buf[0] ? writeCT$wnnzlizzieLet0_1_argbuf_bufchan_buf :
                                                  writeCT$wnnzlizzieLet0_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnzlizzieLet0_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeCT$wnnzlizzieLet0_1_argbuf_rwb_r && writeCT$wnnzlizzieLet0_1_argbuf_bufchan_buf[0]))
        writeCT$wnnzlizzieLet0_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeCT$wnnzlizzieLet0_1_argbuf_rwb_r) && (! writeCT$wnnzlizzieLet0_1_argbuf_bufchan_buf[0])))
        writeCT$wnnzlizzieLet0_1_argbuf_bufchan_buf <= writeCT$wnnzlizzieLet0_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz) : (writeCT$wnnzlizzieLet0_1_argbuf_rwb,Pointer_CT$wnnz) > (lizzieLet39_1_argbuf,Pointer_CT$wnnz) */
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet0_1_argbuf_rwb_bufchan_d;
  logic writeCT$wnnzlizzieLet0_1_argbuf_rwb_bufchan_r;
  assign writeCT$wnnzlizzieLet0_1_argbuf_rwb_r = ((! writeCT$wnnzlizzieLet0_1_argbuf_rwb_bufchan_d[0]) || writeCT$wnnzlizzieLet0_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnzlizzieLet0_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCT$wnnzlizzieLet0_1_argbuf_rwb_r)
        writeCT$wnnzlizzieLet0_1_argbuf_rwb_bufchan_d <= writeCT$wnnzlizzieLet0_1_argbuf_rwb_d;
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet0_1_argbuf_rwb_bufchan_buf;
  assign writeCT$wnnzlizzieLet0_1_argbuf_rwb_bufchan_r = (! writeCT$wnnzlizzieLet0_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet39_1_argbuf_d = (writeCT$wnnzlizzieLet0_1_argbuf_rwb_bufchan_buf[0] ? writeCT$wnnzlizzieLet0_1_argbuf_rwb_bufchan_buf :
                                   writeCT$wnnzlizzieLet0_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnzlizzieLet0_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet39_1_argbuf_r && writeCT$wnnzlizzieLet0_1_argbuf_rwb_bufchan_buf[0]))
        writeCT$wnnzlizzieLet0_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet39_1_argbuf_r) && (! writeCT$wnnzlizzieLet0_1_argbuf_rwb_bufchan_buf[0])))
        writeCT$wnnzlizzieLet0_1_argbuf_rwb_bufchan_buf <= writeCT$wnnzlizzieLet0_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz) : (writeCT$wnnzlizzieLet59_1_argbuf,Pointer_CT$wnnz) > (writeCT$wnnzlizzieLet59_1_argbuf_rwb,Pointer_CT$wnnz) */
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet59_1_argbuf_bufchan_d;
  logic writeCT$wnnzlizzieLet59_1_argbuf_bufchan_r;
  assign writeCT$wnnzlizzieLet59_1_argbuf_r = ((! writeCT$wnnzlizzieLet59_1_argbuf_bufchan_d[0]) || writeCT$wnnzlizzieLet59_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnzlizzieLet59_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCT$wnnzlizzieLet59_1_argbuf_r)
        writeCT$wnnzlizzieLet59_1_argbuf_bufchan_d <= writeCT$wnnzlizzieLet59_1_argbuf_d;
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet59_1_argbuf_bufchan_buf;
  assign writeCT$wnnzlizzieLet59_1_argbuf_bufchan_r = (! writeCT$wnnzlizzieLet59_1_argbuf_bufchan_buf[0]);
  assign writeCT$wnnzlizzieLet59_1_argbuf_rwb_d = (writeCT$wnnzlizzieLet59_1_argbuf_bufchan_buf[0] ? writeCT$wnnzlizzieLet59_1_argbuf_bufchan_buf :
                                                   writeCT$wnnzlizzieLet59_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnzlizzieLet59_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeCT$wnnzlizzieLet59_1_argbuf_rwb_r && writeCT$wnnzlizzieLet59_1_argbuf_bufchan_buf[0]))
        writeCT$wnnzlizzieLet59_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeCT$wnnzlizzieLet59_1_argbuf_rwb_r) && (! writeCT$wnnzlizzieLet59_1_argbuf_bufchan_buf[0])))
        writeCT$wnnzlizzieLet59_1_argbuf_bufchan_buf <= writeCT$wnnzlizzieLet59_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz) : (writeCT$wnnzlizzieLet59_1_argbuf_rwb,Pointer_CT$wnnz) > (sca2_1_argbuf,Pointer_CT$wnnz) */
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet59_1_argbuf_rwb_bufchan_d;
  logic writeCT$wnnzlizzieLet59_1_argbuf_rwb_bufchan_r;
  assign writeCT$wnnzlizzieLet59_1_argbuf_rwb_r = ((! writeCT$wnnzlizzieLet59_1_argbuf_rwb_bufchan_d[0]) || writeCT$wnnzlizzieLet59_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnzlizzieLet59_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCT$wnnzlizzieLet59_1_argbuf_rwb_r)
        writeCT$wnnzlizzieLet59_1_argbuf_rwb_bufchan_d <= writeCT$wnnzlizzieLet59_1_argbuf_rwb_d;
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet59_1_argbuf_rwb_bufchan_buf;
  assign writeCT$wnnzlizzieLet59_1_argbuf_rwb_bufchan_r = (! writeCT$wnnzlizzieLet59_1_argbuf_rwb_bufchan_buf[0]);
  assign sca2_1_argbuf_d = (writeCT$wnnzlizzieLet59_1_argbuf_rwb_bufchan_buf[0] ? writeCT$wnnzlizzieLet59_1_argbuf_rwb_bufchan_buf :
                            writeCT$wnnzlizzieLet59_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnzlizzieLet59_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((sca2_1_argbuf_r && writeCT$wnnzlizzieLet59_1_argbuf_rwb_bufchan_buf[0]))
        writeCT$wnnzlizzieLet59_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
      else if (((! sca2_1_argbuf_r) && (! writeCT$wnnzlizzieLet59_1_argbuf_rwb_bufchan_buf[0])))
        writeCT$wnnzlizzieLet59_1_argbuf_rwb_bufchan_buf <= writeCT$wnnzlizzieLet59_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz) : (writeCT$wnnzlizzieLet5_1_argbuf,Pointer_CT$wnnz) > (writeCT$wnnzlizzieLet5_1_argbuf_rwb,Pointer_CT$wnnz) */
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet5_1_argbuf_bufchan_d;
  logic writeCT$wnnzlizzieLet5_1_argbuf_bufchan_r;
  assign writeCT$wnnzlizzieLet5_1_argbuf_r = ((! writeCT$wnnzlizzieLet5_1_argbuf_bufchan_d[0]) || writeCT$wnnzlizzieLet5_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnzlizzieLet5_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCT$wnnzlizzieLet5_1_argbuf_r)
        writeCT$wnnzlizzieLet5_1_argbuf_bufchan_d <= writeCT$wnnzlizzieLet5_1_argbuf_d;
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet5_1_argbuf_bufchan_buf;
  assign writeCT$wnnzlizzieLet5_1_argbuf_bufchan_r = (! writeCT$wnnzlizzieLet5_1_argbuf_bufchan_buf[0]);
  assign writeCT$wnnzlizzieLet5_1_argbuf_rwb_d = (writeCT$wnnzlizzieLet5_1_argbuf_bufchan_buf[0] ? writeCT$wnnzlizzieLet5_1_argbuf_bufchan_buf :
                                                  writeCT$wnnzlizzieLet5_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnzlizzieLet5_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeCT$wnnzlizzieLet5_1_argbuf_rwb_r && writeCT$wnnzlizzieLet5_1_argbuf_bufchan_buf[0]))
        writeCT$wnnzlizzieLet5_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeCT$wnnzlizzieLet5_1_argbuf_rwb_r) && (! writeCT$wnnzlizzieLet5_1_argbuf_bufchan_buf[0])))
        writeCT$wnnzlizzieLet5_1_argbuf_bufchan_buf <= writeCT$wnnzlizzieLet5_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz) : (writeCT$wnnzlizzieLet5_1_argbuf_rwb,Pointer_CT$wnnz) > (sca3_1_argbuf,Pointer_CT$wnnz) */
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet5_1_argbuf_rwb_bufchan_d;
  logic writeCT$wnnzlizzieLet5_1_argbuf_rwb_bufchan_r;
  assign writeCT$wnnzlizzieLet5_1_argbuf_rwb_r = ((! writeCT$wnnzlizzieLet5_1_argbuf_rwb_bufchan_d[0]) || writeCT$wnnzlizzieLet5_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnzlizzieLet5_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCT$wnnzlizzieLet5_1_argbuf_rwb_r)
        writeCT$wnnzlizzieLet5_1_argbuf_rwb_bufchan_d <= writeCT$wnnzlizzieLet5_1_argbuf_rwb_d;
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet5_1_argbuf_rwb_bufchan_buf;
  assign writeCT$wnnzlizzieLet5_1_argbuf_rwb_bufchan_r = (! writeCT$wnnzlizzieLet5_1_argbuf_rwb_bufchan_buf[0]);
  assign sca3_1_argbuf_d = (writeCT$wnnzlizzieLet5_1_argbuf_rwb_bufchan_buf[0] ? writeCT$wnnzlizzieLet5_1_argbuf_rwb_bufchan_buf :
                            writeCT$wnnzlizzieLet5_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnzlizzieLet5_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((sca3_1_argbuf_r && writeCT$wnnzlizzieLet5_1_argbuf_rwb_bufchan_buf[0]))
        writeCT$wnnzlizzieLet5_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
      else if (((! sca3_1_argbuf_r) && (! writeCT$wnnzlizzieLet5_1_argbuf_rwb_bufchan_buf[0])))
        writeCT$wnnzlizzieLet5_1_argbuf_rwb_bufchan_buf <= writeCT$wnnzlizzieLet5_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz) : (writeCT$wnnzlizzieLet60_1_argbuf,Pointer_CT$wnnz) > (writeCT$wnnzlizzieLet60_1_argbuf_rwb,Pointer_CT$wnnz) */
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet60_1_argbuf_bufchan_d;
  logic writeCT$wnnzlizzieLet60_1_argbuf_bufchan_r;
  assign writeCT$wnnzlizzieLet60_1_argbuf_r = ((! writeCT$wnnzlizzieLet60_1_argbuf_bufchan_d[0]) || writeCT$wnnzlizzieLet60_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnzlizzieLet60_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCT$wnnzlizzieLet60_1_argbuf_r)
        writeCT$wnnzlizzieLet60_1_argbuf_bufchan_d <= writeCT$wnnzlizzieLet60_1_argbuf_d;
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet60_1_argbuf_bufchan_buf;
  assign writeCT$wnnzlizzieLet60_1_argbuf_bufchan_r = (! writeCT$wnnzlizzieLet60_1_argbuf_bufchan_buf[0]);
  assign writeCT$wnnzlizzieLet60_1_argbuf_rwb_d = (writeCT$wnnzlizzieLet60_1_argbuf_bufchan_buf[0] ? writeCT$wnnzlizzieLet60_1_argbuf_bufchan_buf :
                                                   writeCT$wnnzlizzieLet60_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnzlizzieLet60_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeCT$wnnzlizzieLet60_1_argbuf_rwb_r && writeCT$wnnzlizzieLet60_1_argbuf_bufchan_buf[0]))
        writeCT$wnnzlizzieLet60_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeCT$wnnzlizzieLet60_1_argbuf_rwb_r) && (! writeCT$wnnzlizzieLet60_1_argbuf_bufchan_buf[0])))
        writeCT$wnnzlizzieLet60_1_argbuf_bufchan_buf <= writeCT$wnnzlizzieLet60_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz) : (writeCT$wnnzlizzieLet60_1_argbuf_rwb,Pointer_CT$wnnz) > (sca1_1_argbuf,Pointer_CT$wnnz) */
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet60_1_argbuf_rwb_bufchan_d;
  logic writeCT$wnnzlizzieLet60_1_argbuf_rwb_bufchan_r;
  assign writeCT$wnnzlizzieLet60_1_argbuf_rwb_r = ((! writeCT$wnnzlizzieLet60_1_argbuf_rwb_bufchan_d[0]) || writeCT$wnnzlizzieLet60_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnzlizzieLet60_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCT$wnnzlizzieLet60_1_argbuf_rwb_r)
        writeCT$wnnzlizzieLet60_1_argbuf_rwb_bufchan_d <= writeCT$wnnzlizzieLet60_1_argbuf_rwb_d;
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet60_1_argbuf_rwb_bufchan_buf;
  assign writeCT$wnnzlizzieLet60_1_argbuf_rwb_bufchan_r = (! writeCT$wnnzlizzieLet60_1_argbuf_rwb_bufchan_buf[0]);
  assign sca1_1_argbuf_d = (writeCT$wnnzlizzieLet60_1_argbuf_rwb_bufchan_buf[0] ? writeCT$wnnzlizzieLet60_1_argbuf_rwb_bufchan_buf :
                            writeCT$wnnzlizzieLet60_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnzlizzieLet60_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((sca1_1_argbuf_r && writeCT$wnnzlizzieLet60_1_argbuf_rwb_bufchan_buf[0]))
        writeCT$wnnzlizzieLet60_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
      else if (((! sca1_1_argbuf_r) && (! writeCT$wnnzlizzieLet60_1_argbuf_rwb_bufchan_buf[0])))
        writeCT$wnnzlizzieLet60_1_argbuf_rwb_bufchan_buf <= writeCT$wnnzlizzieLet60_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz) : (writeCT$wnnzlizzieLet61_1_argbuf,Pointer_CT$wnnz) > (writeCT$wnnzlizzieLet61_1_argbuf_rwb,Pointer_CT$wnnz) */
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet61_1_argbuf_bufchan_d;
  logic writeCT$wnnzlizzieLet61_1_argbuf_bufchan_r;
  assign writeCT$wnnzlizzieLet61_1_argbuf_r = ((! writeCT$wnnzlizzieLet61_1_argbuf_bufchan_d[0]) || writeCT$wnnzlizzieLet61_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnzlizzieLet61_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCT$wnnzlizzieLet61_1_argbuf_r)
        writeCT$wnnzlizzieLet61_1_argbuf_bufchan_d <= writeCT$wnnzlizzieLet61_1_argbuf_d;
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet61_1_argbuf_bufchan_buf;
  assign writeCT$wnnzlizzieLet61_1_argbuf_bufchan_r = (! writeCT$wnnzlizzieLet61_1_argbuf_bufchan_buf[0]);
  assign writeCT$wnnzlizzieLet61_1_argbuf_rwb_d = (writeCT$wnnzlizzieLet61_1_argbuf_bufchan_buf[0] ? writeCT$wnnzlizzieLet61_1_argbuf_bufchan_buf :
                                                   writeCT$wnnzlizzieLet61_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnzlizzieLet61_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeCT$wnnzlizzieLet61_1_argbuf_rwb_r && writeCT$wnnzlizzieLet61_1_argbuf_bufchan_buf[0]))
        writeCT$wnnzlizzieLet61_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeCT$wnnzlizzieLet61_1_argbuf_rwb_r) && (! writeCT$wnnzlizzieLet61_1_argbuf_bufchan_buf[0])))
        writeCT$wnnzlizzieLet61_1_argbuf_bufchan_buf <= writeCT$wnnzlizzieLet61_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz) : (writeCT$wnnzlizzieLet61_1_argbuf_rwb,Pointer_CT$wnnz) > (sca0_1_argbuf,Pointer_CT$wnnz) */
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet61_1_argbuf_rwb_bufchan_d;
  logic writeCT$wnnzlizzieLet61_1_argbuf_rwb_bufchan_r;
  assign writeCT$wnnzlizzieLet61_1_argbuf_rwb_r = ((! writeCT$wnnzlizzieLet61_1_argbuf_rwb_bufchan_d[0]) || writeCT$wnnzlizzieLet61_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnzlizzieLet61_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCT$wnnzlizzieLet61_1_argbuf_rwb_r)
        writeCT$wnnzlizzieLet61_1_argbuf_rwb_bufchan_d <= writeCT$wnnzlizzieLet61_1_argbuf_rwb_d;
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet61_1_argbuf_rwb_bufchan_buf;
  assign writeCT$wnnzlizzieLet61_1_argbuf_rwb_bufchan_r = (! writeCT$wnnzlizzieLet61_1_argbuf_rwb_bufchan_buf[0]);
  assign sca0_1_argbuf_d = (writeCT$wnnzlizzieLet61_1_argbuf_rwb_bufchan_buf[0] ? writeCT$wnnzlizzieLet61_1_argbuf_rwb_bufchan_buf :
                            writeCT$wnnzlizzieLet61_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnzlizzieLet61_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((sca0_1_argbuf_r && writeCT$wnnzlizzieLet61_1_argbuf_rwb_bufchan_buf[0]))
        writeCT$wnnzlizzieLet61_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
      else if (((! sca0_1_argbuf_r) && (! writeCT$wnnzlizzieLet61_1_argbuf_rwb_bufchan_buf[0])))
        writeCT$wnnzlizzieLet61_1_argbuf_rwb_bufchan_buf <= writeCT$wnnzlizzieLet61_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CTf''''''''''''_f''''''''''''_Int) : (writeCTf''''''''''''_f''''''''''''_IntlizzieLet14_1_argbuf,Pointer_CTf''''''''''''_f''''''''''''_Int) > (writeCTf''''''''''''_f''''''''''''_IntlizzieLet14_1_argbuf_rwb,Pointer_CTf''''''''''''_f''''''''''''_Int) */
  \Pointer_CTf''''''''''''_f''''''''''''_Int_t  \writeCTf''''''''''''_f''''''''''''_IntlizzieLet14_1_argbuf_bufchan_d ;
  logic \writeCTf''''''''''''_f''''''''''''_IntlizzieLet14_1_argbuf_bufchan_r ;
  assign \writeCTf''''''''''''_f''''''''''''_IntlizzieLet14_1_argbuf_r  = ((! \writeCTf''''''''''''_f''''''''''''_IntlizzieLet14_1_argbuf_bufchan_d [0]) || \writeCTf''''''''''''_f''''''''''''_IntlizzieLet14_1_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf''''''''''''_f''''''''''''_IntlizzieLet14_1_argbuf_bufchan_d  <= {16'd0,
                                                                                 1'd0};
    else
      if (\writeCTf''''''''''''_f''''''''''''_IntlizzieLet14_1_argbuf_r )
        \writeCTf''''''''''''_f''''''''''''_IntlizzieLet14_1_argbuf_bufchan_d  <= \writeCTf''''''''''''_f''''''''''''_IntlizzieLet14_1_argbuf_d ;
  \Pointer_CTf''''''''''''_f''''''''''''_Int_t  \writeCTf''''''''''''_f''''''''''''_IntlizzieLet14_1_argbuf_bufchan_buf ;
  assign \writeCTf''''''''''''_f''''''''''''_IntlizzieLet14_1_argbuf_bufchan_r  = (! \writeCTf''''''''''''_f''''''''''''_IntlizzieLet14_1_argbuf_bufchan_buf [0]);
  assign \writeCTf''''''''''''_f''''''''''''_IntlizzieLet14_1_argbuf_rwb_d  = (\writeCTf''''''''''''_f''''''''''''_IntlizzieLet14_1_argbuf_bufchan_buf [0] ? \writeCTf''''''''''''_f''''''''''''_IntlizzieLet14_1_argbuf_bufchan_buf  :
                                                                               \writeCTf''''''''''''_f''''''''''''_IntlizzieLet14_1_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf''''''''''''_f''''''''''''_IntlizzieLet14_1_argbuf_bufchan_buf  <= {16'd0,
                                                                                   1'd0};
    else
      if ((\writeCTf''''''''''''_f''''''''''''_IntlizzieLet14_1_argbuf_rwb_r  && \writeCTf''''''''''''_f''''''''''''_IntlizzieLet14_1_argbuf_bufchan_buf [0]))
        \writeCTf''''''''''''_f''''''''''''_IntlizzieLet14_1_argbuf_bufchan_buf  <= {16'd0,
                                                                                     1'd0};
      else if (((! \writeCTf''''''''''''_f''''''''''''_IntlizzieLet14_1_argbuf_rwb_r ) && (! \writeCTf''''''''''''_f''''''''''''_IntlizzieLet14_1_argbuf_bufchan_buf [0])))
        \writeCTf''''''''''''_f''''''''''''_IntlizzieLet14_1_argbuf_bufchan_buf  <= \writeCTf''''''''''''_f''''''''''''_IntlizzieLet14_1_argbuf_bufchan_d ;
  
  /* buf (Ty Pointer_CTf''''''''''''_f''''''''''''_Int) : (writeCTf''''''''''''_f''''''''''''_IntlizzieLet14_1_argbuf_rwb,Pointer_CTf''''''''''''_f''''''''''''_Int) > (sca3_1_1_argbuf,Pointer_CTf''''''''''''_f''''''''''''_Int) */
  \Pointer_CTf''''''''''''_f''''''''''''_Int_t  \writeCTf''''''''''''_f''''''''''''_IntlizzieLet14_1_argbuf_rwb_bufchan_d ;
  logic \writeCTf''''''''''''_f''''''''''''_IntlizzieLet14_1_argbuf_rwb_bufchan_r ;
  assign \writeCTf''''''''''''_f''''''''''''_IntlizzieLet14_1_argbuf_rwb_r  = ((! \writeCTf''''''''''''_f''''''''''''_IntlizzieLet14_1_argbuf_rwb_bufchan_d [0]) || \writeCTf''''''''''''_f''''''''''''_IntlizzieLet14_1_argbuf_rwb_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf''''''''''''_f''''''''''''_IntlizzieLet14_1_argbuf_rwb_bufchan_d  <= {16'd0,
                                                                                     1'd0};
    else
      if (\writeCTf''''''''''''_f''''''''''''_IntlizzieLet14_1_argbuf_rwb_r )
        \writeCTf''''''''''''_f''''''''''''_IntlizzieLet14_1_argbuf_rwb_bufchan_d  <= \writeCTf''''''''''''_f''''''''''''_IntlizzieLet14_1_argbuf_rwb_d ;
  \Pointer_CTf''''''''''''_f''''''''''''_Int_t  \writeCTf''''''''''''_f''''''''''''_IntlizzieLet14_1_argbuf_rwb_bufchan_buf ;
  assign \writeCTf''''''''''''_f''''''''''''_IntlizzieLet14_1_argbuf_rwb_bufchan_r  = (! \writeCTf''''''''''''_f''''''''''''_IntlizzieLet14_1_argbuf_rwb_bufchan_buf [0]);
  assign sca3_1_1_argbuf_d = (\writeCTf''''''''''''_f''''''''''''_IntlizzieLet14_1_argbuf_rwb_bufchan_buf [0] ? \writeCTf''''''''''''_f''''''''''''_IntlizzieLet14_1_argbuf_rwb_bufchan_buf  :
                              \writeCTf''''''''''''_f''''''''''''_IntlizzieLet14_1_argbuf_rwb_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf''''''''''''_f''''''''''''_IntlizzieLet14_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                                       1'd0};
    else
      if ((sca3_1_1_argbuf_r && \writeCTf''''''''''''_f''''''''''''_IntlizzieLet14_1_argbuf_rwb_bufchan_buf [0]))
        \writeCTf''''''''''''_f''''''''''''_IntlizzieLet14_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                                         1'd0};
      else if (((! sca3_1_1_argbuf_r) && (! \writeCTf''''''''''''_f''''''''''''_IntlizzieLet14_1_argbuf_rwb_bufchan_buf [0])))
        \writeCTf''''''''''''_f''''''''''''_IntlizzieLet14_1_argbuf_rwb_bufchan_buf  <= \writeCTf''''''''''''_f''''''''''''_IntlizzieLet14_1_argbuf_rwb_bufchan_d ;
  
  /* buf (Ty Pointer_CTf''''''''''''_f''''''''''''_Int) : (writeCTf''''''''''''_f''''''''''''_IntlizzieLet56_1_argbuf,Pointer_CTf''''''''''''_f''''''''''''_Int) > (writeCTf''''''''''''_f''''''''''''_IntlizzieLet56_1_argbuf_rwb,Pointer_CTf''''''''''''_f''''''''''''_Int) */
  \Pointer_CTf''''''''''''_f''''''''''''_Int_t  \writeCTf''''''''''''_f''''''''''''_IntlizzieLet56_1_argbuf_bufchan_d ;
  logic \writeCTf''''''''''''_f''''''''''''_IntlizzieLet56_1_argbuf_bufchan_r ;
  assign \writeCTf''''''''''''_f''''''''''''_IntlizzieLet56_1_argbuf_r  = ((! \writeCTf''''''''''''_f''''''''''''_IntlizzieLet56_1_argbuf_bufchan_d [0]) || \writeCTf''''''''''''_f''''''''''''_IntlizzieLet56_1_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf''''''''''''_f''''''''''''_IntlizzieLet56_1_argbuf_bufchan_d  <= {16'd0,
                                                                                 1'd0};
    else
      if (\writeCTf''''''''''''_f''''''''''''_IntlizzieLet56_1_argbuf_r )
        \writeCTf''''''''''''_f''''''''''''_IntlizzieLet56_1_argbuf_bufchan_d  <= \writeCTf''''''''''''_f''''''''''''_IntlizzieLet56_1_argbuf_d ;
  \Pointer_CTf''''''''''''_f''''''''''''_Int_t  \writeCTf''''''''''''_f''''''''''''_IntlizzieLet56_1_argbuf_bufchan_buf ;
  assign \writeCTf''''''''''''_f''''''''''''_IntlizzieLet56_1_argbuf_bufchan_r  = (! \writeCTf''''''''''''_f''''''''''''_IntlizzieLet56_1_argbuf_bufchan_buf [0]);
  assign \writeCTf''''''''''''_f''''''''''''_IntlizzieLet56_1_argbuf_rwb_d  = (\writeCTf''''''''''''_f''''''''''''_IntlizzieLet56_1_argbuf_bufchan_buf [0] ? \writeCTf''''''''''''_f''''''''''''_IntlizzieLet56_1_argbuf_bufchan_buf  :
                                                                               \writeCTf''''''''''''_f''''''''''''_IntlizzieLet56_1_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf''''''''''''_f''''''''''''_IntlizzieLet56_1_argbuf_bufchan_buf  <= {16'd0,
                                                                                   1'd0};
    else
      if ((\writeCTf''''''''''''_f''''''''''''_IntlizzieLet56_1_argbuf_rwb_r  && \writeCTf''''''''''''_f''''''''''''_IntlizzieLet56_1_argbuf_bufchan_buf [0]))
        \writeCTf''''''''''''_f''''''''''''_IntlizzieLet56_1_argbuf_bufchan_buf  <= {16'd0,
                                                                                     1'd0};
      else if (((! \writeCTf''''''''''''_f''''''''''''_IntlizzieLet56_1_argbuf_rwb_r ) && (! \writeCTf''''''''''''_f''''''''''''_IntlizzieLet56_1_argbuf_bufchan_buf [0])))
        \writeCTf''''''''''''_f''''''''''''_IntlizzieLet56_1_argbuf_bufchan_buf  <= \writeCTf''''''''''''_f''''''''''''_IntlizzieLet56_1_argbuf_bufchan_d ;
  
  /* buf (Ty Pointer_CTf''''''''''''_f''''''''''''_Int) : (writeCTf''''''''''''_f''''''''''''_IntlizzieLet56_1_argbuf_rwb,Pointer_CTf''''''''''''_f''''''''''''_Int) > (lizzieLet7_1_1_argbuf,Pointer_CTf''''''''''''_f''''''''''''_Int) */
  \Pointer_CTf''''''''''''_f''''''''''''_Int_t  \writeCTf''''''''''''_f''''''''''''_IntlizzieLet56_1_argbuf_rwb_bufchan_d ;
  logic \writeCTf''''''''''''_f''''''''''''_IntlizzieLet56_1_argbuf_rwb_bufchan_r ;
  assign \writeCTf''''''''''''_f''''''''''''_IntlizzieLet56_1_argbuf_rwb_r  = ((! \writeCTf''''''''''''_f''''''''''''_IntlizzieLet56_1_argbuf_rwb_bufchan_d [0]) || \writeCTf''''''''''''_f''''''''''''_IntlizzieLet56_1_argbuf_rwb_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf''''''''''''_f''''''''''''_IntlizzieLet56_1_argbuf_rwb_bufchan_d  <= {16'd0,
                                                                                     1'd0};
    else
      if (\writeCTf''''''''''''_f''''''''''''_IntlizzieLet56_1_argbuf_rwb_r )
        \writeCTf''''''''''''_f''''''''''''_IntlizzieLet56_1_argbuf_rwb_bufchan_d  <= \writeCTf''''''''''''_f''''''''''''_IntlizzieLet56_1_argbuf_rwb_d ;
  \Pointer_CTf''''''''''''_f''''''''''''_Int_t  \writeCTf''''''''''''_f''''''''''''_IntlizzieLet56_1_argbuf_rwb_bufchan_buf ;
  assign \writeCTf''''''''''''_f''''''''''''_IntlizzieLet56_1_argbuf_rwb_bufchan_r  = (! \writeCTf''''''''''''_f''''''''''''_IntlizzieLet56_1_argbuf_rwb_bufchan_buf [0]);
  assign lizzieLet7_1_1_argbuf_d = (\writeCTf''''''''''''_f''''''''''''_IntlizzieLet56_1_argbuf_rwb_bufchan_buf [0] ? \writeCTf''''''''''''_f''''''''''''_IntlizzieLet56_1_argbuf_rwb_bufchan_buf  :
                                    \writeCTf''''''''''''_f''''''''''''_IntlizzieLet56_1_argbuf_rwb_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf''''''''''''_f''''''''''''_IntlizzieLet56_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                                       1'd0};
    else
      if ((lizzieLet7_1_1_argbuf_r && \writeCTf''''''''''''_f''''''''''''_IntlizzieLet56_1_argbuf_rwb_bufchan_buf [0]))
        \writeCTf''''''''''''_f''''''''''''_IntlizzieLet56_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                                         1'd0};
      else if (((! lizzieLet7_1_1_argbuf_r) && (! \writeCTf''''''''''''_f''''''''''''_IntlizzieLet56_1_argbuf_rwb_bufchan_buf [0])))
        \writeCTf''''''''''''_f''''''''''''_IntlizzieLet56_1_argbuf_rwb_bufchan_buf  <= \writeCTf''''''''''''_f''''''''''''_IntlizzieLet56_1_argbuf_rwb_bufchan_d ;
  
  /* buf (Ty Pointer_CTf''''''''''''_f''''''''''''_Int) : (writeCTf''''''''''''_f''''''''''''_IntlizzieLet63_1_argbuf,Pointer_CTf''''''''''''_f''''''''''''_Int) > (writeCTf''''''''''''_f''''''''''''_IntlizzieLet63_1_argbuf_rwb,Pointer_CTf''''''''''''_f''''''''''''_Int) */
  \Pointer_CTf''''''''''''_f''''''''''''_Int_t  \writeCTf''''''''''''_f''''''''''''_IntlizzieLet63_1_argbuf_bufchan_d ;
  logic \writeCTf''''''''''''_f''''''''''''_IntlizzieLet63_1_argbuf_bufchan_r ;
  assign \writeCTf''''''''''''_f''''''''''''_IntlizzieLet63_1_argbuf_r  = ((! \writeCTf''''''''''''_f''''''''''''_IntlizzieLet63_1_argbuf_bufchan_d [0]) || \writeCTf''''''''''''_f''''''''''''_IntlizzieLet63_1_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf''''''''''''_f''''''''''''_IntlizzieLet63_1_argbuf_bufchan_d  <= {16'd0,
                                                                                 1'd0};
    else
      if (\writeCTf''''''''''''_f''''''''''''_IntlizzieLet63_1_argbuf_r )
        \writeCTf''''''''''''_f''''''''''''_IntlizzieLet63_1_argbuf_bufchan_d  <= \writeCTf''''''''''''_f''''''''''''_IntlizzieLet63_1_argbuf_d ;
  \Pointer_CTf''''''''''''_f''''''''''''_Int_t  \writeCTf''''''''''''_f''''''''''''_IntlizzieLet63_1_argbuf_bufchan_buf ;
  assign \writeCTf''''''''''''_f''''''''''''_IntlizzieLet63_1_argbuf_bufchan_r  = (! \writeCTf''''''''''''_f''''''''''''_IntlizzieLet63_1_argbuf_bufchan_buf [0]);
  assign \writeCTf''''''''''''_f''''''''''''_IntlizzieLet63_1_argbuf_rwb_d  = (\writeCTf''''''''''''_f''''''''''''_IntlizzieLet63_1_argbuf_bufchan_buf [0] ? \writeCTf''''''''''''_f''''''''''''_IntlizzieLet63_1_argbuf_bufchan_buf  :
                                                                               \writeCTf''''''''''''_f''''''''''''_IntlizzieLet63_1_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf''''''''''''_f''''''''''''_IntlizzieLet63_1_argbuf_bufchan_buf  <= {16'd0,
                                                                                   1'd0};
    else
      if ((\writeCTf''''''''''''_f''''''''''''_IntlizzieLet63_1_argbuf_rwb_r  && \writeCTf''''''''''''_f''''''''''''_IntlizzieLet63_1_argbuf_bufchan_buf [0]))
        \writeCTf''''''''''''_f''''''''''''_IntlizzieLet63_1_argbuf_bufchan_buf  <= {16'd0,
                                                                                     1'd0};
      else if (((! \writeCTf''''''''''''_f''''''''''''_IntlizzieLet63_1_argbuf_rwb_r ) && (! \writeCTf''''''''''''_f''''''''''''_IntlizzieLet63_1_argbuf_bufchan_buf [0])))
        \writeCTf''''''''''''_f''''''''''''_IntlizzieLet63_1_argbuf_bufchan_buf  <= \writeCTf''''''''''''_f''''''''''''_IntlizzieLet63_1_argbuf_bufchan_d ;
  
  /* buf (Ty Pointer_CTf''''''''''''_f''''''''''''_Int) : (writeCTf''''''''''''_f''''''''''''_IntlizzieLet63_1_argbuf_rwb,Pointer_CTf''''''''''''_f''''''''''''_Int) > (sca2_1_1_argbuf,Pointer_CTf''''''''''''_f''''''''''''_Int) */
  \Pointer_CTf''''''''''''_f''''''''''''_Int_t  \writeCTf''''''''''''_f''''''''''''_IntlizzieLet63_1_argbuf_rwb_bufchan_d ;
  logic \writeCTf''''''''''''_f''''''''''''_IntlizzieLet63_1_argbuf_rwb_bufchan_r ;
  assign \writeCTf''''''''''''_f''''''''''''_IntlizzieLet63_1_argbuf_rwb_r  = ((! \writeCTf''''''''''''_f''''''''''''_IntlizzieLet63_1_argbuf_rwb_bufchan_d [0]) || \writeCTf''''''''''''_f''''''''''''_IntlizzieLet63_1_argbuf_rwb_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf''''''''''''_f''''''''''''_IntlizzieLet63_1_argbuf_rwb_bufchan_d  <= {16'd0,
                                                                                     1'd0};
    else
      if (\writeCTf''''''''''''_f''''''''''''_IntlizzieLet63_1_argbuf_rwb_r )
        \writeCTf''''''''''''_f''''''''''''_IntlizzieLet63_1_argbuf_rwb_bufchan_d  <= \writeCTf''''''''''''_f''''''''''''_IntlizzieLet63_1_argbuf_rwb_d ;
  \Pointer_CTf''''''''''''_f''''''''''''_Int_t  \writeCTf''''''''''''_f''''''''''''_IntlizzieLet63_1_argbuf_rwb_bufchan_buf ;
  assign \writeCTf''''''''''''_f''''''''''''_IntlizzieLet63_1_argbuf_rwb_bufchan_r  = (! \writeCTf''''''''''''_f''''''''''''_IntlizzieLet63_1_argbuf_rwb_bufchan_buf [0]);
  assign sca2_1_1_argbuf_d = (\writeCTf''''''''''''_f''''''''''''_IntlizzieLet63_1_argbuf_rwb_bufchan_buf [0] ? \writeCTf''''''''''''_f''''''''''''_IntlizzieLet63_1_argbuf_rwb_bufchan_buf  :
                              \writeCTf''''''''''''_f''''''''''''_IntlizzieLet63_1_argbuf_rwb_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf''''''''''''_f''''''''''''_IntlizzieLet63_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                                       1'd0};
    else
      if ((sca2_1_1_argbuf_r && \writeCTf''''''''''''_f''''''''''''_IntlizzieLet63_1_argbuf_rwb_bufchan_buf [0]))
        \writeCTf''''''''''''_f''''''''''''_IntlizzieLet63_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                                         1'd0};
      else if (((! sca2_1_1_argbuf_r) && (! \writeCTf''''''''''''_f''''''''''''_IntlizzieLet63_1_argbuf_rwb_bufchan_buf [0])))
        \writeCTf''''''''''''_f''''''''''''_IntlizzieLet63_1_argbuf_rwb_bufchan_buf  <= \writeCTf''''''''''''_f''''''''''''_IntlizzieLet63_1_argbuf_rwb_bufchan_d ;
  
  /* buf (Ty Pointer_CTf''''''''''''_f''''''''''''_Int) : (writeCTf''''''''''''_f''''''''''''_IntlizzieLet64_1_argbuf,Pointer_CTf''''''''''''_f''''''''''''_Int) > (writeCTf''''''''''''_f''''''''''''_IntlizzieLet64_1_argbuf_rwb,Pointer_CTf''''''''''''_f''''''''''''_Int) */
  \Pointer_CTf''''''''''''_f''''''''''''_Int_t  \writeCTf''''''''''''_f''''''''''''_IntlizzieLet64_1_argbuf_bufchan_d ;
  logic \writeCTf''''''''''''_f''''''''''''_IntlizzieLet64_1_argbuf_bufchan_r ;
  assign \writeCTf''''''''''''_f''''''''''''_IntlizzieLet64_1_argbuf_r  = ((! \writeCTf''''''''''''_f''''''''''''_IntlizzieLet64_1_argbuf_bufchan_d [0]) || \writeCTf''''''''''''_f''''''''''''_IntlizzieLet64_1_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf''''''''''''_f''''''''''''_IntlizzieLet64_1_argbuf_bufchan_d  <= {16'd0,
                                                                                 1'd0};
    else
      if (\writeCTf''''''''''''_f''''''''''''_IntlizzieLet64_1_argbuf_r )
        \writeCTf''''''''''''_f''''''''''''_IntlizzieLet64_1_argbuf_bufchan_d  <= \writeCTf''''''''''''_f''''''''''''_IntlizzieLet64_1_argbuf_d ;
  \Pointer_CTf''''''''''''_f''''''''''''_Int_t  \writeCTf''''''''''''_f''''''''''''_IntlizzieLet64_1_argbuf_bufchan_buf ;
  assign \writeCTf''''''''''''_f''''''''''''_IntlizzieLet64_1_argbuf_bufchan_r  = (! \writeCTf''''''''''''_f''''''''''''_IntlizzieLet64_1_argbuf_bufchan_buf [0]);
  assign \writeCTf''''''''''''_f''''''''''''_IntlizzieLet64_1_argbuf_rwb_d  = (\writeCTf''''''''''''_f''''''''''''_IntlizzieLet64_1_argbuf_bufchan_buf [0] ? \writeCTf''''''''''''_f''''''''''''_IntlizzieLet64_1_argbuf_bufchan_buf  :
                                                                               \writeCTf''''''''''''_f''''''''''''_IntlizzieLet64_1_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf''''''''''''_f''''''''''''_IntlizzieLet64_1_argbuf_bufchan_buf  <= {16'd0,
                                                                                   1'd0};
    else
      if ((\writeCTf''''''''''''_f''''''''''''_IntlizzieLet64_1_argbuf_rwb_r  && \writeCTf''''''''''''_f''''''''''''_IntlizzieLet64_1_argbuf_bufchan_buf [0]))
        \writeCTf''''''''''''_f''''''''''''_IntlizzieLet64_1_argbuf_bufchan_buf  <= {16'd0,
                                                                                     1'd0};
      else if (((! \writeCTf''''''''''''_f''''''''''''_IntlizzieLet64_1_argbuf_rwb_r ) && (! \writeCTf''''''''''''_f''''''''''''_IntlizzieLet64_1_argbuf_bufchan_buf [0])))
        \writeCTf''''''''''''_f''''''''''''_IntlizzieLet64_1_argbuf_bufchan_buf  <= \writeCTf''''''''''''_f''''''''''''_IntlizzieLet64_1_argbuf_bufchan_d ;
  
  /* buf (Ty Pointer_CTf''''''''''''_f''''''''''''_Int) : (writeCTf''''''''''''_f''''''''''''_IntlizzieLet64_1_argbuf_rwb,Pointer_CTf''''''''''''_f''''''''''''_Int) > (sca1_1_1_argbuf,Pointer_CTf''''''''''''_f''''''''''''_Int) */
  \Pointer_CTf''''''''''''_f''''''''''''_Int_t  \writeCTf''''''''''''_f''''''''''''_IntlizzieLet64_1_argbuf_rwb_bufchan_d ;
  logic \writeCTf''''''''''''_f''''''''''''_IntlizzieLet64_1_argbuf_rwb_bufchan_r ;
  assign \writeCTf''''''''''''_f''''''''''''_IntlizzieLet64_1_argbuf_rwb_r  = ((! \writeCTf''''''''''''_f''''''''''''_IntlizzieLet64_1_argbuf_rwb_bufchan_d [0]) || \writeCTf''''''''''''_f''''''''''''_IntlizzieLet64_1_argbuf_rwb_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf''''''''''''_f''''''''''''_IntlizzieLet64_1_argbuf_rwb_bufchan_d  <= {16'd0,
                                                                                     1'd0};
    else
      if (\writeCTf''''''''''''_f''''''''''''_IntlizzieLet64_1_argbuf_rwb_r )
        \writeCTf''''''''''''_f''''''''''''_IntlizzieLet64_1_argbuf_rwb_bufchan_d  <= \writeCTf''''''''''''_f''''''''''''_IntlizzieLet64_1_argbuf_rwb_d ;
  \Pointer_CTf''''''''''''_f''''''''''''_Int_t  \writeCTf''''''''''''_f''''''''''''_IntlizzieLet64_1_argbuf_rwb_bufchan_buf ;
  assign \writeCTf''''''''''''_f''''''''''''_IntlizzieLet64_1_argbuf_rwb_bufchan_r  = (! \writeCTf''''''''''''_f''''''''''''_IntlizzieLet64_1_argbuf_rwb_bufchan_buf [0]);
  assign sca1_1_1_argbuf_d = (\writeCTf''''''''''''_f''''''''''''_IntlizzieLet64_1_argbuf_rwb_bufchan_buf [0] ? \writeCTf''''''''''''_f''''''''''''_IntlizzieLet64_1_argbuf_rwb_bufchan_buf  :
                              \writeCTf''''''''''''_f''''''''''''_IntlizzieLet64_1_argbuf_rwb_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf''''''''''''_f''''''''''''_IntlizzieLet64_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                                       1'd0};
    else
      if ((sca1_1_1_argbuf_r && \writeCTf''''''''''''_f''''''''''''_IntlizzieLet64_1_argbuf_rwb_bufchan_buf [0]))
        \writeCTf''''''''''''_f''''''''''''_IntlizzieLet64_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                                         1'd0};
      else if (((! sca1_1_1_argbuf_r) && (! \writeCTf''''''''''''_f''''''''''''_IntlizzieLet64_1_argbuf_rwb_bufchan_buf [0])))
        \writeCTf''''''''''''_f''''''''''''_IntlizzieLet64_1_argbuf_rwb_bufchan_buf  <= \writeCTf''''''''''''_f''''''''''''_IntlizzieLet64_1_argbuf_rwb_bufchan_d ;
  
  /* buf (Ty Pointer_CTf''''''''''''_f''''''''''''_Int) : (writeCTf''''''''''''_f''''''''''''_IntlizzieLet65_1_argbuf,Pointer_CTf''''''''''''_f''''''''''''_Int) > (writeCTf''''''''''''_f''''''''''''_IntlizzieLet65_1_argbuf_rwb,Pointer_CTf''''''''''''_f''''''''''''_Int) */
  \Pointer_CTf''''''''''''_f''''''''''''_Int_t  \writeCTf''''''''''''_f''''''''''''_IntlizzieLet65_1_argbuf_bufchan_d ;
  logic \writeCTf''''''''''''_f''''''''''''_IntlizzieLet65_1_argbuf_bufchan_r ;
  assign \writeCTf''''''''''''_f''''''''''''_IntlizzieLet65_1_argbuf_r  = ((! \writeCTf''''''''''''_f''''''''''''_IntlizzieLet65_1_argbuf_bufchan_d [0]) || \writeCTf''''''''''''_f''''''''''''_IntlizzieLet65_1_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf''''''''''''_f''''''''''''_IntlizzieLet65_1_argbuf_bufchan_d  <= {16'd0,
                                                                                 1'd0};
    else
      if (\writeCTf''''''''''''_f''''''''''''_IntlizzieLet65_1_argbuf_r )
        \writeCTf''''''''''''_f''''''''''''_IntlizzieLet65_1_argbuf_bufchan_d  <= \writeCTf''''''''''''_f''''''''''''_IntlizzieLet65_1_argbuf_d ;
  \Pointer_CTf''''''''''''_f''''''''''''_Int_t  \writeCTf''''''''''''_f''''''''''''_IntlizzieLet65_1_argbuf_bufchan_buf ;
  assign \writeCTf''''''''''''_f''''''''''''_IntlizzieLet65_1_argbuf_bufchan_r  = (! \writeCTf''''''''''''_f''''''''''''_IntlizzieLet65_1_argbuf_bufchan_buf [0]);
  assign \writeCTf''''''''''''_f''''''''''''_IntlizzieLet65_1_argbuf_rwb_d  = (\writeCTf''''''''''''_f''''''''''''_IntlizzieLet65_1_argbuf_bufchan_buf [0] ? \writeCTf''''''''''''_f''''''''''''_IntlizzieLet65_1_argbuf_bufchan_buf  :
                                                                               \writeCTf''''''''''''_f''''''''''''_IntlizzieLet65_1_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf''''''''''''_f''''''''''''_IntlizzieLet65_1_argbuf_bufchan_buf  <= {16'd0,
                                                                                   1'd0};
    else
      if ((\writeCTf''''''''''''_f''''''''''''_IntlizzieLet65_1_argbuf_rwb_r  && \writeCTf''''''''''''_f''''''''''''_IntlizzieLet65_1_argbuf_bufchan_buf [0]))
        \writeCTf''''''''''''_f''''''''''''_IntlizzieLet65_1_argbuf_bufchan_buf  <= {16'd0,
                                                                                     1'd0};
      else if (((! \writeCTf''''''''''''_f''''''''''''_IntlizzieLet65_1_argbuf_rwb_r ) && (! \writeCTf''''''''''''_f''''''''''''_IntlizzieLet65_1_argbuf_bufchan_buf [0])))
        \writeCTf''''''''''''_f''''''''''''_IntlizzieLet65_1_argbuf_bufchan_buf  <= \writeCTf''''''''''''_f''''''''''''_IntlizzieLet65_1_argbuf_bufchan_d ;
  
  /* buf (Ty Pointer_CTf''''''''''''_f''''''''''''_Int) : (writeCTf''''''''''''_f''''''''''''_IntlizzieLet65_1_argbuf_rwb,Pointer_CTf''''''''''''_f''''''''''''_Int) > (sca0_1_1_argbuf,Pointer_CTf''''''''''''_f''''''''''''_Int) */
  \Pointer_CTf''''''''''''_f''''''''''''_Int_t  \writeCTf''''''''''''_f''''''''''''_IntlizzieLet65_1_argbuf_rwb_bufchan_d ;
  logic \writeCTf''''''''''''_f''''''''''''_IntlizzieLet65_1_argbuf_rwb_bufchan_r ;
  assign \writeCTf''''''''''''_f''''''''''''_IntlizzieLet65_1_argbuf_rwb_r  = ((! \writeCTf''''''''''''_f''''''''''''_IntlizzieLet65_1_argbuf_rwb_bufchan_d [0]) || \writeCTf''''''''''''_f''''''''''''_IntlizzieLet65_1_argbuf_rwb_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf''''''''''''_f''''''''''''_IntlizzieLet65_1_argbuf_rwb_bufchan_d  <= {16'd0,
                                                                                     1'd0};
    else
      if (\writeCTf''''''''''''_f''''''''''''_IntlizzieLet65_1_argbuf_rwb_r )
        \writeCTf''''''''''''_f''''''''''''_IntlizzieLet65_1_argbuf_rwb_bufchan_d  <= \writeCTf''''''''''''_f''''''''''''_IntlizzieLet65_1_argbuf_rwb_d ;
  \Pointer_CTf''''''''''''_f''''''''''''_Int_t  \writeCTf''''''''''''_f''''''''''''_IntlizzieLet65_1_argbuf_rwb_bufchan_buf ;
  assign \writeCTf''''''''''''_f''''''''''''_IntlizzieLet65_1_argbuf_rwb_bufchan_r  = (! \writeCTf''''''''''''_f''''''''''''_IntlizzieLet65_1_argbuf_rwb_bufchan_buf [0]);
  assign sca0_1_1_argbuf_d = (\writeCTf''''''''''''_f''''''''''''_IntlizzieLet65_1_argbuf_rwb_bufchan_buf [0] ? \writeCTf''''''''''''_f''''''''''''_IntlizzieLet65_1_argbuf_rwb_bufchan_buf  :
                              \writeCTf''''''''''''_f''''''''''''_IntlizzieLet65_1_argbuf_rwb_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf''''''''''''_f''''''''''''_IntlizzieLet65_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                                       1'd0};
    else
      if ((sca0_1_1_argbuf_r && \writeCTf''''''''''''_f''''''''''''_IntlizzieLet65_1_argbuf_rwb_bufchan_buf [0]))
        \writeCTf''''''''''''_f''''''''''''_IntlizzieLet65_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                                         1'd0};
      else if (((! sca0_1_1_argbuf_r) && (! \writeCTf''''''''''''_f''''''''''''_IntlizzieLet65_1_argbuf_rwb_bufchan_buf [0])))
        \writeCTf''''''''''''_f''''''''''''_IntlizzieLet65_1_argbuf_rwb_bufchan_buf  <= \writeCTf''''''''''''_f''''''''''''_IntlizzieLet65_1_argbuf_rwb_bufchan_d ;
  
  /* buf (Ty Pointer_CTf_f_Int) : (writeCTf_f_IntlizzieLet52_1_argbuf,Pointer_CTf_f_Int) > (writeCTf_f_IntlizzieLet52_1_argbuf_rwb,Pointer_CTf_f_Int) */
  Pointer_CTf_f_Int_t writeCTf_f_IntlizzieLet52_1_argbuf_bufchan_d;
  logic writeCTf_f_IntlizzieLet52_1_argbuf_bufchan_r;
  assign writeCTf_f_IntlizzieLet52_1_argbuf_r = ((! writeCTf_f_IntlizzieLet52_1_argbuf_bufchan_d[0]) || writeCTf_f_IntlizzieLet52_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTf_f_IntlizzieLet52_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCTf_f_IntlizzieLet52_1_argbuf_r)
        writeCTf_f_IntlizzieLet52_1_argbuf_bufchan_d <= writeCTf_f_IntlizzieLet52_1_argbuf_d;
  Pointer_CTf_f_Int_t writeCTf_f_IntlizzieLet52_1_argbuf_bufchan_buf;
  assign writeCTf_f_IntlizzieLet52_1_argbuf_bufchan_r = (! writeCTf_f_IntlizzieLet52_1_argbuf_bufchan_buf[0]);
  assign writeCTf_f_IntlizzieLet52_1_argbuf_rwb_d = (writeCTf_f_IntlizzieLet52_1_argbuf_bufchan_buf[0] ? writeCTf_f_IntlizzieLet52_1_argbuf_bufchan_buf :
                                                     writeCTf_f_IntlizzieLet52_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTf_f_IntlizzieLet52_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeCTf_f_IntlizzieLet52_1_argbuf_rwb_r && writeCTf_f_IntlizzieLet52_1_argbuf_bufchan_buf[0]))
        writeCTf_f_IntlizzieLet52_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeCTf_f_IntlizzieLet52_1_argbuf_rwb_r) && (! writeCTf_f_IntlizzieLet52_1_argbuf_bufchan_buf[0])))
        writeCTf_f_IntlizzieLet52_1_argbuf_bufchan_buf <= writeCTf_f_IntlizzieLet52_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CTf_f_Int) : (writeCTf_f_IntlizzieLet52_1_argbuf_rwb,Pointer_CTf_f_Int) > (sca3_2_1_argbuf,Pointer_CTf_f_Int) */
  Pointer_CTf_f_Int_t writeCTf_f_IntlizzieLet52_1_argbuf_rwb_bufchan_d;
  logic writeCTf_f_IntlizzieLet52_1_argbuf_rwb_bufchan_r;
  assign writeCTf_f_IntlizzieLet52_1_argbuf_rwb_r = ((! writeCTf_f_IntlizzieLet52_1_argbuf_rwb_bufchan_d[0]) || writeCTf_f_IntlizzieLet52_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTf_f_IntlizzieLet52_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCTf_f_IntlizzieLet52_1_argbuf_rwb_r)
        writeCTf_f_IntlizzieLet52_1_argbuf_rwb_bufchan_d <= writeCTf_f_IntlizzieLet52_1_argbuf_rwb_d;
  Pointer_CTf_f_Int_t writeCTf_f_IntlizzieLet52_1_argbuf_rwb_bufchan_buf;
  assign writeCTf_f_IntlizzieLet52_1_argbuf_rwb_bufchan_r = (! writeCTf_f_IntlizzieLet52_1_argbuf_rwb_bufchan_buf[0]);
  assign sca3_2_1_argbuf_d = (writeCTf_f_IntlizzieLet52_1_argbuf_rwb_bufchan_buf[0] ? writeCTf_f_IntlizzieLet52_1_argbuf_rwb_bufchan_buf :
                              writeCTf_f_IntlizzieLet52_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTf_f_IntlizzieLet52_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((sca3_2_1_argbuf_r && writeCTf_f_IntlizzieLet52_1_argbuf_rwb_bufchan_buf[0]))
        writeCTf_f_IntlizzieLet52_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! sca3_2_1_argbuf_r) && (! writeCTf_f_IntlizzieLet52_1_argbuf_rwb_bufchan_buf[0])))
        writeCTf_f_IntlizzieLet52_1_argbuf_rwb_bufchan_buf <= writeCTf_f_IntlizzieLet52_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CTf_f_Int) : (writeCTf_f_IntlizzieLet57_1_argbuf,Pointer_CTf_f_Int) > (writeCTf_f_IntlizzieLet57_1_argbuf_rwb,Pointer_CTf_f_Int) */
  Pointer_CTf_f_Int_t writeCTf_f_IntlizzieLet57_1_argbuf_bufchan_d;
  logic writeCTf_f_IntlizzieLet57_1_argbuf_bufchan_r;
  assign writeCTf_f_IntlizzieLet57_1_argbuf_r = ((! writeCTf_f_IntlizzieLet57_1_argbuf_bufchan_d[0]) || writeCTf_f_IntlizzieLet57_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTf_f_IntlizzieLet57_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCTf_f_IntlizzieLet57_1_argbuf_r)
        writeCTf_f_IntlizzieLet57_1_argbuf_bufchan_d <= writeCTf_f_IntlizzieLet57_1_argbuf_d;
  Pointer_CTf_f_Int_t writeCTf_f_IntlizzieLet57_1_argbuf_bufchan_buf;
  assign writeCTf_f_IntlizzieLet57_1_argbuf_bufchan_r = (! writeCTf_f_IntlizzieLet57_1_argbuf_bufchan_buf[0]);
  assign writeCTf_f_IntlizzieLet57_1_argbuf_rwb_d = (writeCTf_f_IntlizzieLet57_1_argbuf_bufchan_buf[0] ? writeCTf_f_IntlizzieLet57_1_argbuf_bufchan_buf :
                                                     writeCTf_f_IntlizzieLet57_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTf_f_IntlizzieLet57_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeCTf_f_IntlizzieLet57_1_argbuf_rwb_r && writeCTf_f_IntlizzieLet57_1_argbuf_bufchan_buf[0]))
        writeCTf_f_IntlizzieLet57_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeCTf_f_IntlizzieLet57_1_argbuf_rwb_r) && (! writeCTf_f_IntlizzieLet57_1_argbuf_bufchan_buf[0])))
        writeCTf_f_IntlizzieLet57_1_argbuf_bufchan_buf <= writeCTf_f_IntlizzieLet57_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CTf_f_Int) : (writeCTf_f_IntlizzieLet57_1_argbuf_rwb,Pointer_CTf_f_Int) > (lizzieLet36_1_1_argbuf,Pointer_CTf_f_Int) */
  Pointer_CTf_f_Int_t writeCTf_f_IntlizzieLet57_1_argbuf_rwb_bufchan_d;
  logic writeCTf_f_IntlizzieLet57_1_argbuf_rwb_bufchan_r;
  assign writeCTf_f_IntlizzieLet57_1_argbuf_rwb_r = ((! writeCTf_f_IntlizzieLet57_1_argbuf_rwb_bufchan_d[0]) || writeCTf_f_IntlizzieLet57_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTf_f_IntlizzieLet57_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCTf_f_IntlizzieLet57_1_argbuf_rwb_r)
        writeCTf_f_IntlizzieLet57_1_argbuf_rwb_bufchan_d <= writeCTf_f_IntlizzieLet57_1_argbuf_rwb_d;
  Pointer_CTf_f_Int_t writeCTf_f_IntlizzieLet57_1_argbuf_rwb_bufchan_buf;
  assign writeCTf_f_IntlizzieLet57_1_argbuf_rwb_bufchan_r = (! writeCTf_f_IntlizzieLet57_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet36_1_1_argbuf_d = (writeCTf_f_IntlizzieLet57_1_argbuf_rwb_bufchan_buf[0] ? writeCTf_f_IntlizzieLet57_1_argbuf_rwb_bufchan_buf :
                                     writeCTf_f_IntlizzieLet57_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTf_f_IntlizzieLet57_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((lizzieLet36_1_1_argbuf_r && writeCTf_f_IntlizzieLet57_1_argbuf_rwb_bufchan_buf[0]))
        writeCTf_f_IntlizzieLet57_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! lizzieLet36_1_1_argbuf_r) && (! writeCTf_f_IntlizzieLet57_1_argbuf_rwb_bufchan_buf[0])))
        writeCTf_f_IntlizzieLet57_1_argbuf_rwb_bufchan_buf <= writeCTf_f_IntlizzieLet57_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CTf_f_Int) : (writeCTf_f_IntlizzieLet68_1_argbuf,Pointer_CTf_f_Int) > (writeCTf_f_IntlizzieLet68_1_argbuf_rwb,Pointer_CTf_f_Int) */
  Pointer_CTf_f_Int_t writeCTf_f_IntlizzieLet68_1_argbuf_bufchan_d;
  logic writeCTf_f_IntlizzieLet68_1_argbuf_bufchan_r;
  assign writeCTf_f_IntlizzieLet68_1_argbuf_r = ((! writeCTf_f_IntlizzieLet68_1_argbuf_bufchan_d[0]) || writeCTf_f_IntlizzieLet68_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTf_f_IntlizzieLet68_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCTf_f_IntlizzieLet68_1_argbuf_r)
        writeCTf_f_IntlizzieLet68_1_argbuf_bufchan_d <= writeCTf_f_IntlizzieLet68_1_argbuf_d;
  Pointer_CTf_f_Int_t writeCTf_f_IntlizzieLet68_1_argbuf_bufchan_buf;
  assign writeCTf_f_IntlizzieLet68_1_argbuf_bufchan_r = (! writeCTf_f_IntlizzieLet68_1_argbuf_bufchan_buf[0]);
  assign writeCTf_f_IntlizzieLet68_1_argbuf_rwb_d = (writeCTf_f_IntlizzieLet68_1_argbuf_bufchan_buf[0] ? writeCTf_f_IntlizzieLet68_1_argbuf_bufchan_buf :
                                                     writeCTf_f_IntlizzieLet68_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTf_f_IntlizzieLet68_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeCTf_f_IntlizzieLet68_1_argbuf_rwb_r && writeCTf_f_IntlizzieLet68_1_argbuf_bufchan_buf[0]))
        writeCTf_f_IntlizzieLet68_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeCTf_f_IntlizzieLet68_1_argbuf_rwb_r) && (! writeCTf_f_IntlizzieLet68_1_argbuf_bufchan_buf[0])))
        writeCTf_f_IntlizzieLet68_1_argbuf_bufchan_buf <= writeCTf_f_IntlizzieLet68_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CTf_f_Int) : (writeCTf_f_IntlizzieLet68_1_argbuf_rwb,Pointer_CTf_f_Int) > (sca2_2_1_argbuf,Pointer_CTf_f_Int) */
  Pointer_CTf_f_Int_t writeCTf_f_IntlizzieLet68_1_argbuf_rwb_bufchan_d;
  logic writeCTf_f_IntlizzieLet68_1_argbuf_rwb_bufchan_r;
  assign writeCTf_f_IntlizzieLet68_1_argbuf_rwb_r = ((! writeCTf_f_IntlizzieLet68_1_argbuf_rwb_bufchan_d[0]) || writeCTf_f_IntlizzieLet68_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTf_f_IntlizzieLet68_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCTf_f_IntlizzieLet68_1_argbuf_rwb_r)
        writeCTf_f_IntlizzieLet68_1_argbuf_rwb_bufchan_d <= writeCTf_f_IntlizzieLet68_1_argbuf_rwb_d;
  Pointer_CTf_f_Int_t writeCTf_f_IntlizzieLet68_1_argbuf_rwb_bufchan_buf;
  assign writeCTf_f_IntlizzieLet68_1_argbuf_rwb_bufchan_r = (! writeCTf_f_IntlizzieLet68_1_argbuf_rwb_bufchan_buf[0]);
  assign sca2_2_1_argbuf_d = (writeCTf_f_IntlizzieLet68_1_argbuf_rwb_bufchan_buf[0] ? writeCTf_f_IntlizzieLet68_1_argbuf_rwb_bufchan_buf :
                              writeCTf_f_IntlizzieLet68_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTf_f_IntlizzieLet68_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((sca2_2_1_argbuf_r && writeCTf_f_IntlizzieLet68_1_argbuf_rwb_bufchan_buf[0]))
        writeCTf_f_IntlizzieLet68_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! sca2_2_1_argbuf_r) && (! writeCTf_f_IntlizzieLet68_1_argbuf_rwb_bufchan_buf[0])))
        writeCTf_f_IntlizzieLet68_1_argbuf_rwb_bufchan_buf <= writeCTf_f_IntlizzieLet68_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CTf_f_Int) : (writeCTf_f_IntlizzieLet69_1_argbuf,Pointer_CTf_f_Int) > (writeCTf_f_IntlizzieLet69_1_argbuf_rwb,Pointer_CTf_f_Int) */
  Pointer_CTf_f_Int_t writeCTf_f_IntlizzieLet69_1_argbuf_bufchan_d;
  logic writeCTf_f_IntlizzieLet69_1_argbuf_bufchan_r;
  assign writeCTf_f_IntlizzieLet69_1_argbuf_r = ((! writeCTf_f_IntlizzieLet69_1_argbuf_bufchan_d[0]) || writeCTf_f_IntlizzieLet69_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTf_f_IntlizzieLet69_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCTf_f_IntlizzieLet69_1_argbuf_r)
        writeCTf_f_IntlizzieLet69_1_argbuf_bufchan_d <= writeCTf_f_IntlizzieLet69_1_argbuf_d;
  Pointer_CTf_f_Int_t writeCTf_f_IntlizzieLet69_1_argbuf_bufchan_buf;
  assign writeCTf_f_IntlizzieLet69_1_argbuf_bufchan_r = (! writeCTf_f_IntlizzieLet69_1_argbuf_bufchan_buf[0]);
  assign writeCTf_f_IntlizzieLet69_1_argbuf_rwb_d = (writeCTf_f_IntlizzieLet69_1_argbuf_bufchan_buf[0] ? writeCTf_f_IntlizzieLet69_1_argbuf_bufchan_buf :
                                                     writeCTf_f_IntlizzieLet69_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTf_f_IntlizzieLet69_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeCTf_f_IntlizzieLet69_1_argbuf_rwb_r && writeCTf_f_IntlizzieLet69_1_argbuf_bufchan_buf[0]))
        writeCTf_f_IntlizzieLet69_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeCTf_f_IntlizzieLet69_1_argbuf_rwb_r) && (! writeCTf_f_IntlizzieLet69_1_argbuf_bufchan_buf[0])))
        writeCTf_f_IntlizzieLet69_1_argbuf_bufchan_buf <= writeCTf_f_IntlizzieLet69_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CTf_f_Int) : (writeCTf_f_IntlizzieLet69_1_argbuf_rwb,Pointer_CTf_f_Int) > (sca1_2_1_argbuf,Pointer_CTf_f_Int) */
  Pointer_CTf_f_Int_t writeCTf_f_IntlizzieLet69_1_argbuf_rwb_bufchan_d;
  logic writeCTf_f_IntlizzieLet69_1_argbuf_rwb_bufchan_r;
  assign writeCTf_f_IntlizzieLet69_1_argbuf_rwb_r = ((! writeCTf_f_IntlizzieLet69_1_argbuf_rwb_bufchan_d[0]) || writeCTf_f_IntlizzieLet69_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTf_f_IntlizzieLet69_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCTf_f_IntlizzieLet69_1_argbuf_rwb_r)
        writeCTf_f_IntlizzieLet69_1_argbuf_rwb_bufchan_d <= writeCTf_f_IntlizzieLet69_1_argbuf_rwb_d;
  Pointer_CTf_f_Int_t writeCTf_f_IntlizzieLet69_1_argbuf_rwb_bufchan_buf;
  assign writeCTf_f_IntlizzieLet69_1_argbuf_rwb_bufchan_r = (! writeCTf_f_IntlizzieLet69_1_argbuf_rwb_bufchan_buf[0]);
  assign sca1_2_1_argbuf_d = (writeCTf_f_IntlizzieLet69_1_argbuf_rwb_bufchan_buf[0] ? writeCTf_f_IntlizzieLet69_1_argbuf_rwb_bufchan_buf :
                              writeCTf_f_IntlizzieLet69_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTf_f_IntlizzieLet69_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((sca1_2_1_argbuf_r && writeCTf_f_IntlizzieLet69_1_argbuf_rwb_bufchan_buf[0]))
        writeCTf_f_IntlizzieLet69_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! sca1_2_1_argbuf_r) && (! writeCTf_f_IntlizzieLet69_1_argbuf_rwb_bufchan_buf[0])))
        writeCTf_f_IntlizzieLet69_1_argbuf_rwb_bufchan_buf <= writeCTf_f_IntlizzieLet69_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CTf_f_Int) : (writeCTf_f_IntlizzieLet70_1_argbuf,Pointer_CTf_f_Int) > (writeCTf_f_IntlizzieLet70_1_argbuf_rwb,Pointer_CTf_f_Int) */
  Pointer_CTf_f_Int_t writeCTf_f_IntlizzieLet70_1_argbuf_bufchan_d;
  logic writeCTf_f_IntlizzieLet70_1_argbuf_bufchan_r;
  assign writeCTf_f_IntlizzieLet70_1_argbuf_r = ((! writeCTf_f_IntlizzieLet70_1_argbuf_bufchan_d[0]) || writeCTf_f_IntlizzieLet70_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTf_f_IntlizzieLet70_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCTf_f_IntlizzieLet70_1_argbuf_r)
        writeCTf_f_IntlizzieLet70_1_argbuf_bufchan_d <= writeCTf_f_IntlizzieLet70_1_argbuf_d;
  Pointer_CTf_f_Int_t writeCTf_f_IntlizzieLet70_1_argbuf_bufchan_buf;
  assign writeCTf_f_IntlizzieLet70_1_argbuf_bufchan_r = (! writeCTf_f_IntlizzieLet70_1_argbuf_bufchan_buf[0]);
  assign writeCTf_f_IntlizzieLet70_1_argbuf_rwb_d = (writeCTf_f_IntlizzieLet70_1_argbuf_bufchan_buf[0] ? writeCTf_f_IntlizzieLet70_1_argbuf_bufchan_buf :
                                                     writeCTf_f_IntlizzieLet70_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTf_f_IntlizzieLet70_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeCTf_f_IntlizzieLet70_1_argbuf_rwb_r && writeCTf_f_IntlizzieLet70_1_argbuf_bufchan_buf[0]))
        writeCTf_f_IntlizzieLet70_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeCTf_f_IntlizzieLet70_1_argbuf_rwb_r) && (! writeCTf_f_IntlizzieLet70_1_argbuf_bufchan_buf[0])))
        writeCTf_f_IntlizzieLet70_1_argbuf_bufchan_buf <= writeCTf_f_IntlizzieLet70_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CTf_f_Int) : (writeCTf_f_IntlizzieLet70_1_argbuf_rwb,Pointer_CTf_f_Int) > (sca0_2_1_argbuf,Pointer_CTf_f_Int) */
  Pointer_CTf_f_Int_t writeCTf_f_IntlizzieLet70_1_argbuf_rwb_bufchan_d;
  logic writeCTf_f_IntlizzieLet70_1_argbuf_rwb_bufchan_r;
  assign writeCTf_f_IntlizzieLet70_1_argbuf_rwb_r = ((! writeCTf_f_IntlizzieLet70_1_argbuf_rwb_bufchan_d[0]) || writeCTf_f_IntlizzieLet70_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTf_f_IntlizzieLet70_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCTf_f_IntlizzieLet70_1_argbuf_rwb_r)
        writeCTf_f_IntlizzieLet70_1_argbuf_rwb_bufchan_d <= writeCTf_f_IntlizzieLet70_1_argbuf_rwb_d;
  Pointer_CTf_f_Int_t writeCTf_f_IntlizzieLet70_1_argbuf_rwb_bufchan_buf;
  assign writeCTf_f_IntlizzieLet70_1_argbuf_rwb_bufchan_r = (! writeCTf_f_IntlizzieLet70_1_argbuf_rwb_bufchan_buf[0]);
  assign sca0_2_1_argbuf_d = (writeCTf_f_IntlizzieLet70_1_argbuf_rwb_bufchan_buf[0] ? writeCTf_f_IntlizzieLet70_1_argbuf_rwb_bufchan_buf :
                              writeCTf_f_IntlizzieLet70_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTf_f_IntlizzieLet70_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((sca0_2_1_argbuf_r && writeCTf_f_IntlizzieLet70_1_argbuf_rwb_bufchan_buf[0]))
        writeCTf_f_IntlizzieLet70_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! sca0_2_1_argbuf_r) && (! writeCTf_f_IntlizzieLet70_1_argbuf_rwb_bufchan_buf[0])))
        writeCTf_f_IntlizzieLet70_1_argbuf_rwb_bufchan_buf <= writeCTf_f_IntlizzieLet70_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet10_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet10_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet10_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet10_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet10_1_argbuf_r = ((! writeQTree_IntlizzieLet10_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet10_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet10_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet10_1_argbuf_r)
        writeQTree_IntlizzieLet10_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet10_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet10_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet10_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet10_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet10_1_argbuf_rwb_d = (writeQTree_IntlizzieLet10_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet10_1_argbuf_bufchan_buf :
                                                     writeQTree_IntlizzieLet10_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet10_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet10_1_argbuf_rwb_r && writeQTree_IntlizzieLet10_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet10_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet10_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet10_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet10_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet10_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet10_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet2_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet10_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet10_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet10_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet10_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet10_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet10_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet10_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet10_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet10_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet10_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet10_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet10_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet2_1_1_argbuf_d = (writeQTree_IntlizzieLet10_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet10_1_argbuf_rwb_bufchan_buf :
                                    writeQTree_IntlizzieLet10_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet10_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((lizzieLet2_1_1_argbuf_r && writeQTree_IntlizzieLet10_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet10_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! lizzieLet2_1_1_argbuf_r) && (! writeQTree_IntlizzieLet10_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet10_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet10_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet11_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet11_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet11_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet11_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet11_1_argbuf_r = ((! writeQTree_IntlizzieLet11_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet11_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet11_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet11_1_argbuf_r)
        writeQTree_IntlizzieLet11_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet11_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet11_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet11_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet11_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet11_1_argbuf_rwb_d = (writeQTree_IntlizzieLet11_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet11_1_argbuf_bufchan_buf :
                                                     writeQTree_IntlizzieLet11_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet11_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet11_1_argbuf_rwb_r && writeQTree_IntlizzieLet11_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet11_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet11_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet11_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet11_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet11_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet11_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet3_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet11_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet11_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet11_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet11_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet11_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet11_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet11_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet11_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet11_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet11_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet11_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet11_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet3_1_1_argbuf_d = (writeQTree_IntlizzieLet11_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet11_1_argbuf_rwb_bufchan_buf :
                                    writeQTree_IntlizzieLet11_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet11_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((lizzieLet3_1_1_argbuf_r && writeQTree_IntlizzieLet11_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet11_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! lizzieLet3_1_1_argbuf_r) && (! writeQTree_IntlizzieLet11_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet11_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet11_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet13_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet13_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet13_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet13_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet13_1_argbuf_r = ((! writeQTree_IntlizzieLet13_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet13_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet13_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet13_1_argbuf_r)
        writeQTree_IntlizzieLet13_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet13_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet13_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet13_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet13_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet13_1_argbuf_rwb_d = (writeQTree_IntlizzieLet13_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet13_1_argbuf_bufchan_buf :
                                                     writeQTree_IntlizzieLet13_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet13_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet13_1_argbuf_rwb_r && writeQTree_IntlizzieLet13_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet13_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet13_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet13_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet13_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet13_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet13_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet4_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet13_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet13_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet13_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet13_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet13_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet13_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet13_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet13_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet13_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet13_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet13_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet13_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet4_1_1_argbuf_d = (writeQTree_IntlizzieLet13_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet13_1_argbuf_rwb_bufchan_buf :
                                    writeQTree_IntlizzieLet13_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet13_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((lizzieLet4_1_1_argbuf_r && writeQTree_IntlizzieLet13_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet13_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! lizzieLet4_1_1_argbuf_r) && (! writeQTree_IntlizzieLet13_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet13_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet13_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet15_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet15_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet15_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet15_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet15_1_argbuf_r = ((! writeQTree_IntlizzieLet15_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet15_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet15_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet15_1_argbuf_r)
        writeQTree_IntlizzieLet15_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet15_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet15_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet15_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet15_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet15_1_argbuf_rwb_d = (writeQTree_IntlizzieLet15_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet15_1_argbuf_bufchan_buf :
                                                     writeQTree_IntlizzieLet15_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet15_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet15_1_argbuf_rwb_r && writeQTree_IntlizzieLet15_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet15_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet15_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet15_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet15_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet15_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet15_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet5_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet15_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet15_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet15_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet15_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet15_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet15_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet15_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet15_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet15_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet15_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet15_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet15_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet5_1_1_argbuf_d = (writeQTree_IntlizzieLet15_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet15_1_argbuf_rwb_bufchan_buf :
                                    writeQTree_IntlizzieLet15_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet15_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((lizzieLet5_1_1_argbuf_r && writeQTree_IntlizzieLet15_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet15_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! lizzieLet5_1_1_argbuf_r) && (! writeQTree_IntlizzieLet15_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet15_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet15_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet16_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet16_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet16_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet16_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet16_1_argbuf_r = ((! writeQTree_IntlizzieLet16_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet16_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet16_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet16_1_argbuf_r)
        writeQTree_IntlizzieLet16_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet16_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet16_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet16_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet16_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet16_1_argbuf_rwb_d = (writeQTree_IntlizzieLet16_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet16_1_argbuf_bufchan_buf :
                                                     writeQTree_IntlizzieLet16_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet16_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet16_1_argbuf_rwb_r && writeQTree_IntlizzieLet16_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet16_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet16_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet16_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet16_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet16_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet16_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet6_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet16_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet16_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet16_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet16_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet16_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet16_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet16_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet16_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet16_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet16_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet16_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet16_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet6_1_1_argbuf_d = (writeQTree_IntlizzieLet16_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet16_1_argbuf_rwb_bufchan_buf :
                                    writeQTree_IntlizzieLet16_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet16_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((lizzieLet6_1_1_argbuf_r && writeQTree_IntlizzieLet16_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet16_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! lizzieLet6_1_1_argbuf_r) && (! writeQTree_IntlizzieLet16_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet16_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet16_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet20_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet20_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet20_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet20_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet20_1_argbuf_r = ((! writeQTree_IntlizzieLet20_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet20_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet20_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet20_1_argbuf_r)
        writeQTree_IntlizzieLet20_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet20_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet20_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet20_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet20_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet20_1_argbuf_rwb_d = (writeQTree_IntlizzieLet20_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet20_1_argbuf_bufchan_buf :
                                                     writeQTree_IntlizzieLet20_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet20_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet20_1_argbuf_rwb_r && writeQTree_IntlizzieLet20_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet20_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet20_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet20_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet20_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet20_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet20_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet8_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet20_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet20_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet20_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet20_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet20_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet20_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet20_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet20_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet20_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet20_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet20_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet20_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet8_1_1_argbuf_d = (writeQTree_IntlizzieLet20_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet20_1_argbuf_rwb_bufchan_buf :
                                    writeQTree_IntlizzieLet20_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet20_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((lizzieLet8_1_1_argbuf_r && writeQTree_IntlizzieLet20_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet20_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! lizzieLet8_1_1_argbuf_r) && (! writeQTree_IntlizzieLet20_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet20_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet20_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet21_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet21_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet21_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet21_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet21_1_argbuf_r = ((! writeQTree_IntlizzieLet21_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet21_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet21_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet21_1_argbuf_r)
        writeQTree_IntlizzieLet21_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet21_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet21_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet21_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet21_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet21_1_argbuf_rwb_d = (writeQTree_IntlizzieLet21_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet21_1_argbuf_bufchan_buf :
                                                     writeQTree_IntlizzieLet21_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet21_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet21_1_argbuf_rwb_r && writeQTree_IntlizzieLet21_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet21_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet21_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet21_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet21_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet21_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet21_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet9_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet21_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet21_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet21_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet21_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet21_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet21_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet21_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet21_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet21_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet21_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet21_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet21_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet9_1_1_argbuf_d = (writeQTree_IntlizzieLet21_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet21_1_argbuf_rwb_bufchan_buf :
                                    writeQTree_IntlizzieLet21_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet21_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((lizzieLet9_1_1_argbuf_r && writeQTree_IntlizzieLet21_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet21_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! lizzieLet9_1_1_argbuf_r) && (! writeQTree_IntlizzieLet21_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet21_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet21_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet22_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet22_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet22_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet22_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet22_1_argbuf_r = ((! writeQTree_IntlizzieLet22_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet22_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet22_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet22_1_argbuf_r)
        writeQTree_IntlizzieLet22_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet22_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet22_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet22_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet22_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet22_1_argbuf_rwb_d = (writeQTree_IntlizzieLet22_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet22_1_argbuf_bufchan_buf :
                                                     writeQTree_IntlizzieLet22_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet22_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet22_1_argbuf_rwb_r && writeQTree_IntlizzieLet22_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet22_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet22_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet22_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet22_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet22_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet22_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet10_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet22_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet22_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet22_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet22_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet22_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet22_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet22_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet22_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet22_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet22_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet22_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet22_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet10_1_1_argbuf_d = (writeQTree_IntlizzieLet22_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet22_1_argbuf_rwb_bufchan_buf :
                                     writeQTree_IntlizzieLet22_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet22_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((lizzieLet10_1_1_argbuf_r && writeQTree_IntlizzieLet22_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet22_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! lizzieLet10_1_1_argbuf_r) && (! writeQTree_IntlizzieLet22_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet22_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet22_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet23_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet23_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet23_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet23_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet23_1_argbuf_r = ((! writeQTree_IntlizzieLet23_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet23_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet23_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet23_1_argbuf_r)
        writeQTree_IntlizzieLet23_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet23_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet23_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet23_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet23_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet23_1_argbuf_rwb_d = (writeQTree_IntlizzieLet23_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet23_1_argbuf_bufchan_buf :
                                                     writeQTree_IntlizzieLet23_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet23_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet23_1_argbuf_rwb_r && writeQTree_IntlizzieLet23_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet23_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet23_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet23_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet23_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet23_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet23_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet11_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet23_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet23_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet23_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet23_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet23_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet23_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet23_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet23_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet23_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet23_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet23_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet23_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet11_1_1_argbuf_d = (writeQTree_IntlizzieLet23_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet23_1_argbuf_rwb_bufchan_buf :
                                     writeQTree_IntlizzieLet23_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet23_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((lizzieLet11_1_1_argbuf_r && writeQTree_IntlizzieLet23_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet23_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! lizzieLet11_1_1_argbuf_r) && (! writeQTree_IntlizzieLet23_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet23_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet23_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet25_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet25_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet25_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet25_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet25_1_argbuf_r = ((! writeQTree_IntlizzieLet25_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet25_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet25_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet25_1_argbuf_r)
        writeQTree_IntlizzieLet25_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet25_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet25_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet25_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet25_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet25_1_argbuf_rwb_d = (writeQTree_IntlizzieLet25_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet25_1_argbuf_bufchan_buf :
                                                     writeQTree_IntlizzieLet25_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet25_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet25_1_argbuf_rwb_r && writeQTree_IntlizzieLet25_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet25_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet25_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet25_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet25_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet25_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet25_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet12_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet25_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet25_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet25_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet25_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet25_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet25_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet25_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet25_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet25_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet25_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet25_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet25_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet12_1_argbuf_d = (writeQTree_IntlizzieLet25_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet25_1_argbuf_rwb_bufchan_buf :
                                   writeQTree_IntlizzieLet25_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet25_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((lizzieLet12_1_argbuf_r && writeQTree_IntlizzieLet25_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet25_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! lizzieLet12_1_argbuf_r) && (! writeQTree_IntlizzieLet25_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet25_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet25_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet26_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet26_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet26_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet26_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet26_1_argbuf_r = ((! writeQTree_IntlizzieLet26_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet26_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet26_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet26_1_argbuf_r)
        writeQTree_IntlizzieLet26_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet26_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet26_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet26_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet26_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet26_1_argbuf_rwb_d = (writeQTree_IntlizzieLet26_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet26_1_argbuf_bufchan_buf :
                                                     writeQTree_IntlizzieLet26_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet26_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet26_1_argbuf_rwb_r && writeQTree_IntlizzieLet26_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet26_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet26_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet26_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet26_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet26_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet26_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet13_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet26_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet26_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet26_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet26_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet26_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet26_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet26_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet26_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet26_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet26_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet26_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet26_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet13_1_1_argbuf_d = (writeQTree_IntlizzieLet26_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet26_1_argbuf_rwb_bufchan_buf :
                                     writeQTree_IntlizzieLet26_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet26_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((lizzieLet13_1_1_argbuf_r && writeQTree_IntlizzieLet26_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet26_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! lizzieLet13_1_1_argbuf_r) && (! writeQTree_IntlizzieLet26_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet26_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet26_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet27_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet27_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet27_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet27_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet27_1_argbuf_r = ((! writeQTree_IntlizzieLet27_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet27_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet27_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet27_1_argbuf_r)
        writeQTree_IntlizzieLet27_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet27_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet27_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet27_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet27_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet27_1_argbuf_rwb_d = (writeQTree_IntlizzieLet27_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet27_1_argbuf_bufchan_buf :
                                                     writeQTree_IntlizzieLet27_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet27_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet27_1_argbuf_rwb_r && writeQTree_IntlizzieLet27_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet27_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet27_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet27_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet27_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet27_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet27_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet14_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet27_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet27_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet27_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet27_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet27_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet27_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet27_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet27_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet27_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet27_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet27_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet27_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet14_1_1_argbuf_d = (writeQTree_IntlizzieLet27_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet27_1_argbuf_rwb_bufchan_buf :
                                     writeQTree_IntlizzieLet27_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet27_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((lizzieLet14_1_1_argbuf_r && writeQTree_IntlizzieLet27_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet27_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! lizzieLet14_1_1_argbuf_r) && (! writeQTree_IntlizzieLet27_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet27_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet27_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet28_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet28_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet28_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet28_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet28_1_argbuf_r = ((! writeQTree_IntlizzieLet28_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet28_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet28_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet28_1_argbuf_r)
        writeQTree_IntlizzieLet28_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet28_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet28_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet28_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet28_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet28_1_argbuf_rwb_d = (writeQTree_IntlizzieLet28_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet28_1_argbuf_bufchan_buf :
                                                     writeQTree_IntlizzieLet28_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet28_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet28_1_argbuf_rwb_r && writeQTree_IntlizzieLet28_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet28_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet28_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet28_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet28_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet28_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet28_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet15_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet28_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet28_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet28_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet28_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet28_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet28_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet28_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet28_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet28_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet28_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet28_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet28_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet15_1_1_argbuf_d = (writeQTree_IntlizzieLet28_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet28_1_argbuf_rwb_bufchan_buf :
                                     writeQTree_IntlizzieLet28_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet28_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((lizzieLet15_1_1_argbuf_r && writeQTree_IntlizzieLet28_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet28_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! lizzieLet15_1_1_argbuf_r) && (! writeQTree_IntlizzieLet28_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet28_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet28_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet31_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet31_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet31_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet31_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet31_1_argbuf_r = ((! writeQTree_IntlizzieLet31_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet31_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet31_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet31_1_argbuf_r)
        writeQTree_IntlizzieLet31_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet31_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet31_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet31_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet31_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet31_1_argbuf_rwb_d = (writeQTree_IntlizzieLet31_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet31_1_argbuf_bufchan_buf :
                                                     writeQTree_IntlizzieLet31_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet31_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet31_1_argbuf_rwb_r && writeQTree_IntlizzieLet31_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet31_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet31_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet31_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet31_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet31_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet31_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet16_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet31_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet31_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet31_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet31_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet31_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet31_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet31_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet31_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet31_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet31_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet31_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet31_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet16_1_1_argbuf_d = (writeQTree_IntlizzieLet31_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet31_1_argbuf_rwb_bufchan_buf :
                                     writeQTree_IntlizzieLet31_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet31_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((lizzieLet16_1_1_argbuf_r && writeQTree_IntlizzieLet31_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet31_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! lizzieLet16_1_1_argbuf_r) && (! writeQTree_IntlizzieLet31_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet31_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet31_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet32_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet32_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet32_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet32_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet32_1_argbuf_r = ((! writeQTree_IntlizzieLet32_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet32_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet32_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet32_1_argbuf_r)
        writeQTree_IntlizzieLet32_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet32_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet32_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet32_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet32_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet32_1_argbuf_rwb_d = (writeQTree_IntlizzieLet32_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet32_1_argbuf_bufchan_buf :
                                                     writeQTree_IntlizzieLet32_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet32_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet32_1_argbuf_rwb_r && writeQTree_IntlizzieLet32_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet32_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet32_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet32_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet32_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet32_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet32_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet17_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet32_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet32_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet32_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet32_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet32_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet32_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet32_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet32_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet32_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet32_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet32_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet32_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet17_1_1_argbuf_d = (writeQTree_IntlizzieLet32_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet32_1_argbuf_rwb_bufchan_buf :
                                     writeQTree_IntlizzieLet32_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet32_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((lizzieLet17_1_1_argbuf_r && writeQTree_IntlizzieLet32_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet32_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! lizzieLet17_1_1_argbuf_r) && (! writeQTree_IntlizzieLet32_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet32_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet32_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet33_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet33_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet33_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet33_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet33_1_argbuf_r = ((! writeQTree_IntlizzieLet33_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet33_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet33_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet33_1_argbuf_r)
        writeQTree_IntlizzieLet33_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet33_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet33_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet33_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet33_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet33_1_argbuf_rwb_d = (writeQTree_IntlizzieLet33_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet33_1_argbuf_bufchan_buf :
                                                     writeQTree_IntlizzieLet33_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet33_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet33_1_argbuf_rwb_r && writeQTree_IntlizzieLet33_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet33_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet33_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet33_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet33_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet33_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet33_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet18_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet33_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet33_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet33_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet33_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet33_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet33_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet33_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet33_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet33_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet33_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet33_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet33_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet18_1_1_argbuf_d = (writeQTree_IntlizzieLet33_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet33_1_argbuf_rwb_bufchan_buf :
                                     writeQTree_IntlizzieLet33_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet33_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((lizzieLet18_1_1_argbuf_r && writeQTree_IntlizzieLet33_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet33_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! lizzieLet18_1_1_argbuf_r) && (! writeQTree_IntlizzieLet33_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet33_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet33_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet34_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet34_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet34_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet34_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet34_1_argbuf_r = ((! writeQTree_IntlizzieLet34_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet34_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet34_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet34_1_argbuf_r)
        writeQTree_IntlizzieLet34_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet34_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet34_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet34_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet34_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet34_1_argbuf_rwb_d = (writeQTree_IntlizzieLet34_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet34_1_argbuf_bufchan_buf :
                                                     writeQTree_IntlizzieLet34_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet34_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet34_1_argbuf_rwb_r && writeQTree_IntlizzieLet34_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet34_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet34_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet34_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet34_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet34_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet34_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet19_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet34_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet34_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet34_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet34_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet34_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet34_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet34_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet34_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet34_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet34_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet34_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet34_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet19_1_1_argbuf_d = (writeQTree_IntlizzieLet34_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet34_1_argbuf_rwb_bufchan_buf :
                                     writeQTree_IntlizzieLet34_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet34_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((lizzieLet19_1_1_argbuf_r && writeQTree_IntlizzieLet34_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet34_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! lizzieLet19_1_1_argbuf_r) && (! writeQTree_IntlizzieLet34_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet34_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet34_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet36_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet36_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet36_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet36_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet36_1_argbuf_r = ((! writeQTree_IntlizzieLet36_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet36_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet36_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet36_1_argbuf_r)
        writeQTree_IntlizzieLet36_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet36_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet36_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet36_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet36_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet36_1_argbuf_rwb_d = (writeQTree_IntlizzieLet36_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet36_1_argbuf_bufchan_buf :
                                                     writeQTree_IntlizzieLet36_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet36_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet36_1_argbuf_rwb_r && writeQTree_IntlizzieLet36_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet36_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet36_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet36_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet36_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet36_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet36_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet20_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet36_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet36_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet36_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet36_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet36_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet36_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet36_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet36_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet36_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet36_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet36_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet36_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet20_1_1_argbuf_d = (writeQTree_IntlizzieLet36_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet36_1_argbuf_rwb_bufchan_buf :
                                     writeQTree_IntlizzieLet36_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet36_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((lizzieLet20_1_1_argbuf_r && writeQTree_IntlizzieLet36_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet36_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! lizzieLet20_1_1_argbuf_r) && (! writeQTree_IntlizzieLet36_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet36_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet36_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet37_2_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet37_2_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet37_2_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet37_2_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet37_2_1_argbuf_r = ((! writeQTree_IntlizzieLet37_2_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet37_2_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet37_2_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet37_2_1_argbuf_r)
        writeQTree_IntlizzieLet37_2_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet37_2_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet37_2_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet37_2_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet37_2_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet37_2_1_argbuf_rwb_d = (writeQTree_IntlizzieLet37_2_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet37_2_1_argbuf_bufchan_buf :
                                                       writeQTree_IntlizzieLet37_2_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet37_2_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet37_2_1_argbuf_rwb_r && writeQTree_IntlizzieLet37_2_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet37_2_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet37_2_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet37_2_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet37_2_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet37_2_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet37_2_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet21_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet37_2_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet37_2_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet37_2_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet37_2_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet37_2_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet37_2_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                             1'd0};
    else
      if (writeQTree_IntlizzieLet37_2_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet37_2_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet37_2_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet37_2_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet37_2_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet37_2_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet21_1_1_argbuf_d = (writeQTree_IntlizzieLet37_2_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet37_2_1_argbuf_rwb_bufchan_buf :
                                     writeQTree_IntlizzieLet37_2_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet37_2_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
    else
      if ((lizzieLet21_1_1_argbuf_r && writeQTree_IntlizzieLet37_2_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet37_2_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                 1'd0};
      else if (((! lizzieLet21_1_1_argbuf_r) && (! writeQTree_IntlizzieLet37_2_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet37_2_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet37_2_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet38_1_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet38_1_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet38_1_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet38_1_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet38_1_1_argbuf_r = ((! writeQTree_IntlizzieLet38_1_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet38_1_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet38_1_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet38_1_1_argbuf_r)
        writeQTree_IntlizzieLet38_1_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet38_1_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet38_1_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet38_1_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet38_1_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet38_1_1_argbuf_rwb_d = (writeQTree_IntlizzieLet38_1_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet38_1_1_argbuf_bufchan_buf :
                                                       writeQTree_IntlizzieLet38_1_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet38_1_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet38_1_1_argbuf_rwb_r && writeQTree_IntlizzieLet38_1_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet38_1_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet38_1_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet38_1_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet38_1_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet38_1_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet38_1_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet22_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet38_1_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet38_1_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet38_1_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet38_1_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet38_1_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet38_1_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                             1'd0};
    else
      if (writeQTree_IntlizzieLet38_1_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet38_1_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet38_1_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet38_1_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet38_1_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet38_1_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet22_1_1_argbuf_d = (writeQTree_IntlizzieLet38_1_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet38_1_1_argbuf_rwb_bufchan_buf :
                                     writeQTree_IntlizzieLet38_1_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet38_1_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
    else
      if ((lizzieLet22_1_1_argbuf_r && writeQTree_IntlizzieLet38_1_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet38_1_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                 1'd0};
      else if (((! lizzieLet22_1_1_argbuf_r) && (! writeQTree_IntlizzieLet38_1_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet38_1_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet38_1_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet39_1_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet39_1_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet39_1_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet39_1_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet39_1_1_argbuf_r = ((! writeQTree_IntlizzieLet39_1_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet39_1_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet39_1_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet39_1_1_argbuf_r)
        writeQTree_IntlizzieLet39_1_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet39_1_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet39_1_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet39_1_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet39_1_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet39_1_1_argbuf_rwb_d = (writeQTree_IntlizzieLet39_1_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet39_1_1_argbuf_bufchan_buf :
                                                       writeQTree_IntlizzieLet39_1_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet39_1_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet39_1_1_argbuf_rwb_r && writeQTree_IntlizzieLet39_1_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet39_1_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet39_1_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet39_1_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet39_1_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet39_1_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet39_1_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet23_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet39_1_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet39_1_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet39_1_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet39_1_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet39_1_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet39_1_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                             1'd0};
    else
      if (writeQTree_IntlizzieLet39_1_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet39_1_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet39_1_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet39_1_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet39_1_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet39_1_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet23_1_1_argbuf_d = (writeQTree_IntlizzieLet39_1_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet39_1_1_argbuf_rwb_bufchan_buf :
                                     writeQTree_IntlizzieLet39_1_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet39_1_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
    else
      if ((lizzieLet23_1_1_argbuf_r && writeQTree_IntlizzieLet39_1_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet39_1_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                 1'd0};
      else if (((! lizzieLet23_1_1_argbuf_r) && (! writeQTree_IntlizzieLet39_1_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet39_1_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet39_1_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet40_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet40_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet40_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet40_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet40_1_argbuf_r = ((! writeQTree_IntlizzieLet40_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet40_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet40_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet40_1_argbuf_r)
        writeQTree_IntlizzieLet40_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet40_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet40_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet40_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet40_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet40_1_argbuf_rwb_d = (writeQTree_IntlizzieLet40_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet40_1_argbuf_bufchan_buf :
                                                     writeQTree_IntlizzieLet40_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet40_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet40_1_argbuf_rwb_r && writeQTree_IntlizzieLet40_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet40_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet40_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet40_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet40_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet40_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet40_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet24_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet40_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet40_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet40_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet40_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet40_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet40_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet40_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet40_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet40_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet40_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet40_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet40_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet24_1_argbuf_d = (writeQTree_IntlizzieLet40_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet40_1_argbuf_rwb_bufchan_buf :
                                   writeQTree_IntlizzieLet40_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet40_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((lizzieLet24_1_argbuf_r && writeQTree_IntlizzieLet40_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet40_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! lizzieLet24_1_argbuf_r) && (! writeQTree_IntlizzieLet40_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet40_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet40_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet41_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet41_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet41_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet41_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet41_1_argbuf_r = ((! writeQTree_IntlizzieLet41_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet41_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet41_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet41_1_argbuf_r)
        writeQTree_IntlizzieLet41_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet41_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet41_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet41_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet41_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet41_1_argbuf_rwb_d = (writeQTree_IntlizzieLet41_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet41_1_argbuf_bufchan_buf :
                                                     writeQTree_IntlizzieLet41_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet41_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet41_1_argbuf_rwb_r && writeQTree_IntlizzieLet41_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet41_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet41_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet41_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet41_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet41_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet41_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet25_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet41_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet41_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet41_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet41_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet41_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet41_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet41_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet41_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet41_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet41_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet41_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet41_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet25_1_1_argbuf_d = (writeQTree_IntlizzieLet41_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet41_1_argbuf_rwb_bufchan_buf :
                                     writeQTree_IntlizzieLet41_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet41_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((lizzieLet25_1_1_argbuf_r && writeQTree_IntlizzieLet41_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet41_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! lizzieLet25_1_1_argbuf_r) && (! writeQTree_IntlizzieLet41_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet41_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet41_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet42_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet42_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet42_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet42_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet42_1_argbuf_r = ((! writeQTree_IntlizzieLet42_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet42_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet42_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet42_1_argbuf_r)
        writeQTree_IntlizzieLet42_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet42_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet42_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet42_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet42_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet42_1_argbuf_rwb_d = (writeQTree_IntlizzieLet42_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet42_1_argbuf_bufchan_buf :
                                                     writeQTree_IntlizzieLet42_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet42_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet42_1_argbuf_rwb_r && writeQTree_IntlizzieLet42_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet42_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet42_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet42_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet42_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet42_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet42_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet26_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet42_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet42_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet42_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet42_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet42_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet42_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet42_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet42_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet42_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet42_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet42_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet42_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet26_1_1_argbuf_d = (writeQTree_IntlizzieLet42_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet42_1_argbuf_rwb_bufchan_buf :
                                     writeQTree_IntlizzieLet42_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet42_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((lizzieLet26_1_1_argbuf_r && writeQTree_IntlizzieLet42_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet42_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! lizzieLet26_1_1_argbuf_r) && (! writeQTree_IntlizzieLet42_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet42_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet42_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet45_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet45_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet45_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet45_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet45_1_argbuf_r = ((! writeQTree_IntlizzieLet45_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet45_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet45_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet45_1_argbuf_r)
        writeQTree_IntlizzieLet45_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet45_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet45_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet45_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet45_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet45_1_argbuf_rwb_d = (writeQTree_IntlizzieLet45_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet45_1_argbuf_bufchan_buf :
                                                     writeQTree_IntlizzieLet45_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet45_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet45_1_argbuf_rwb_r && writeQTree_IntlizzieLet45_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet45_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet45_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet45_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet45_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet45_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet45_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet27_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet45_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet45_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet45_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet45_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet45_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet45_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet45_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet45_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet45_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet45_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet45_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet45_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet27_1_1_argbuf_d = (writeQTree_IntlizzieLet45_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet45_1_argbuf_rwb_bufchan_buf :
                                     writeQTree_IntlizzieLet45_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet45_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((lizzieLet27_1_1_argbuf_r && writeQTree_IntlizzieLet45_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet45_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! lizzieLet27_1_1_argbuf_r) && (! writeQTree_IntlizzieLet45_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet45_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet45_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet46_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet46_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet46_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet46_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet46_1_argbuf_r = ((! writeQTree_IntlizzieLet46_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet46_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet46_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet46_1_argbuf_r)
        writeQTree_IntlizzieLet46_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet46_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet46_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet46_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet46_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet46_1_argbuf_rwb_d = (writeQTree_IntlizzieLet46_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet46_1_argbuf_bufchan_buf :
                                                     writeQTree_IntlizzieLet46_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet46_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet46_1_argbuf_rwb_r && writeQTree_IntlizzieLet46_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet46_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet46_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet46_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet46_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet46_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet46_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet28_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet46_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet46_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet46_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet46_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet46_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet46_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet46_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet46_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet46_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet46_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet46_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet46_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet28_1_1_argbuf_d = (writeQTree_IntlizzieLet46_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet46_1_argbuf_rwb_bufchan_buf :
                                     writeQTree_IntlizzieLet46_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet46_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((lizzieLet28_1_1_argbuf_r && writeQTree_IntlizzieLet46_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet46_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! lizzieLet28_1_1_argbuf_r) && (! writeQTree_IntlizzieLet46_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet46_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet46_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet47_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet47_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet47_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet47_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet47_1_argbuf_r = ((! writeQTree_IntlizzieLet47_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet47_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet47_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet47_1_argbuf_r)
        writeQTree_IntlizzieLet47_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet47_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet47_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet47_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet47_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet47_1_argbuf_rwb_d = (writeQTree_IntlizzieLet47_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet47_1_argbuf_bufchan_buf :
                                                     writeQTree_IntlizzieLet47_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet47_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet47_1_argbuf_rwb_r && writeQTree_IntlizzieLet47_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet47_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet47_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet47_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet47_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet47_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet47_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet29_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet47_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet47_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet47_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet47_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet47_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet47_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet47_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet47_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet47_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet47_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet47_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet47_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet29_1_argbuf_d = (writeQTree_IntlizzieLet47_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet47_1_argbuf_rwb_bufchan_buf :
                                   writeQTree_IntlizzieLet47_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet47_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((lizzieLet29_1_argbuf_r && writeQTree_IntlizzieLet47_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet47_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! lizzieLet29_1_argbuf_r) && (! writeQTree_IntlizzieLet47_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet47_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet47_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet48_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet48_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet48_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet48_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet48_1_argbuf_r = ((! writeQTree_IntlizzieLet48_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet48_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet48_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet48_1_argbuf_r)
        writeQTree_IntlizzieLet48_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet48_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet48_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet48_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet48_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet48_1_argbuf_rwb_d = (writeQTree_IntlizzieLet48_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet48_1_argbuf_bufchan_buf :
                                                     writeQTree_IntlizzieLet48_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet48_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet48_1_argbuf_rwb_r && writeQTree_IntlizzieLet48_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet48_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet48_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet48_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet48_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet48_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet48_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet30_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet48_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet48_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet48_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet48_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet48_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet48_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet48_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet48_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet48_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet48_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet48_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet48_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet30_1_argbuf_d = (writeQTree_IntlizzieLet48_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet48_1_argbuf_rwb_bufchan_buf :
                                   writeQTree_IntlizzieLet48_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet48_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((lizzieLet30_1_argbuf_r && writeQTree_IntlizzieLet48_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet48_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! lizzieLet30_1_argbuf_r) && (! writeQTree_IntlizzieLet48_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet48_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet48_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet50_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet50_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet50_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet50_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet50_1_argbuf_r = ((! writeQTree_IntlizzieLet50_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet50_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet50_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet50_1_argbuf_r)
        writeQTree_IntlizzieLet50_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet50_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet50_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet50_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet50_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet50_1_argbuf_rwb_d = (writeQTree_IntlizzieLet50_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet50_1_argbuf_bufchan_buf :
                                                     writeQTree_IntlizzieLet50_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet50_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet50_1_argbuf_rwb_r && writeQTree_IntlizzieLet50_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet50_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet50_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet50_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet50_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet50_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet50_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet31_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet50_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet50_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet50_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet50_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet50_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet50_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet50_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet50_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet50_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet50_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet50_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet50_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet31_1_1_argbuf_d = (writeQTree_IntlizzieLet50_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet50_1_argbuf_rwb_bufchan_buf :
                                     writeQTree_IntlizzieLet50_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet50_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((lizzieLet31_1_1_argbuf_r && writeQTree_IntlizzieLet50_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet50_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! lizzieLet31_1_1_argbuf_r) && (! writeQTree_IntlizzieLet50_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet50_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet50_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet51_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet51_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet51_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet51_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet51_1_argbuf_r = ((! writeQTree_IntlizzieLet51_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet51_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet51_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet51_1_argbuf_r)
        writeQTree_IntlizzieLet51_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet51_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet51_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet51_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet51_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet51_1_argbuf_rwb_d = (writeQTree_IntlizzieLet51_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet51_1_argbuf_bufchan_buf :
                                                     writeQTree_IntlizzieLet51_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet51_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet51_1_argbuf_rwb_r && writeQTree_IntlizzieLet51_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet51_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet51_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet51_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet51_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet51_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet51_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet32_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet51_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet51_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet51_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet51_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet51_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet51_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet51_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet51_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet51_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet51_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet51_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet51_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet32_1_1_argbuf_d = (writeQTree_IntlizzieLet51_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet51_1_argbuf_rwb_bufchan_buf :
                                     writeQTree_IntlizzieLet51_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet51_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((lizzieLet32_1_1_argbuf_r && writeQTree_IntlizzieLet51_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet51_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! lizzieLet32_1_1_argbuf_r) && (! writeQTree_IntlizzieLet51_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet51_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet51_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet53_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet53_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet53_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet53_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet53_1_argbuf_r = ((! writeQTree_IntlizzieLet53_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet53_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet53_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet53_1_argbuf_r)
        writeQTree_IntlizzieLet53_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet53_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet53_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet53_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet53_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet53_1_argbuf_rwb_d = (writeQTree_IntlizzieLet53_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet53_1_argbuf_bufchan_buf :
                                                     writeQTree_IntlizzieLet53_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet53_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet53_1_argbuf_rwb_r && writeQTree_IntlizzieLet53_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet53_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet53_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet53_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet53_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet53_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet53_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet33_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet53_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet53_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet53_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet53_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet53_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet53_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet53_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet53_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet53_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet53_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet53_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet53_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet33_1_1_argbuf_d = (writeQTree_IntlizzieLet53_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet53_1_argbuf_rwb_bufchan_buf :
                                     writeQTree_IntlizzieLet53_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet53_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((lizzieLet33_1_1_argbuf_r && writeQTree_IntlizzieLet53_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet53_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! lizzieLet33_1_1_argbuf_r) && (! writeQTree_IntlizzieLet53_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet53_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet53_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet54_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet54_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet54_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet54_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet54_1_argbuf_r = ((! writeQTree_IntlizzieLet54_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet54_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet54_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet54_1_argbuf_r)
        writeQTree_IntlizzieLet54_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet54_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet54_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet54_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet54_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet54_1_argbuf_rwb_d = (writeQTree_IntlizzieLet54_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet54_1_argbuf_bufchan_buf :
                                                     writeQTree_IntlizzieLet54_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet54_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet54_1_argbuf_rwb_r && writeQTree_IntlizzieLet54_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet54_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet54_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet54_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet54_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet54_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet54_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet34_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet54_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet54_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet54_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet54_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet54_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet54_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet54_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet54_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet54_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet54_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet54_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet54_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet34_1_1_argbuf_d = (writeQTree_IntlizzieLet54_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet54_1_argbuf_rwb_bufchan_buf :
                                     writeQTree_IntlizzieLet54_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet54_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((lizzieLet34_1_1_argbuf_r && writeQTree_IntlizzieLet54_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet54_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! lizzieLet34_1_1_argbuf_r) && (! writeQTree_IntlizzieLet54_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet54_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet54_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet55_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet55_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet55_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet55_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet55_1_argbuf_r = ((! writeQTree_IntlizzieLet55_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet55_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet55_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet55_1_argbuf_r)
        writeQTree_IntlizzieLet55_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet55_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet55_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet55_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet55_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet55_1_argbuf_rwb_d = (writeQTree_IntlizzieLet55_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet55_1_argbuf_bufchan_buf :
                                                     writeQTree_IntlizzieLet55_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet55_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet55_1_argbuf_rwb_r && writeQTree_IntlizzieLet55_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet55_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet55_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet55_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet55_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet55_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet55_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet35_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet55_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet55_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet55_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet55_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet55_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet55_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet55_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet55_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet55_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet55_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet55_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet55_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet35_1_argbuf_d = (writeQTree_IntlizzieLet55_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet55_1_argbuf_rwb_bufchan_buf :
                                   writeQTree_IntlizzieLet55_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet55_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((lizzieLet35_1_argbuf_r && writeQTree_IntlizzieLet55_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet55_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! lizzieLet35_1_argbuf_r) && (! writeQTree_IntlizzieLet55_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet55_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet55_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet66_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet66_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet66_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet66_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet66_1_argbuf_r = ((! writeQTree_IntlizzieLet66_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet66_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet66_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet66_1_argbuf_r)
        writeQTree_IntlizzieLet66_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet66_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet66_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet66_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet66_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet66_1_argbuf_rwb_d = (writeQTree_IntlizzieLet66_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet66_1_argbuf_bufchan_buf :
                                                     writeQTree_IntlizzieLet66_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet66_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet66_1_argbuf_rwb_r && writeQTree_IntlizzieLet66_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet66_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet66_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet66_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet66_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet66_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet66_1_argbuf_rwb,Pointer_QTree_Int) > (contRet_0_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet66_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet66_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet66_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet66_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet66_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet66_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet66_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet66_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet66_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet66_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet66_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet66_1_argbuf_rwb_bufchan_buf[0]);
  assign contRet_0_1_1_argbuf_d = (writeQTree_IntlizzieLet66_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet66_1_argbuf_rwb_bufchan_buf :
                                   writeQTree_IntlizzieLet66_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet66_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((contRet_0_1_1_argbuf_r && writeQTree_IntlizzieLet66_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet66_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! contRet_0_1_1_argbuf_r) && (! writeQTree_IntlizzieLet66_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet66_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet66_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet71_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet71_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet71_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet71_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet71_1_argbuf_r = ((! writeQTree_IntlizzieLet71_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet71_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet71_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet71_1_argbuf_r)
        writeQTree_IntlizzieLet71_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet71_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet71_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet71_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet71_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet71_1_argbuf_rwb_d = (writeQTree_IntlizzieLet71_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet71_1_argbuf_bufchan_buf :
                                                     writeQTree_IntlizzieLet71_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet71_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet71_1_argbuf_rwb_r && writeQTree_IntlizzieLet71_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet71_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet71_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet71_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet71_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet71_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet71_1_argbuf_rwb,Pointer_QTree_Int) > (contRet_0_2_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet71_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet71_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet71_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet71_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet71_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet71_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet71_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet71_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet71_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet71_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet71_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet71_1_argbuf_rwb_bufchan_buf[0]);
  assign contRet_0_2_1_argbuf_d = (writeQTree_IntlizzieLet71_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet71_1_argbuf_rwb_bufchan_buf :
                                   writeQTree_IntlizzieLet71_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet71_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((contRet_0_2_1_argbuf_r && writeQTree_IntlizzieLet71_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet71_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! contRet_0_2_1_argbuf_r) && (! writeQTree_IntlizzieLet71_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet71_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet71_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet8_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet8_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet8_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet8_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet8_1_argbuf_r = ((! writeQTree_IntlizzieLet8_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet8_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet8_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet8_1_argbuf_r)
        writeQTree_IntlizzieLet8_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet8_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet8_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet8_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet8_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet8_1_argbuf_rwb_d = (writeQTree_IntlizzieLet8_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet8_1_argbuf_bufchan_buf :
                                                    writeQTree_IntlizzieLet8_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet8_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet8_1_argbuf_rwb_r && writeQTree_IntlizzieLet8_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet8_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet8_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet8_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet8_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet8_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet8_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet0_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet8_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet8_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet8_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet8_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet8_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet8_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet8_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet8_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet8_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet8_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet8_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet8_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet0_1_1_argbuf_d = (writeQTree_IntlizzieLet8_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet8_1_argbuf_rwb_bufchan_buf :
                                    writeQTree_IntlizzieLet8_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet8_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet0_1_1_argbuf_r && writeQTree_IntlizzieLet8_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet8_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet0_1_1_argbuf_r) && (! writeQTree_IntlizzieLet8_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet8_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet8_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet9_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet9_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet9_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet9_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet9_1_argbuf_r = ((! writeQTree_IntlizzieLet9_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet9_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet9_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet9_1_argbuf_r)
        writeQTree_IntlizzieLet9_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet9_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet9_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet9_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet9_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet9_1_argbuf_rwb_d = (writeQTree_IntlizzieLet9_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet9_1_argbuf_bufchan_buf :
                                                    writeQTree_IntlizzieLet9_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet9_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet9_1_argbuf_rwb_r && writeQTree_IntlizzieLet9_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet9_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet9_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet9_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet9_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet9_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet9_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet1_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet9_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet9_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet9_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet9_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet9_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet9_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet9_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet9_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet9_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet9_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet9_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet9_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet1_1_1_argbuf_d = (writeQTree_IntlizzieLet9_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet9_1_argbuf_rwb_bufchan_buf :
                                    writeQTree_IntlizzieLet9_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet9_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet1_1_1_argbuf_r && writeQTree_IntlizzieLet9_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet9_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet1_1_1_argbuf_r) && (! writeQTree_IntlizzieLet9_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet9_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet9_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (wsmk_1_goMux_mux,Pointer_QTree_Int) > (wsmk_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t wsmk_1_goMux_mux_bufchan_d;
  logic wsmk_1_goMux_mux_bufchan_r;
  assign wsmk_1_goMux_mux_r = ((! wsmk_1_goMux_mux_bufchan_d[0]) || wsmk_1_goMux_mux_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) wsmk_1_goMux_mux_bufchan_d <= {16'd0, 1'd0};
    else
      if (wsmk_1_goMux_mux_r)
        wsmk_1_goMux_mux_bufchan_d <= wsmk_1_goMux_mux_d;
  Pointer_QTree_Int_t wsmk_1_goMux_mux_bufchan_buf;
  assign wsmk_1_goMux_mux_bufchan_r = (! wsmk_1_goMux_mux_bufchan_buf[0]);
  assign wsmk_1_1_argbuf_d = (wsmk_1_goMux_mux_bufchan_buf[0] ? wsmk_1_goMux_mux_bufchan_buf :
                              wsmk_1_goMux_mux_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) wsmk_1_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((wsmk_1_1_argbuf_r && wsmk_1_goMux_mux_bufchan_buf[0]))
        wsmk_1_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
      else if (((! wsmk_1_1_argbuf_r) && (! wsmk_1_goMux_mux_bufchan_buf[0])))
        wsmk_1_goMux_mux_bufchan_buf <= wsmk_1_goMux_mux_bufchan_d;
  
  /* buf (Ty CT$wnnz) : (wwsmn_2_1lizzieLet58_4Lcall_$wnnz2_1sc_0_4_1q4a8u_2_1Lcall_$wnnz1,CT$wnnz) > (lizzieLet60_1_argbuf,CT$wnnz) */
  CT$wnnz_t wwsmn_2_1lizzieLet58_4Lcall_$wnnz2_1sc_0_4_1q4a8u_2_1Lcall_$wnnz1_bufchan_d;
  logic wwsmn_2_1lizzieLet58_4Lcall_$wnnz2_1sc_0_4_1q4a8u_2_1Lcall_$wnnz1_bufchan_r;
  assign wwsmn_2_1lizzieLet58_4Lcall_$wnnz2_1sc_0_4_1q4a8u_2_1Lcall_$wnnz1_r = ((! wwsmn_2_1lizzieLet58_4Lcall_$wnnz2_1sc_0_4_1q4a8u_2_1Lcall_$wnnz1_bufchan_d[0]) || wwsmn_2_1lizzieLet58_4Lcall_$wnnz2_1sc_0_4_1q4a8u_2_1Lcall_$wnnz1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      wwsmn_2_1lizzieLet58_4Lcall_$wnnz2_1sc_0_4_1q4a8u_2_1Lcall_$wnnz1_bufchan_d <= {115'd0,
                                                                                      1'd0};
    else
      if (wwsmn_2_1lizzieLet58_4Lcall_$wnnz2_1sc_0_4_1q4a8u_2_1Lcall_$wnnz1_r)
        wwsmn_2_1lizzieLet58_4Lcall_$wnnz2_1sc_0_4_1q4a8u_2_1Lcall_$wnnz1_bufchan_d <= wwsmn_2_1lizzieLet58_4Lcall_$wnnz2_1sc_0_4_1q4a8u_2_1Lcall_$wnnz1_d;
  CT$wnnz_t wwsmn_2_1lizzieLet58_4Lcall_$wnnz2_1sc_0_4_1q4a8u_2_1Lcall_$wnnz1_bufchan_buf;
  assign wwsmn_2_1lizzieLet58_4Lcall_$wnnz2_1sc_0_4_1q4a8u_2_1Lcall_$wnnz1_bufchan_r = (! wwsmn_2_1lizzieLet58_4Lcall_$wnnz2_1sc_0_4_1q4a8u_2_1Lcall_$wnnz1_bufchan_buf[0]);
  assign lizzieLet60_1_argbuf_d = (wwsmn_2_1lizzieLet58_4Lcall_$wnnz2_1sc_0_4_1q4a8u_2_1Lcall_$wnnz1_bufchan_buf[0] ? wwsmn_2_1lizzieLet58_4Lcall_$wnnz2_1sc_0_4_1q4a8u_2_1Lcall_$wnnz1_bufchan_buf :
                                   wwsmn_2_1lizzieLet58_4Lcall_$wnnz2_1sc_0_4_1q4a8u_2_1Lcall_$wnnz1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      wwsmn_2_1lizzieLet58_4Lcall_$wnnz2_1sc_0_4_1q4a8u_2_1Lcall_$wnnz1_bufchan_buf <= {115'd0,
                                                                                        1'd0};
    else
      if ((lizzieLet60_1_argbuf_r && wwsmn_2_1lizzieLet58_4Lcall_$wnnz2_1sc_0_4_1q4a8u_2_1Lcall_$wnnz1_bufchan_buf[0]))
        wwsmn_2_1lizzieLet58_4Lcall_$wnnz2_1sc_0_4_1q4a8u_2_1Lcall_$wnnz1_bufchan_buf <= {115'd0,
                                                                                          1'd0};
      else if (((! lizzieLet60_1_argbuf_r) && (! wwsmn_2_1lizzieLet58_4Lcall_$wnnz2_1sc_0_4_1q4a8u_2_1Lcall_$wnnz1_bufchan_buf[0])))
        wwsmn_2_1lizzieLet58_4Lcall_$wnnz2_1sc_0_4_1q4a8u_2_1Lcall_$wnnz1_bufchan_buf <= wwsmn_2_1lizzieLet58_4Lcall_$wnnz2_1sc_0_4_1q4a8u_2_1Lcall_$wnnz1_bufchan_d;
  
  /* dcon (Ty CT$wnnz,Dcon Lcall_$wnnz1) : [(wwsmn_2_destruct,Int#),
                                       (lizzieLet58_4Lcall_$wnnz2,Int#),
                                       (sc_0_4_destruct,Pointer_CT$wnnz),
                                       (q4a8u_2_destruct,Pointer_QTree_Int)] > (wwsmn_2_1lizzieLet58_4Lcall_$wnnz2_1sc_0_4_1q4a8u_2_1Lcall_$wnnz1,CT$wnnz) */
  assign wwsmn_2_1lizzieLet58_4Lcall_$wnnz2_1sc_0_4_1q4a8u_2_1Lcall_$wnnz1_d = Lcall_$wnnz1_dc((& {wwsmn_2_destruct_d[0],
                                                                                                   lizzieLet58_4Lcall_$wnnz2_d[0],
                                                                                                   sc_0_4_destruct_d[0],
                                                                                                   q4a8u_2_destruct_d[0]}), wwsmn_2_destruct_d, lizzieLet58_4Lcall_$wnnz2_d, sc_0_4_destruct_d, q4a8u_2_destruct_d);
  assign {wwsmn_2_destruct_r,
          lizzieLet58_4Lcall_$wnnz2_r,
          sc_0_4_destruct_r,
          q4a8u_2_destruct_r} = {4 {(wwsmn_2_1lizzieLet58_4Lcall_$wnnz2_1sc_0_4_1q4a8u_2_1Lcall_$wnnz1_r && wwsmn_2_1lizzieLet58_4Lcall_$wnnz2_1sc_0_4_1q4a8u_2_1Lcall_$wnnz1_d[0])}};
  
  /* buf (Ty CT$wnnz) : (wwsmn_3_1ww1XmW_1_1lizzieLet58_4Lcall_$wnnz1_1sc_0_5_1Lcall_$wnnz0,CT$wnnz) > (lizzieLet61_1_argbuf,CT$wnnz) */
  CT$wnnz_t wwsmn_3_1ww1XmW_1_1lizzieLet58_4Lcall_$wnnz1_1sc_0_5_1Lcall_$wnnz0_bufchan_d;
  logic wwsmn_3_1ww1XmW_1_1lizzieLet58_4Lcall_$wnnz1_1sc_0_5_1Lcall_$wnnz0_bufchan_r;
  assign wwsmn_3_1ww1XmW_1_1lizzieLet58_4Lcall_$wnnz1_1sc_0_5_1Lcall_$wnnz0_r = ((! wwsmn_3_1ww1XmW_1_1lizzieLet58_4Lcall_$wnnz1_1sc_0_5_1Lcall_$wnnz0_bufchan_d[0]) || wwsmn_3_1ww1XmW_1_1lizzieLet58_4Lcall_$wnnz1_1sc_0_5_1Lcall_$wnnz0_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      wwsmn_3_1ww1XmW_1_1lizzieLet58_4Lcall_$wnnz1_1sc_0_5_1Lcall_$wnnz0_bufchan_d <= {115'd0,
                                                                                       1'd0};
    else
      if (wwsmn_3_1ww1XmW_1_1lizzieLet58_4Lcall_$wnnz1_1sc_0_5_1Lcall_$wnnz0_r)
        wwsmn_3_1ww1XmW_1_1lizzieLet58_4Lcall_$wnnz1_1sc_0_5_1Lcall_$wnnz0_bufchan_d <= wwsmn_3_1ww1XmW_1_1lizzieLet58_4Lcall_$wnnz1_1sc_0_5_1Lcall_$wnnz0_d;
  CT$wnnz_t wwsmn_3_1ww1XmW_1_1lizzieLet58_4Lcall_$wnnz1_1sc_0_5_1Lcall_$wnnz0_bufchan_buf;
  assign wwsmn_3_1ww1XmW_1_1lizzieLet58_4Lcall_$wnnz1_1sc_0_5_1Lcall_$wnnz0_bufchan_r = (! wwsmn_3_1ww1XmW_1_1lizzieLet58_4Lcall_$wnnz1_1sc_0_5_1Lcall_$wnnz0_bufchan_buf[0]);
  assign lizzieLet61_1_argbuf_d = (wwsmn_3_1ww1XmW_1_1lizzieLet58_4Lcall_$wnnz1_1sc_0_5_1Lcall_$wnnz0_bufchan_buf[0] ? wwsmn_3_1ww1XmW_1_1lizzieLet58_4Lcall_$wnnz1_1sc_0_5_1Lcall_$wnnz0_bufchan_buf :
                                   wwsmn_3_1ww1XmW_1_1lizzieLet58_4Lcall_$wnnz1_1sc_0_5_1Lcall_$wnnz0_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      wwsmn_3_1ww1XmW_1_1lizzieLet58_4Lcall_$wnnz1_1sc_0_5_1Lcall_$wnnz0_bufchan_buf <= {115'd0,
                                                                                         1'd0};
    else
      if ((lizzieLet61_1_argbuf_r && wwsmn_3_1ww1XmW_1_1lizzieLet58_4Lcall_$wnnz1_1sc_0_5_1Lcall_$wnnz0_bufchan_buf[0]))
        wwsmn_3_1ww1XmW_1_1lizzieLet58_4Lcall_$wnnz1_1sc_0_5_1Lcall_$wnnz0_bufchan_buf <= {115'd0,
                                                                                           1'd0};
      else if (((! lizzieLet61_1_argbuf_r) && (! wwsmn_3_1ww1XmW_1_1lizzieLet58_4Lcall_$wnnz1_1sc_0_5_1Lcall_$wnnz0_bufchan_buf[0])))
        wwsmn_3_1ww1XmW_1_1lizzieLet58_4Lcall_$wnnz1_1sc_0_5_1Lcall_$wnnz0_bufchan_buf <= wwsmn_3_1ww1XmW_1_1lizzieLet58_4Lcall_$wnnz1_1sc_0_5_1Lcall_$wnnz0_bufchan_d;
  
  /* dcon (Ty CT$wnnz,Dcon Lcall_$wnnz0) : [(wwsmn_3_destruct,Int#),
                                       (ww1XmW_1_destruct,Int#),
                                       (lizzieLet58_4Lcall_$wnnz1,Int#),
                                       (sc_0_5_destruct,Pointer_CT$wnnz)] > (wwsmn_3_1ww1XmW_1_1lizzieLet58_4Lcall_$wnnz1_1sc_0_5_1Lcall_$wnnz0,CT$wnnz) */
  assign wwsmn_3_1ww1XmW_1_1lizzieLet58_4Lcall_$wnnz1_1sc_0_5_1Lcall_$wnnz0_d = Lcall_$wnnz0_dc((& {wwsmn_3_destruct_d[0],
                                                                                                    ww1XmW_1_destruct_d[0],
                                                                                                    lizzieLet58_4Lcall_$wnnz1_d[0],
                                                                                                    sc_0_5_destruct_d[0]}), wwsmn_3_destruct_d, ww1XmW_1_destruct_d, lizzieLet58_4Lcall_$wnnz1_d, sc_0_5_destruct_d);
  assign {wwsmn_3_destruct_r,
          ww1XmW_1_destruct_r,
          lizzieLet58_4Lcall_$wnnz1_r,
          sc_0_5_destruct_r} = {4 {(wwsmn_3_1ww1XmW_1_1lizzieLet58_4Lcall_$wnnz1_1sc_0_5_1Lcall_$wnnz0_r && wwsmn_3_1ww1XmW_1_1lizzieLet58_4Lcall_$wnnz1_1sc_0_5_1Lcall_$wnnz0_d[0])}};
  
  /* op_add (Ty Int#) : (wwsmn_4_1ww1XmW_2_1_Add32,Int#) (ww2XmZ_1_destruct,Int#) > (es_6_2_1ww2XmZ_1_1_Add32,Int#) */
  assign es_6_2_1ww2XmZ_1_1_Add32_d = {(wwsmn_4_1ww1XmW_2_1_Add32_d[32:1] + ww2XmZ_1_destruct_d[32:1]),
                                       (wwsmn_4_1ww1XmW_2_1_Add32_d[0] && ww2XmZ_1_destruct_d[0])};
  assign {wwsmn_4_1ww1XmW_2_1_Add32_r,
          ww2XmZ_1_destruct_r} = {2 {(es_6_2_1ww2XmZ_1_1_Add32_r && es_6_2_1ww2XmZ_1_1_Add32_d[0])}};
  
  /* op_add (Ty Int#) : (wwsmn_4_destruct,Int#) (ww1XmW_2_destruct,Int#) > (wwsmn_4_1ww1XmW_2_1_Add32,Int#) */
  assign wwsmn_4_1ww1XmW_2_1_Add32_d = {(wwsmn_4_destruct_d[32:1] + ww1XmW_2_destruct_d[32:1]),
                                        (wwsmn_4_destruct_d[0] && ww1XmW_2_destruct_d[0])};
  assign {wwsmn_4_destruct_r,
          ww1XmW_2_destruct_r} = {2 {(wwsmn_4_1ww1XmW_2_1_Add32_r && wwsmn_4_1ww1XmW_2_1_Add32_d[0])}};
endmodule