`timescale 1ns/1ns
import mAddAdd_package::*;

module mAddAdd(
  input logic clk,
  input logic reset,
  input Go_t \\QTree_Bool_src_d ,
  output logic \\QTree_Bool_src_r ,
  input QTree_Bool_t dummy_write_QTree_Bool_d,
  output logic dummy_write_QTree_Bool_r,
  input Go_t sourceGo_d,
  output logic sourceGo_r,
  input Pointer_QTree_Bool_t m1a81_0_d,
  output logic m1a81_0_r,
  input Pointer_QTree_Bool_t m2a82_1_d,
  output logic m2a82_1_r,
  input Pointer_QTree_Bool_t m3a83_2_d,
  output logic m3a83_2_r,
  output \Word16#_t  forkHP1_QTree_Bool_snk_dout,
  input logic forkHP1_QTree_Bool_snk_rout,
  output Pointer_QTree_Bool_t dummy_write_QTree_Bool_sink_dout,
  input logic dummy_write_QTree_Bool_sink_rout,
  output Pointer_QTree_Bool_t f_resbuf_dout,
  input logic f_resbuf_rout
  );
  /* --define=INPUTS=((__05CQTree_Bool_src, 0, 1, Go), (dummy_write_QTree_Bool, 66, 73786976294838206464, QTree_Bool), (sourceGo, 0, 1, Go), (m1a81_0, 16, 65536, Pointer_QTree_Bool), (m2a82_1, 16, 65536, Pointer_QTree_Bool), (m3a83_2, 16, 65536, Pointer_QTree_Bool)) */
  /* --define=TAPS=() */
  /* --define=OUTPUTS=((forkHP1_QTree_Bool_snk, 16, 65536, Word16__023), (dummy_write_QTree_Bool_sink, 16, 65536, Pointer_QTree_Bool), (f_resbuf, 16, 65536, Pointer_QTree_Bool)) */
  /* TYPE_START
QTree_Bool 16 2 (0,[0]) (1,[1]) (2,[16p,16p,16p,16p]) (3,[0])
CTf 16 3 (0,[0]) (1,[16p,16p,16p,16p,16p,16p,16p,16p,16p,16p]) (2,[16p,16p,16p,16p,16p,16p,16p,16p]) (3,[16p,16p,16p,16p,16p,16p]) (4,[16p,16p,16p,16p])
CTf__027__027__027__027__027__027__027__027__027__027__027__027 16 3 (0,[0]) (1,[16p,16p,16p,16p,16p,16p,16p]) (2,[16p,16p,16p,16p,16p,16p]) (3,[16p,16p,16p,16p,16p]) (4,[16p,16p,16p,16p])
TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf__027__027__027__027__027__027__027__027__027__027__027__027 16 0 (0,[0,16p,16p,16p])
TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf 16 0 (0,[0,16p,16p,16p,16p])
TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool 16 0 (0,[0,16p,16p])
TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool 16 0 (0,[0,16p,16p,16p])
TYPE_END */
  /*  */
  /*  */
  Go_t goFork_d;
  logic goFork_r;
  Go_t goFor_2_d;
  logic goFor_2_r;
  Go_t goFor_3_d;
  logic goFor_3_r;
  Go_t goFor_4_d;
  logic goFor_4_r;
  Go_t goFor_5_d;
  logic goFor_5_r;
  \Word16#_t  initHP_QTree_Bool_d;
  logic initHP_QTree_Bool_r;
  \Word16#_t  incrHP_QTree_Bool_d;
  logic incrHP_QTree_Bool_r;
  Go_t incrHP_mergeQTree_Bool_d;
  logic incrHP_mergeQTree_Bool_r;
  Go_t incrHP_QTree_Bool1_d;
  logic incrHP_QTree_Bool1_r;
  Go_t incrHP_QTree_Bool2_d;
  logic incrHP_QTree_Bool2_r;
  \Word16#_t  addHP_QTree_Bool_d;
  logic addHP_QTree_Bool_r;
  \Word16#_t  mergeHP_QTree_Bool_d;
  logic mergeHP_QTree_Bool_r;
  Go_t incrHP_mergeQTree_Bool_buf_d;
  logic incrHP_mergeQTree_Bool_buf_r;
  \Word16#_t  mergeHP_QTree_Bool_buf_d;
  logic mergeHP_QTree_Bool_buf_r;
  Go_t go_1_dummy_write_QTree_Bool_d;
  logic go_1_dummy_write_QTree_Bool_r;
  Go_t go_2_dummy_write_QTree_Bool_d;
  logic go_2_dummy_write_QTree_Bool_r;
  \Word16#_t  forkHP1_QTree_Bool_d;
  logic forkHP1_QTree_Bool_r;
  \Word16#_t  forkHP1_QTree_Bool_snk_d;
  logic forkHP1_QTree_Bool_snk_r;
  \Word16#_t  forkHP1_QTree_Boo3_d;
  logic forkHP1_QTree_Boo3_r;
  \Word16#_t  forkHP1_QTree_Boo4_d;
  logic forkHP1_QTree_Boo4_r;
  C2_t memMergeChoice_QTree_Bool_d;
  logic memMergeChoice_QTree_Bool_r;
  MemIn_QTree_Bool_t memMergeIn_QTree_Bool_d;
  logic memMergeIn_QTree_Bool_r;
  MemOut_QTree_Bool_t memOut_QTree_Bool_d;
  logic memOut_QTree_Bool_r;
  MemOut_QTree_Bool_t memReadOut_QTree_Bool_d;
  logic memReadOut_QTree_Bool_r;
  MemOut_QTree_Bool_t memWriteOut_QTree_Bool_d;
  logic memWriteOut_QTree_Bool_r;
  MemIn_QTree_Bool_t memMergeIn_QTree_Bool_dbuf_d;
  logic memMergeIn_QTree_Bool_dbuf_r;
  MemIn_QTree_Bool_t memMergeIn_QTree_Bool_rbuf_d;
  logic memMergeIn_QTree_Bool_rbuf_r;
  MemOut_QTree_Bool_t memOut_QTree_Bool_dbuf_d;
  logic memOut_QTree_Bool_dbuf_r;
  MemOut_QTree_Bool_t memOut_QTree_Bool_rbuf_d;
  logic memOut_QTree_Bool_rbuf_r;
  C5_t readMerge_choice_QTree_Bool_d;
  logic readMerge_choice_QTree_Bool_r;
  Pointer_QTree_Bool_t readMerge_data_QTree_Bool_d;
  logic readMerge_data_QTree_Bool_r;
  QTree_Bool_t readPointer_QTree_Boolm1a84_1_argbuf_d;
  logic readPointer_QTree_Boolm1a84_1_argbuf_r;
  QTree_Bool_t readPointer_QTree_Boolm2a85_1_argbuf_d;
  logic readPointer_QTree_Boolm2a85_1_argbuf_r;
  QTree_Bool_t readPointer_QTree_Boolm3a86_1_argbuf_d;
  logic readPointer_QTree_Boolm3a86_1_argbuf_r;
  QTree_Bool_t readPointer_QTree_Boolq4a90_1_argbuf_d;
  logic readPointer_QTree_Boolq4a90_1_argbuf_r;
  QTree_Bool_t readPointer_QTree_Boolt4a91_1_argbuf_d;
  logic readPointer_QTree_Boolt4a91_1_argbuf_r;
  \Word16#_t  destructReadIn_QTree_Bool_d;
  logic destructReadIn_QTree_Bool_r;
  MemIn_QTree_Bool_t dconReadIn_QTree_Bool_d;
  logic dconReadIn_QTree_Bool_r;
  QTree_Bool_t destructReadOut_QTree_Bool_d;
  logic destructReadOut_QTree_Bool_r;
  C35_t writeMerge_choice_QTree_Bool_d;
  logic writeMerge_choice_QTree_Bool_r;
  QTree_Bool_t writeMerge_data_QTree_Bool_d;
  logic writeMerge_data_QTree_Bool_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet10_1_1_argbuf_d;
  logic writeQTree_BoollizzieLet10_1_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet11_1_1_argbuf_d;
  logic writeQTree_BoollizzieLet11_1_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet12_1_1_argbuf_d;
  logic writeQTree_BoollizzieLet12_1_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet15_1_1_argbuf_d;
  logic writeQTree_BoollizzieLet15_1_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet18_1_argbuf_d;
  logic writeQTree_BoollizzieLet18_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet19_1_argbuf_d;
  logic writeQTree_BoollizzieLet19_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet23_1_argbuf_d;
  logic writeQTree_BoollizzieLet23_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet24_1_argbuf_d;
  logic writeQTree_BoollizzieLet24_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet28_1_argbuf_d;
  logic writeQTree_BoollizzieLet28_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet29_1_argbuf_d;
  logic writeQTree_BoollizzieLet29_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet30_1_argbuf_d;
  logic writeQTree_BoollizzieLet30_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet31_1_argbuf_d;
  logic writeQTree_BoollizzieLet31_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet34_1_argbuf_d;
  logic writeQTree_BoollizzieLet34_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet35_1_argbuf_d;
  logic writeQTree_BoollizzieLet35_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet36_1_argbuf_d;
  logic writeQTree_BoollizzieLet36_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet37_1_argbuf_d;
  logic writeQTree_BoollizzieLet37_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet39_1_argbuf_d;
  logic writeQTree_BoollizzieLet39_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet3_1_argbuf_d;
  logic writeQTree_BoollizzieLet3_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet40_1_argbuf_d;
  logic writeQTree_BoollizzieLet40_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet42_1_argbuf_d;
  logic writeQTree_BoollizzieLet42_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet43_1_argbuf_d;
  logic writeQTree_BoollizzieLet43_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet44_1_argbuf_d;
  logic writeQTree_BoollizzieLet44_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet47_1_argbuf_d;
  logic writeQTree_BoollizzieLet47_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet50_1_argbuf_d;
  logic writeQTree_BoollizzieLet50_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet51_1_argbuf_d;
  logic writeQTree_BoollizzieLet51_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet53_1_argbuf_d;
  logic writeQTree_BoollizzieLet53_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet55_1_argbuf_d;
  logic writeQTree_BoollizzieLet55_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet56_1_argbuf_d;
  logic writeQTree_BoollizzieLet56_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet59_1_argbuf_d;
  logic writeQTree_BoollizzieLet59_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet64_1_argbuf_d;
  logic writeQTree_BoollizzieLet64_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet69_1_argbuf_d;
  logic writeQTree_BoollizzieLet69_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet6_1_argbuf_d;
  logic writeQTree_BoollizzieLet6_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet7_1_argbuf_d;
  logic writeQTree_BoollizzieLet7_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet9_1_1_argbuf_d;
  logic writeQTree_BoollizzieLet9_1_1_argbuf_r;
  Pointer_QTree_Bool_t dummy_write_QTree_Bool_sink_d;
  logic dummy_write_QTree_Bool_sink_r;
  MemIn_QTree_Bool_t dconWriteIn_QTree_Bool_d;
  logic dconWriteIn_QTree_Bool_r;
  Pointer_QTree_Bool_t dconPtr_QTree_Bool_d;
  logic dconPtr_QTree_Bool_r;
  Pointer_QTree_Bool_t _171_d;
  logic _171_r;
  assign _171_r = 1'd1;
  Pointer_QTree_Bool_t demuxWriteResult_QTree_Bool_d;
  logic demuxWriteResult_QTree_Bool_r;
  \Word16#_t  initHP_CTf_d;
  logic initHP_CTf_r;
  \Word16#_t  incrHP_CTf_d;
  logic incrHP_CTf_r;
  Go_t incrHP_mergeCTf_d;
  logic incrHP_mergeCTf_r;
  Go_t incrHP_CTf1_d;
  logic incrHP_CTf1_r;
  Go_t incrHP_CTf2_d;
  logic incrHP_CTf2_r;
  \Word16#_t  addHP_CTf_d;
  logic addHP_CTf_r;
  \Word16#_t  mergeHP_CTf_d;
  logic mergeHP_CTf_r;
  Go_t incrHP_mergeCTf_buf_d;
  logic incrHP_mergeCTf_buf_r;
  \Word16#_t  mergeHP_CTf_buf_d;
  logic mergeHP_CTf_buf_r;
  \Word16#_t  forkHP1_CTf_d;
  logic forkHP1_CTf_r;
  \Word16#_t  forkHP1_CT2_d;
  logic forkHP1_CT2_r;
  \Word16#_t  forkHP1_CT3_d;
  logic forkHP1_CT3_r;
  C2_t memMergeChoice_CTf_d;
  logic memMergeChoice_CTf_r;
  MemIn_CTf_t memMergeIn_CTf_d;
  logic memMergeIn_CTf_r;
  MemOut_CTf_t memOut_CTf_d;
  logic memOut_CTf_r;
  MemOut_CTf_t memReadOut_CTf_d;
  logic memReadOut_CTf_r;
  MemOut_CTf_t memWriteOut_CTf_d;
  logic memWriteOut_CTf_r;
  MemIn_CTf_t memMergeIn_CTf_dbuf_d;
  logic memMergeIn_CTf_dbuf_r;
  MemIn_CTf_t memMergeIn_CTf_rbuf_d;
  logic memMergeIn_CTf_rbuf_r;
  MemOut_CTf_t memOut_CTf_dbuf_d;
  logic memOut_CTf_dbuf_r;
  MemOut_CTf_t memOut_CTf_rbuf_d;
  logic memOut_CTf_rbuf_r;
  \Word16#_t  destructReadIn_CTf_d;
  logic destructReadIn_CTf_r;
  MemIn_CTf_t dconReadIn_CTf_d;
  logic dconReadIn_CTf_r;
  CTf_t readPointer_CTfscfarg_0_1_argbuf_d;
  logic readPointer_CTfscfarg_0_1_argbuf_r;
  C5_t writeMerge_choice_CTf_d;
  logic writeMerge_choice_CTf_r;
  CTf_t writeMerge_data_CTf_d;
  logic writeMerge_data_CTf_r;
  Pointer_CTf_t writeCTflizzieLet41_1_argbuf_d;
  logic writeCTflizzieLet41_1_argbuf_r;
  Pointer_CTf_t writeCTflizzieLet57_1_argbuf_d;
  logic writeCTflizzieLet57_1_argbuf_r;
  Pointer_CTf_t writeCTflizzieLet61_1_argbuf_d;
  logic writeCTflizzieLet61_1_argbuf_r;
  Pointer_CTf_t writeCTflizzieLet62_1_argbuf_d;
  logic writeCTflizzieLet62_1_argbuf_r;
  Pointer_CTf_t writeCTflizzieLet63_1_argbuf_d;
  logic writeCTflizzieLet63_1_argbuf_r;
  MemIn_CTf_t dconWriteIn_CTf_d;
  logic dconWriteIn_CTf_r;
  Pointer_CTf_t dconPtr_CTf_d;
  logic dconPtr_CTf_r;
  Pointer_CTf_t _170_d;
  logic _170_r;
  assign _170_r = 1'd1;
  Pointer_CTf_t demuxWriteResult_CTf_d;
  logic demuxWriteResult_CTf_r;
  \Word16#_t  \initHP_CTf''''''''''''_d ;
  logic \initHP_CTf''''''''''''_r ;
  \Word16#_t  \incrHP_CTf''''''''''''_d ;
  logic \incrHP_CTf''''''''''''_r ;
  Go_t \incrHP_mergeCTf''''''''''''_d ;
  logic \incrHP_mergeCTf''''''''''''_r ;
  Go_t \incrHP_CTf''''''''''''1_d ;
  logic \incrHP_CTf''''''''''''1_r ;
  Go_t \incrHP_CTf''''''''''''2_d ;
  logic \incrHP_CTf''''''''''''2_r ;
  \Word16#_t  \addHP_CTf''''''''''''_d ;
  logic \addHP_CTf''''''''''''_r ;
  \Word16#_t  \mergeHP_CTf''''''''''''_d ;
  logic \mergeHP_CTf''''''''''''_r ;
  Go_t \incrHP_mergeCTf''''''''''''_buf_d ;
  logic \incrHP_mergeCTf''''''''''''_buf_r ;
  \Word16#_t  \mergeHP_CTf''''''''''''_buf_d ;
  logic \mergeHP_CTf''''''''''''_buf_r ;
  \Word16#_t  \forkHP1_CTf''''''''''''_d ;
  logic \forkHP1_CTf''''''''''''_r ;
  \Word16#_t  \forkHP1_CTf'''''''''''2_d ;
  logic \forkHP1_CTf'''''''''''2_r ;
  \Word16#_t  \forkHP1_CTf'''''''''''3_d ;
  logic \forkHP1_CTf'''''''''''3_r ;
  C2_t \memMergeChoice_CTf''''''''''''_d ;
  logic \memMergeChoice_CTf''''''''''''_r ;
  \MemIn_CTf''''''''''''_t  \memMergeIn_CTf''''''''''''_d ;
  logic \memMergeIn_CTf''''''''''''_r ;
  \MemOut_CTf''''''''''''_t  \memOut_CTf''''''''''''_d ;
  logic \memOut_CTf''''''''''''_r ;
  \MemOut_CTf''''''''''''_t  \memReadOut_CTf''''''''''''_d ;
  logic \memReadOut_CTf''''''''''''_r ;
  \MemOut_CTf''''''''''''_t  \memWriteOut_CTf''''''''''''_d ;
  logic \memWriteOut_CTf''''''''''''_r ;
  \MemIn_CTf''''''''''''_t  \memMergeIn_CTf''''''''''''_dbuf_d ;
  logic \memMergeIn_CTf''''''''''''_dbuf_r ;
  \MemIn_CTf''''''''''''_t  \memMergeIn_CTf''''''''''''_rbuf_d ;
  logic \memMergeIn_CTf''''''''''''_rbuf_r ;
  \MemOut_CTf''''''''''''_t  \memOut_CTf''''''''''''_dbuf_d ;
  logic \memOut_CTf''''''''''''_dbuf_r ;
  \MemOut_CTf''''''''''''_t  \memOut_CTf''''''''''''_rbuf_d ;
  logic \memOut_CTf''''''''''''_rbuf_r ;
  \Word16#_t  \destructReadIn_CTf''''''''''''_d ;
  logic \destructReadIn_CTf''''''''''''_r ;
  \MemIn_CTf''''''''''''_t  \dconReadIn_CTf''''''''''''_d ;
  logic \dconReadIn_CTf''''''''''''_r ;
  \CTf''''''''''''_t  \readPointer_CTf''''''''''''scfarg_0_1_1_argbuf_d ;
  logic \readPointer_CTf''''''''''''scfarg_0_1_1_argbuf_r ;
  C5_t \writeMerge_choice_CTf''''''''''''_d ;
  logic \writeMerge_choice_CTf''''''''''''_r ;
  \CTf''''''''''''_t  \writeMerge_data_CTf''''''''''''_d ;
  logic \writeMerge_data_CTf''''''''''''_r ;
  \Pointer_CTf''''''''''''_t  \writeCTf''''''''''''lizzieLet54_1_argbuf_d ;
  logic \writeCTf''''''''''''lizzieLet54_1_argbuf_r ;
  \Pointer_CTf''''''''''''_t  \writeCTf''''''''''''lizzieLet58_1_argbuf_d ;
  logic \writeCTf''''''''''''lizzieLet58_1_argbuf_r ;
  \Pointer_CTf''''''''''''_t  \writeCTf''''''''''''lizzieLet66_1_argbuf_d ;
  logic \writeCTf''''''''''''lizzieLet66_1_argbuf_r ;
  \Pointer_CTf''''''''''''_t  \writeCTf''''''''''''lizzieLet67_1_argbuf_d ;
  logic \writeCTf''''''''''''lizzieLet67_1_argbuf_r ;
  \Pointer_CTf''''''''''''_t  \writeCTf''''''''''''lizzieLet68_1_argbuf_d ;
  logic \writeCTf''''''''''''lizzieLet68_1_argbuf_r ;
  \MemIn_CTf''''''''''''_t  \dconWriteIn_CTf''''''''''''_d ;
  logic \dconWriteIn_CTf''''''''''''_r ;
  \Pointer_CTf''''''''''''_t  \dconPtr_CTf''''''''''''_d ;
  logic \dconPtr_CTf''''''''''''_r ;
  \Pointer_CTf''''''''''''_t  _169_d;
  logic _169_r;
  assign _169_r = 1'd1;
  \Pointer_CTf''''''''''''_t  \demuxWriteResult_CTf''''''''''''_d ;
  logic \demuxWriteResult_CTf''''''''''''_r ;
  Go_t go_1_argbuf_d;
  logic go_1_argbuf_r;
  Go_t \call_f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf''''''''''''go_3_d ;
  logic \call_f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf''''''''''''go_3_r ;
  Pointer_QTree_Bool_t \call_f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf''''''''''''q4a90_d ;
  logic \call_f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf''''''''''''q4a90_r ;
  Pointer_QTree_Bool_t \call_f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf''''''''''''t4a91_d ;
  logic \call_f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf''''''''''''t4a91_r ;
  \Pointer_CTf''''''''''''_t  \call_f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf''''''''''''sc_0_1_d ;
  logic \call_f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf''''''''''''sc_0_1_r ;
  Go_t \call_f''''''''''''_initBufi_d ;
  logic \call_f''''''''''''_initBufi_r ;
  C5_t go_3_goMux_choice_d;
  logic go_3_goMux_choice_r;
  Go_t go_3_goMux_data_d;
  logic go_3_goMux_data_r;
  Go_t \call_f''''''''''''_unlockFork1_d ;
  logic \call_f''''''''''''_unlockFork1_r ;
  Go_t \call_f''''''''''''_unlockFork2_d ;
  logic \call_f''''''''''''_unlockFork2_r ;
  Go_t \call_f''''''''''''_unlockFork3_d ;
  logic \call_f''''''''''''_unlockFork3_r ;
  Go_t \call_f''''''''''''_unlockFork4_d ;
  logic \call_f''''''''''''_unlockFork4_r ;
  Go_t \call_f''''''''''''_initBuf_d ;
  logic \call_f''''''''''''_initBuf_r ;
  Go_t \call_f''''''''''''_goMux1_d ;
  logic \call_f''''''''''''_goMux1_r ;
  Pointer_QTree_Bool_t \call_f''''''''''''_goMux2_d ;
  logic \call_f''''''''''''_goMux2_r ;
  Pointer_QTree_Bool_t \call_f''''''''''''_goMux3_d ;
  logic \call_f''''''''''''_goMux3_r ;
  \Pointer_CTf''''''''''''_t  \call_f''''''''''''_goMux4_d ;
  logic \call_f''''''''''''_goMux4_r ;
  Go_t call_fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfgo_2_d;
  logic call_fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfgo_2_r;
  Pointer_QTree_Bool_t call_fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfm1a84_d;
  logic call_fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfm1a84_r;
  Pointer_QTree_Bool_t call_fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfm2a85_d;
  logic call_fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfm2a85_r;
  Pointer_QTree_Bool_t call_fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfm3a86_d;
  logic call_fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfm3a86_r;
  Pointer_CTf_t call_fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfsc_0_d;
  logic call_fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfsc_0_r;
  Go_t call_f_initBufi_d;
  logic call_f_initBufi_r;
  C5_t go_2_goMux_choice_d;
  logic go_2_goMux_choice_r;
  Go_t go_2_goMux_data_d;
  logic go_2_goMux_data_r;
  Go_t call_f_unlockFork1_d;
  logic call_f_unlockFork1_r;
  Go_t call_f_unlockFork2_d;
  logic call_f_unlockFork2_r;
  Go_t call_f_unlockFork3_d;
  logic call_f_unlockFork3_r;
  Go_t call_f_unlockFork4_d;
  logic call_f_unlockFork4_r;
  Go_t call_f_unlockFork5_d;
  logic call_f_unlockFork5_r;
  Go_t call_f_initBuf_d;
  logic call_f_initBuf_r;
  Go_t call_f_goMux1_d;
  logic call_f_goMux1_r;
  Pointer_QTree_Bool_t call_f_goMux2_d;
  logic call_f_goMux2_r;
  Pointer_QTree_Bool_t call_f_goMux3_d;
  logic call_f_goMux3_r;
  Pointer_QTree_Bool_t call_f_goMux4_d;
  logic call_f_goMux4_r;
  Pointer_CTf_t call_f_goMux5_d;
  logic call_f_goMux5_r;
  QTree_Bool_t lizzieLet10_1_1_argbuf_d;
  logic lizzieLet10_1_1_argbuf_r;
  QTree_Bool_t lizzieLet35_1_argbuf_d;
  logic lizzieLet35_1_argbuf_r;
  QTree_Bool_t lizzieLet39_1_argbuf_d;
  logic lizzieLet39_1_argbuf_r;
  C12_t \f''''''''''''_choice_d ;
  logic \f''''''''''''_choice_r ;
  TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_t \f''''''''''''_data_d ;
  logic \f''''''''''''_data_r ;
  Go_t go_5_1_d;
  logic go_5_1_r;
  Go_t go_5_2_d;
  logic go_5_2_r;
  Pointer_QTree_Bool_t q4a90_1_1_argbuf_d;
  logic q4a90_1_1_argbuf_r;
  Pointer_QTree_Bool_t t4a91_1_1_argbuf_d;
  logic t4a91_1_1_argbuf_r;
  Pointer_QTree_Bool_t \f''''''''''''_resbuf_d ;
  logic \f''''''''''''_resbuf_r ;
  Pointer_QTree_Bool_t \f''''''''''''_10_argbuf_d ;
  logic \f''''''''''''_10_argbuf_r ;
  Pointer_QTree_Bool_t \f''''''''''''_11_argbuf_d ;
  logic \f''''''''''''_11_argbuf_r ;
  Pointer_QTree_Bool_t \f''''''''''''_12_argbuf_d ;
  logic \f''''''''''''_12_argbuf_r ;
  QTree_Bool_t es_8_1es_9_1es_10_1es_11_1QNode_Bool_d;
  logic es_8_1es_9_1es_10_1es_11_1QNode_Bool_r;
  Pointer_QTree_Bool_t \f''''''''''''_2_argbuf_d ;
  logic \f''''''''''''_2_argbuf_r ;
  Pointer_QTree_Bool_t \f''''''''''''_3_argbuf_d ;
  logic \f''''''''''''_3_argbuf_r ;
  Pointer_QTree_Bool_t \f''''''''''''_4_argbuf_d ;
  logic \f''''''''''''_4_argbuf_r ;
  QTree_Bool_t es_0_1es_1_1es_2_1es_3_1QNode_Bool_d;
  logic es_0_1es_1_1es_2_1es_3_1QNode_Bool_r;
  Pointer_QTree_Bool_t \f''''''''''''_5_argbuf_d ;
  logic \f''''''''''''_5_argbuf_r ;
  Pointer_QTree_Bool_t \f''''''''''''_6_argbuf_d ;
  logic \f''''''''''''_6_argbuf_r ;
  Pointer_QTree_Bool_t \f''''''''''''_7_argbuf_d ;
  logic \f''''''''''''_7_argbuf_r ;
  Pointer_QTree_Bool_t \f''''''''''''_8_argbuf_d ;
  logic \f''''''''''''_8_argbuf_r ;
  QTree_Bool_t es_4_1es_5_1es_6_1es_7_1QNode_Bool_d;
  logic es_4_1es_5_1es_6_1es_7_1QNode_Bool_r;
  Pointer_QTree_Bool_t \f''''''''''''_9_argbuf_d ;
  logic \f''''''''''''_9_argbuf_r ;
  Pointer_QTree_Bool_t \f''''''''''''_1_d ;
  logic \f''''''''''''_1_r ;
  Pointer_QTree_Bool_t \f''''''''''''_2_d ;
  logic \f''''''''''''_2_r ;
  Pointer_QTree_Bool_t \f''''''''''''_3_d ;
  logic \f''''''''''''_3_r ;
  Pointer_QTree_Bool_t \f''''''''''''_4_d ;
  logic \f''''''''''''_4_r ;
  Pointer_QTree_Bool_t \f''''''''''''_5_d ;
  logic \f''''''''''''_5_r ;
  Pointer_QTree_Bool_t \f''''''''''''_6_d ;
  logic \f''''''''''''_6_r ;
  Pointer_QTree_Bool_t \f''''''''''''_7_d ;
  logic \f''''''''''''_7_r ;
  Pointer_QTree_Bool_t \f''''''''''''_8_d ;
  logic \f''''''''''''_8_r ;
  Pointer_QTree_Bool_t \f''''''''''''_9_d ;
  logic \f''''''''''''_9_r ;
  Pointer_QTree_Bool_t \f''''''''''''_10_d ;
  logic \f''''''''''''_10_r ;
  Pointer_QTree_Bool_t \f''''''''''''_11_d ;
  logic \f''''''''''''_11_r ;
  Pointer_QTree_Bool_t \f''''''''''''_12_d ;
  logic \f''''''''''''_12_r ;
  Go_t \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolgo_5_d ;
  logic \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolgo_5_r ;
  Pointer_QTree_Bool_t \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolq4a90_1_d ;
  logic \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolq4a90_1_r ;
  Pointer_QTree_Bool_t \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolt4a91_1_d ;
  logic \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolt4a91_1_r ;
  Go_t fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgo_4_d;
  logic fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgo_4_r;
  Pointer_QTree_Bool_t fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm1a84_1_d;
  logic fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm1a84_1_r;
  Pointer_QTree_Bool_t fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm2a85_1_d;
  logic fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm2a85_1_r;
  Pointer_QTree_Bool_t fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm3a86_1_d;
  logic fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm3a86_1_r;
  Go_t go_4_1_d;
  logic go_4_1_r;
  Go_t go_4_2_d;
  logic go_4_2_r;
  Pointer_QTree_Bool_t m1a84_1_1_argbuf_d;
  logic m1a84_1_1_argbuf_r;
  Pointer_QTree_Bool_t m2a85_1_1_argbuf_d;
  logic m2a85_1_1_argbuf_r;
  Pointer_QTree_Bool_t m3a86_1_1_argbuf_d;
  logic m3a86_1_1_argbuf_r;
  TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_t fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1_d;
  logic fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1_r;
  C5_t go_2_goMux_choice_1_d;
  logic go_2_goMux_choice_1_r;
  C5_t go_2_goMux_choice_2_d;
  logic go_2_goMux_choice_2_r;
  C5_t go_2_goMux_choice_3_d;
  logic go_2_goMux_choice_3_r;
  C5_t go_2_goMux_choice_4_d;
  logic go_2_goMux_choice_4_r;
  Pointer_QTree_Bool_t m1a84_goMux_mux_d;
  logic m1a84_goMux_mux_r;
  Pointer_QTree_Bool_t m2a85_goMux_mux_d;
  logic m2a85_goMux_mux_r;
  Pointer_QTree_Bool_t m3a86_goMux_mux_d;
  logic m3a86_goMux_mux_r;
  Pointer_CTf_t sc_0_goMux_mux_d;
  logic sc_0_goMux_mux_r;
  C5_t go_3_goMux_choice_1_d;
  logic go_3_goMux_choice_1_r;
  C5_t go_3_goMux_choice_2_d;
  logic go_3_goMux_choice_2_r;
  C5_t go_3_goMux_choice_3_d;
  logic go_3_goMux_choice_3_r;
  Pointer_QTree_Bool_t q4a90_goMux_mux_d;
  logic q4a90_goMux_mux_r;
  Pointer_QTree_Bool_t t4a91_goMux_mux_d;
  logic t4a91_goMux_mux_r;
  \Pointer_CTf''''''''''''_t  sc_0_1_goMux_mux_d;
  logic sc_0_1_goMux_mux_r;
  CTf_t go_4_1Lfsbos_d;
  logic go_4_1Lfsbos_r;
  CTf_t lizzieLet57_1_argbuf_d;
  logic lizzieLet57_1_argbuf_r;
  Go_t go_4_2_argbuf_d;
  logic go_4_2_argbuf_r;
  TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf_t call_fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf_1_d;
  logic call_fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf_1_r;
  \CTf''''''''''''_t  \go_5_1Lf''''''''''''sbos_d ;
  logic \go_5_1Lf''''''''''''sbos_r ;
  \CTf''''''''''''_t  lizzieLet58_1_argbuf_d;
  logic lizzieLet58_1_argbuf_r;
  Go_t go_5_2_argbuf_d;
  logic go_5_2_argbuf_r;
  \TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf''''''''''''_t  \call_f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf''''''''''''_1_d ;
  logic \call_f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf''''''''''''_1_r ;
  QTree_Bool_t lizzieLet0_1_1QVal_Bool_d;
  logic lizzieLet0_1_1QVal_Bool_r;
  C40_t go_7_goMux_choice_1_d;
  logic go_7_goMux_choice_1_r;
  C40_t go_7_goMux_choice_2_d;
  logic go_7_goMux_choice_2_r;
  Pointer_QTree_Bool_t srtarg_0_goMux_mux_d;
  logic srtarg_0_goMux_mux_r;
  Pointer_CTf_t scfarg_0_goMux_mux_d;
  logic scfarg_0_goMux_mux_r;
  C12_t go_8_goMux_choice_1_d;
  logic go_8_goMux_choice_1_r;
  C12_t go_8_goMux_choice_2_d;
  logic go_8_goMux_choice_2_r;
  Pointer_QTree_Bool_t srtarg_0_1_goMux_mux_d;
  logic srtarg_0_1_goMux_mux_r;
  \Pointer_CTf''''''''''''_t  scfarg_0_1_goMux_mux_d;
  logic scfarg_0_1_goMux_mux_r;
  Pointer_QTree_Bool_t q1a8H_destruct_d;
  logic q1a8H_destruct_r;
  Pointer_QTree_Bool_t q2a8I_destruct_d;
  logic q2a8I_destruct_r;
  Pointer_QTree_Bool_t q3a8J_destruct_d;
  logic q3a8J_destruct_r;
  Pointer_QTree_Bool_t q4a8K_destruct_d;
  logic q4a8K_destruct_r;
  MyBool_t v1a8m_destruct_d;
  logic v1a8m_destruct_r;
  QTree_Bool_t lizzieLet59_1_argbuf_d;
  logic lizzieLet59_1_argbuf_r;
  QTree_Bool_t _168_d;
  logic _168_r;
  assign _168_r = 1'd1;
  QTree_Bool_t lizzieLet0_1QVal_Bool_d;
  logic lizzieLet0_1QVal_Bool_r;
  QTree_Bool_t lizzieLet0_1QNode_Bool_d;
  logic lizzieLet0_1QNode_Bool_r;
  QTree_Bool_t _167_d;
  logic _167_r;
  assign _167_r = 1'd1;
  Go_t lizzieLet0_3QNone_Bool_d;
  logic lizzieLet0_3QNone_Bool_r;
  Go_t lizzieLet0_3QVal_Bool_d;
  logic lizzieLet0_3QVal_Bool_r;
  Go_t lizzieLet0_3QNode_Bool_d;
  logic lizzieLet0_3QNode_Bool_r;
  Go_t lizzieLet0_3QError_Bool_d;
  logic lizzieLet0_3QError_Bool_r;
  Go_t lizzieLet0_3QError_Bool_1_d;
  logic lizzieLet0_3QError_Bool_1_r;
  Go_t lizzieLet0_3QError_Bool_2_d;
  logic lizzieLet0_3QError_Bool_2_r;
  QTree_Bool_t lizzieLet0_3QError_Bool_1QError_Bool_d;
  logic lizzieLet0_3QError_Bool_1QError_Bool_r;
  QTree_Bool_t lizzieLet44_1_argbuf_d;
  logic lizzieLet44_1_argbuf_r;
  Go_t lizzieLet0_3QError_Bool_2_argbuf_d;
  logic lizzieLet0_3QError_Bool_2_argbuf_r;
  QTree_Bool_t lizzieLet0_4QNone_Bool_d;
  logic lizzieLet0_4QNone_Bool_r;
  QTree_Bool_t lizzieLet0_4QVal_Bool_d;
  logic lizzieLet0_4QVal_Bool_r;
  QTree_Bool_t lizzieLet0_4QNode_Bool_d;
  logic lizzieLet0_4QNode_Bool_r;
  QTree_Bool_t _166_d;
  logic _166_r;
  assign _166_r = 1'd1;
  QTree_Bool_t lizzieLet0_4QNode_Bool_1_d;
  logic lizzieLet0_4QNode_Bool_1_r;
  QTree_Bool_t lizzieLet0_4QNode_Bool_2_d;
  logic lizzieLet0_4QNode_Bool_2_r;
  QTree_Bool_t lizzieLet0_4QNode_Bool_3_d;
  logic lizzieLet0_4QNode_Bool_3_r;
  QTree_Bool_t lizzieLet0_4QNode_Bool_4_d;
  logic lizzieLet0_4QNode_Bool_4_r;
  QTree_Bool_t lizzieLet0_4QNode_Bool_5_d;
  logic lizzieLet0_4QNode_Bool_5_r;
  QTree_Bool_t lizzieLet0_4QNode_Bool_6_d;
  logic lizzieLet0_4QNode_Bool_6_r;
  QTree_Bool_t lizzieLet0_4QNode_Bool_7_d;
  logic lizzieLet0_4QNode_Bool_7_r;
  QTree_Bool_t lizzieLet0_4QNode_Bool_8_d;
  logic lizzieLet0_4QNode_Bool_8_r;
  QTree_Bool_t lizzieLet0_4QNode_Bool_9_d;
  logic lizzieLet0_4QNode_Bool_9_r;
  QTree_Bool_t lizzieLet0_4QNode_Bool_10_d;
  logic lizzieLet0_4QNode_Bool_10_r;
  Pointer_QTree_Bool_t lizzieLet0_4QNode_Bool_10QNone_Bool_d;
  logic lizzieLet0_4QNode_Bool_10QNone_Bool_r;
  Pointer_QTree_Bool_t _165_d;
  logic _165_r;
  assign _165_r = 1'd1;
  Pointer_QTree_Bool_t lizzieLet0_4QNode_Bool_10QNode_Bool_d;
  logic lizzieLet0_4QNode_Bool_10QNode_Bool_r;
  Pointer_QTree_Bool_t _164_d;
  logic _164_r;
  assign _164_r = 1'd1;
  Pointer_QTree_Bool_t t1a8R_destruct_d;
  logic t1a8R_destruct_r;
  Pointer_QTree_Bool_t t2a8S_destruct_d;
  logic t2a8S_destruct_r;
  Pointer_QTree_Bool_t t3a8T_destruct_d;
  logic t3a8T_destruct_r;
  Pointer_QTree_Bool_t t4a8U_destruct_d;
  logic t4a8U_destruct_r;
  QTree_Bool_t _163_d;
  logic _163_r;
  assign _163_r = 1'd1;
  QTree_Bool_t _162_d;
  logic _162_r;
  assign _162_r = 1'd1;
  QTree_Bool_t lizzieLet0_4QNode_Bool_1QNode_Bool_d;
  logic lizzieLet0_4QNode_Bool_1QNode_Bool_r;
  QTree_Bool_t _161_d;
  logic _161_r;
  assign _161_r = 1'd1;
  Go_t lizzieLet0_4QNode_Bool_3QNone_Bool_d;
  logic lizzieLet0_4QNode_Bool_3QNone_Bool_r;
  Go_t lizzieLet0_4QNode_Bool_3QVal_Bool_d;
  logic lizzieLet0_4QNode_Bool_3QVal_Bool_r;
  Go_t lizzieLet0_4QNode_Bool_3QNode_Bool_d;
  logic lizzieLet0_4QNode_Bool_3QNode_Bool_r;
  Go_t lizzieLet0_4QNode_Bool_3QError_Bool_d;
  logic lizzieLet0_4QNode_Bool_3QError_Bool_r;
  Go_t lizzieLet0_4QNode_Bool_3QError_Bool_1_d;
  logic lizzieLet0_4QNode_Bool_3QError_Bool_1_r;
  Go_t lizzieLet0_4QNode_Bool_3QError_Bool_2_d;
  logic lizzieLet0_4QNode_Bool_3QError_Bool_2_r;
  QTree_Bool_t lizzieLet0_4QNode_Bool_3QError_Bool_1QError_Bool_d;
  logic lizzieLet0_4QNode_Bool_3QError_Bool_1QError_Bool_r;
  QTree_Bool_t lizzieLet43_1_argbuf_d;
  logic lizzieLet43_1_argbuf_r;
  Go_t lizzieLet0_4QNode_Bool_3QError_Bool_2_argbuf_d;
  logic lizzieLet0_4QNode_Bool_3QError_Bool_2_argbuf_r;
  Go_t lizzieLet0_4QNode_Bool_3QVal_Bool_1_d;
  logic lizzieLet0_4QNode_Bool_3QVal_Bool_1_r;
  Go_t lizzieLet0_4QNode_Bool_3QVal_Bool_2_d;
  logic lizzieLet0_4QNode_Bool_3QVal_Bool_2_r;
  QTree_Bool_t lizzieLet0_4QNode_Bool_3QVal_Bool_1QError_Bool_d;
  logic lizzieLet0_4QNode_Bool_3QVal_Bool_1QError_Bool_r;
  QTree_Bool_t lizzieLet37_1_argbuf_d;
  logic lizzieLet37_1_argbuf_r;
  Go_t lizzieLet0_4QNode_Bool_3QVal_Bool_2_argbuf_d;
  logic lizzieLet0_4QNode_Bool_3QVal_Bool_2_argbuf_r;
  QTree_Bool_t lizzieLet0_4QNode_Bool_4QNone_Bool_d;
  logic lizzieLet0_4QNode_Bool_4QNone_Bool_r;
  QTree_Bool_t _160_d;
  logic _160_r;
  assign _160_r = 1'd1;
  QTree_Bool_t lizzieLet0_4QNode_Bool_4QNode_Bool_d;
  logic lizzieLet0_4QNode_Bool_4QNode_Bool_r;
  QTree_Bool_t _159_d;
  logic _159_r;
  assign _159_r = 1'd1;
  QTree_Bool_t lizzieLet0_4QNode_Bool_4QNode_Bool_1_d;
  logic lizzieLet0_4QNode_Bool_4QNode_Bool_1_r;
  QTree_Bool_t lizzieLet0_4QNode_Bool_4QNode_Bool_2_d;
  logic lizzieLet0_4QNode_Bool_4QNode_Bool_2_r;
  QTree_Bool_t lizzieLet0_4QNode_Bool_4QNode_Bool_3_d;
  logic lizzieLet0_4QNode_Bool_4QNode_Bool_3_r;
  QTree_Bool_t lizzieLet0_4QNode_Bool_4QNode_Bool_4_d;
  logic lizzieLet0_4QNode_Bool_4QNode_Bool_4_r;
  QTree_Bool_t lizzieLet0_4QNode_Bool_4QNode_Bool_5_d;
  logic lizzieLet0_4QNode_Bool_4QNode_Bool_5_r;
  QTree_Bool_t lizzieLet0_4QNode_Bool_4QNode_Bool_6_d;
  logic lizzieLet0_4QNode_Bool_4QNode_Bool_6_r;
  QTree_Bool_t lizzieLet0_4QNode_Bool_4QNode_Bool_7_d;
  logic lizzieLet0_4QNode_Bool_4QNode_Bool_7_r;
  QTree_Bool_t lizzieLet0_4QNode_Bool_4QNode_Bool_8_d;
  logic lizzieLet0_4QNode_Bool_4QNode_Bool_8_r;
  QTree_Bool_t lizzieLet0_4QNode_Bool_4QNode_Bool_9_d;
  logic lizzieLet0_4QNode_Bool_4QNode_Bool_9_r;
  QTree_Bool_t lizzieLet0_4QNode_Bool_4QNode_Bool_10_d;
  logic lizzieLet0_4QNode_Bool_4QNode_Bool_10_r;
  QTree_Bool_t lizzieLet0_4QNode_Bool_4QNode_Bool_11_d;
  logic lizzieLet0_4QNode_Bool_4QNode_Bool_11_r;
  QTree_Bool_t lizzieLet0_4QNode_Bool_4QNode_Bool_12_d;
  logic lizzieLet0_4QNode_Bool_4QNode_Bool_12_r;
  Pointer_QTree_Bool_t lizzieLet0_4QNode_Bool_4QNode_Bool_10QNone_Bool_d;
  logic lizzieLet0_4QNode_Bool_4QNode_Bool_10QNone_Bool_r;
  Pointer_QTree_Bool_t _158_d;
  logic _158_r;
  assign _158_r = 1'd1;
  Pointer_QTree_Bool_t lizzieLet0_4QNode_Bool_4QNode_Bool_10QNode_Bool_d;
  logic lizzieLet0_4QNode_Bool_4QNode_Bool_10QNode_Bool_r;
  Pointer_QTree_Bool_t _157_d;
  logic _157_r;
  assign _157_r = 1'd1;
  Pointer_QTree_Bool_t lizzieLet0_4QNode_Bool_4QNode_Bool_10QNone_Bool_1_argbuf_d;
  logic lizzieLet0_4QNode_Bool_4QNode_Bool_10QNone_Bool_1_argbuf_r;
  Pointer_QTree_Bool_t lizzieLet0_4QNode_Bool_4QNode_Bool_11QNone_Bool_d;
  logic lizzieLet0_4QNode_Bool_4QNode_Bool_11QNone_Bool_r;
  Pointer_QTree_Bool_t _156_d;
  logic _156_r;
  assign _156_r = 1'd1;
  Pointer_QTree_Bool_t lizzieLet0_4QNode_Bool_4QNode_Bool_11QNode_Bool_d;
  logic lizzieLet0_4QNode_Bool_4QNode_Bool_11QNode_Bool_r;
  Pointer_QTree_Bool_t _155_d;
  logic _155_r;
  assign _155_r = 1'd1;
  Pointer_QTree_Bool_t lizzieLet0_4QNode_Bool_4QNode_Bool_11QNone_Bool_1_argbuf_d;
  logic lizzieLet0_4QNode_Bool_4QNode_Bool_11QNone_Bool_1_argbuf_r;
  Pointer_QTree_Bool_t lizzieLet0_4QNode_Bool_4QNode_Bool_12QNone_Bool_d;
  logic lizzieLet0_4QNode_Bool_4QNode_Bool_12QNone_Bool_r;
  Pointer_QTree_Bool_t _154_d;
  logic _154_r;
  assign _154_r = 1'd1;
  Pointer_QTree_Bool_t lizzieLet0_4QNode_Bool_4QNode_Bool_12QNode_Bool_d;
  logic lizzieLet0_4QNode_Bool_4QNode_Bool_12QNode_Bool_r;
  Pointer_QTree_Bool_t _153_d;
  logic _153_r;
  assign _153_r = 1'd1;
  Pointer_QTree_Bool_t lizzieLet0_4QNode_Bool_4QNode_Bool_12QNode_Bool_1_argbuf_d;
  logic lizzieLet0_4QNode_Bool_4QNode_Bool_12QNode_Bool_1_argbuf_r;
  Pointer_QTree_Bool_t lizzieLet0_4QNode_Bool_4QNode_Bool_12QNone_Bool_1_argbuf_d;
  logic lizzieLet0_4QNode_Bool_4QNode_Bool_12QNone_Bool_1_argbuf_r;
  Pointer_QTree_Bool_t \t1'a8W_destruct_d ;
  logic \t1'a8W_destruct_r ;
  Pointer_QTree_Bool_t \t2'a8X_destruct_d ;
  logic \t2'a8X_destruct_r ;
  Pointer_QTree_Bool_t \t3'a8Y_destruct_d ;
  logic \t3'a8Y_destruct_r ;
  Pointer_QTree_Bool_t \t4'a8Z_destruct_d ;
  logic \t4'a8Z_destruct_r ;
  QTree_Bool_t _152_d;
  logic _152_r;
  assign _152_r = 1'd1;
  QTree_Bool_t _151_d;
  logic _151_r;
  assign _151_r = 1'd1;
  QTree_Bool_t lizzieLet0_4QNode_Bool_4QNode_Bool_1QNode_Bool_d;
  logic lizzieLet0_4QNode_Bool_4QNode_Bool_1QNode_Bool_r;
  QTree_Bool_t _150_d;
  logic _150_r;
  assign _150_r = 1'd1;
  Pointer_QTree_Bool_t lizzieLet0_4QNode_Bool_4QNode_Bool_3QNone_Bool_d;
  logic lizzieLet0_4QNode_Bool_4QNode_Bool_3QNone_Bool_r;
  Pointer_QTree_Bool_t _149_d;
  logic _149_r;
  assign _149_r = 1'd1;
  Pointer_QTree_Bool_t lizzieLet0_4QNode_Bool_4QNode_Bool_3QNode_Bool_d;
  logic lizzieLet0_4QNode_Bool_4QNode_Bool_3QNode_Bool_r;
  Pointer_QTree_Bool_t _148_d;
  logic _148_r;
  assign _148_r = 1'd1;
  Pointer_QTree_Bool_t lizzieLet0_4QNode_Bool_4QNode_Bool_3QNode_Bool_1_argbuf_d;
  logic lizzieLet0_4QNode_Bool_4QNode_Bool_3QNode_Bool_1_argbuf_r;
  Pointer_QTree_Bool_t lizzieLet0_4QNode_Bool_4QNode_Bool_3QNone_Bool_1_argbuf_d;
  logic lizzieLet0_4QNode_Bool_4QNode_Bool_3QNone_Bool_1_argbuf_r;
  Go_t lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_d;
  logic lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_r;
  Go_t lizzieLet0_4QNode_Bool_4QNode_Bool_4QVal_Bool_d;
  logic lizzieLet0_4QNode_Bool_4QNode_Bool_4QVal_Bool_r;
  Go_t lizzieLet0_4QNode_Bool_4QNode_Bool_4QNode_Bool_d;
  logic lizzieLet0_4QNode_Bool_4QNode_Bool_4QNode_Bool_r;
  Go_t lizzieLet0_4QNode_Bool_4QNode_Bool_4QError_Bool_d;
  logic lizzieLet0_4QNode_Bool_4QNode_Bool_4QError_Bool_r;
  Go_t lizzieLet0_4QNode_Bool_4QNode_Bool_4QError_Bool_1_d;
  logic lizzieLet0_4QNode_Bool_4QNode_Bool_4QError_Bool_1_r;
  Go_t lizzieLet0_4QNode_Bool_4QNode_Bool_4QError_Bool_2_d;
  logic lizzieLet0_4QNode_Bool_4QNode_Bool_4QError_Bool_2_r;
  QTree_Bool_t lizzieLet0_4QNode_Bool_4QNode_Bool_4QError_Bool_1QError_Bool_d;
  logic lizzieLet0_4QNode_Bool_4QNode_Bool_4QError_Bool_1QError_Bool_r;
  QTree_Bool_t lizzieLet42_1_argbuf_d;
  logic lizzieLet42_1_argbuf_r;
  Go_t lizzieLet0_4QNode_Bool_4QNode_Bool_4QError_Bool_2_argbuf_d;
  logic lizzieLet0_4QNode_Bool_4QNode_Bool_4QError_Bool_2_argbuf_r;
  Go_t lizzieLet0_4QNode_Bool_4QNode_Bool_4QNode_Bool_1_argbuf_d;
  logic lizzieLet0_4QNode_Bool_4QNode_Bool_4QNode_Bool_1_argbuf_r;
  Go_t lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_1_d;
  logic lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_1_r;
  Go_t lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_2_d;
  logic lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_2_r;
  Go_t lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_3_d;
  logic lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_3_r;
  Go_t lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_4_d;
  logic lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_4_r;
  Go_t lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_5_d;
  logic lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_5_r;
  Go_t lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_1_argbuf_d;
  logic lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_1_argbuf_r;
  TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_t \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool9_d ;
  logic \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool9_r ;
  Go_t lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_2_argbuf_d;
  logic lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_2_argbuf_r;
  TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_t \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool10_d ;
  logic \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool10_r ;
  Go_t lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_3_argbuf_d;
  logic lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_3_argbuf_r;
  TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_t \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool11_d ;
  logic \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool11_r ;
  Go_t lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_4_argbuf_d;
  logic lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_4_argbuf_r;
  TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_t \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool12_d ;
  logic \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool12_r ;
  Go_t lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_5_argbuf_d;
  logic lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_5_argbuf_r;
  Go_t lizzieLet0_4QNode_Bool_4QNode_Bool_4QVal_Bool_1_d;
  logic lizzieLet0_4QNode_Bool_4QNode_Bool_4QVal_Bool_1_r;
  Go_t lizzieLet0_4QNode_Bool_4QNode_Bool_4QVal_Bool_2_d;
  logic lizzieLet0_4QNode_Bool_4QNode_Bool_4QVal_Bool_2_r;
  QTree_Bool_t lizzieLet0_4QNode_Bool_4QNode_Bool_4QVal_Bool_1QError_Bool_d;
  logic lizzieLet0_4QNode_Bool_4QNode_Bool_4QVal_Bool_1QError_Bool_r;
  QTree_Bool_t lizzieLet40_1_argbuf_d;
  logic lizzieLet40_1_argbuf_r;
  Go_t lizzieLet0_4QNode_Bool_4QNode_Bool_4QVal_Bool_2_argbuf_d;
  logic lizzieLet0_4QNode_Bool_4QNode_Bool_4QVal_Bool_2_argbuf_r;
  Pointer_CTf_t lizzieLet0_4QNode_Bool_4QNode_Bool_5QNone_Bool_d;
  logic lizzieLet0_4QNode_Bool_4QNode_Bool_5QNone_Bool_r;
  Pointer_CTf_t lizzieLet0_4QNode_Bool_4QNode_Bool_5QVal_Bool_d;
  logic lizzieLet0_4QNode_Bool_4QNode_Bool_5QVal_Bool_r;
  Pointer_CTf_t lizzieLet0_4QNode_Bool_4QNode_Bool_5QNode_Bool_d;
  logic lizzieLet0_4QNode_Bool_4QNode_Bool_5QNode_Bool_r;
  Pointer_CTf_t lizzieLet0_4QNode_Bool_4QNode_Bool_5QError_Bool_d;
  logic lizzieLet0_4QNode_Bool_4QNode_Bool_5QError_Bool_r;
  Pointer_CTf_t lizzieLet0_4QNode_Bool_4QNode_Bool_5QError_Bool_1_argbuf_d;
  logic lizzieLet0_4QNode_Bool_4QNode_Bool_5QError_Bool_1_argbuf_r;
  CTf_t \lizzieLet0_4QNode_Bool_4QNode_Bool_5QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_6QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_9QNode_Bool_1t1'a8W_1lizzieLet0_4QNode_Bool_4QNode_Bool_7QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_10QNode_Bool_1t2'a8X_1lizzieLet0_4QNode_Bool_4QNode_Bool_8QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_11QNode_Bool_1t3'a8Y_1Lcall_f3_d ;
  logic \lizzieLet0_4QNode_Bool_4QNode_Bool_5QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_6QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_9QNode_Bool_1t1'a8W_1lizzieLet0_4QNode_Bool_4QNode_Bool_7QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_10QNode_Bool_1t2'a8X_1lizzieLet0_4QNode_Bool_4QNode_Bool_8QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_11QNode_Bool_1t3'a8Y_1Lcall_f3_r ;
  CTf_t lizzieLet41_1_argbuf_d;
  logic lizzieLet41_1_argbuf_r;
  Pointer_CTf_t lizzieLet0_4QNode_Bool_4QNode_Bool_5QNone_Bool_1_argbuf_d;
  logic lizzieLet0_4QNode_Bool_4QNode_Bool_5QNone_Bool_1_argbuf_r;
  Pointer_CTf_t lizzieLet0_4QNode_Bool_4QNode_Bool_5QVal_Bool_1_argbuf_d;
  logic lizzieLet0_4QNode_Bool_4QNode_Bool_5QVal_Bool_1_argbuf_r;
  Pointer_QTree_Bool_t lizzieLet0_4QNode_Bool_4QNode_Bool_6QNone_Bool_d;
  logic lizzieLet0_4QNode_Bool_4QNode_Bool_6QNone_Bool_r;
  Pointer_QTree_Bool_t _147_d;
  logic _147_r;
  assign _147_r = 1'd1;
  Pointer_QTree_Bool_t lizzieLet0_4QNode_Bool_4QNode_Bool_6QNode_Bool_d;
  logic lizzieLet0_4QNode_Bool_4QNode_Bool_6QNode_Bool_r;
  Pointer_QTree_Bool_t _146_d;
  logic _146_r;
  assign _146_r = 1'd1;
  Pointer_QTree_Bool_t lizzieLet0_4QNode_Bool_4QNode_Bool_6QNone_Bool_1_argbuf_d;
  logic lizzieLet0_4QNode_Bool_4QNode_Bool_6QNone_Bool_1_argbuf_r;
  Pointer_QTree_Bool_t lizzieLet0_4QNode_Bool_4QNode_Bool_7QNone_Bool_d;
  logic lizzieLet0_4QNode_Bool_4QNode_Bool_7QNone_Bool_r;
  Pointer_QTree_Bool_t _145_d;
  logic _145_r;
  assign _145_r = 1'd1;
  Pointer_QTree_Bool_t lizzieLet0_4QNode_Bool_4QNode_Bool_7QNode_Bool_d;
  logic lizzieLet0_4QNode_Bool_4QNode_Bool_7QNode_Bool_r;
  Pointer_QTree_Bool_t _144_d;
  logic _144_r;
  assign _144_r = 1'd1;
  Pointer_QTree_Bool_t lizzieLet0_4QNode_Bool_4QNode_Bool_7QNone_Bool_1_argbuf_d;
  logic lizzieLet0_4QNode_Bool_4QNode_Bool_7QNone_Bool_1_argbuf_r;
  Pointer_QTree_Bool_t lizzieLet0_4QNode_Bool_4QNode_Bool_8QNone_Bool_d;
  logic lizzieLet0_4QNode_Bool_4QNode_Bool_8QNone_Bool_r;
  Pointer_QTree_Bool_t _143_d;
  logic _143_r;
  assign _143_r = 1'd1;
  Pointer_QTree_Bool_t lizzieLet0_4QNode_Bool_4QNode_Bool_8QNode_Bool_d;
  logic lizzieLet0_4QNode_Bool_4QNode_Bool_8QNode_Bool_r;
  Pointer_QTree_Bool_t _142_d;
  logic _142_r;
  assign _142_r = 1'd1;
  Pointer_QTree_Bool_t lizzieLet0_4QNode_Bool_4QNode_Bool_8QNone_Bool_1_argbuf_d;
  logic lizzieLet0_4QNode_Bool_4QNode_Bool_8QNone_Bool_1_argbuf_r;
  Pointer_QTree_Bool_t lizzieLet0_4QNode_Bool_4QNode_Bool_9QNone_Bool_d;
  logic lizzieLet0_4QNode_Bool_4QNode_Bool_9QNone_Bool_r;
  Pointer_QTree_Bool_t _141_d;
  logic _141_r;
  assign _141_r = 1'd1;
  Pointer_QTree_Bool_t lizzieLet0_4QNode_Bool_4QNode_Bool_9QNode_Bool_d;
  logic lizzieLet0_4QNode_Bool_4QNode_Bool_9QNode_Bool_r;
  Pointer_QTree_Bool_t _140_d;
  logic _140_r;
  assign _140_r = 1'd1;
  Pointer_QTree_Bool_t lizzieLet0_4QNode_Bool_4QNode_Bool_9QNone_Bool_1_argbuf_d;
  logic lizzieLet0_4QNode_Bool_4QNode_Bool_9QNone_Bool_1_argbuf_r;
  QTree_Bool_t lizzieLet0_4QNode_Bool_4QNone_Bool_1_d;
  logic lizzieLet0_4QNode_Bool_4QNone_Bool_1_r;
  QTree_Bool_t lizzieLet0_4QNode_Bool_4QNone_Bool_2_d;
  logic lizzieLet0_4QNode_Bool_4QNone_Bool_2_r;
  QTree_Bool_t lizzieLet0_4QNode_Bool_4QNone_Bool_3_d;
  logic lizzieLet0_4QNode_Bool_4QNone_Bool_3_r;
  QTree_Bool_t lizzieLet0_4QNode_Bool_4QNone_Bool_4_d;
  logic lizzieLet0_4QNode_Bool_4QNone_Bool_4_r;
  QTree_Bool_t lizzieLet0_4QNode_Bool_4QNone_Bool_5_d;
  logic lizzieLet0_4QNode_Bool_4QNone_Bool_5_r;
  QTree_Bool_t lizzieLet0_4QNode_Bool_4QNone_Bool_6_d;
  logic lizzieLet0_4QNode_Bool_4QNone_Bool_6_r;
  QTree_Bool_t lizzieLet0_4QNode_Bool_4QNone_Bool_7_d;
  logic lizzieLet0_4QNode_Bool_4QNone_Bool_7_r;
  QTree_Bool_t lizzieLet0_4QNode_Bool_4QNone_Bool_8_d;
  logic lizzieLet0_4QNode_Bool_4QNone_Bool_8_r;
  QTree_Bool_t lizzieLet0_4QNode_Bool_4QNone_Bool_9_d;
  logic lizzieLet0_4QNode_Bool_4QNone_Bool_9_r;
  Pointer_QTree_Bool_t t1a8M_destruct_d;
  logic t1a8M_destruct_r;
  Pointer_QTree_Bool_t t2a8N_destruct_d;
  logic t2a8N_destruct_r;
  Pointer_QTree_Bool_t t3a8O_destruct_d;
  logic t3a8O_destruct_r;
  Pointer_QTree_Bool_t t4a8P_destruct_d;
  logic t4a8P_destruct_r;
  QTree_Bool_t _139_d;
  logic _139_r;
  assign _139_r = 1'd1;
  QTree_Bool_t _138_d;
  logic _138_r;
  assign _138_r = 1'd1;
  QTree_Bool_t lizzieLet0_4QNode_Bool_4QNone_Bool_1QNode_Bool_d;
  logic lizzieLet0_4QNode_Bool_4QNone_Bool_1QNode_Bool_r;
  QTree_Bool_t _137_d;
  logic _137_r;
  assign _137_r = 1'd1;
  Pointer_QTree_Bool_t _136_d;
  logic _136_r;
  assign _136_r = 1'd1;
  Pointer_QTree_Bool_t _135_d;
  logic _135_r;
  assign _135_r = 1'd1;
  Pointer_QTree_Bool_t lizzieLet0_4QNode_Bool_4QNone_Bool_3QNode_Bool_d;
  logic lizzieLet0_4QNode_Bool_4QNone_Bool_3QNode_Bool_r;
  Pointer_QTree_Bool_t _134_d;
  logic _134_r;
  assign _134_r = 1'd1;
  Pointer_QTree_Bool_t lizzieLet0_4QNode_Bool_4QNone_Bool_3QNode_Bool_1_argbuf_d;
  logic lizzieLet0_4QNode_Bool_4QNone_Bool_3QNode_Bool_1_argbuf_r;
  Go_t lizzieLet0_4QNode_Bool_4QNone_Bool_4QNone_Bool_d;
  logic lizzieLet0_4QNode_Bool_4QNone_Bool_4QNone_Bool_r;
  Go_t lizzieLet0_4QNode_Bool_4QNone_Bool_4QVal_Bool_d;
  logic lizzieLet0_4QNode_Bool_4QNone_Bool_4QVal_Bool_r;
  Go_t lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_d;
  logic lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_r;
  Go_t lizzieLet0_4QNode_Bool_4QNone_Bool_4QError_Bool_d;
  logic lizzieLet0_4QNode_Bool_4QNone_Bool_4QError_Bool_r;
  Go_t lizzieLet0_4QNode_Bool_4QNone_Bool_4QError_Bool_1_d;
  logic lizzieLet0_4QNode_Bool_4QNone_Bool_4QError_Bool_1_r;
  Go_t lizzieLet0_4QNode_Bool_4QNone_Bool_4QError_Bool_2_d;
  logic lizzieLet0_4QNode_Bool_4QNone_Bool_4QError_Bool_2_r;
  QTree_Bool_t lizzieLet0_4QNode_Bool_4QNone_Bool_4QError_Bool_1QError_Bool_d;
  logic lizzieLet0_4QNode_Bool_4QNone_Bool_4QError_Bool_1QError_Bool_r;
  QTree_Bool_t lizzieLet36_1_argbuf_d;
  logic lizzieLet36_1_argbuf_r;
  Go_t lizzieLet0_4QNode_Bool_4QNone_Bool_4QError_Bool_2_argbuf_d;
  logic lizzieLet0_4QNode_Bool_4QNone_Bool_4QError_Bool_2_argbuf_r;
  Go_t lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_1_d;
  logic lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_1_r;
  Go_t lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_2_d;
  logic lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_2_r;
  Go_t lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_3_d;
  logic lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_3_r;
  Go_t lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_4_d;
  logic lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_4_r;
  Go_t lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_5_d;
  logic lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_5_r;
  Go_t lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_1_argbuf_d;
  logic lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_1_argbuf_r;
  TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_t \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool5_d ;
  logic \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool5_r ;
  Go_t lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_2_argbuf_d;
  logic lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_2_argbuf_r;
  TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_t \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool6_d ;
  logic \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool6_r ;
  Go_t lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_3_argbuf_d;
  logic lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_3_argbuf_r;
  TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_t \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool7_d ;
  logic \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool7_r ;
  Go_t lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_4_argbuf_d;
  logic lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_4_argbuf_r;
  TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_t \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool8_d ;
  logic \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool8_r ;
  Go_t lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_5_argbuf_d;
  logic lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_5_argbuf_r;
  Go_t lizzieLet0_4QNode_Bool_4QNone_Bool_4QNone_Bool_1_argbuf_d;
  logic lizzieLet0_4QNode_Bool_4QNone_Bool_4QNone_Bool_1_argbuf_r;
  Go_t lizzieLet0_4QNode_Bool_4QNone_Bool_4QVal_Bool_1_d;
  logic lizzieLet0_4QNode_Bool_4QNone_Bool_4QVal_Bool_1_r;
  Go_t lizzieLet0_4QNode_Bool_4QNone_Bool_4QVal_Bool_2_d;
  logic lizzieLet0_4QNode_Bool_4QNone_Bool_4QVal_Bool_2_r;
  QTree_Bool_t lizzieLet0_4QNode_Bool_4QNone_Bool_4QVal_Bool_1QError_Bool_d;
  logic lizzieLet0_4QNode_Bool_4QNone_Bool_4QVal_Bool_1QError_Bool_r;
  QTree_Bool_t lizzieLet34_1_argbuf_d;
  logic lizzieLet34_1_argbuf_r;
  Go_t lizzieLet0_4QNode_Bool_4QNone_Bool_4QVal_Bool_2_argbuf_d;
  logic lizzieLet0_4QNode_Bool_4QNone_Bool_4QVal_Bool_2_argbuf_r;
  Pointer_QTree_Bool_t lizzieLet0_4QNode_Bool_4QNone_Bool_5QNone_Bool_d;
  logic lizzieLet0_4QNode_Bool_4QNone_Bool_5QNone_Bool_r;
  Pointer_QTree_Bool_t _133_d;
  logic _133_r;
  assign _133_r = 1'd1;
  Pointer_QTree_Bool_t _132_d;
  logic _132_r;
  assign _132_r = 1'd1;
  Pointer_QTree_Bool_t _131_d;
  logic _131_r;
  assign _131_r = 1'd1;
  Pointer_QTree_Bool_t lizzieLet0_4QNode_Bool_4QNone_Bool_5QNone_Bool_1_argbuf_d;
  logic lizzieLet0_4QNode_Bool_4QNone_Bool_5QNone_Bool_1_argbuf_r;
  Pointer_CTf_t lizzieLet0_4QNode_Bool_4QNone_Bool_6QNone_Bool_d;
  logic lizzieLet0_4QNode_Bool_4QNone_Bool_6QNone_Bool_r;
  Pointer_CTf_t lizzieLet0_4QNode_Bool_4QNone_Bool_6QVal_Bool_d;
  logic lizzieLet0_4QNode_Bool_4QNone_Bool_6QVal_Bool_r;
  Pointer_CTf_t lizzieLet0_4QNode_Bool_4QNone_Bool_6QNode_Bool_d;
  logic lizzieLet0_4QNode_Bool_4QNone_Bool_6QNode_Bool_r;
  Pointer_CTf_t lizzieLet0_4QNode_Bool_4QNone_Bool_6QError_Bool_d;
  logic lizzieLet0_4QNode_Bool_4QNone_Bool_6QError_Bool_r;
  Pointer_CTf_t lizzieLet0_4QNode_Bool_4QNone_Bool_6QError_Bool_1_argbuf_d;
  logic lizzieLet0_4QNode_Bool_4QNone_Bool_6QError_Bool_1_argbuf_r;
  Pointer_CTf_t lizzieLet0_4QNode_Bool_4QNone_Bool_6QNode_Bool_1_argbuf_d;
  logic lizzieLet0_4QNode_Bool_4QNone_Bool_6QNode_Bool_1_argbuf_r;
  Pointer_CTf_t lizzieLet0_4QNode_Bool_4QNone_Bool_6QNone_Bool_1_argbuf_d;
  logic lizzieLet0_4QNode_Bool_4QNone_Bool_6QNone_Bool_1_argbuf_r;
  Pointer_CTf_t lizzieLet0_4QNode_Bool_4QNone_Bool_6QVal_Bool_1_argbuf_d;
  logic lizzieLet0_4QNode_Bool_4QNone_Bool_6QVal_Bool_1_argbuf_r;
  Pointer_QTree_Bool_t _130_d;
  logic _130_r;
  assign _130_r = 1'd1;
  Pointer_QTree_Bool_t _129_d;
  logic _129_r;
  assign _129_r = 1'd1;
  Pointer_QTree_Bool_t lizzieLet0_4QNode_Bool_4QNone_Bool_7QNode_Bool_d;
  logic lizzieLet0_4QNode_Bool_4QNone_Bool_7QNode_Bool_r;
  Pointer_QTree_Bool_t _128_d;
  logic _128_r;
  assign _128_r = 1'd1;
  Pointer_QTree_Bool_t lizzieLet0_4QNode_Bool_4QNone_Bool_7QNode_Bool_1_argbuf_d;
  logic lizzieLet0_4QNode_Bool_4QNone_Bool_7QNode_Bool_1_argbuf_r;
  Pointer_QTree_Bool_t _127_d;
  logic _127_r;
  assign _127_r = 1'd1;
  Pointer_QTree_Bool_t _126_d;
  logic _126_r;
  assign _126_r = 1'd1;
  Pointer_QTree_Bool_t lizzieLet0_4QNode_Bool_4QNone_Bool_8QNode_Bool_d;
  logic lizzieLet0_4QNode_Bool_4QNone_Bool_8QNode_Bool_r;
  Pointer_QTree_Bool_t _125_d;
  logic _125_r;
  assign _125_r = 1'd1;
  Pointer_QTree_Bool_t lizzieLet0_4QNode_Bool_4QNone_Bool_8QNode_Bool_1_argbuf_d;
  logic lizzieLet0_4QNode_Bool_4QNone_Bool_8QNode_Bool_1_argbuf_r;
  Pointer_QTree_Bool_t _124_d;
  logic _124_r;
  assign _124_r = 1'd1;
  Pointer_QTree_Bool_t _123_d;
  logic _123_r;
  assign _123_r = 1'd1;
  Pointer_QTree_Bool_t lizzieLet0_4QNode_Bool_4QNone_Bool_9QNode_Bool_d;
  logic lizzieLet0_4QNode_Bool_4QNone_Bool_9QNode_Bool_r;
  Pointer_QTree_Bool_t _122_d;
  logic _122_r;
  assign _122_r = 1'd1;
  Pointer_QTree_Bool_t lizzieLet0_4QNode_Bool_4QNone_Bool_9QNode_Bool_1_argbuf_d;
  logic lizzieLet0_4QNode_Bool_4QNone_Bool_9QNode_Bool_1_argbuf_r;
  Pointer_QTree_Bool_t lizzieLet0_4QNode_Bool_5QNone_Bool_d;
  logic lizzieLet0_4QNode_Bool_5QNone_Bool_r;
  Pointer_QTree_Bool_t _121_d;
  logic _121_r;
  assign _121_r = 1'd1;
  Pointer_QTree_Bool_t _120_d;
  logic _120_r;
  assign _120_r = 1'd1;
  Pointer_QTree_Bool_t _119_d;
  logic _119_r;
  assign _119_r = 1'd1;
  Pointer_CTf_t lizzieLet0_4QNode_Bool_6QNone_Bool_d;
  logic lizzieLet0_4QNode_Bool_6QNone_Bool_r;
  Pointer_CTf_t lizzieLet0_4QNode_Bool_6QVal_Bool_d;
  logic lizzieLet0_4QNode_Bool_6QVal_Bool_r;
  Pointer_CTf_t lizzieLet0_4QNode_Bool_6QNode_Bool_d;
  logic lizzieLet0_4QNode_Bool_6QNode_Bool_r;
  Pointer_CTf_t lizzieLet0_4QNode_Bool_6QError_Bool_d;
  logic lizzieLet0_4QNode_Bool_6QError_Bool_r;
  Pointer_CTf_t lizzieLet0_4QNode_Bool_6QError_Bool_1_argbuf_d;
  logic lizzieLet0_4QNode_Bool_6QError_Bool_1_argbuf_r;
  Pointer_CTf_t lizzieLet0_4QNode_Bool_6QVal_Bool_1_argbuf_d;
  logic lizzieLet0_4QNode_Bool_6QVal_Bool_1_argbuf_r;
  Pointer_QTree_Bool_t lizzieLet0_4QNode_Bool_7QNone_Bool_d;
  logic lizzieLet0_4QNode_Bool_7QNone_Bool_r;
  Pointer_QTree_Bool_t _118_d;
  logic _118_r;
  assign _118_r = 1'd1;
  Pointer_QTree_Bool_t lizzieLet0_4QNode_Bool_7QNode_Bool_d;
  logic lizzieLet0_4QNode_Bool_7QNode_Bool_r;
  Pointer_QTree_Bool_t _117_d;
  logic _117_r;
  assign _117_r = 1'd1;
  Pointer_QTree_Bool_t lizzieLet0_4QNode_Bool_8QNone_Bool_d;
  logic lizzieLet0_4QNode_Bool_8QNone_Bool_r;
  Pointer_QTree_Bool_t _116_d;
  logic _116_r;
  assign _116_r = 1'd1;
  Pointer_QTree_Bool_t lizzieLet0_4QNode_Bool_8QNode_Bool_d;
  logic lizzieLet0_4QNode_Bool_8QNode_Bool_r;
  Pointer_QTree_Bool_t _115_d;
  logic _115_r;
  assign _115_r = 1'd1;
  Pointer_QTree_Bool_t lizzieLet0_4QNode_Bool_9QNone_Bool_d;
  logic lizzieLet0_4QNode_Bool_9QNone_Bool_r;
  Pointer_QTree_Bool_t _114_d;
  logic _114_r;
  assign _114_r = 1'd1;
  Pointer_QTree_Bool_t lizzieLet0_4QNode_Bool_9QNode_Bool_d;
  logic lizzieLet0_4QNode_Bool_9QNode_Bool_r;
  Pointer_QTree_Bool_t _113_d;
  logic _113_r;
  assign _113_r = 1'd1;
  QTree_Bool_t lizzieLet0_4QNone_Bool_1_d;
  logic lizzieLet0_4QNone_Bool_1_r;
  QTree_Bool_t lizzieLet0_4QNone_Bool_2_d;
  logic lizzieLet0_4QNone_Bool_2_r;
  QTree_Bool_t lizzieLet0_4QNone_Bool_3_d;
  logic lizzieLet0_4QNone_Bool_3_r;
  QTree_Bool_t lizzieLet0_4QNone_Bool_4_d;
  logic lizzieLet0_4QNone_Bool_4_r;
  QTree_Bool_t lizzieLet0_4QNone_Bool_5_d;
  logic lizzieLet0_4QNone_Bool_5_r;
  QTree_Bool_t lizzieLet0_4QNone_Bool_6_d;
  logic lizzieLet0_4QNone_Bool_6_r;
  QTree_Bool_t lizzieLet0_4QNone_Bool_7_d;
  logic lizzieLet0_4QNone_Bool_7_r;
  Pointer_QTree_Bool_t q1a8d_destruct_d;
  logic q1a8d_destruct_r;
  Pointer_QTree_Bool_t q2a8e_destruct_d;
  logic q2a8e_destruct_r;
  Pointer_QTree_Bool_t q3a8f_destruct_d;
  logic q3a8f_destruct_r;
  Pointer_QTree_Bool_t q4a8g_destruct_d;
  logic q4a8g_destruct_r;
  MyBool_t v1a87_destruct_d;
  logic v1a87_destruct_r;
  QTree_Bool_t _112_d;
  logic _112_r;
  assign _112_r = 1'd1;
  QTree_Bool_t lizzieLet0_4QNone_Bool_1QVal_Bool_d;
  logic lizzieLet0_4QNone_Bool_1QVal_Bool_r;
  QTree_Bool_t lizzieLet0_4QNone_Bool_1QNode_Bool_d;
  logic lizzieLet0_4QNone_Bool_1QNode_Bool_r;
  QTree_Bool_t _111_d;
  logic _111_r;
  assign _111_r = 1'd1;
  Go_t lizzieLet0_4QNone_Bool_3QNone_Bool_d;
  logic lizzieLet0_4QNone_Bool_3QNone_Bool_r;
  Go_t lizzieLet0_4QNone_Bool_3QVal_Bool_d;
  logic lizzieLet0_4QNone_Bool_3QVal_Bool_r;
  Go_t lizzieLet0_4QNone_Bool_3QNode_Bool_d;
  logic lizzieLet0_4QNone_Bool_3QNode_Bool_r;
  Go_t lizzieLet0_4QNone_Bool_3QError_Bool_d;
  logic lizzieLet0_4QNone_Bool_3QError_Bool_r;
  Go_t lizzieLet0_4QNone_Bool_3QError_Bool_1_d;
  logic lizzieLet0_4QNone_Bool_3QError_Bool_1_r;
  Go_t lizzieLet0_4QNone_Bool_3QError_Bool_2_d;
  logic lizzieLet0_4QNone_Bool_3QError_Bool_2_r;
  QTree_Bool_t lizzieLet0_4QNone_Bool_3QError_Bool_1QError_Bool_d;
  logic lizzieLet0_4QNone_Bool_3QError_Bool_1QError_Bool_r;
  QTree_Bool_t lizzieLet12_1_1_argbuf_d;
  logic lizzieLet12_1_1_argbuf_r;
  Go_t lizzieLet0_4QNone_Bool_3QError_Bool_2_argbuf_d;
  logic lizzieLet0_4QNone_Bool_3QError_Bool_2_argbuf_r;
  Go_t lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_d;
  logic lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_r;
  C40_t go_7_goMux_choice_d;
  logic go_7_goMux_choice_r;
  Go_t go_7_goMux_data_d;
  logic go_7_goMux_data_r;
  QTree_Bool_t _110_d;
  logic _110_r;
  assign _110_r = 1'd1;
  QTree_Bool_t lizzieLet0_4QNone_Bool_4QVal_Bool_d;
  logic lizzieLet0_4QNone_Bool_4QVal_Bool_r;
  QTree_Bool_t lizzieLet0_4QNone_Bool_4QNode_Bool_d;
  logic lizzieLet0_4QNone_Bool_4QNode_Bool_r;
  QTree_Bool_t _109_d;
  logic _109_r;
  assign _109_r = 1'd1;
  QTree_Bool_t lizzieLet0_4QNone_Bool_4QNode_Bool_1_d;
  logic lizzieLet0_4QNone_Bool_4QNode_Bool_1_r;
  QTree_Bool_t lizzieLet0_4QNone_Bool_4QNode_Bool_2_d;
  logic lizzieLet0_4QNone_Bool_4QNode_Bool_2_r;
  QTree_Bool_t lizzieLet0_4QNone_Bool_4QNode_Bool_3_d;
  logic lizzieLet0_4QNone_Bool_4QNode_Bool_3_r;
  QTree_Bool_t lizzieLet0_4QNone_Bool_4QNode_Bool_4_d;
  logic lizzieLet0_4QNone_Bool_4QNode_Bool_4_r;
  QTree_Bool_t lizzieLet0_4QNone_Bool_4QNode_Bool_5_d;
  logic lizzieLet0_4QNone_Bool_4QNode_Bool_5_r;
  QTree_Bool_t lizzieLet0_4QNone_Bool_4QNode_Bool_6_d;
  logic lizzieLet0_4QNone_Bool_4QNode_Bool_6_r;
  QTree_Bool_t lizzieLet0_4QNone_Bool_4QNode_Bool_7_d;
  logic lizzieLet0_4QNone_Bool_4QNode_Bool_7_r;
  QTree_Bool_t lizzieLet0_4QNone_Bool_4QNode_Bool_8_d;
  logic lizzieLet0_4QNone_Bool_4QNode_Bool_8_r;
  QTree_Bool_t lizzieLet0_4QNone_Bool_4QNode_Bool_9_d;
  logic lizzieLet0_4QNone_Bool_4QNode_Bool_9_r;
  Pointer_QTree_Bool_t t1a8i_destruct_d;
  logic t1a8i_destruct_r;
  Pointer_QTree_Bool_t t2a8j_destruct_d;
  logic t2a8j_destruct_r;
  Pointer_QTree_Bool_t t3a8k_destruct_d;
  logic t3a8k_destruct_r;
  Pointer_QTree_Bool_t t4a8l_destruct_d;
  logic t4a8l_destruct_r;
  QTree_Bool_t _108_d;
  logic _108_r;
  assign _108_r = 1'd1;
  QTree_Bool_t _107_d;
  logic _107_r;
  assign _107_r = 1'd1;
  QTree_Bool_t lizzieLet0_4QNone_Bool_4QNode_Bool_1QNode_Bool_d;
  logic lizzieLet0_4QNone_Bool_4QNode_Bool_1QNode_Bool_r;
  QTree_Bool_t _106_d;
  logic _106_r;
  assign _106_r = 1'd1;
  Go_t lizzieLet0_4QNone_Bool_4QNode_Bool_3QNone_Bool_d;
  logic lizzieLet0_4QNone_Bool_4QNode_Bool_3QNone_Bool_r;
  Go_t lizzieLet0_4QNone_Bool_4QNode_Bool_3QVal_Bool_d;
  logic lizzieLet0_4QNone_Bool_4QNode_Bool_3QVal_Bool_r;
  Go_t lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_d;
  logic lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_r;
  Go_t lizzieLet0_4QNone_Bool_4QNode_Bool_3QError_Bool_d;
  logic lizzieLet0_4QNone_Bool_4QNode_Bool_3QError_Bool_r;
  Go_t lizzieLet0_4QNone_Bool_4QNode_Bool_3QError_Bool_1_d;
  logic lizzieLet0_4QNone_Bool_4QNode_Bool_3QError_Bool_1_r;
  Go_t lizzieLet0_4QNone_Bool_4QNode_Bool_3QError_Bool_2_d;
  logic lizzieLet0_4QNone_Bool_4QNode_Bool_3QError_Bool_2_r;
  QTree_Bool_t lizzieLet0_4QNone_Bool_4QNode_Bool_3QError_Bool_1QError_Bool_d;
  logic lizzieLet0_4QNone_Bool_4QNode_Bool_3QError_Bool_1QError_Bool_r;
  QTree_Bool_t lizzieLet11_1_1_argbuf_d;
  logic lizzieLet11_1_1_argbuf_r;
  Go_t lizzieLet0_4QNone_Bool_4QNode_Bool_3QError_Bool_2_argbuf_d;
  logic lizzieLet0_4QNone_Bool_4QNode_Bool_3QError_Bool_2_argbuf_r;
  Go_t lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_1_d;
  logic lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_1_r;
  Go_t lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_2_d;
  logic lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_2_r;
  Go_t lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_3_d;
  logic lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_3_r;
  Go_t lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_4_d;
  logic lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_4_r;
  Go_t lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_5_d;
  logic lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_5_r;
  Go_t lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_1_argbuf_d;
  logic lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_1_argbuf_r;
  TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_t \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_1_d ;
  logic \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_1_r ;
  Go_t lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_2_argbuf_d;
  logic lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_2_argbuf_r;
  TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_t \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool2_d ;
  logic \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool2_r ;
  Go_t lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_3_argbuf_d;
  logic lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_3_argbuf_r;
  TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_t \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool3_d ;
  logic \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool3_r ;
  Go_t lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_4_argbuf_d;
  logic lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_4_argbuf_r;
  TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_t \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool4_d ;
  logic \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool4_r ;
  Go_t lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_5_argbuf_d;
  logic lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_5_argbuf_r;
  Go_t lizzieLet0_4QNone_Bool_4QNode_Bool_3QNone_Bool_1_argbuf_d;
  logic lizzieLet0_4QNone_Bool_4QNode_Bool_3QNone_Bool_1_argbuf_r;
  Go_t lizzieLet0_4QNone_Bool_4QNode_Bool_3QVal_Bool_1_d;
  logic lizzieLet0_4QNone_Bool_4QNode_Bool_3QVal_Bool_1_r;
  Go_t lizzieLet0_4QNone_Bool_4QNode_Bool_3QVal_Bool_2_d;
  logic lizzieLet0_4QNone_Bool_4QNode_Bool_3QVal_Bool_2_r;
  QTree_Bool_t lizzieLet0_4QNone_Bool_4QNode_Bool_3QVal_Bool_1QError_Bool_d;
  logic lizzieLet0_4QNone_Bool_4QNode_Bool_3QVal_Bool_1QError_Bool_r;
  QTree_Bool_t lizzieLet9_1_1_argbuf_d;
  logic lizzieLet9_1_1_argbuf_r;
  Go_t lizzieLet0_4QNone_Bool_4QNode_Bool_3QVal_Bool_2_argbuf_d;
  logic lizzieLet0_4QNone_Bool_4QNode_Bool_3QVal_Bool_2_argbuf_r;
  Pointer_QTree_Bool_t lizzieLet0_4QNone_Bool_4QNode_Bool_4QNone_Bool_d;
  logic lizzieLet0_4QNone_Bool_4QNode_Bool_4QNone_Bool_r;
  Pointer_QTree_Bool_t _105_d;
  logic _105_r;
  assign _105_r = 1'd1;
  Pointer_QTree_Bool_t _104_d;
  logic _104_r;
  assign _104_r = 1'd1;
  Pointer_QTree_Bool_t _103_d;
  logic _103_r;
  assign _103_r = 1'd1;
  Pointer_QTree_Bool_t lizzieLet0_4QNone_Bool_4QNode_Bool_4QNone_Bool_1_argbuf_d;
  logic lizzieLet0_4QNone_Bool_4QNode_Bool_4QNone_Bool_1_argbuf_r;
  Pointer_CTf_t lizzieLet0_4QNone_Bool_4QNode_Bool_5QNone_Bool_d;
  logic lizzieLet0_4QNone_Bool_4QNode_Bool_5QNone_Bool_r;
  Pointer_CTf_t lizzieLet0_4QNone_Bool_4QNode_Bool_5QVal_Bool_d;
  logic lizzieLet0_4QNone_Bool_4QNode_Bool_5QVal_Bool_r;
  Pointer_CTf_t lizzieLet0_4QNone_Bool_4QNode_Bool_5QNode_Bool_d;
  logic lizzieLet0_4QNone_Bool_4QNode_Bool_5QNode_Bool_r;
  Pointer_CTf_t lizzieLet0_4QNone_Bool_4QNode_Bool_5QError_Bool_d;
  logic lizzieLet0_4QNone_Bool_4QNode_Bool_5QError_Bool_r;
  Pointer_CTf_t lizzieLet0_4QNone_Bool_4QNode_Bool_5QError_Bool_1_argbuf_d;
  logic lizzieLet0_4QNone_Bool_4QNode_Bool_5QError_Bool_1_argbuf_r;
  Pointer_CTf_t lizzieLet0_4QNone_Bool_4QNode_Bool_5QNode_Bool_1_argbuf_d;
  logic lizzieLet0_4QNone_Bool_4QNode_Bool_5QNode_Bool_1_argbuf_r;
  Pointer_CTf_t lizzieLet0_4QNone_Bool_4QNode_Bool_5QNone_Bool_1_argbuf_d;
  logic lizzieLet0_4QNone_Bool_4QNode_Bool_5QNone_Bool_1_argbuf_r;
  Pointer_CTf_t lizzieLet0_4QNone_Bool_4QNode_Bool_5QVal_Bool_1_argbuf_d;
  logic lizzieLet0_4QNone_Bool_4QNode_Bool_5QVal_Bool_1_argbuf_r;
  Pointer_QTree_Bool_t _102_d;
  logic _102_r;
  assign _102_r = 1'd1;
  Pointer_QTree_Bool_t _101_d;
  logic _101_r;
  assign _101_r = 1'd1;
  Pointer_QTree_Bool_t lizzieLet0_4QNone_Bool_4QNode_Bool_6QNode_Bool_d;
  logic lizzieLet0_4QNone_Bool_4QNode_Bool_6QNode_Bool_r;
  Pointer_QTree_Bool_t _100_d;
  logic _100_r;
  assign _100_r = 1'd1;
  Pointer_QTree_Bool_t lizzieLet0_4QNone_Bool_4QNode_Bool_6QNode_Bool_1_argbuf_d;
  logic lizzieLet0_4QNone_Bool_4QNode_Bool_6QNode_Bool_1_argbuf_r;
  Pointer_QTree_Bool_t _99_d;
  logic _99_r;
  assign _99_r = 1'd1;
  Pointer_QTree_Bool_t _98_d;
  logic _98_r;
  assign _98_r = 1'd1;
  Pointer_QTree_Bool_t lizzieLet0_4QNone_Bool_4QNode_Bool_7QNode_Bool_d;
  logic lizzieLet0_4QNone_Bool_4QNode_Bool_7QNode_Bool_r;
  Pointer_QTree_Bool_t _97_d;
  logic _97_r;
  assign _97_r = 1'd1;
  Pointer_QTree_Bool_t lizzieLet0_4QNone_Bool_4QNode_Bool_7QNode_Bool_1_argbuf_d;
  logic lizzieLet0_4QNone_Bool_4QNode_Bool_7QNode_Bool_1_argbuf_r;
  Pointer_QTree_Bool_t _96_d;
  logic _96_r;
  assign _96_r = 1'd1;
  Pointer_QTree_Bool_t _95_d;
  logic _95_r;
  assign _95_r = 1'd1;
  Pointer_QTree_Bool_t lizzieLet0_4QNone_Bool_4QNode_Bool_8QNode_Bool_d;
  logic lizzieLet0_4QNone_Bool_4QNode_Bool_8QNode_Bool_r;
  Pointer_QTree_Bool_t _94_d;
  logic _94_r;
  assign _94_r = 1'd1;
  Pointer_QTree_Bool_t lizzieLet0_4QNone_Bool_4QNode_Bool_8QNode_Bool_1_argbuf_d;
  logic lizzieLet0_4QNone_Bool_4QNode_Bool_8QNode_Bool_1_argbuf_r;
  Pointer_QTree_Bool_t _93_d;
  logic _93_r;
  assign _93_r = 1'd1;
  Pointer_QTree_Bool_t _92_d;
  logic _92_r;
  assign _92_r = 1'd1;
  Pointer_QTree_Bool_t lizzieLet0_4QNone_Bool_4QNode_Bool_9QNode_Bool_d;
  logic lizzieLet0_4QNone_Bool_4QNode_Bool_9QNode_Bool_r;
  Pointer_QTree_Bool_t _91_d;
  logic _91_r;
  assign _91_r = 1'd1;
  Pointer_QTree_Bool_t lizzieLet0_4QNone_Bool_4QNode_Bool_9QNode_Bool_1_argbuf_d;
  logic lizzieLet0_4QNone_Bool_4QNode_Bool_9QNode_Bool_1_argbuf_r;
  QTree_Bool_t lizzieLet0_4QNone_Bool_4QVal_Bool_1_d;
  logic lizzieLet0_4QNone_Bool_4QVal_Bool_1_r;
  QTree_Bool_t lizzieLet0_4QNone_Bool_4QVal_Bool_2_d;
  logic lizzieLet0_4QNone_Bool_4QVal_Bool_2_r;
  QTree_Bool_t lizzieLet0_4QNone_Bool_4QVal_Bool_3_d;
  logic lizzieLet0_4QNone_Bool_4QVal_Bool_3_r;
  QTree_Bool_t lizzieLet0_4QNone_Bool_4QVal_Bool_4_d;
  logic lizzieLet0_4QNone_Bool_4QVal_Bool_4_r;
  QTree_Bool_t lizzieLet0_4QNone_Bool_4QVal_Bool_5_d;
  logic lizzieLet0_4QNone_Bool_4QVal_Bool_5_r;
  QTree_Bool_t lizzieLet0_4QNone_Bool_4QVal_Bool_6_d;
  logic lizzieLet0_4QNone_Bool_4QVal_Bool_6_r;
  MyBool_t va88_destruct_d;
  logic va88_destruct_r;
  QTree_Bool_t _90_d;
  logic _90_r;
  assign _90_r = 1'd1;
  QTree_Bool_t lizzieLet0_4QNone_Bool_4QVal_Bool_1QVal_Bool_d;
  logic lizzieLet0_4QNone_Bool_4QVal_Bool_1QVal_Bool_r;
  QTree_Bool_t _89_d;
  logic _89_r;
  assign _89_r = 1'd1;
  QTree_Bool_t _88_d;
  logic _88_r;
  assign _88_r = 1'd1;
  Go_t lizzieLet0_4QNone_Bool_4QVal_Bool_3QNone_Bool_d;
  logic lizzieLet0_4QNone_Bool_4QVal_Bool_3QNone_Bool_r;
  Go_t lizzieLet0_4QNone_Bool_4QVal_Bool_3QVal_Bool_d;
  logic lizzieLet0_4QNone_Bool_4QVal_Bool_3QVal_Bool_r;
  Go_t lizzieLet0_4QNone_Bool_4QVal_Bool_3QNode_Bool_d;
  logic lizzieLet0_4QNone_Bool_4QVal_Bool_3QNode_Bool_r;
  Go_t lizzieLet0_4QNone_Bool_4QVal_Bool_3QError_Bool_d;
  logic lizzieLet0_4QNone_Bool_4QVal_Bool_3QError_Bool_r;
  Go_t lizzieLet0_4QNone_Bool_4QVal_Bool_3QError_Bool_1_d;
  logic lizzieLet0_4QNone_Bool_4QVal_Bool_3QError_Bool_1_r;
  Go_t lizzieLet0_4QNone_Bool_4QVal_Bool_3QError_Bool_2_d;
  logic lizzieLet0_4QNone_Bool_4QVal_Bool_3QError_Bool_2_r;
  QTree_Bool_t lizzieLet0_4QNone_Bool_4QVal_Bool_3QError_Bool_1QError_Bool_d;
  logic lizzieLet0_4QNone_Bool_4QVal_Bool_3QError_Bool_1QError_Bool_r;
  QTree_Bool_t lizzieLet7_1_argbuf_d;
  logic lizzieLet7_1_argbuf_r;
  Go_t lizzieLet0_4QNone_Bool_4QVal_Bool_3QError_Bool_2_argbuf_d;
  logic lizzieLet0_4QNone_Bool_4QVal_Bool_3QError_Bool_2_argbuf_r;
  Go_t lizzieLet0_4QNone_Bool_4QVal_Bool_3QNode_Bool_1_d;
  logic lizzieLet0_4QNone_Bool_4QVal_Bool_3QNode_Bool_1_r;
  Go_t lizzieLet0_4QNone_Bool_4QVal_Bool_3QNode_Bool_2_d;
  logic lizzieLet0_4QNone_Bool_4QVal_Bool_3QNode_Bool_2_r;
  QTree_Bool_t lizzieLet0_4QNone_Bool_4QVal_Bool_3QNode_Bool_1QError_Bool_d;
  logic lizzieLet0_4QNone_Bool_4QVal_Bool_3QNode_Bool_1QError_Bool_r;
  QTree_Bool_t lizzieLet6_1_argbuf_d;
  logic lizzieLet6_1_argbuf_r;
  Go_t lizzieLet0_4QNone_Bool_4QVal_Bool_3QNode_Bool_2_argbuf_d;
  logic lizzieLet0_4QNone_Bool_4QVal_Bool_3QNode_Bool_2_argbuf_r;
  Go_t lizzieLet0_4QNone_Bool_4QVal_Bool_3QNone_Bool_1_argbuf_d;
  logic lizzieLet0_4QNone_Bool_4QVal_Bool_3QNone_Bool_1_argbuf_r;
  Pointer_QTree_Bool_t lizzieLet0_4QNone_Bool_4QVal_Bool_4QNone_Bool_d;
  logic lizzieLet0_4QNone_Bool_4QVal_Bool_4QNone_Bool_r;
  Pointer_QTree_Bool_t _87_d;
  logic _87_r;
  assign _87_r = 1'd1;
  Pointer_QTree_Bool_t _86_d;
  logic _86_r;
  assign _86_r = 1'd1;
  Pointer_QTree_Bool_t _85_d;
  logic _85_r;
  assign _85_r = 1'd1;
  Pointer_QTree_Bool_t lizzieLet0_4QNone_Bool_4QVal_Bool_4QNone_Bool_1_argbuf_d;
  logic lizzieLet0_4QNone_Bool_4QVal_Bool_4QNone_Bool_1_argbuf_r;
  Pointer_CTf_t lizzieLet0_4QNone_Bool_4QVal_Bool_5QNone_Bool_d;
  logic lizzieLet0_4QNone_Bool_4QVal_Bool_5QNone_Bool_r;
  Pointer_CTf_t lizzieLet0_4QNone_Bool_4QVal_Bool_5QVal_Bool_d;
  logic lizzieLet0_4QNone_Bool_4QVal_Bool_5QVal_Bool_r;
  Pointer_CTf_t lizzieLet0_4QNone_Bool_4QVal_Bool_5QNode_Bool_d;
  logic lizzieLet0_4QNone_Bool_4QVal_Bool_5QNode_Bool_r;
  Pointer_CTf_t lizzieLet0_4QNone_Bool_4QVal_Bool_5QError_Bool_d;
  logic lizzieLet0_4QNone_Bool_4QVal_Bool_5QError_Bool_r;
  Pointer_CTf_t lizzieLet0_4QNone_Bool_4QVal_Bool_5QError_Bool_1_argbuf_d;
  logic lizzieLet0_4QNone_Bool_4QVal_Bool_5QError_Bool_1_argbuf_r;
  Pointer_CTf_t lizzieLet0_4QNone_Bool_4QVal_Bool_5QNode_Bool_1_argbuf_d;
  logic lizzieLet0_4QNone_Bool_4QVal_Bool_5QNode_Bool_1_argbuf_r;
  Pointer_CTf_t lizzieLet0_4QNone_Bool_4QVal_Bool_5QNone_Bool_1_argbuf_d;
  logic lizzieLet0_4QNone_Bool_4QVal_Bool_5QNone_Bool_1_argbuf_r;
  MyBool_t _84_d;
  logic _84_r;
  assign _84_r = 1'd1;
  MyBool_t lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_d;
  logic lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_r;
  MyBool_t _83_d;
  logic _83_r;
  assign _83_r = 1'd1;
  MyBool_t _82_d;
  logic _82_r;
  assign _82_r = 1'd1;
  MyBool_t lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1_d;
  logic lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1_r;
  MyBool_t lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_2_d;
  logic lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_2_r;
  MyBool_t lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3_d;
  logic lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3_r;
  Go_t lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyFalse_d;
  logic lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyFalse_r;
  Go_t lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyTrue_d;
  logic lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyTrue_r;
  Go_t lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyTrue_1_d;
  logic lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyTrue_1_r;
  Go_t lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyTrue_2_d;
  logic lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyTrue_2_r;
  Go_t lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyTrue_1_argbuf_d;
  logic lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyTrue_1_argbuf_r;
  TupGo_t \lvlrf2-0TupGo2_d ;
  logic \lvlrf2-0TupGo2_r ;
  Go_t lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyTrue_2_argbuf_d;
  logic lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyTrue_2_argbuf_r;
  Pointer_CTf_t lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_2MyFalse_d;
  logic lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_2MyFalse_r;
  Pointer_CTf_t lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_2MyTrue_d;
  logic lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_2MyTrue_r;
  Pointer_CTf_t lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_2MyTrue_1_argbuf_d;
  logic lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_2MyTrue_1_argbuf_r;
  MyBool_t lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_d;
  logic lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_r;
  MyBool_t _81_d;
  logic _81_r;
  assign _81_r = 1'd1;
  MyBool_t lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1_d;
  logic lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1_r;
  MyBool_t lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_2_d;
  logic lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_2_r;
  Go_t lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_d;
  logic lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_r;
  Go_t lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_d;
  logic lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_r;
  Go_t lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1_d;
  logic lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1_r;
  Go_t lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_d;
  logic lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_r;
  QTree_Bool_t lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_d;
  logic lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_r;
  QTree_Bool_t lizzieLet3_1_argbuf_d;
  logic lizzieLet3_1_argbuf_r;
  Go_t lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_argbuf_d;
  logic lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_argbuf_r;
  Go_t lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_d;
  logic lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_r;
  Go_t lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_d;
  logic lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_r;
  Go_t lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_argbuf_d;
  logic lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_argbuf_r;
  TupGo_t \lvlrf2-0TupGo_1_d ;
  logic \lvlrf2-0TupGo_1_r ;
  Go_t lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_argbuf_d;
  logic lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_argbuf_r;
  Pointer_CTf_t lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_2MyFalse_d;
  logic lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_2MyFalse_r;
  Pointer_CTf_t lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_2MyTrue_d;
  logic lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_2MyTrue_r;
  Pointer_CTf_t lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_2MyFalse_1_argbuf_d;
  logic lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_2MyFalse_1_argbuf_r;
  Pointer_CTf_t lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_2MyTrue_1_argbuf_d;
  logic lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_2MyTrue_1_argbuf_r;
  Pointer_QTree_Bool_t _80_d;
  logic _80_r;
  assign _80_r = 1'd1;
  Pointer_QTree_Bool_t lizzieLet0_4QNone_Bool_5QVal_Bool_d;
  logic lizzieLet0_4QNone_Bool_5QVal_Bool_r;
  Pointer_QTree_Bool_t lizzieLet0_4QNone_Bool_5QNode_Bool_d;
  logic lizzieLet0_4QNone_Bool_5QNode_Bool_r;
  Pointer_QTree_Bool_t _79_d;
  logic _79_r;
  assign _79_r = 1'd1;
  Pointer_QTree_Bool_t lizzieLet0_4QNone_Bool_6QNone_Bool_d;
  logic lizzieLet0_4QNone_Bool_6QNone_Bool_r;
  Pointer_QTree_Bool_t _78_d;
  logic _78_r;
  assign _78_r = 1'd1;
  Pointer_QTree_Bool_t _77_d;
  logic _77_r;
  assign _77_r = 1'd1;
  Pointer_QTree_Bool_t _76_d;
  logic _76_r;
  assign _76_r = 1'd1;
  Pointer_QTree_Bool_t lizzieLet0_4QNone_Bool_6QNone_Bool_1_argbuf_d;
  logic lizzieLet0_4QNone_Bool_6QNone_Bool_1_argbuf_r;
  Pointer_CTf_t lizzieLet0_4QNone_Bool_7QNone_Bool_d;
  logic lizzieLet0_4QNone_Bool_7QNone_Bool_r;
  Pointer_CTf_t lizzieLet0_4QNone_Bool_7QVal_Bool_d;
  logic lizzieLet0_4QNone_Bool_7QVal_Bool_r;
  Pointer_CTf_t lizzieLet0_4QNone_Bool_7QNode_Bool_d;
  logic lizzieLet0_4QNone_Bool_7QNode_Bool_r;
  Pointer_CTf_t lizzieLet0_4QNone_Bool_7QError_Bool_d;
  logic lizzieLet0_4QNone_Bool_7QError_Bool_r;
  Pointer_CTf_t lizzieLet0_4QNone_Bool_7QError_Bool_1_argbuf_d;
  logic lizzieLet0_4QNone_Bool_7QError_Bool_1_argbuf_r;
  Pointer_CTf_t lizzieLet0_4QNone_Bool_7QNone_Bool_1_argbuf_d;
  logic lizzieLet0_4QNone_Bool_7QNone_Bool_1_argbuf_r;
  QTree_Bool_t lizzieLet0_4QVal_Bool_1_d;
  logic lizzieLet0_4QVal_Bool_1_r;
  QTree_Bool_t lizzieLet0_4QVal_Bool_2_d;
  logic lizzieLet0_4QVal_Bool_2_r;
  QTree_Bool_t lizzieLet0_4QVal_Bool_3_d;
  logic lizzieLet0_4QVal_Bool_3_r;
  QTree_Bool_t lizzieLet0_4QVal_Bool_4_d;
  logic lizzieLet0_4QVal_Bool_4_r;
  QTree_Bool_t lizzieLet0_4QVal_Bool_5_d;
  logic lizzieLet0_4QVal_Bool_5_r;
  QTree_Bool_t lizzieLet0_4QVal_Bool_6_d;
  logic lizzieLet0_4QVal_Bool_6_r;
  QTree_Bool_t lizzieLet0_4QVal_Bool_7_d;
  logic lizzieLet0_4QVal_Bool_7_r;
  QTree_Bool_t lizzieLet0_4QVal_Bool_8_d;
  logic lizzieLet0_4QVal_Bool_8_r;
  MyBool_t va8s_destruct_d;
  logic va8s_destruct_r;
  QTree_Bool_t _75_d;
  logic _75_r;
  assign _75_r = 1'd1;
  QTree_Bool_t lizzieLet0_4QVal_Bool_1QVal_Bool_d;
  logic lizzieLet0_4QVal_Bool_1QVal_Bool_r;
  QTree_Bool_t _74_d;
  logic _74_r;
  assign _74_r = 1'd1;
  QTree_Bool_t _73_d;
  logic _73_r;
  assign _73_r = 1'd1;
  Go_t lizzieLet0_4QVal_Bool_3QNone_Bool_d;
  logic lizzieLet0_4QVal_Bool_3QNone_Bool_r;
  Go_t lizzieLet0_4QVal_Bool_3QVal_Bool_d;
  logic lizzieLet0_4QVal_Bool_3QVal_Bool_r;
  Go_t lizzieLet0_4QVal_Bool_3QNode_Bool_d;
  logic lizzieLet0_4QVal_Bool_3QNode_Bool_r;
  Go_t lizzieLet0_4QVal_Bool_3QError_Bool_d;
  logic lizzieLet0_4QVal_Bool_3QError_Bool_r;
  Go_t lizzieLet0_4QVal_Bool_3QError_Bool_1_d;
  logic lizzieLet0_4QVal_Bool_3QError_Bool_1_r;
  Go_t lizzieLet0_4QVal_Bool_3QError_Bool_2_d;
  logic lizzieLet0_4QVal_Bool_3QError_Bool_2_r;
  QTree_Bool_t lizzieLet0_4QVal_Bool_3QError_Bool_1QError_Bool_d;
  logic lizzieLet0_4QVal_Bool_3QError_Bool_1QError_Bool_r;
  QTree_Bool_t lizzieLet31_1_argbuf_d;
  logic lizzieLet31_1_argbuf_r;
  Go_t lizzieLet0_4QVal_Bool_3QError_Bool_2_argbuf_d;
  logic lizzieLet0_4QVal_Bool_3QError_Bool_2_argbuf_r;
  Go_t lizzieLet0_4QVal_Bool_3QNode_Bool_1_d;
  logic lizzieLet0_4QVal_Bool_3QNode_Bool_1_r;
  Go_t lizzieLet0_4QVal_Bool_3QNode_Bool_2_d;
  logic lizzieLet0_4QVal_Bool_3QNode_Bool_2_r;
  QTree_Bool_t lizzieLet0_4QVal_Bool_3QNode_Bool_1QError_Bool_d;
  logic lizzieLet0_4QVal_Bool_3QNode_Bool_1QError_Bool_r;
  QTree_Bool_t lizzieLet30_1_argbuf_d;
  logic lizzieLet30_1_argbuf_r;
  Go_t lizzieLet0_4QVal_Bool_3QNode_Bool_2_argbuf_d;
  logic lizzieLet0_4QVal_Bool_3QNode_Bool_2_argbuf_r;
  QTree_Bool_t lizzieLet0_4QVal_Bool_4QNone_Bool_d;
  logic lizzieLet0_4QVal_Bool_4QNone_Bool_r;
  QTree_Bool_t lizzieLet0_4QVal_Bool_4QVal_Bool_d;
  logic lizzieLet0_4QVal_Bool_4QVal_Bool_r;
  QTree_Bool_t _72_d;
  logic _72_r;
  assign _72_r = 1'd1;
  QTree_Bool_t _71_d;
  logic _71_r;
  assign _71_r = 1'd1;
  QTree_Bool_t lizzieLet0_4QVal_Bool_4QNone_Bool_1_d;
  logic lizzieLet0_4QVal_Bool_4QNone_Bool_1_r;
  QTree_Bool_t lizzieLet0_4QVal_Bool_4QNone_Bool_2_d;
  logic lizzieLet0_4QVal_Bool_4QNone_Bool_2_r;
  QTree_Bool_t lizzieLet0_4QVal_Bool_4QNone_Bool_3_d;
  logic lizzieLet0_4QVal_Bool_4QNone_Bool_3_r;
  QTree_Bool_t lizzieLet0_4QVal_Bool_4QNone_Bool_4_d;
  logic lizzieLet0_4QVal_Bool_4QNone_Bool_4_r;
  QTree_Bool_t lizzieLet0_4QVal_Bool_4QNone_Bool_5_d;
  logic lizzieLet0_4QVal_Bool_4QNone_Bool_5_r;
  QTree_Bool_t lizzieLet0_4QVal_Bool_4QNone_Bool_6_d;
  logic lizzieLet0_4QVal_Bool_4QNone_Bool_6_r;
  MyBool_t va8n_destruct_d;
  logic va8n_destruct_r;
  QTree_Bool_t _70_d;
  logic _70_r;
  assign _70_r = 1'd1;
  QTree_Bool_t lizzieLet0_4QVal_Bool_4QNone_Bool_1QVal_Bool_d;
  logic lizzieLet0_4QVal_Bool_4QNone_Bool_1QVal_Bool_r;
  QTree_Bool_t _69_d;
  logic _69_r;
  assign _69_r = 1'd1;
  QTree_Bool_t _68_d;
  logic _68_r;
  assign _68_r = 1'd1;
  Go_t lizzieLet0_4QVal_Bool_4QNone_Bool_3QNone_Bool_d;
  logic lizzieLet0_4QVal_Bool_4QNone_Bool_3QNone_Bool_r;
  Go_t lizzieLet0_4QVal_Bool_4QNone_Bool_3QVal_Bool_d;
  logic lizzieLet0_4QVal_Bool_4QNone_Bool_3QVal_Bool_r;
  Go_t lizzieLet0_4QVal_Bool_4QNone_Bool_3QNode_Bool_d;
  logic lizzieLet0_4QVal_Bool_4QNone_Bool_3QNode_Bool_r;
  Go_t lizzieLet0_4QVal_Bool_4QNone_Bool_3QError_Bool_d;
  logic lizzieLet0_4QVal_Bool_4QNone_Bool_3QError_Bool_r;
  Go_t lizzieLet0_4QVal_Bool_4QNone_Bool_3QError_Bool_1_d;
  logic lizzieLet0_4QVal_Bool_4QNone_Bool_3QError_Bool_1_r;
  Go_t lizzieLet0_4QVal_Bool_4QNone_Bool_3QError_Bool_2_d;
  logic lizzieLet0_4QVal_Bool_4QNone_Bool_3QError_Bool_2_r;
  QTree_Bool_t lizzieLet0_4QVal_Bool_4QNone_Bool_3QError_Bool_1QError_Bool_d;
  logic lizzieLet0_4QVal_Bool_4QNone_Bool_3QError_Bool_1QError_Bool_r;
  QTree_Bool_t lizzieLet19_1_argbuf_d;
  logic lizzieLet19_1_argbuf_r;
  Go_t lizzieLet0_4QVal_Bool_4QNone_Bool_3QError_Bool_2_argbuf_d;
  logic lizzieLet0_4QVal_Bool_4QNone_Bool_3QError_Bool_2_argbuf_r;
  Go_t lizzieLet0_4QVal_Bool_4QNone_Bool_3QNode_Bool_1_d;
  logic lizzieLet0_4QVal_Bool_4QNone_Bool_3QNode_Bool_1_r;
  Go_t lizzieLet0_4QVal_Bool_4QNone_Bool_3QNode_Bool_2_d;
  logic lizzieLet0_4QVal_Bool_4QNone_Bool_3QNode_Bool_2_r;
  QTree_Bool_t lizzieLet0_4QVal_Bool_4QNone_Bool_3QNode_Bool_1QError_Bool_d;
  logic lizzieLet0_4QVal_Bool_4QNone_Bool_3QNode_Bool_1QError_Bool_r;
  QTree_Bool_t lizzieLet18_1_argbuf_d;
  logic lizzieLet18_1_argbuf_r;
  Go_t lizzieLet0_4QVal_Bool_4QNone_Bool_3QNode_Bool_2_argbuf_d;
  logic lizzieLet0_4QVal_Bool_4QNone_Bool_3QNode_Bool_2_argbuf_r;
  Go_t lizzieLet0_4QVal_Bool_4QNone_Bool_3QNone_Bool_1_argbuf_d;
  logic lizzieLet0_4QVal_Bool_4QNone_Bool_3QNone_Bool_1_argbuf_r;
  Pointer_QTree_Bool_t lizzieLet0_4QVal_Bool_4QNone_Bool_4QNone_Bool_d;
  logic lizzieLet0_4QVal_Bool_4QNone_Bool_4QNone_Bool_r;
  Pointer_QTree_Bool_t _67_d;
  logic _67_r;
  assign _67_r = 1'd1;
  Pointer_QTree_Bool_t _66_d;
  logic _66_r;
  assign _66_r = 1'd1;
  Pointer_QTree_Bool_t _65_d;
  logic _65_r;
  assign _65_r = 1'd1;
  Pointer_QTree_Bool_t lizzieLet0_4QVal_Bool_4QNone_Bool_4QNone_Bool_1_argbuf_d;
  logic lizzieLet0_4QVal_Bool_4QNone_Bool_4QNone_Bool_1_argbuf_r;
  Pointer_CTf_t lizzieLet0_4QVal_Bool_4QNone_Bool_5QNone_Bool_d;
  logic lizzieLet0_4QVal_Bool_4QNone_Bool_5QNone_Bool_r;
  Pointer_CTf_t lizzieLet0_4QVal_Bool_4QNone_Bool_5QVal_Bool_d;
  logic lizzieLet0_4QVal_Bool_4QNone_Bool_5QVal_Bool_r;
  Pointer_CTf_t lizzieLet0_4QVal_Bool_4QNone_Bool_5QNode_Bool_d;
  logic lizzieLet0_4QVal_Bool_4QNone_Bool_5QNode_Bool_r;
  Pointer_CTf_t lizzieLet0_4QVal_Bool_4QNone_Bool_5QError_Bool_d;
  logic lizzieLet0_4QVal_Bool_4QNone_Bool_5QError_Bool_r;
  Pointer_CTf_t lizzieLet0_4QVal_Bool_4QNone_Bool_5QError_Bool_1_argbuf_d;
  logic lizzieLet0_4QVal_Bool_4QNone_Bool_5QError_Bool_1_argbuf_r;
  Pointer_CTf_t lizzieLet0_4QVal_Bool_4QNone_Bool_5QNode_Bool_1_argbuf_d;
  logic lizzieLet0_4QVal_Bool_4QNone_Bool_5QNode_Bool_1_argbuf_r;
  Pointer_CTf_t lizzieLet0_4QVal_Bool_4QNone_Bool_5QNone_Bool_1_argbuf_d;
  logic lizzieLet0_4QVal_Bool_4QNone_Bool_5QNone_Bool_1_argbuf_r;
  MyBool_t _64_d;
  logic _64_r;
  assign _64_r = 1'd1;
  MyBool_t lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_d;
  logic lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_r;
  MyBool_t _63_d;
  logic _63_r;
  assign _63_r = 1'd1;
  MyBool_t _62_d;
  logic _62_r;
  assign _62_r = 1'd1;
  MyBool_t lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1_d;
  logic lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1_r;
  MyBool_t lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_2_d;
  logic lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_2_r;
  MyBool_t lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3_d;
  logic lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3_r;
  Go_t lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyFalse_d;
  logic lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyFalse_r;
  Go_t lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyTrue_d;
  logic lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyTrue_r;
  Go_t lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyTrue_1_d;
  logic lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyTrue_1_r;
  Go_t lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyTrue_2_d;
  logic lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyTrue_2_r;
  Go_t lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyTrue_1_argbuf_d;
  logic lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyTrue_1_argbuf_r;
  TupGo_t \lvlrf2-0TupGo6_d ;
  logic \lvlrf2-0TupGo6_r ;
  Go_t lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyTrue_2_argbuf_d;
  logic lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyTrue_2_argbuf_r;
  Pointer_CTf_t lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_2MyFalse_d;
  logic lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_2MyFalse_r;
  Pointer_CTf_t lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_2MyTrue_d;
  logic lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_2MyTrue_r;
  Pointer_CTf_t lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_2MyTrue_1_argbuf_d;
  logic lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_2MyTrue_1_argbuf_r;
  MyBool_t lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_d;
  logic lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_r;
  MyBool_t _61_d;
  logic _61_r;
  assign _61_r = 1'd1;
  MyBool_t lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1_d;
  logic lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1_r;
  MyBool_t lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_2_d;
  logic lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_2_r;
  Go_t lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyFalse_d;
  logic lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyFalse_r;
  Go_t lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyTrue_d;
  logic lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyTrue_r;
  Go_t lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyFalse_1_d;
  logic lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyFalse_1_r;
  Go_t lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_d;
  logic lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_r;
  QTree_Bool_t lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_d;
  logic lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_r;
  QTree_Bool_t lizzieLet15_1_1_argbuf_d;
  logic lizzieLet15_1_1_argbuf_r;
  Go_t lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_argbuf_d;
  logic lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_argbuf_r;
  Go_t lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_d;
  logic lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_r;
  Go_t lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_d;
  logic lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_r;
  Go_t lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_argbuf_d;
  logic lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_argbuf_r;
  TupGo_t \lvlrf2-0TupGo5_d ;
  logic \lvlrf2-0TupGo5_r ;
  Go_t lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_argbuf_d;
  logic lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_argbuf_r;
  Pointer_CTf_t lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_2MyFalse_d;
  logic lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_2MyFalse_r;
  Pointer_CTf_t lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_2MyTrue_d;
  logic lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_2MyTrue_r;
  Pointer_CTf_t lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_2MyFalse_1_argbuf_d;
  logic lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_2MyFalse_1_argbuf_r;
  Pointer_CTf_t lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_2MyTrue_1_argbuf_d;
  logic lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_2MyTrue_1_argbuf_r;
  Pointer_QTree_Bool_t lizzieLet0_4QVal_Bool_5QNone_Bool_d;
  logic lizzieLet0_4QVal_Bool_5QNone_Bool_r;
  Pointer_QTree_Bool_t _60_d;
  logic _60_r;
  assign _60_r = 1'd1;
  Pointer_QTree_Bool_t _59_d;
  logic _59_r;
  assign _59_r = 1'd1;
  Pointer_QTree_Bool_t _58_d;
  logic _58_r;
  assign _58_r = 1'd1;
  Pointer_QTree_Bool_t _57_d;
  logic _57_r;
  assign _57_r = 1'd1;
  Pointer_QTree_Bool_t lizzieLet0_4QVal_Bool_6QVal_Bool_d;
  logic lizzieLet0_4QVal_Bool_6QVal_Bool_r;
  Pointer_QTree_Bool_t _56_d;
  logic _56_r;
  assign _56_r = 1'd1;
  Pointer_QTree_Bool_t _55_d;
  logic _55_r;
  assign _55_r = 1'd1;
  Pointer_CTf_t lizzieLet0_4QVal_Bool_7QNone_Bool_d;
  logic lizzieLet0_4QVal_Bool_7QNone_Bool_r;
  Pointer_CTf_t lizzieLet0_4QVal_Bool_7QVal_Bool_d;
  logic lizzieLet0_4QVal_Bool_7QVal_Bool_r;
  Pointer_CTf_t lizzieLet0_4QVal_Bool_7QNode_Bool_d;
  logic lizzieLet0_4QVal_Bool_7QNode_Bool_r;
  Pointer_CTf_t lizzieLet0_4QVal_Bool_7QError_Bool_d;
  logic lizzieLet0_4QVal_Bool_7QError_Bool_r;
  Pointer_CTf_t lizzieLet0_4QVal_Bool_7QError_Bool_1_argbuf_d;
  logic lizzieLet0_4QVal_Bool_7QError_Bool_1_argbuf_r;
  Pointer_CTf_t lizzieLet0_4QVal_Bool_7QNode_Bool_1_argbuf_d;
  logic lizzieLet0_4QVal_Bool_7QNode_Bool_1_argbuf_r;
  MyBool_t lizzieLet0_4QVal_Bool_8QNone_Bool_d;
  logic lizzieLet0_4QVal_Bool_8QNone_Bool_r;
  MyBool_t lizzieLet0_4QVal_Bool_8QVal_Bool_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_r;
  MyBool_t _54_d;
  logic _54_r;
  assign _54_r = 1'd1;
  MyBool_t _53_d;
  logic _53_r;
  assign _53_r = 1'd1;
  MyBool_t lizzieLet0_4QVal_Bool_8QVal_Bool_1_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_1_r;
  MyBool_t lizzieLet0_4QVal_Bool_8QVal_Bool_2_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_2_r;
  MyBool_t lizzieLet0_4QVal_Bool_8QVal_Bool_3_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_3_r;
  MyBool_t lizzieLet0_4QVal_Bool_8QVal_Bool_4_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_4_r;
  MyBool_t lizzieLet0_4QVal_Bool_8QVal_Bool_5_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_5_r;
  Go_t lizzieLet0_4QVal_Bool_8QVal_Bool_1MyFalse_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_1MyFalse_r;
  Go_t lizzieLet0_4QVal_Bool_8QVal_Bool_1MyTrue_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_1MyTrue_r;
  QTree_Bool_t lizzieLet0_4QVal_Bool_8QVal_Bool_2MyFalse_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_2MyFalse_r;
  QTree_Bool_t lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_r;
  QTree_Bool_t lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1_r;
  QTree_Bool_t lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2_r;
  Go_t lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNone_Bool_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNone_Bool_r;
  Go_t lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QVal_Bool_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QVal_Bool_r;
  Go_t lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNode_Bool_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNode_Bool_r;
  Go_t lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QError_Bool_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QError_Bool_r;
  Go_t lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QError_Bool_1_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QError_Bool_1_r;
  Go_t lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QError_Bool_2_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QError_Bool_2_r;
  QTree_Bool_t lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QError_Bool_1QError_Bool_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QError_Bool_1QError_Bool_r;
  QTree_Bool_t lizzieLet29_1_argbuf_d;
  logic lizzieLet29_1_argbuf_r;
  Go_t lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QError_Bool_2_argbuf_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QError_Bool_2_argbuf_r;
  Go_t lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNode_Bool_1_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNode_Bool_1_r;
  Go_t lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNode_Bool_2_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNode_Bool_2_r;
  QTree_Bool_t lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNode_Bool_1QError_Bool_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNode_Bool_1QError_Bool_r;
  QTree_Bool_t lizzieLet28_1_argbuf_d;
  logic lizzieLet28_1_argbuf_r;
  Go_t lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNode_Bool_2_argbuf_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNode_Bool_2_argbuf_r;
  Go_t lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNone_Bool_1_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNone_Bool_1_r;
  Go_t lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNone_Bool_2_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNone_Bool_2_r;
  Go_t lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNone_Bool_1_argbuf_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNone_Bool_1_argbuf_r;
  TupGo_t \lvlrf2-0TupGo9_d ;
  logic \lvlrf2-0TupGo9_r ;
  Go_t lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNone_Bool_2_argbuf_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNone_Bool_2_argbuf_r;
  Go_t lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QVal_Bool_1_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QVal_Bool_1_r;
  Go_t lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QVal_Bool_2_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QVal_Bool_2_r;
  Go_t lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QVal_Bool_1_argbuf_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QVal_Bool_1_argbuf_r;
  TupGo_t \lvlrf2-0TupGo10_d ;
  logic \lvlrf2-0TupGo10_r ;
  Go_t lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QVal_Bool_2_argbuf_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QVal_Bool_2_argbuf_r;
  Pointer_CTf_t lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QNone_Bool_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QNone_Bool_r;
  Pointer_CTf_t lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QVal_Bool_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QVal_Bool_r;
  Pointer_CTf_t lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QNode_Bool_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QNode_Bool_r;
  Pointer_CTf_t lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QError_Bool_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QError_Bool_r;
  Pointer_CTf_t lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QError_Bool_1_argbuf_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QError_Bool_1_argbuf_r;
  Pointer_CTf_t lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QNode_Bool_1_argbuf_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QNode_Bool_1_argbuf_r;
  Pointer_CTf_t lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QNone_Bool_1_argbuf_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QNone_Bool_1_argbuf_r;
  Pointer_CTf_t lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QVal_Bool_1_argbuf_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QVal_Bool_1_argbuf_r;
  Pointer_QTree_Bool_t lizzieLet0_4QVal_Bool_8QVal_Bool_3MyFalse_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_3MyFalse_r;
  Pointer_QTree_Bool_t _52_d;
  logic _52_r;
  assign _52_r = 1'd1;
  Pointer_CTf_t lizzieLet0_4QVal_Bool_8QVal_Bool_4MyFalse_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_4MyFalse_r;
  Pointer_CTf_t lizzieLet0_4QVal_Bool_8QVal_Bool_4MyTrue_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_4MyTrue_r;
  MyBool_t lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_r;
  MyBool_t _51_d;
  logic _51_r;
  assign _51_r = 1'd1;
  MyBool_t lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_1_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_1_r;
  MyBool_t lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2_r;
  MyBool_t lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_3_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_3_r;
  MyBool_t lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_4_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_4_r;
  Go_t lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_1MyFalse_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_1MyFalse_r;
  Go_t lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_1MyTrue_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_1MyTrue_r;
  Go_t lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_1MyFalse_1_argbuf_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_1MyFalse_1_argbuf_r;
  QTree_Bool_t _50_d;
  logic _50_r;
  assign _50_r = 1'd1;
  QTree_Bool_t lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_r;
  QTree_Bool_t lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1_r;
  QTree_Bool_t lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2_r;
  Go_t lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNone_Bool_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNone_Bool_r;
  Go_t lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QVal_Bool_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QVal_Bool_r;
  Go_t lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNode_Bool_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNode_Bool_r;
  Go_t lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QError_Bool_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QError_Bool_r;
  Go_t lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QError_Bool_1_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QError_Bool_1_r;
  Go_t lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QError_Bool_2_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QError_Bool_2_r;
  QTree_Bool_t lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QError_Bool_1QError_Bool_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QError_Bool_1QError_Bool_r;
  QTree_Bool_t lizzieLet24_1_argbuf_d;
  logic lizzieLet24_1_argbuf_r;
  Go_t lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QError_Bool_2_argbuf_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QError_Bool_2_argbuf_r;
  Go_t lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNode_Bool_1_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNode_Bool_1_r;
  Go_t lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNode_Bool_2_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNode_Bool_2_r;
  QTree_Bool_t lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNode_Bool_1QError_Bool_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNode_Bool_1QError_Bool_r;
  QTree_Bool_t lizzieLet23_1_argbuf_d;
  logic lizzieLet23_1_argbuf_r;
  Go_t lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNode_Bool_2_argbuf_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNode_Bool_2_argbuf_r;
  Go_t lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNone_Bool_1_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNone_Bool_1_r;
  Go_t lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNone_Bool_2_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNone_Bool_2_r;
  Go_t lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNone_Bool_1_argbuf_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNone_Bool_1_argbuf_r;
  TupGo_t \lvlrf2-0TupGo7_d ;
  logic \lvlrf2-0TupGo7_r ;
  Go_t lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNone_Bool_2_argbuf_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNone_Bool_2_argbuf_r;
  Go_t lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QVal_Bool_1_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QVal_Bool_1_r;
  Go_t lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QVal_Bool_2_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QVal_Bool_2_r;
  Go_t lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QVal_Bool_1_argbuf_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QVal_Bool_1_argbuf_r;
  TupGo_t \lvlrf2-0TupGo8_d ;
  logic \lvlrf2-0TupGo8_r ;
  Go_t lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QVal_Bool_2_argbuf_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QVal_Bool_2_argbuf_r;
  Pointer_CTf_t lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QNone_Bool_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QNone_Bool_r;
  Pointer_CTf_t lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QVal_Bool_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QVal_Bool_r;
  Pointer_CTf_t lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QNode_Bool_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QNode_Bool_r;
  Pointer_CTf_t lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QError_Bool_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QError_Bool_r;
  Pointer_CTf_t lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QError_Bool_1_argbuf_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QError_Bool_1_argbuf_r;
  Pointer_CTf_t lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QNode_Bool_1_argbuf_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QNode_Bool_1_argbuf_r;
  Pointer_CTf_t lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QNone_Bool_1_argbuf_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QNone_Bool_1_argbuf_r;
  Pointer_CTf_t lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QVal_Bool_1_argbuf_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QVal_Bool_1_argbuf_r;
  Pointer_QTree_Bool_t lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_3MyFalse_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_3MyFalse_r;
  Pointer_QTree_Bool_t _49_d;
  logic _49_r;
  assign _49_r = 1'd1;
  Pointer_QTree_Bool_t lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_3MyFalse_1_argbuf_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_3MyFalse_1_argbuf_r;
  Pointer_CTf_t lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_4MyFalse_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_4MyFalse_r;
  Pointer_CTf_t lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_4MyTrue_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_4MyTrue_r;
  Pointer_CTf_t lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_4MyFalse_1_argbuf_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_4MyFalse_1_argbuf_r;
  QTree_Bool_t lizzieLet0_5QNone_Bool_d;
  logic lizzieLet0_5QNone_Bool_r;
  QTree_Bool_t lizzieLet0_5QVal_Bool_d;
  logic lizzieLet0_5QVal_Bool_r;
  QTree_Bool_t lizzieLet0_5QNode_Bool_d;
  logic lizzieLet0_5QNode_Bool_r;
  QTree_Bool_t _48_d;
  logic _48_r;
  assign _48_r = 1'd1;
  Pointer_QTree_Bool_t _47_d;
  logic _47_r;
  assign _47_r = 1'd1;
  Pointer_QTree_Bool_t lizzieLet0_6QVal_Bool_d;
  logic lizzieLet0_6QVal_Bool_r;
  Pointer_QTree_Bool_t lizzieLet0_6QNode_Bool_d;
  logic lizzieLet0_6QNode_Bool_r;
  Pointer_QTree_Bool_t _46_d;
  logic _46_r;
  assign _46_r = 1'd1;
  Pointer_QTree_Bool_t lizzieLet0_7QNone_Bool_d;
  logic lizzieLet0_7QNone_Bool_r;
  Pointer_QTree_Bool_t _45_d;
  logic _45_r;
  assign _45_r = 1'd1;
  Pointer_QTree_Bool_t _44_d;
  logic _44_r;
  assign _44_r = 1'd1;
  Pointer_QTree_Bool_t _43_d;
  logic _43_r;
  assign _43_r = 1'd1;
  Pointer_QTree_Bool_t lizzieLet0_8QNone_Bool_d;
  logic lizzieLet0_8QNone_Bool_r;
  Pointer_QTree_Bool_t lizzieLet0_8QVal_Bool_d;
  logic lizzieLet0_8QVal_Bool_r;
  Pointer_QTree_Bool_t _42_d;
  logic _42_r;
  assign _42_r = 1'd1;
  Pointer_QTree_Bool_t _41_d;
  logic _41_r;
  assign _41_r = 1'd1;
  Pointer_CTf_t lizzieLet0_9QNone_Bool_d;
  logic lizzieLet0_9QNone_Bool_r;
  Pointer_CTf_t lizzieLet0_9QVal_Bool_d;
  logic lizzieLet0_9QVal_Bool_r;
  Pointer_CTf_t lizzieLet0_9QNode_Bool_d;
  logic lizzieLet0_9QNode_Bool_r;
  Pointer_CTf_t lizzieLet0_9QError_Bool_d;
  logic lizzieLet0_9QError_Bool_r;
  Pointer_CTf_t lizzieLet0_9QError_Bool_1_argbuf_d;
  logic lizzieLet0_9QError_Bool_1_argbuf_r;
  Pointer_QTree_Bool_t q1a98_destruct_d;
  logic q1a98_destruct_r;
  Pointer_QTree_Bool_t q2a99_destruct_d;
  logic q2a99_destruct_r;
  Pointer_QTree_Bool_t q3a9a_destruct_d;
  logic q3a9a_destruct_r;
  Pointer_QTree_Bool_t q5a9b_destruct_d;
  logic q5a9b_destruct_r;
  MyBool_t v1a92_destruct_d;
  logic v1a92_destruct_r;
  QTree_Bool_t _40_d;
  logic _40_r;
  assign _40_r = 1'd1;
  QTree_Bool_t lizzieLet45_1QVal_Bool_d;
  logic lizzieLet45_1QVal_Bool_r;
  QTree_Bool_t lizzieLet45_1QNode_Bool_d;
  logic lizzieLet45_1QNode_Bool_r;
  QTree_Bool_t _39_d;
  logic _39_r;
  assign _39_r = 1'd1;
  Go_t lizzieLet45_3QNone_Bool_d;
  logic lizzieLet45_3QNone_Bool_r;
  Go_t lizzieLet45_3QVal_Bool_d;
  logic lizzieLet45_3QVal_Bool_r;
  Go_t lizzieLet45_3QNode_Bool_d;
  logic lizzieLet45_3QNode_Bool_r;
  Go_t lizzieLet45_3QError_Bool_d;
  logic lizzieLet45_3QError_Bool_r;
  Go_t lizzieLet45_3QError_Bool_1_d;
  logic lizzieLet45_3QError_Bool_1_r;
  Go_t lizzieLet45_3QError_Bool_2_d;
  logic lizzieLet45_3QError_Bool_2_r;
  QTree_Bool_t lizzieLet45_3QError_Bool_1QError_Bool_d;
  logic lizzieLet45_3QError_Bool_1QError_Bool_r;
  QTree_Bool_t lizzieLet56_1_argbuf_d;
  logic lizzieLet56_1_argbuf_r;
  Go_t lizzieLet45_3QError_Bool_2_argbuf_d;
  logic lizzieLet45_3QError_Bool_2_argbuf_r;
  Go_t lizzieLet45_3QNone_Bool_1_argbuf_d;
  logic lizzieLet45_3QNone_Bool_1_argbuf_r;
  C12_t go_8_goMux_choice_d;
  logic go_8_goMux_choice_r;
  Go_t go_8_goMux_data_d;
  logic go_8_goMux_data_r;
  QTree_Bool_t _38_d;
  logic _38_r;
  assign _38_r = 1'd1;
  QTree_Bool_t lizzieLet45_4QVal_Bool_d;
  logic lizzieLet45_4QVal_Bool_r;
  QTree_Bool_t lizzieLet45_4QNode_Bool_d;
  logic lizzieLet45_4QNode_Bool_r;
  QTree_Bool_t _37_d;
  logic _37_r;
  assign _37_r = 1'd1;
  QTree_Bool_t lizzieLet45_4QNode_Bool_1_d;
  logic lizzieLet45_4QNode_Bool_1_r;
  QTree_Bool_t lizzieLet45_4QNode_Bool_2_d;
  logic lizzieLet45_4QNode_Bool_2_r;
  QTree_Bool_t lizzieLet45_4QNode_Bool_3_d;
  logic lizzieLet45_4QNode_Bool_3_r;
  QTree_Bool_t lizzieLet45_4QNode_Bool_4_d;
  logic lizzieLet45_4QNode_Bool_4_r;
  QTree_Bool_t lizzieLet45_4QNode_Bool_5_d;
  logic lizzieLet45_4QNode_Bool_5_r;
  QTree_Bool_t lizzieLet45_4QNode_Bool_6_d;
  logic lizzieLet45_4QNode_Bool_6_r;
  QTree_Bool_t lizzieLet45_4QNode_Bool_7_d;
  logic lizzieLet45_4QNode_Bool_7_r;
  QTree_Bool_t lizzieLet45_4QNode_Bool_8_d;
  logic lizzieLet45_4QNode_Bool_8_r;
  QTree_Bool_t lizzieLet45_4QNode_Bool_9_d;
  logic lizzieLet45_4QNode_Bool_9_r;
  Pointer_QTree_Bool_t t1a9d_destruct_d;
  logic t1a9d_destruct_r;
  Pointer_QTree_Bool_t t2a9e_destruct_d;
  logic t2a9e_destruct_r;
  Pointer_QTree_Bool_t t3a9f_destruct_d;
  logic t3a9f_destruct_r;
  Pointer_QTree_Bool_t t5a9g_destruct_d;
  logic t5a9g_destruct_r;
  QTree_Bool_t _36_d;
  logic _36_r;
  assign _36_r = 1'd1;
  QTree_Bool_t _35_d;
  logic _35_r;
  assign _35_r = 1'd1;
  QTree_Bool_t lizzieLet45_4QNode_Bool_1QNode_Bool_d;
  logic lizzieLet45_4QNode_Bool_1QNode_Bool_r;
  QTree_Bool_t _34_d;
  logic _34_r;
  assign _34_r = 1'd1;
  Go_t lizzieLet45_4QNode_Bool_3QNone_Bool_d;
  logic lizzieLet45_4QNode_Bool_3QNone_Bool_r;
  Go_t lizzieLet45_4QNode_Bool_3QVal_Bool_d;
  logic lizzieLet45_4QNode_Bool_3QVal_Bool_r;
  Go_t lizzieLet45_4QNode_Bool_3QNode_Bool_d;
  logic lizzieLet45_4QNode_Bool_3QNode_Bool_r;
  Go_t lizzieLet45_4QNode_Bool_3QError_Bool_d;
  logic lizzieLet45_4QNode_Bool_3QError_Bool_r;
  Go_t lizzieLet45_4QNode_Bool_3QError_Bool_1_d;
  logic lizzieLet45_4QNode_Bool_3QError_Bool_1_r;
  Go_t lizzieLet45_4QNode_Bool_3QError_Bool_2_d;
  logic lizzieLet45_4QNode_Bool_3QError_Bool_2_r;
  QTree_Bool_t lizzieLet45_4QNode_Bool_3QError_Bool_1QError_Bool_d;
  logic lizzieLet45_4QNode_Bool_3QError_Bool_1QError_Bool_r;
  QTree_Bool_t lizzieLet55_1_argbuf_d;
  logic lizzieLet55_1_argbuf_r;
  Go_t lizzieLet45_4QNode_Bool_3QError_Bool_2_argbuf_d;
  logic lizzieLet45_4QNode_Bool_3QError_Bool_2_argbuf_r;
  Go_t lizzieLet45_4QNode_Bool_3QNode_Bool_1_argbuf_d;
  logic lizzieLet45_4QNode_Bool_3QNode_Bool_1_argbuf_r;
  Go_t lizzieLet45_4QNode_Bool_3QNone_Bool_1_argbuf_d;
  logic lizzieLet45_4QNode_Bool_3QNone_Bool_1_argbuf_r;
  Go_t lizzieLet45_4QNode_Bool_3QVal_Bool_1_d;
  logic lizzieLet45_4QNode_Bool_3QVal_Bool_1_r;
  Go_t lizzieLet45_4QNode_Bool_3QVal_Bool_2_d;
  logic lizzieLet45_4QNode_Bool_3QVal_Bool_2_r;
  QTree_Bool_t lizzieLet45_4QNode_Bool_3QVal_Bool_1QError_Bool_d;
  logic lizzieLet45_4QNode_Bool_3QVal_Bool_1QError_Bool_r;
  QTree_Bool_t lizzieLet53_1_argbuf_d;
  logic lizzieLet53_1_argbuf_r;
  Go_t lizzieLet45_4QNode_Bool_3QVal_Bool_2_argbuf_d;
  logic lizzieLet45_4QNode_Bool_3QVal_Bool_2_argbuf_r;
  Pointer_QTree_Bool_t lizzieLet45_4QNode_Bool_4QNone_Bool_d;
  logic lizzieLet45_4QNode_Bool_4QNone_Bool_r;
  Pointer_QTree_Bool_t _33_d;
  logic _33_r;
  assign _33_r = 1'd1;
  Pointer_QTree_Bool_t _32_d;
  logic _32_r;
  assign _32_r = 1'd1;
  Pointer_QTree_Bool_t _31_d;
  logic _31_r;
  assign _31_r = 1'd1;
  Pointer_QTree_Bool_t lizzieLet45_4QNode_Bool_4QNone_Bool_1_argbuf_d;
  logic lizzieLet45_4QNode_Bool_4QNone_Bool_1_argbuf_r;
  \Pointer_CTf''''''''''''_t  lizzieLet45_4QNode_Bool_5QNone_Bool_d;
  logic lizzieLet45_4QNode_Bool_5QNone_Bool_r;
  \Pointer_CTf''''''''''''_t  lizzieLet45_4QNode_Bool_5QVal_Bool_d;
  logic lizzieLet45_4QNode_Bool_5QVal_Bool_r;
  \Pointer_CTf''''''''''''_t  lizzieLet45_4QNode_Bool_5QNode_Bool_d;
  logic lizzieLet45_4QNode_Bool_5QNode_Bool_r;
  \Pointer_CTf''''''''''''_t  lizzieLet45_4QNode_Bool_5QError_Bool_d;
  logic lizzieLet45_4QNode_Bool_5QError_Bool_r;
  \Pointer_CTf''''''''''''_t  lizzieLet45_4QNode_Bool_5QError_Bool_1_argbuf_d;
  logic lizzieLet45_4QNode_Bool_5QError_Bool_1_argbuf_r;
  \CTf''''''''''''_t  \lizzieLet45_4QNode_Bool_5QNode_Bool_1lizzieLet45_4QNode_Bool_6QNode_Bool_1t1a9d_1lizzieLet45_4QNode_Bool_7QNode_Bool_1t2a9e_1lizzieLet45_4QNode_Bool_8QNode_Bool_1t3a9f_1Lcall_f''''''''''''3_d ;
  logic \lizzieLet45_4QNode_Bool_5QNode_Bool_1lizzieLet45_4QNode_Bool_6QNode_Bool_1t1a9d_1lizzieLet45_4QNode_Bool_7QNode_Bool_1t2a9e_1lizzieLet45_4QNode_Bool_8QNode_Bool_1t3a9f_1Lcall_f''''''''''''3_r ;
  \CTf''''''''''''_t  lizzieLet54_1_argbuf_d;
  logic lizzieLet54_1_argbuf_r;
  \Pointer_CTf''''''''''''_t  lizzieLet45_4QNode_Bool_5QNone_Bool_1_argbuf_d;
  logic lizzieLet45_4QNode_Bool_5QNone_Bool_1_argbuf_r;
  \Pointer_CTf''''''''''''_t  lizzieLet45_4QNode_Bool_5QVal_Bool_1_argbuf_d;
  logic lizzieLet45_4QNode_Bool_5QVal_Bool_1_argbuf_r;
  Pointer_QTree_Bool_t _30_d;
  logic _30_r;
  assign _30_r = 1'd1;
  Pointer_QTree_Bool_t _29_d;
  logic _29_r;
  assign _29_r = 1'd1;
  Pointer_QTree_Bool_t lizzieLet45_4QNode_Bool_6QNode_Bool_d;
  logic lizzieLet45_4QNode_Bool_6QNode_Bool_r;
  Pointer_QTree_Bool_t _28_d;
  logic _28_r;
  assign _28_r = 1'd1;
  Pointer_QTree_Bool_t _27_d;
  logic _27_r;
  assign _27_r = 1'd1;
  Pointer_QTree_Bool_t _26_d;
  logic _26_r;
  assign _26_r = 1'd1;
  Pointer_QTree_Bool_t lizzieLet45_4QNode_Bool_7QNode_Bool_d;
  logic lizzieLet45_4QNode_Bool_7QNode_Bool_r;
  Pointer_QTree_Bool_t _25_d;
  logic _25_r;
  assign _25_r = 1'd1;
  Pointer_QTree_Bool_t _24_d;
  logic _24_r;
  assign _24_r = 1'd1;
  Pointer_QTree_Bool_t _23_d;
  logic _23_r;
  assign _23_r = 1'd1;
  Pointer_QTree_Bool_t lizzieLet45_4QNode_Bool_8QNode_Bool_d;
  logic lizzieLet45_4QNode_Bool_8QNode_Bool_r;
  Pointer_QTree_Bool_t _22_d;
  logic _22_r;
  assign _22_r = 1'd1;
  Pointer_QTree_Bool_t _21_d;
  logic _21_r;
  assign _21_r = 1'd1;
  Pointer_QTree_Bool_t _20_d;
  logic _20_r;
  assign _20_r = 1'd1;
  Pointer_QTree_Bool_t lizzieLet45_4QNode_Bool_9QNode_Bool_d;
  logic lizzieLet45_4QNode_Bool_9QNode_Bool_r;
  Pointer_QTree_Bool_t _19_d;
  logic _19_r;
  assign _19_r = 1'd1;
  Pointer_QTree_Bool_t lizzieLet45_4QNode_Bool_9QNode_Bool_1_argbuf_d;
  logic lizzieLet45_4QNode_Bool_9QNode_Bool_1_argbuf_r;
  QTree_Bool_t lizzieLet45_4QVal_Bool_1_d;
  logic lizzieLet45_4QVal_Bool_1_r;
  QTree_Bool_t lizzieLet45_4QVal_Bool_2_d;
  logic lizzieLet45_4QVal_Bool_2_r;
  QTree_Bool_t lizzieLet45_4QVal_Bool_3_d;
  logic lizzieLet45_4QVal_Bool_3_r;
  QTree_Bool_t lizzieLet45_4QVal_Bool_4_d;
  logic lizzieLet45_4QVal_Bool_4_r;
  QTree_Bool_t lizzieLet45_4QVal_Bool_5_d;
  logic lizzieLet45_4QVal_Bool_5_r;
  QTree_Bool_t lizzieLet45_4QVal_Bool_6_d;
  logic lizzieLet45_4QVal_Bool_6_r;
  MyBool_t va93_destruct_d;
  logic va93_destruct_r;
  QTree_Bool_t _18_d;
  logic _18_r;
  assign _18_r = 1'd1;
  QTree_Bool_t lizzieLet45_4QVal_Bool_1QVal_Bool_d;
  logic lizzieLet45_4QVal_Bool_1QVal_Bool_r;
  QTree_Bool_t _17_d;
  logic _17_r;
  assign _17_r = 1'd1;
  QTree_Bool_t _16_d;
  logic _16_r;
  assign _16_r = 1'd1;
  Go_t lizzieLet45_4QVal_Bool_3QNone_Bool_d;
  logic lizzieLet45_4QVal_Bool_3QNone_Bool_r;
  Go_t lizzieLet45_4QVal_Bool_3QVal_Bool_d;
  logic lizzieLet45_4QVal_Bool_3QVal_Bool_r;
  Go_t lizzieLet45_4QVal_Bool_3QNode_Bool_d;
  logic lizzieLet45_4QVal_Bool_3QNode_Bool_r;
  Go_t lizzieLet45_4QVal_Bool_3QError_Bool_d;
  logic lizzieLet45_4QVal_Bool_3QError_Bool_r;
  Go_t lizzieLet45_4QVal_Bool_3QError_Bool_1_d;
  logic lizzieLet45_4QVal_Bool_3QError_Bool_1_r;
  Go_t lizzieLet45_4QVal_Bool_3QError_Bool_2_d;
  logic lizzieLet45_4QVal_Bool_3QError_Bool_2_r;
  QTree_Bool_t lizzieLet45_4QVal_Bool_3QError_Bool_1QError_Bool_d;
  logic lizzieLet45_4QVal_Bool_3QError_Bool_1QError_Bool_r;
  QTree_Bool_t lizzieLet51_1_argbuf_d;
  logic lizzieLet51_1_argbuf_r;
  Go_t lizzieLet45_4QVal_Bool_3QError_Bool_2_argbuf_d;
  logic lizzieLet45_4QVal_Bool_3QError_Bool_2_argbuf_r;
  Go_t lizzieLet45_4QVal_Bool_3QNode_Bool_1_d;
  logic lizzieLet45_4QVal_Bool_3QNode_Bool_1_r;
  Go_t lizzieLet45_4QVal_Bool_3QNode_Bool_2_d;
  logic lizzieLet45_4QVal_Bool_3QNode_Bool_2_r;
  QTree_Bool_t lizzieLet45_4QVal_Bool_3QNode_Bool_1QError_Bool_d;
  logic lizzieLet45_4QVal_Bool_3QNode_Bool_1QError_Bool_r;
  QTree_Bool_t lizzieLet50_1_argbuf_d;
  logic lizzieLet50_1_argbuf_r;
  Go_t lizzieLet45_4QVal_Bool_3QNode_Bool_2_argbuf_d;
  logic lizzieLet45_4QVal_Bool_3QNode_Bool_2_argbuf_r;
  Go_t lizzieLet45_4QVal_Bool_3QNone_Bool_1_argbuf_d;
  logic lizzieLet45_4QVal_Bool_3QNone_Bool_1_argbuf_r;
  Pointer_QTree_Bool_t lizzieLet45_4QVal_Bool_4QNone_Bool_d;
  logic lizzieLet45_4QVal_Bool_4QNone_Bool_r;
  Pointer_QTree_Bool_t _15_d;
  logic _15_r;
  assign _15_r = 1'd1;
  Pointer_QTree_Bool_t _14_d;
  logic _14_r;
  assign _14_r = 1'd1;
  Pointer_QTree_Bool_t _13_d;
  logic _13_r;
  assign _13_r = 1'd1;
  Pointer_QTree_Bool_t lizzieLet45_4QVal_Bool_4QNone_Bool_1_argbuf_d;
  logic lizzieLet45_4QVal_Bool_4QNone_Bool_1_argbuf_r;
  \Pointer_CTf''''''''''''_t  lizzieLet45_4QVal_Bool_5QNone_Bool_d;
  logic lizzieLet45_4QVal_Bool_5QNone_Bool_r;
  \Pointer_CTf''''''''''''_t  lizzieLet45_4QVal_Bool_5QVal_Bool_d;
  logic lizzieLet45_4QVal_Bool_5QVal_Bool_r;
  \Pointer_CTf''''''''''''_t  lizzieLet45_4QVal_Bool_5QNode_Bool_d;
  logic lizzieLet45_4QVal_Bool_5QNode_Bool_r;
  \Pointer_CTf''''''''''''_t  lizzieLet45_4QVal_Bool_5QError_Bool_d;
  logic lizzieLet45_4QVal_Bool_5QError_Bool_r;
  \Pointer_CTf''''''''''''_t  lizzieLet45_4QVal_Bool_5QError_Bool_1_argbuf_d;
  logic lizzieLet45_4QVal_Bool_5QError_Bool_1_argbuf_r;
  \Pointer_CTf''''''''''''_t  lizzieLet45_4QVal_Bool_5QNode_Bool_1_argbuf_d;
  logic lizzieLet45_4QVal_Bool_5QNode_Bool_1_argbuf_r;
  \Pointer_CTf''''''''''''_t  lizzieLet45_4QVal_Bool_5QNone_Bool_1_argbuf_d;
  logic lizzieLet45_4QVal_Bool_5QNone_Bool_1_argbuf_r;
  MyBool_t _12_d;
  logic _12_r;
  assign _12_r = 1'd1;
  MyBool_t lizzieLet45_4QVal_Bool_6QVal_Bool_d;
  logic lizzieLet45_4QVal_Bool_6QVal_Bool_r;
  MyBool_t _11_d;
  logic _11_r;
  assign _11_r = 1'd1;
  MyBool_t _10_d;
  logic _10_r;
  assign _10_r = 1'd1;
  MyBool_t lizzieLet45_4QVal_Bool_6QVal_Bool_1_d;
  logic lizzieLet45_4QVal_Bool_6QVal_Bool_1_r;
  MyBool_t lizzieLet45_4QVal_Bool_6QVal_Bool_2_d;
  logic lizzieLet45_4QVal_Bool_6QVal_Bool_2_r;
  MyBool_t lizzieLet45_4QVal_Bool_6QVal_Bool_3_d;
  logic lizzieLet45_4QVal_Bool_6QVal_Bool_3_r;
  Go_t lizzieLet45_4QVal_Bool_6QVal_Bool_1MyFalse_d;
  logic lizzieLet45_4QVal_Bool_6QVal_Bool_1MyFalse_r;
  Go_t lizzieLet45_4QVal_Bool_6QVal_Bool_1MyTrue_d;
  logic lizzieLet45_4QVal_Bool_6QVal_Bool_1MyTrue_r;
  Go_t lizzieLet45_4QVal_Bool_6QVal_Bool_1MyTrue_1_d;
  logic lizzieLet45_4QVal_Bool_6QVal_Bool_1MyTrue_1_r;
  Go_t lizzieLet45_4QVal_Bool_6QVal_Bool_1MyTrue_2_d;
  logic lizzieLet45_4QVal_Bool_6QVal_Bool_1MyTrue_2_r;
  Go_t lizzieLet45_4QVal_Bool_6QVal_Bool_1MyTrue_1_argbuf_d;
  logic lizzieLet45_4QVal_Bool_6QVal_Bool_1MyTrue_1_argbuf_r;
  TupGo_t \lvlrf2-0TupGo4_d ;
  logic \lvlrf2-0TupGo4_r ;
  Go_t lizzieLet45_4QVal_Bool_6QVal_Bool_1MyTrue_2_argbuf_d;
  logic lizzieLet45_4QVal_Bool_6QVal_Bool_1MyTrue_2_argbuf_r;
  \Pointer_CTf''''''''''''_t  lizzieLet45_4QVal_Bool_6QVal_Bool_2MyFalse_d;
  logic lizzieLet45_4QVal_Bool_6QVal_Bool_2MyFalse_r;
  \Pointer_CTf''''''''''''_t  lizzieLet45_4QVal_Bool_6QVal_Bool_2MyTrue_d;
  logic lizzieLet45_4QVal_Bool_6QVal_Bool_2MyTrue_r;
  \Pointer_CTf''''''''''''_t  lizzieLet45_4QVal_Bool_6QVal_Bool_2MyTrue_1_argbuf_d;
  logic lizzieLet45_4QVal_Bool_6QVal_Bool_2MyTrue_1_argbuf_r;
  MyBool_t lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_d;
  logic lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_r;
  MyBool_t _9_d;
  logic _9_r;
  assign _9_r = 1'd1;
  MyBool_t lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1_d;
  logic lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1_r;
  MyBool_t lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_2_d;
  logic lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_2_r;
  Go_t lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_d;
  logic lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_r;
  Go_t lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_d;
  logic lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_r;
  Go_t lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1_d;
  logic lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1_r;
  Go_t lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_d;
  logic lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_r;
  QTree_Bool_t lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_d;
  logic lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_r;
  QTree_Bool_t lizzieLet47_1_argbuf_d;
  logic lizzieLet47_1_argbuf_r;
  Go_t lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_argbuf_d;
  logic lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_argbuf_r;
  Go_t lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_d;
  logic lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_r;
  Go_t lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_d;
  logic lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_r;
  Go_t lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_argbuf_d;
  logic lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_argbuf_r;
  TupGo_t \lvlrf2-0TupGo3_d ;
  logic \lvlrf2-0TupGo3_r ;
  Go_t lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_argbuf_d;
  logic lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_argbuf_r;
  \Pointer_CTf''''''''''''_t  lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_2MyFalse_d;
  logic lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_2MyFalse_r;
  \Pointer_CTf''''''''''''_t  lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_2MyTrue_d;
  logic lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_2MyTrue_r;
  \Pointer_CTf''''''''''''_t  lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_2MyFalse_1_argbuf_d;
  logic lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_2MyFalse_1_argbuf_r;
  \Pointer_CTf''''''''''''_t  lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_2MyTrue_1_argbuf_d;
  logic lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_2MyTrue_1_argbuf_r;
  Pointer_QTree_Bool_t _8_d;
  logic _8_r;
  assign _8_r = 1'd1;
  Pointer_QTree_Bool_t lizzieLet45_5QVal_Bool_d;
  logic lizzieLet45_5QVal_Bool_r;
  Pointer_QTree_Bool_t lizzieLet45_5QNode_Bool_d;
  logic lizzieLet45_5QNode_Bool_r;
  Pointer_QTree_Bool_t _7_d;
  logic _7_r;
  assign _7_r = 1'd1;
  \Pointer_CTf''''''''''''_t  lizzieLet45_6QNone_Bool_d;
  logic lizzieLet45_6QNone_Bool_r;
  \Pointer_CTf''''''''''''_t  lizzieLet45_6QVal_Bool_d;
  logic lizzieLet45_6QVal_Bool_r;
  \Pointer_CTf''''''''''''_t  lizzieLet45_6QNode_Bool_d;
  logic lizzieLet45_6QNode_Bool_r;
  \Pointer_CTf''''''''''''_t  lizzieLet45_6QError_Bool_d;
  logic lizzieLet45_6QError_Bool_r;
  \Pointer_CTf''''''''''''_t  lizzieLet45_6QError_Bool_1_argbuf_d;
  logic lizzieLet45_6QError_Bool_1_argbuf_r;
  \Pointer_CTf''''''''''''_t  lizzieLet45_6QNone_Bool_1_argbuf_d;
  logic lizzieLet45_6QNone_Bool_1_argbuf_r;
  Pointer_QTree_Bool_t lizzieLet45_7QNone_Bool_d;
  logic lizzieLet45_7QNone_Bool_r;
  Pointer_QTree_Bool_t _6_d;
  logic _6_r;
  assign _6_r = 1'd1;
  Pointer_QTree_Bool_t _5_d;
  logic _5_r;
  assign _5_r = 1'd1;
  Pointer_QTree_Bool_t _4_d;
  logic _4_r;
  assign _4_r = 1'd1;
  Pointer_QTree_Bool_t lizzieLet45_7QNone_Bool_1_argbuf_d;
  logic lizzieLet45_7QNone_Bool_1_argbuf_r;
  Pointer_QTree_Bool_t es_13_destruct_d;
  logic es_13_destruct_r;
  Pointer_QTree_Bool_t es_14_1_destruct_d;
  logic es_14_1_destruct_r;
  Pointer_QTree_Bool_t es_15_2_destruct_d;
  logic es_15_2_destruct_r;
  Pointer_CTf_t sc_0_5_destruct_d;
  logic sc_0_5_destruct_r;
  Pointer_QTree_Bool_t es_14_destruct_d;
  logic es_14_destruct_r;
  Pointer_QTree_Bool_t es_15_1_destruct_d;
  logic es_15_1_destruct_r;
  Pointer_CTf_t sc_0_4_destruct_d;
  logic sc_0_4_destruct_r;
  Pointer_QTree_Bool_t q1a8H_3_destruct_d;
  logic q1a8H_3_destruct_r;
  Pointer_QTree_Bool_t t1a8R_3_destruct_d;
  logic t1a8R_3_destruct_r;
  Pointer_QTree_Bool_t \t1'a8W_3_destruct_d ;
  logic \t1'a8W_3_destruct_r ;
  Pointer_QTree_Bool_t es_15_destruct_d;
  logic es_15_destruct_r;
  Pointer_CTf_t sc_0_3_destruct_d;
  logic sc_0_3_destruct_r;
  Pointer_QTree_Bool_t q1a8H_2_destruct_d;
  logic q1a8H_2_destruct_r;
  Pointer_QTree_Bool_t t1a8R_2_destruct_d;
  logic t1a8R_2_destruct_r;
  Pointer_QTree_Bool_t \t1'a8W_2_destruct_d ;
  logic \t1'a8W_2_destruct_r ;
  Pointer_QTree_Bool_t q2a8I_2_destruct_d;
  logic q2a8I_2_destruct_r;
  Pointer_QTree_Bool_t t2a8S_2_destruct_d;
  logic t2a8S_2_destruct_r;
  Pointer_QTree_Bool_t \t2'a8X_2_destruct_d ;
  logic \t2'a8X_2_destruct_r ;
  Pointer_CTf_t sc_0_2_destruct_d;
  logic sc_0_2_destruct_r;
  Pointer_QTree_Bool_t q1a8H_1_destruct_d;
  logic q1a8H_1_destruct_r;
  Pointer_QTree_Bool_t t1a8R_1_destruct_d;
  logic t1a8R_1_destruct_r;
  Pointer_QTree_Bool_t \t1'a8W_1_destruct_d ;
  logic \t1'a8W_1_destruct_r ;
  Pointer_QTree_Bool_t q2a8I_1_destruct_d;
  logic q2a8I_1_destruct_r;
  Pointer_QTree_Bool_t t2a8S_1_destruct_d;
  logic t2a8S_1_destruct_r;
  Pointer_QTree_Bool_t \t2'a8X_1_destruct_d ;
  logic \t2'a8X_1_destruct_r ;
  Pointer_QTree_Bool_t q3a8J_1_destruct_d;
  logic q3a8J_1_destruct_r;
  Pointer_QTree_Bool_t t3a8T_1_destruct_d;
  logic t3a8T_1_destruct_r;
  Pointer_QTree_Bool_t \t3'a8Y_1_destruct_d ;
  logic \t3'a8Y_1_destruct_r ;
  CTf_t _3_d;
  logic _3_r;
  assign _3_r = 1'd1;
  CTf_t lizzieLet60_1Lcall_f3_d;
  logic lizzieLet60_1Lcall_f3_r;
  CTf_t lizzieLet60_1Lcall_f2_d;
  logic lizzieLet60_1Lcall_f2_r;
  CTf_t lizzieLet60_1Lcall_f1_d;
  logic lizzieLet60_1Lcall_f1_r;
  CTf_t lizzieLet60_1Lcall_f0_d;
  logic lizzieLet60_1Lcall_f0_r;
  Go_t _2_d;
  logic _2_r;
  assign _2_r = 1'd1;
  Go_t lizzieLet60_3Lcall_f3_d;
  logic lizzieLet60_3Lcall_f3_r;
  Go_t lizzieLet60_3Lcall_f2_d;
  logic lizzieLet60_3Lcall_f2_r;
  Go_t lizzieLet60_3Lcall_f1_d;
  logic lizzieLet60_3Lcall_f1_r;
  Go_t lizzieLet60_3Lcall_f0_d;
  logic lizzieLet60_3Lcall_f0_r;
  Go_t lizzieLet60_3Lcall_f0_1_argbuf_d;
  logic lizzieLet60_3Lcall_f0_1_argbuf_r;
  Go_t lizzieLet60_3Lcall_f1_1_argbuf_d;
  logic lizzieLet60_3Lcall_f1_1_argbuf_r;
  Go_t lizzieLet60_3Lcall_f2_1_argbuf_d;
  logic lizzieLet60_3Lcall_f2_1_argbuf_r;
  Go_t lizzieLet60_3Lcall_f3_1_argbuf_d;
  logic lizzieLet60_3Lcall_f3_1_argbuf_r;
  Pointer_QTree_Bool_t lizzieLet60_4Lfsbos_d;
  logic lizzieLet60_4Lfsbos_r;
  Pointer_QTree_Bool_t lizzieLet60_4Lcall_f3_d;
  logic lizzieLet60_4Lcall_f3_r;
  Pointer_QTree_Bool_t lizzieLet60_4Lcall_f2_d;
  logic lizzieLet60_4Lcall_f2_r;
  Pointer_QTree_Bool_t lizzieLet60_4Lcall_f1_d;
  logic lizzieLet60_4Lcall_f1_r;
  Pointer_QTree_Bool_t lizzieLet60_4Lcall_f0_d;
  logic lizzieLet60_4Lcall_f0_r;
  QTree_Bool_t lizzieLet60_4Lcall_f0_1es_13_1es_14_1_1es_15_2_1QNode_Bool_d;
  logic lizzieLet60_4Lcall_f0_1es_13_1es_14_1_1es_15_2_1QNode_Bool_r;
  QTree_Bool_t lizzieLet64_1_argbuf_d;
  logic lizzieLet64_1_argbuf_r;
  CTf_t lizzieLet60_4Lcall_f1_1es_14_1es_15_1_1sc_0_4_1Lcall_f0_d;
  logic lizzieLet60_4Lcall_f1_1es_14_1es_15_1_1sc_0_4_1Lcall_f0_r;
  CTf_t lizzieLet63_1_argbuf_d;
  logic lizzieLet63_1_argbuf_r;
  CTf_t \lizzieLet60_4Lcall_f2_1es_15_1sc_0_3_1q1a8H_2_1t1a8R_2_1t1'a8W_2_1Lcall_f1_d ;
  logic \lizzieLet60_4Lcall_f2_1es_15_1sc_0_3_1q1a8H_2_1t1a8R_2_1t1'a8W_2_1Lcall_f1_r ;
  CTf_t lizzieLet62_1_argbuf_d;
  logic lizzieLet62_1_argbuf_r;
  CTf_t \lizzieLet60_4Lcall_f3_1sc_0_2_1q1a8H_1_1t1a8R_1_1t1'a8W_1_1q2a8I_1_1t2a8S_1_1t2'a8X_1_1Lcall_f2_d ;
  logic \lizzieLet60_4Lcall_f3_1sc_0_2_1q1a8H_1_1t1a8R_1_1t1'a8W_1_1q2a8I_1_1t2a8S_1_1t2'a8X_1_1Lcall_f2_r ;
  CTf_t lizzieLet61_1_argbuf_d;
  logic lizzieLet61_1_argbuf_r;
  Pointer_QTree_Bool_t lizzieLet60_4Lfsbos_1_merge_merge_merge_fork_1_d;
  logic lizzieLet60_4Lfsbos_1_merge_merge_merge_fork_1_r;
  Pointer_QTree_Bool_t lizzieLet60_4Lfsbos_1_merge_merge_merge_fork_2_d;
  logic lizzieLet60_4Lfsbos_1_merge_merge_merge_fork_2_r;
  Go_t call_f_goConst_d;
  logic call_f_goConst_r;
  Pointer_QTree_Bool_t f_resbuf_d;
  logic f_resbuf_r;
  Pointer_QTree_Bool_t es_1_1_destruct_d;
  logic es_1_1_destruct_r;
  Pointer_QTree_Bool_t es_2_2_destruct_d;
  logic es_2_2_destruct_r;
  Pointer_QTree_Bool_t es_3_3_destruct_d;
  logic es_3_3_destruct_r;
  \Pointer_CTf''''''''''''_t  sc_0_9_destruct_d;
  logic sc_0_9_destruct_r;
  Pointer_QTree_Bool_t es_2_1_destruct_d;
  logic es_2_1_destruct_r;
  Pointer_QTree_Bool_t es_3_2_destruct_d;
  logic es_3_2_destruct_r;
  \Pointer_CTf''''''''''''_t  sc_0_8_destruct_d;
  logic sc_0_8_destruct_r;
  Pointer_QTree_Bool_t q1a98_3_destruct_d;
  logic q1a98_3_destruct_r;
  Pointer_QTree_Bool_t t1a9d_3_destruct_d;
  logic t1a9d_3_destruct_r;
  Pointer_QTree_Bool_t es_3_1_destruct_d;
  logic es_3_1_destruct_r;
  \Pointer_CTf''''''''''''_t  sc_0_7_destruct_d;
  logic sc_0_7_destruct_r;
  Pointer_QTree_Bool_t q1a98_2_destruct_d;
  logic q1a98_2_destruct_r;
  Pointer_QTree_Bool_t t1a9d_2_destruct_d;
  logic t1a9d_2_destruct_r;
  Pointer_QTree_Bool_t q2a99_2_destruct_d;
  logic q2a99_2_destruct_r;
  Pointer_QTree_Bool_t t2a9e_2_destruct_d;
  logic t2a9e_2_destruct_r;
  \Pointer_CTf''''''''''''_t  sc_0_6_destruct_d;
  logic sc_0_6_destruct_r;
  Pointer_QTree_Bool_t q1a98_1_destruct_d;
  logic q1a98_1_destruct_r;
  Pointer_QTree_Bool_t t1a9d_1_destruct_d;
  logic t1a9d_1_destruct_r;
  Pointer_QTree_Bool_t q2a99_1_destruct_d;
  logic q2a99_1_destruct_r;
  Pointer_QTree_Bool_t t2a9e_1_destruct_d;
  logic t2a9e_1_destruct_r;
  Pointer_QTree_Bool_t q3a9a_1_destruct_d;
  logic q3a9a_1_destruct_r;
  Pointer_QTree_Bool_t t3a9f_1_destruct_d;
  logic t3a9f_1_destruct_r;
  \CTf''''''''''''_t  _1_d;
  logic _1_r;
  assign _1_r = 1'd1;
  \CTf''''''''''''_t  \lizzieLet65_1Lcall_f''''''''''''3_d ;
  logic \lizzieLet65_1Lcall_f''''''''''''3_r ;
  \CTf''''''''''''_t  \lizzieLet65_1Lcall_f''''''''''''2_d ;
  logic \lizzieLet65_1Lcall_f''''''''''''2_r ;
  \CTf''''''''''''_t  \lizzieLet65_1Lcall_f''''''''''''1_d ;
  logic \lizzieLet65_1Lcall_f''''''''''''1_r ;
  \CTf''''''''''''_t  \lizzieLet65_1Lcall_f''''''''''''0_d ;
  logic \lizzieLet65_1Lcall_f''''''''''''0_r ;
  Go_t _0_d;
  logic _0_r;
  assign _0_r = 1'd1;
  Go_t \lizzieLet65_3Lcall_f''''''''''''3_d ;
  logic \lizzieLet65_3Lcall_f''''''''''''3_r ;
  Go_t \lizzieLet65_3Lcall_f''''''''''''2_d ;
  logic \lizzieLet65_3Lcall_f''''''''''''2_r ;
  Go_t \lizzieLet65_3Lcall_f''''''''''''1_d ;
  logic \lizzieLet65_3Lcall_f''''''''''''1_r ;
  Go_t \lizzieLet65_3Lcall_f''''''''''''0_d ;
  logic \lizzieLet65_3Lcall_f''''''''''''0_r ;
  Go_t \lizzieLet65_3Lcall_f''''''''''''0_1_argbuf_d ;
  logic \lizzieLet65_3Lcall_f''''''''''''0_1_argbuf_r ;
  Go_t \lizzieLet65_3Lcall_f''''''''''''1_1_argbuf_d ;
  logic \lizzieLet65_3Lcall_f''''''''''''1_1_argbuf_r ;
  Go_t \lizzieLet65_3Lcall_f''''''''''''2_1_argbuf_d ;
  logic \lizzieLet65_3Lcall_f''''''''''''2_1_argbuf_r ;
  Go_t \lizzieLet65_3Lcall_f''''''''''''3_1_argbuf_d ;
  logic \lizzieLet65_3Lcall_f''''''''''''3_1_argbuf_r ;
  Pointer_QTree_Bool_t \lizzieLet65_4Lf''''''''''''sbos_d ;
  logic \lizzieLet65_4Lf''''''''''''sbos_r ;
  Pointer_QTree_Bool_t \lizzieLet65_4Lcall_f''''''''''''3_d ;
  logic \lizzieLet65_4Lcall_f''''''''''''3_r ;
  Pointer_QTree_Bool_t \lizzieLet65_4Lcall_f''''''''''''2_d ;
  logic \lizzieLet65_4Lcall_f''''''''''''2_r ;
  Pointer_QTree_Bool_t \lizzieLet65_4Lcall_f''''''''''''1_d ;
  logic \lizzieLet65_4Lcall_f''''''''''''1_r ;
  Pointer_QTree_Bool_t \lizzieLet65_4Lcall_f''''''''''''0_d ;
  logic \lizzieLet65_4Lcall_f''''''''''''0_r ;
  QTree_Bool_t \lizzieLet65_4Lcall_f''''''''''''0_1es_1_1_1es_2_2_1es_3_3_1QNode_Bool_d ;
  logic \lizzieLet65_4Lcall_f''''''''''''0_1es_1_1_1es_2_2_1es_3_3_1QNode_Bool_r ;
  QTree_Bool_t lizzieLet69_1_argbuf_d;
  logic lizzieLet69_1_argbuf_r;
  \CTf''''''''''''_t  \lizzieLet65_4Lcall_f''''''''''''1_1es_2_1_1es_3_2_1sc_0_8_1Lcall_f''''''''''''0_d ;
  logic \lizzieLet65_4Lcall_f''''''''''''1_1es_2_1_1es_3_2_1sc_0_8_1Lcall_f''''''''''''0_r ;
  \CTf''''''''''''_t  lizzieLet68_1_argbuf_d;
  logic lizzieLet68_1_argbuf_r;
  \CTf''''''''''''_t  \lizzieLet65_4Lcall_f''''''''''''2_1es_3_1_1sc_0_7_1q1a98_2_1t1a9d_2_1Lcall_f''''''''''''1_d ;
  logic \lizzieLet65_4Lcall_f''''''''''''2_1es_3_1_1sc_0_7_1q1a98_2_1t1a9d_2_1Lcall_f''''''''''''1_r ;
  \CTf''''''''''''_t  lizzieLet67_1_argbuf_d;
  logic lizzieLet67_1_argbuf_r;
  \CTf''''''''''''_t  \lizzieLet65_4Lcall_f''''''''''''3_1sc_0_6_1q1a98_1_1t1a9d_1_1q2a99_1_1t2a9e_1_1Lcall_f''''''''''''2_d ;
  logic \lizzieLet65_4Lcall_f''''''''''''3_1sc_0_6_1q1a98_1_1t1a9d_1_1q2a99_1_1t2a9e_1_1Lcall_f''''''''''''2_r ;
  \CTf''''''''''''_t  lizzieLet66_1_argbuf_d;
  logic lizzieLet66_1_argbuf_r;
  Pointer_QTree_Bool_t \lizzieLet65_4Lf''''''''''''sbos_1_merge_merge_fork_1_d ;
  logic \lizzieLet65_4Lf''''''''''''sbos_1_merge_merge_fork_1_r ;
  Pointer_QTree_Bool_t \lizzieLet65_4Lf''''''''''''sbos_1_merge_merge_fork_2_d ;
  logic \lizzieLet65_4Lf''''''''''''sbos_1_merge_merge_fork_2_r ;
  Go_t \call_f''''''''''''_goConst_d ;
  logic \call_f''''''''''''_goConst_r ;
  C10_t \lvlrf2-0_choice_d ;
  logic \lvlrf2-0_choice_r ;
  TupGo_t \lvlrf2-0_data_d ;
  logic \lvlrf2-0_data_r ;
  MyBool_t go_6_1MyTrue_d;
  logic go_6_1MyTrue_r;
  Pointer_QTree_Bool_t \lvlrf2-0_resbuf_d ;
  logic \lvlrf2-0_resbuf_r ;
  Pointer_QTree_Bool_t \lvlrf2-0_10_argbuf_d ;
  logic \lvlrf2-0_10_argbuf_r ;
  Pointer_QTree_Bool_t lizzieLet27_1_argbuf_d;
  logic lizzieLet27_1_argbuf_r;
  Pointer_QTree_Bool_t \lvlrf2-0_2_argbuf_d ;
  logic \lvlrf2-0_2_argbuf_r ;
  Pointer_QTree_Bool_t lizzieLet5_1_argbuf_d;
  logic lizzieLet5_1_argbuf_r;
  Pointer_QTree_Bool_t \lvlrf2-0_3_argbuf_d ;
  logic \lvlrf2-0_3_argbuf_r ;
  Pointer_QTree_Bool_t lizzieLet48_1_argbuf_d;
  logic lizzieLet48_1_argbuf_r;
  Pointer_QTree_Bool_t \lvlrf2-0_4_argbuf_d ;
  logic \lvlrf2-0_4_argbuf_r ;
  Pointer_QTree_Bool_t lizzieLet49_1_argbuf_d;
  logic lizzieLet49_1_argbuf_r;
  Pointer_QTree_Bool_t \lvlrf2-0_5_argbuf_d ;
  logic \lvlrf2-0_5_argbuf_r ;
  Pointer_QTree_Bool_t lizzieLet16_1_argbuf_d;
  logic lizzieLet16_1_argbuf_r;
  Pointer_QTree_Bool_t \lvlrf2-0_6_argbuf_d ;
  logic \lvlrf2-0_6_argbuf_r ;
  Pointer_QTree_Bool_t lizzieLet17_1_argbuf_d;
  logic lizzieLet17_1_argbuf_r;
  Pointer_QTree_Bool_t \lvlrf2-0_7_argbuf_d ;
  logic \lvlrf2-0_7_argbuf_r ;
  Pointer_QTree_Bool_t lizzieLet21_1_argbuf_d;
  logic lizzieLet21_1_argbuf_r;
  Pointer_QTree_Bool_t \lvlrf2-0_8_argbuf_d ;
  logic \lvlrf2-0_8_argbuf_r ;
  Pointer_QTree_Bool_t lizzieLet22_1_argbuf_d;
  logic lizzieLet22_1_argbuf_r;
  Pointer_QTree_Bool_t \lvlrf2-0_9_argbuf_d ;
  logic \lvlrf2-0_9_argbuf_r ;
  Pointer_QTree_Bool_t lizzieLet26_1_argbuf_d;
  logic lizzieLet26_1_argbuf_r;
  Pointer_QTree_Bool_t \lvlrf2-0_1_d ;
  logic \lvlrf2-0_1_r ;
  Pointer_QTree_Bool_t \lvlrf2-0_2_d ;
  logic \lvlrf2-0_2_r ;
  Pointer_QTree_Bool_t \lvlrf2-0_3_d ;
  logic \lvlrf2-0_3_r ;
  Pointer_QTree_Bool_t \lvlrf2-0_4_d ;
  logic \lvlrf2-0_4_r ;
  Pointer_QTree_Bool_t \lvlrf2-0_5_d ;
  logic \lvlrf2-0_5_r ;
  Pointer_QTree_Bool_t \lvlrf2-0_6_d ;
  logic \lvlrf2-0_6_r ;
  Pointer_QTree_Bool_t \lvlrf2-0_7_d ;
  logic \lvlrf2-0_7_r ;
  Pointer_QTree_Bool_t \lvlrf2-0_8_d ;
  logic \lvlrf2-0_8_r ;
  Pointer_QTree_Bool_t \lvlrf2-0_9_d ;
  logic \lvlrf2-0_9_r ;
  Pointer_QTree_Bool_t \lvlrf2-0_10_d ;
  logic \lvlrf2-0_10_r ;
  Go_t \lvlrf2-0TupGogo_6_d ;
  logic \lvlrf2-0TupGogo_6_r ;
  Pointer_QTree_Bool_t lizzieLet4_1_argbuf_d;
  logic lizzieLet4_1_argbuf_r;
  Pointer_QTree_Bool_t m1a84_1_argbuf_d;
  logic m1a84_1_argbuf_r;
  Pointer_QTree_Bool_t m1a84_1_d;
  logic m1a84_1_r;
  Pointer_QTree_Bool_t m1a84_2_d;
  logic m1a84_2_r;
  Pointer_QTree_Bool_t m2a85_1_argbuf_d;
  logic m2a85_1_argbuf_r;
  Pointer_QTree_Bool_t m2a85_1_d;
  logic m2a85_1_r;
  Pointer_QTree_Bool_t m2a85_2_d;
  logic m2a85_2_r;
  Pointer_QTree_Bool_t m3a86_1_argbuf_d;
  logic m3a86_1_argbuf_r;
  Pointer_QTree_Bool_t m3a86_1_d;
  logic m3a86_1_r;
  Pointer_QTree_Bool_t m3a86_2_d;
  logic m3a86_2_r;
  Pointer_QTree_Bool_t q1a8H_3_1_argbuf_d;
  logic q1a8H_3_1_argbuf_r;
  Pointer_QTree_Bool_t q1a98_3_1_argbuf_d;
  logic q1a98_3_1_argbuf_r;
  Pointer_QTree_Bool_t q2a8I_2_1_argbuf_d;
  logic q2a8I_2_1_argbuf_r;
  Pointer_QTree_Bool_t q2a99_2_1_argbuf_d;
  logic q2a99_2_1_argbuf_r;
  Pointer_QTree_Bool_t q3a8J_1_1_argbuf_d;
  logic q3a8J_1_1_argbuf_r;
  Pointer_QTree_Bool_t q3a9a_1_1_argbuf_d;
  logic q3a9a_1_1_argbuf_r;
  Pointer_QTree_Bool_t q4a90_1_argbuf_d;
  logic q4a90_1_argbuf_r;
  Pointer_QTree_Bool_t q4a90_1_d;
  logic q4a90_1_r;
  Pointer_QTree_Bool_t q4a90_2_d;
  logic q4a90_2_r;
  \CTf''''''''''''_t  \readPointer_CTf''''''''''''scfarg_0_1_1_argbuf_rwb_d ;
  logic \readPointer_CTf''''''''''''scfarg_0_1_1_argbuf_rwb_r ;
  \CTf''''''''''''_t  lizzieLet65_1_d;
  logic lizzieLet65_1_r;
  \CTf''''''''''''_t  lizzieLet65_2_d;
  logic lizzieLet65_2_r;
  \CTf''''''''''''_t  lizzieLet65_3_d;
  logic lizzieLet65_3_r;
  \CTf''''''''''''_t  lizzieLet65_4_d;
  logic lizzieLet65_4_r;
  CTf_t readPointer_CTfscfarg_0_1_argbuf_rwb_d;
  logic readPointer_CTfscfarg_0_1_argbuf_rwb_r;
  CTf_t lizzieLet60_1_d;
  logic lizzieLet60_1_r;
  CTf_t lizzieLet60_2_d;
  logic lizzieLet60_2_r;
  CTf_t lizzieLet60_3_d;
  logic lizzieLet60_3_r;
  CTf_t lizzieLet60_4_d;
  logic lizzieLet60_4_r;
  QTree_Bool_t readPointer_QTree_Boolm1a84_1_argbuf_rwb_d;
  logic readPointer_QTree_Boolm1a84_1_argbuf_rwb_r;
  QTree_Bool_t lizzieLet0_1_d;
  logic lizzieLet0_1_r;
  QTree_Bool_t lizzieLet0_2_d;
  logic lizzieLet0_2_r;
  QTree_Bool_t lizzieLet0_3_d;
  logic lizzieLet0_3_r;
  QTree_Bool_t lizzieLet0_4_d;
  logic lizzieLet0_4_r;
  QTree_Bool_t lizzieLet0_5_d;
  logic lizzieLet0_5_r;
  QTree_Bool_t lizzieLet0_6_d;
  logic lizzieLet0_6_r;
  QTree_Bool_t lizzieLet0_7_d;
  logic lizzieLet0_7_r;
  QTree_Bool_t lizzieLet0_8_d;
  logic lizzieLet0_8_r;
  QTree_Bool_t lizzieLet0_9_d;
  logic lizzieLet0_9_r;
  QTree_Bool_t readPointer_QTree_Boolm2a85_1_argbuf_rwb_d;
  logic readPointer_QTree_Boolm2a85_1_argbuf_rwb_r;
  QTree_Bool_t readPointer_QTree_Boolm3a86_1_argbuf_rwb_d;
  logic readPointer_QTree_Boolm3a86_1_argbuf_rwb_r;
  QTree_Bool_t readPointer_QTree_Boolq4a90_1_argbuf_rwb_d;
  logic readPointer_QTree_Boolq4a90_1_argbuf_rwb_r;
  QTree_Bool_t lizzieLet45_1_d;
  logic lizzieLet45_1_r;
  QTree_Bool_t lizzieLet45_2_d;
  logic lizzieLet45_2_r;
  QTree_Bool_t lizzieLet45_3_d;
  logic lizzieLet45_3_r;
  QTree_Bool_t lizzieLet45_4_d;
  logic lizzieLet45_4_r;
  QTree_Bool_t lizzieLet45_5_d;
  logic lizzieLet45_5_r;
  QTree_Bool_t lizzieLet45_6_d;
  logic lizzieLet45_6_r;
  QTree_Bool_t lizzieLet45_7_d;
  logic lizzieLet45_7_r;
  QTree_Bool_t readPointer_QTree_Boolt4a91_1_argbuf_rwb_d;
  logic readPointer_QTree_Boolt4a91_1_argbuf_rwb_r;
  Pointer_CTf_t sc_0_5_1_argbuf_d;
  logic sc_0_5_1_argbuf_r;
  \Pointer_CTf''''''''''''_t  sc_0_9_1_argbuf_d;
  logic sc_0_9_1_argbuf_r;
  \Pointer_CTf''''''''''''_t  scfarg_0_1_1_argbuf_d;
  logic scfarg_0_1_1_argbuf_r;
  Pointer_CTf_t scfarg_0_1_argbuf_d;
  logic scfarg_0_1_argbuf_r;
  Pointer_QTree_Bool_t \t1'a8W_3_1_argbuf_d ;
  logic \t1'a8W_3_1_argbuf_r ;
  Pointer_QTree_Bool_t t1a8M_1_argbuf_d;
  logic t1a8M_1_argbuf_r;
  Pointer_QTree_Bool_t t1a8R_3_1_argbuf_d;
  logic t1a8R_3_1_argbuf_r;
  Pointer_QTree_Bool_t t1a8i_1_argbuf_d;
  logic t1a8i_1_argbuf_r;
  Pointer_QTree_Bool_t t1a9d_3_1_argbuf_d;
  logic t1a9d_3_1_argbuf_r;
  Pointer_QTree_Bool_t \t2'a8X_2_1_argbuf_d ;
  logic \t2'a8X_2_1_argbuf_r ;
  Pointer_QTree_Bool_t t2a8N_1_argbuf_d;
  logic t2a8N_1_argbuf_r;
  Pointer_QTree_Bool_t t2a8S_2_1_argbuf_d;
  logic t2a8S_2_1_argbuf_r;
  Pointer_QTree_Bool_t t2a8j_1_argbuf_d;
  logic t2a8j_1_argbuf_r;
  Pointer_QTree_Bool_t t2a9e_2_1_argbuf_d;
  logic t2a9e_2_1_argbuf_r;
  Pointer_QTree_Bool_t \t3'a8Y_1_1_argbuf_d ;
  logic \t3'a8Y_1_1_argbuf_r ;
  Pointer_QTree_Bool_t t3a8O_1_argbuf_d;
  logic t3a8O_1_argbuf_r;
  Pointer_QTree_Bool_t t3a8T_1_1_argbuf_d;
  logic t3a8T_1_1_argbuf_r;
  Pointer_QTree_Bool_t t3a8k_1_argbuf_d;
  logic t3a8k_1_argbuf_r;
  Pointer_QTree_Bool_t t3a9f_1_1_argbuf_d;
  logic t3a9f_1_1_argbuf_r;
  Pointer_QTree_Bool_t \t4'a8Z_1_argbuf_d ;
  logic \t4'a8Z_1_argbuf_r ;
  Pointer_QTree_Bool_t t4a8P_1_argbuf_d;
  logic t4a8P_1_argbuf_r;
  Pointer_QTree_Bool_t t4a8l_1_argbuf_d;
  logic t4a8l_1_argbuf_r;
  Pointer_QTree_Bool_t t4a91_1_argbuf_d;
  logic t4a91_1_argbuf_r;
  Pointer_QTree_Bool_t t4a91_1_d;
  logic t4a91_1_r;
  Pointer_QTree_Bool_t t4a91_2_d;
  logic t4a91_2_r;
  Pointer_QTree_Bool_t t5a9g_1_argbuf_d;
  logic t5a9g_1_argbuf_r;
  \Pointer_CTf''''''''''''_t  \writeCTf''''''''''''lizzieLet54_1_argbuf_rwb_d ;
  logic \writeCTf''''''''''''lizzieLet54_1_argbuf_rwb_r ;
  \Pointer_CTf''''''''''''_t  sca3_1_1_argbuf_d;
  logic sca3_1_1_argbuf_r;
  \Pointer_CTf''''''''''''_t  \writeCTf''''''''''''lizzieLet58_1_argbuf_rwb_d ;
  logic \writeCTf''''''''''''lizzieLet58_1_argbuf_rwb_r ;
  \Pointer_CTf''''''''''''_t  lizzieLet7_1_1_argbuf_d;
  logic lizzieLet7_1_1_argbuf_r;
  \Pointer_CTf''''''''''''_t  \writeCTf''''''''''''lizzieLet66_1_argbuf_rwb_d ;
  logic \writeCTf''''''''''''lizzieLet66_1_argbuf_rwb_r ;
  \Pointer_CTf''''''''''''_t  sca2_1_1_argbuf_d;
  logic sca2_1_1_argbuf_r;
  \Pointer_CTf''''''''''''_t  \writeCTf''''''''''''lizzieLet67_1_argbuf_rwb_d ;
  logic \writeCTf''''''''''''lizzieLet67_1_argbuf_rwb_r ;
  \Pointer_CTf''''''''''''_t  sca1_1_1_argbuf_d;
  logic sca1_1_1_argbuf_r;
  \Pointer_CTf''''''''''''_t  \writeCTf''''''''''''lizzieLet68_1_argbuf_rwb_d ;
  logic \writeCTf''''''''''''lizzieLet68_1_argbuf_rwb_r ;
  \Pointer_CTf''''''''''''_t  sca0_1_1_argbuf_d;
  logic sca0_1_1_argbuf_r;
  Pointer_CTf_t writeCTflizzieLet41_1_argbuf_rwb_d;
  logic writeCTflizzieLet41_1_argbuf_rwb_r;
  Pointer_CTf_t sca3_1_argbuf_d;
  logic sca3_1_argbuf_r;
  Pointer_CTf_t writeCTflizzieLet57_1_argbuf_rwb_d;
  logic writeCTflizzieLet57_1_argbuf_rwb_r;
  Pointer_CTf_t lizzieLet33_1_argbuf_d;
  logic lizzieLet33_1_argbuf_r;
  Pointer_CTf_t writeCTflizzieLet61_1_argbuf_rwb_d;
  logic writeCTflizzieLet61_1_argbuf_rwb_r;
  Pointer_CTf_t sca2_1_argbuf_d;
  logic sca2_1_argbuf_r;
  Pointer_CTf_t writeCTflizzieLet62_1_argbuf_rwb_d;
  logic writeCTflizzieLet62_1_argbuf_rwb_r;
  Pointer_CTf_t sca1_1_argbuf_d;
  logic sca1_1_argbuf_r;
  Pointer_CTf_t writeCTflizzieLet63_1_argbuf_rwb_d;
  logic writeCTflizzieLet63_1_argbuf_rwb_r;
  Pointer_CTf_t sca0_1_argbuf_d;
  logic sca0_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet10_1_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet10_1_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t lizzieLet12_1_argbuf_d;
  logic lizzieLet12_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet11_1_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet11_1_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t lizzieLet13_1_argbuf_d;
  logic lizzieLet13_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet12_1_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet12_1_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t lizzieLet14_1_argbuf_d;
  logic lizzieLet14_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet15_1_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet15_1_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t lizzieLet15_1_argbuf_d;
  logic lizzieLet15_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet18_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet18_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t lizzieLet16_1_1_argbuf_d;
  logic lizzieLet16_1_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet19_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet19_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t lizzieLet17_1_1_argbuf_d;
  logic lizzieLet17_1_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet23_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet23_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t lizzieLet18_1_1_argbuf_d;
  logic lizzieLet18_1_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet24_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet24_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t lizzieLet19_1_1_argbuf_d;
  logic lizzieLet19_1_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet28_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet28_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t lizzieLet20_1_argbuf_d;
  logic lizzieLet20_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet29_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet29_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t lizzieLet21_1_1_argbuf_d;
  logic lizzieLet21_1_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet30_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet30_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t lizzieLet22_1_1_argbuf_d;
  logic lizzieLet22_1_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet31_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet31_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t lizzieLet23_1_1_argbuf_d;
  logic lizzieLet23_1_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet34_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet34_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t lizzieLet24_1_1_argbuf_d;
  logic lizzieLet24_1_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet35_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet35_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t lizzieLet25_1_argbuf_d;
  logic lizzieLet25_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet36_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet36_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t lizzieLet26_1_1_argbuf_d;
  logic lizzieLet26_1_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet37_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet37_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t lizzieLet27_1_1_argbuf_d;
  logic lizzieLet27_1_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet39_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet39_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t lizzieLet28_1_1_argbuf_d;
  logic lizzieLet28_1_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet3_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet3_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t lizzieLet8_1_argbuf_d;
  logic lizzieLet8_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet40_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet40_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t lizzieLet29_1_1_argbuf_d;
  logic lizzieLet29_1_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet42_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet42_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t lizzieLet30_1_1_argbuf_d;
  logic lizzieLet30_1_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet43_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet43_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t lizzieLet31_1_1_argbuf_d;
  logic lizzieLet31_1_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet44_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet44_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t lizzieLet32_1_argbuf_d;
  logic lizzieLet32_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet47_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet47_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t lizzieLet1_1_1_argbuf_d;
  logic lizzieLet1_1_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet50_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet50_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t lizzieLet2_1_1_argbuf_d;
  logic lizzieLet2_1_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet51_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet51_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t lizzieLet3_1_1_argbuf_d;
  logic lizzieLet3_1_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet53_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet53_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t lizzieLet4_1_1_argbuf_d;
  logic lizzieLet4_1_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet55_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet55_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t lizzieLet5_1_1_argbuf_d;
  logic lizzieLet5_1_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet56_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet56_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t lizzieLet6_1_1_argbuf_d;
  logic lizzieLet6_1_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet59_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet59_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet64_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet64_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t contRet_0_1_argbuf_d;
  logic contRet_0_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet69_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet69_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t contRet_0_1_1_argbuf_d;
  logic contRet_0_1_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet6_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet6_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t lizzieLet9_1_argbuf_d;
  logic lizzieLet9_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet7_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet7_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t lizzieLet10_1_argbuf_d;
  logic lizzieLet10_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet9_1_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet9_1_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t lizzieLet11_1_argbuf_d;
  logic lizzieLet11_1_argbuf_r;
  
  /* fork (Ty Go) : (sourceGo,Go) > [(goFork,Go),
                                (goFor_2,Go),
                                (goFor_3,Go),
                                (goFor_4,Go),
                                (goFor_5,Go)] */
  logic [4:0] sourceGo_emitted;
  logic [4:0] sourceGo_done;
  assign goFork_d = (sourceGo_d[0] && (! sourceGo_emitted[0]));
  assign goFor_2_d = (sourceGo_d[0] && (! sourceGo_emitted[1]));
  assign goFor_3_d = (sourceGo_d[0] && (! sourceGo_emitted[2]));
  assign goFor_4_d = (sourceGo_d[0] && (! sourceGo_emitted[3]));
  assign goFor_5_d = (sourceGo_d[0] && (! sourceGo_emitted[4]));
  assign sourceGo_done = (sourceGo_emitted | ({goFor_5_d[0],
                                               goFor_4_d[0],
                                               goFor_3_d[0],
                                               goFor_2_d[0],
                                               goFork_d[0]} & {goFor_5_r,
                                                               goFor_4_r,
                                                               goFor_3_r,
                                                               goFor_2_r,
                                                               goFork_r}));
  assign sourceGo_r = (& sourceGo_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) sourceGo_emitted <= 5'd0;
    else
      sourceGo_emitted <= (sourceGo_r ? 5'd0 :
                           sourceGo_done);
  
  /* const (Ty Word16#,
       Lit 0) : (go_1_dummy_write_QTree_Bool,Go) > (initHP_QTree_Bool,Word16#) */
  assign initHP_QTree_Bool_d = {16'd0,
                                go_1_dummy_write_QTree_Bool_d[0]};
  assign go_1_dummy_write_QTree_Bool_r = initHP_QTree_Bool_r;
  
  /* const (Ty Word16#,
       Lit 1) : (incrHP_QTree_Bool1,Go) > (incrHP_QTree_Bool,Word16#) */
  assign incrHP_QTree_Bool_d = {16'd1, incrHP_QTree_Bool1_d[0]};
  assign incrHP_QTree_Bool1_r = incrHP_QTree_Bool_r;
  
  /* merge (Ty Go) : [(go_2_dummy_write_QTree_Bool,Go),
                 (incrHP_QTree_Bool2,Go)] > (incrHP_mergeQTree_Bool,Go) */
  logic [1:0] incrHP_mergeQTree_Bool_selected;
  logic [1:0] incrHP_mergeQTree_Bool_select;
  always_comb
    begin
      incrHP_mergeQTree_Bool_selected = 2'd0;
      if ((| incrHP_mergeQTree_Bool_select))
        incrHP_mergeQTree_Bool_selected = incrHP_mergeQTree_Bool_select;
      else
        if (go_2_dummy_write_QTree_Bool_d[0])
          incrHP_mergeQTree_Bool_selected[0] = 1'd1;
        else if (incrHP_QTree_Bool2_d[0])
          incrHP_mergeQTree_Bool_selected[1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeQTree_Bool_select <= 2'd0;
    else
      incrHP_mergeQTree_Bool_select <= (incrHP_mergeQTree_Bool_r ? 2'd0 :
                                        incrHP_mergeQTree_Bool_selected);
  always_comb
    if (incrHP_mergeQTree_Bool_selected[0])
      incrHP_mergeQTree_Bool_d = go_2_dummy_write_QTree_Bool_d;
    else if (incrHP_mergeQTree_Bool_selected[1])
      incrHP_mergeQTree_Bool_d = incrHP_QTree_Bool2_d;
    else incrHP_mergeQTree_Bool_d = 1'd0;
  assign {incrHP_QTree_Bool2_r,
          go_2_dummy_write_QTree_Bool_r} = (incrHP_mergeQTree_Bool_r ? incrHP_mergeQTree_Bool_selected :
                                            2'd0);
  
  /* fork (Ty Go) : (incrHP_mergeQTree_Bool_buf,Go) > [(incrHP_QTree_Bool1,Go),
                                                  (incrHP_QTree_Bool2,Go)] */
  logic [1:0] incrHP_mergeQTree_Bool_buf_emitted;
  logic [1:0] incrHP_mergeQTree_Bool_buf_done;
  assign incrHP_QTree_Bool1_d = (incrHP_mergeQTree_Bool_buf_d[0] && (! incrHP_mergeQTree_Bool_buf_emitted[0]));
  assign incrHP_QTree_Bool2_d = (incrHP_mergeQTree_Bool_buf_d[0] && (! incrHP_mergeQTree_Bool_buf_emitted[1]));
  assign incrHP_mergeQTree_Bool_buf_done = (incrHP_mergeQTree_Bool_buf_emitted | ({incrHP_QTree_Bool2_d[0],
                                                                                   incrHP_QTree_Bool1_d[0]} & {incrHP_QTree_Bool2_r,
                                                                                                               incrHP_QTree_Bool1_r}));
  assign incrHP_mergeQTree_Bool_buf_r = (& incrHP_mergeQTree_Bool_buf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeQTree_Bool_buf_emitted <= 2'd0;
    else
      incrHP_mergeQTree_Bool_buf_emitted <= (incrHP_mergeQTree_Bool_buf_r ? 2'd0 :
                                             incrHP_mergeQTree_Bool_buf_done);
  
  /* op_add (Ty Word16#) : (incrHP_QTree_Bool,Word16#) (forkHP1_QTree_Bool,Word16#) > (addHP_QTree_Bool,Word16#) */
  assign addHP_QTree_Bool_d = {(incrHP_QTree_Bool_d[16:1] + forkHP1_QTree_Bool_d[16:1]),
                               (incrHP_QTree_Bool_d[0] && forkHP1_QTree_Bool_d[0])};
  assign {incrHP_QTree_Bool_r,
          forkHP1_QTree_Bool_r} = {2 {(addHP_QTree_Bool_r && addHP_QTree_Bool_d[0])}};
  
  /* merge (Ty Word16#) : [(initHP_QTree_Bool,Word16#),
                      (addHP_QTree_Bool,Word16#)] > (mergeHP_QTree_Bool,Word16#) */
  logic [1:0] mergeHP_QTree_Bool_selected;
  logic [1:0] mergeHP_QTree_Bool_select;
  always_comb
    begin
      mergeHP_QTree_Bool_selected = 2'd0;
      if ((| mergeHP_QTree_Bool_select))
        mergeHP_QTree_Bool_selected = mergeHP_QTree_Bool_select;
      else
        if (initHP_QTree_Bool_d[0]) mergeHP_QTree_Bool_selected[0] = 1'd1;
        else if (addHP_QTree_Bool_d[0])
          mergeHP_QTree_Bool_selected[1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_QTree_Bool_select <= 2'd0;
    else
      mergeHP_QTree_Bool_select <= (mergeHP_QTree_Bool_r ? 2'd0 :
                                    mergeHP_QTree_Bool_selected);
  always_comb
    if (mergeHP_QTree_Bool_selected[0])
      mergeHP_QTree_Bool_d = initHP_QTree_Bool_d;
    else if (mergeHP_QTree_Bool_selected[1])
      mergeHP_QTree_Bool_d = addHP_QTree_Bool_d;
    else mergeHP_QTree_Bool_d = {16'd0, 1'd0};
  assign {addHP_QTree_Bool_r,
          initHP_QTree_Bool_r} = (mergeHP_QTree_Bool_r ? mergeHP_QTree_Bool_selected :
                                  2'd0);
  
  /* buf (Ty Go) : (incrHP_mergeQTree_Bool,Go) > (incrHP_mergeQTree_Bool_buf,Go) */
  Go_t incrHP_mergeQTree_Bool_bufchan_d;
  logic incrHP_mergeQTree_Bool_bufchan_r;
  assign incrHP_mergeQTree_Bool_r = ((! incrHP_mergeQTree_Bool_bufchan_d[0]) || incrHP_mergeQTree_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeQTree_Bool_bufchan_d <= 1'd0;
    else
      if (incrHP_mergeQTree_Bool_r)
        incrHP_mergeQTree_Bool_bufchan_d <= incrHP_mergeQTree_Bool_d;
  Go_t incrHP_mergeQTree_Bool_bufchan_buf;
  assign incrHP_mergeQTree_Bool_bufchan_r = (! incrHP_mergeQTree_Bool_bufchan_buf[0]);
  assign incrHP_mergeQTree_Bool_buf_d = (incrHP_mergeQTree_Bool_bufchan_buf[0] ? incrHP_mergeQTree_Bool_bufchan_buf :
                                         incrHP_mergeQTree_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeQTree_Bool_bufchan_buf <= 1'd0;
    else
      if ((incrHP_mergeQTree_Bool_buf_r && incrHP_mergeQTree_Bool_bufchan_buf[0]))
        incrHP_mergeQTree_Bool_bufchan_buf <= 1'd0;
      else if (((! incrHP_mergeQTree_Bool_buf_r) && (! incrHP_mergeQTree_Bool_bufchan_buf[0])))
        incrHP_mergeQTree_Bool_bufchan_buf <= incrHP_mergeQTree_Bool_bufchan_d;
  
  /* buf (Ty Word16#) : (mergeHP_QTree_Bool,Word16#) > (mergeHP_QTree_Bool_buf,Word16#) */
  \Word16#_t  mergeHP_QTree_Bool_bufchan_d;
  logic mergeHP_QTree_Bool_bufchan_r;
  assign mergeHP_QTree_Bool_r = ((! mergeHP_QTree_Bool_bufchan_d[0]) || mergeHP_QTree_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_QTree_Bool_bufchan_d <= {16'd0, 1'd0};
    else
      if (mergeHP_QTree_Bool_r)
        mergeHP_QTree_Bool_bufchan_d <= mergeHP_QTree_Bool_d;
  \Word16#_t  mergeHP_QTree_Bool_bufchan_buf;
  assign mergeHP_QTree_Bool_bufchan_r = (! mergeHP_QTree_Bool_bufchan_buf[0]);
  assign mergeHP_QTree_Bool_buf_d = (mergeHP_QTree_Bool_bufchan_buf[0] ? mergeHP_QTree_Bool_bufchan_buf :
                                     mergeHP_QTree_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      mergeHP_QTree_Bool_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((mergeHP_QTree_Bool_buf_r && mergeHP_QTree_Bool_bufchan_buf[0]))
        mergeHP_QTree_Bool_bufchan_buf <= {16'd0, 1'd0};
      else if (((! mergeHP_QTree_Bool_buf_r) && (! mergeHP_QTree_Bool_bufchan_buf[0])))
        mergeHP_QTree_Bool_bufchan_buf <= mergeHP_QTree_Bool_bufchan_d;
  
  /* sink (Ty Word16#) : (forkHP1_QTree_Bool_snk,Word16#) > */
  assign {forkHP1_QTree_Bool_snk_r,
          forkHP1_QTree_Bool_snk_dout} = {forkHP1_QTree_Bool_snk_rout,
                                          forkHP1_QTree_Bool_snk_d};
  
  /* source (Ty Go) : > (\QTree_Bool_src,Go) */
  
  /* fork (Ty Go) : (\QTree_Bool_src,Go) > [(go_1_dummy_write_QTree_Bool,Go),
                                       (go_2_dummy_write_QTree_Bool,Go)] */
  logic [1:0] \\QTree_Bool_src_emitted ;
  logic [1:0] \\QTree_Bool_src_done ;
  assign go_1_dummy_write_QTree_Bool_d = (\\QTree_Bool_src_d [0] && (! \\QTree_Bool_src_emitted [0]));
  assign go_2_dummy_write_QTree_Bool_d = (\\QTree_Bool_src_d [0] && (! \\QTree_Bool_src_emitted [1]));
  assign \\QTree_Bool_src_done  = (\\QTree_Bool_src_emitted  | ({go_2_dummy_write_QTree_Bool_d[0],
                                                                 go_1_dummy_write_QTree_Bool_d[0]} & {go_2_dummy_write_QTree_Bool_r,
                                                                                                      go_1_dummy_write_QTree_Bool_r}));
  assign \\QTree_Bool_src_r  = (& \\QTree_Bool_src_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \\QTree_Bool_src_emitted  <= 2'd0;
    else
      \\QTree_Bool_src_emitted  <= (\\QTree_Bool_src_r  ? 2'd0 :
                                    \\QTree_Bool_src_done );
  
  /* source (Ty QTree_Bool) : > (dummy_write_QTree_Bool,QTree_Bool) */
  
  /* sink (Ty Pointer_QTree_Bool) : (dummy_write_QTree_Bool_sink,Pointer_QTree_Bool) > */
  assign {dummy_write_QTree_Bool_sink_r,
          dummy_write_QTree_Bool_sink_dout} = {dummy_write_QTree_Bool_sink_rout,
                                               dummy_write_QTree_Bool_sink_d};
  
  /* fork (Ty Word16#) : (mergeHP_QTree_Bool_buf,Word16#) > [(forkHP1_QTree_Bool,Word16#),
                                                        (forkHP1_QTree_Bool_snk,Word16#),
                                                        (forkHP1_QTree_Boo3,Word16#),
                                                        (forkHP1_QTree_Boo4,Word16#)] */
  logic [3:0] mergeHP_QTree_Bool_buf_emitted;
  logic [3:0] mergeHP_QTree_Bool_buf_done;
  assign forkHP1_QTree_Bool_d = {mergeHP_QTree_Bool_buf_d[16:1],
                                 (mergeHP_QTree_Bool_buf_d[0] && (! mergeHP_QTree_Bool_buf_emitted[0]))};
  assign forkHP1_QTree_Bool_snk_d = {mergeHP_QTree_Bool_buf_d[16:1],
                                     (mergeHP_QTree_Bool_buf_d[0] && (! mergeHP_QTree_Bool_buf_emitted[1]))};
  assign forkHP1_QTree_Boo3_d = {mergeHP_QTree_Bool_buf_d[16:1],
                                 (mergeHP_QTree_Bool_buf_d[0] && (! mergeHP_QTree_Bool_buf_emitted[2]))};
  assign forkHP1_QTree_Boo4_d = {mergeHP_QTree_Bool_buf_d[16:1],
                                 (mergeHP_QTree_Bool_buf_d[0] && (! mergeHP_QTree_Bool_buf_emitted[3]))};
  assign mergeHP_QTree_Bool_buf_done = (mergeHP_QTree_Bool_buf_emitted | ({forkHP1_QTree_Boo4_d[0],
                                                                           forkHP1_QTree_Boo3_d[0],
                                                                           forkHP1_QTree_Bool_snk_d[0],
                                                                           forkHP1_QTree_Bool_d[0]} & {forkHP1_QTree_Boo4_r,
                                                                                                       forkHP1_QTree_Boo3_r,
                                                                                                       forkHP1_QTree_Bool_snk_r,
                                                                                                       forkHP1_QTree_Bool_r}));
  assign mergeHP_QTree_Bool_buf_r = (& mergeHP_QTree_Bool_buf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_QTree_Bool_buf_emitted <= 4'd0;
    else
      mergeHP_QTree_Bool_buf_emitted <= (mergeHP_QTree_Bool_buf_r ? 4'd0 :
                                         mergeHP_QTree_Bool_buf_done);
  
  /* mergectrl (Ty C2,
           Ty MemIn_QTree_Bool) : [(dconReadIn_QTree_Bool,MemIn_QTree_Bool),
                                   (dconWriteIn_QTree_Bool,MemIn_QTree_Bool)] > (memMergeChoice_QTree_Bool,C2) (memMergeIn_QTree_Bool,MemIn_QTree_Bool) */
  logic [1:0] dconReadIn_QTree_Bool_select_d;
  assign dconReadIn_QTree_Bool_select_d = ((| dconReadIn_QTree_Bool_select_q) ? dconReadIn_QTree_Bool_select_q :
                                           (dconReadIn_QTree_Bool_d[0] ? 2'd1 :
                                            (dconWriteIn_QTree_Bool_d[0] ? 2'd2 :
                                             2'd0)));
  logic [1:0] dconReadIn_QTree_Bool_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) dconReadIn_QTree_Bool_select_q <= 2'd0;
    else
      dconReadIn_QTree_Bool_select_q <= (dconReadIn_QTree_Bool_done ? 2'd0 :
                                         dconReadIn_QTree_Bool_select_d);
  logic [1:0] dconReadIn_QTree_Bool_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) dconReadIn_QTree_Bool_emit_q <= 2'd0;
    else
      dconReadIn_QTree_Bool_emit_q <= (dconReadIn_QTree_Bool_done ? 2'd0 :
                                       dconReadIn_QTree_Bool_emit_d);
  logic [1:0] dconReadIn_QTree_Bool_emit_d;
  assign dconReadIn_QTree_Bool_emit_d = (dconReadIn_QTree_Bool_emit_q | ({memMergeChoice_QTree_Bool_d[0],
                                                                          memMergeIn_QTree_Bool_d[0]} & {memMergeChoice_QTree_Bool_r,
                                                                                                         memMergeIn_QTree_Bool_r}));
  logic dconReadIn_QTree_Bool_done;
  assign dconReadIn_QTree_Bool_done = (& dconReadIn_QTree_Bool_emit_d);
  assign {dconWriteIn_QTree_Bool_r,
          dconReadIn_QTree_Bool_r} = (dconReadIn_QTree_Bool_done ? dconReadIn_QTree_Bool_select_d :
                                      2'd0);
  assign memMergeIn_QTree_Bool_d = ((dconReadIn_QTree_Bool_select_d[0] && (! dconReadIn_QTree_Bool_emit_q[0])) ? dconReadIn_QTree_Bool_d :
                                    ((dconReadIn_QTree_Bool_select_d[1] && (! dconReadIn_QTree_Bool_emit_q[0])) ? dconWriteIn_QTree_Bool_d :
                                     {83'd0, 1'd0}));
  assign memMergeChoice_QTree_Bool_d = ((dconReadIn_QTree_Bool_select_d[0] && (! dconReadIn_QTree_Bool_emit_q[1])) ? C1_2_dc(1'd1) :
                                        ((dconReadIn_QTree_Bool_select_d[1] && (! dconReadIn_QTree_Bool_emit_q[1])) ? C2_2_dc(1'd1) :
                                         {1'd0, 1'd0}));
  
  /* bram (Ty MemIn_QTree_Bool,
      Ty MemOut_QTree_Bool) : (memMergeIn_QTree_Bool_dbuf,MemIn_QTree_Bool) > (memOut_QTree_Bool,MemOut_QTree_Bool) */
  logic [65:0] memMergeIn_QTree_Bool_dbuf_mem[65535:0];
  logic [15:0] memMergeIn_QTree_Bool_dbuf_address;
  logic [65:0] memMergeIn_QTree_Bool_dbuf_din;
  logic [65:0] memOut_QTree_Bool_q;
  logic memOut_QTree_Bool_valid;
  logic memMergeIn_QTree_Bool_dbuf_we;
  logic memOut_QTree_Bool_we;
  assign memMergeIn_QTree_Bool_dbuf_din = memMergeIn_QTree_Bool_dbuf_d[83:18];
  assign memMergeIn_QTree_Bool_dbuf_address = memMergeIn_QTree_Bool_dbuf_d[17:2];
  assign memMergeIn_QTree_Bool_dbuf_we = (memMergeIn_QTree_Bool_dbuf_d[1:1] && memMergeIn_QTree_Bool_dbuf_d[0]);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        memOut_QTree_Bool_we <= 1'd0;
        memOut_QTree_Bool_valid <= 1'd0;
      end
    else
      begin
        memOut_QTree_Bool_we <= memMergeIn_QTree_Bool_dbuf_we;
        memOut_QTree_Bool_valid <= memMergeIn_QTree_Bool_dbuf_d[0];
        if (memMergeIn_QTree_Bool_dbuf_we)
          begin
            memMergeIn_QTree_Bool_dbuf_mem[memMergeIn_QTree_Bool_dbuf_address] <= memMergeIn_QTree_Bool_dbuf_din;
            memOut_QTree_Bool_q <= memMergeIn_QTree_Bool_dbuf_din;
          end
        else
          memOut_QTree_Bool_q <= memMergeIn_QTree_Bool_dbuf_mem[memMergeIn_QTree_Bool_dbuf_address];
      end
  assign memOut_QTree_Bool_d = {memOut_QTree_Bool_q,
                                memOut_QTree_Bool_we,
                                memOut_QTree_Bool_valid};
  assign memMergeIn_QTree_Bool_dbuf_r = ((! memOut_QTree_Bool_valid) || memOut_QTree_Bool_r);
  logic [31:0] profiling_MemIn_QTree_Bool_read;
  logic [31:0] profiling_MemIn_QTree_Bool_write;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        profiling_MemIn_QTree_Bool_write <= 0;
        profiling_MemIn_QTree_Bool_read <= 0;
      end
    else
      if ((memMergeIn_QTree_Bool_dbuf_we == 1'd1))
        profiling_MemIn_QTree_Bool_write <= (profiling_MemIn_QTree_Bool_write + 1);
      else
        if ((memOut_QTree_Bool_valid == 1'd1))
          profiling_MemIn_QTree_Bool_read <= (profiling_MemIn_QTree_Bool_read + 1);
  
  /* demux (Ty C2,
       Ty MemOut_QTree_Bool) : (memMergeChoice_QTree_Bool,C2) (memOut_QTree_Bool_dbuf,MemOut_QTree_Bool) > [(memReadOut_QTree_Bool,MemOut_QTree_Bool),
                                                                                                            (memWriteOut_QTree_Bool,MemOut_QTree_Bool)] */
  logic [1:0] memOut_QTree_Bool_dbuf_onehotd;
  always_comb
    if ((memMergeChoice_QTree_Bool_d[0] && memOut_QTree_Bool_dbuf_d[0]))
      unique case (memMergeChoice_QTree_Bool_d[1:1])
        1'd0: memOut_QTree_Bool_dbuf_onehotd = 2'd1;
        1'd1: memOut_QTree_Bool_dbuf_onehotd = 2'd2;
        default: memOut_QTree_Bool_dbuf_onehotd = 2'd0;
      endcase
    else memOut_QTree_Bool_dbuf_onehotd = 2'd0;
  assign memReadOut_QTree_Bool_d = {memOut_QTree_Bool_dbuf_d[67:1],
                                    memOut_QTree_Bool_dbuf_onehotd[0]};
  assign memWriteOut_QTree_Bool_d = {memOut_QTree_Bool_dbuf_d[67:1],
                                     memOut_QTree_Bool_dbuf_onehotd[1]};
  assign memOut_QTree_Bool_dbuf_r = (| (memOut_QTree_Bool_dbuf_onehotd & {memWriteOut_QTree_Bool_r,
                                                                          memReadOut_QTree_Bool_r}));
  assign memMergeChoice_QTree_Bool_r = memOut_QTree_Bool_dbuf_r;
  
  /* dbuf (Ty MemIn_QTree_Bool) : (memMergeIn_QTree_Bool_rbuf,MemIn_QTree_Bool) > (memMergeIn_QTree_Bool_dbuf,MemIn_QTree_Bool) */
  assign memMergeIn_QTree_Bool_rbuf_r = ((! memMergeIn_QTree_Bool_dbuf_d[0]) || memMergeIn_QTree_Bool_dbuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memMergeIn_QTree_Bool_dbuf_d <= {83'd0, 1'd0};
    else
      if (memMergeIn_QTree_Bool_rbuf_r)
        memMergeIn_QTree_Bool_dbuf_d <= memMergeIn_QTree_Bool_rbuf_d;
  
  /* rbuf (Ty MemIn_QTree_Bool) : (memMergeIn_QTree_Bool,MemIn_QTree_Bool) > (memMergeIn_QTree_Bool_rbuf,MemIn_QTree_Bool) */
  MemIn_QTree_Bool_t memMergeIn_QTree_Bool_buf;
  assign memMergeIn_QTree_Bool_r = (! memMergeIn_QTree_Bool_buf[0]);
  assign memMergeIn_QTree_Bool_rbuf_d = (memMergeIn_QTree_Bool_buf[0] ? memMergeIn_QTree_Bool_buf :
                                         memMergeIn_QTree_Bool_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memMergeIn_QTree_Bool_buf <= {83'd0, 1'd0};
    else
      if ((memMergeIn_QTree_Bool_rbuf_r && memMergeIn_QTree_Bool_buf[0]))
        memMergeIn_QTree_Bool_buf <= {83'd0, 1'd0};
      else if (((! memMergeIn_QTree_Bool_rbuf_r) && (! memMergeIn_QTree_Bool_buf[0])))
        memMergeIn_QTree_Bool_buf <= memMergeIn_QTree_Bool_d;
  
  /* dbuf (Ty MemOut_QTree_Bool) : (memOut_QTree_Bool_rbuf,MemOut_QTree_Bool) > (memOut_QTree_Bool_dbuf,MemOut_QTree_Bool) */
  assign memOut_QTree_Bool_rbuf_r = ((! memOut_QTree_Bool_dbuf_d[0]) || memOut_QTree_Bool_dbuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memOut_QTree_Bool_dbuf_d <= {67'd0, 1'd0};
    else
      if (memOut_QTree_Bool_rbuf_r)
        memOut_QTree_Bool_dbuf_d <= memOut_QTree_Bool_rbuf_d;
  
  /* rbuf (Ty MemOut_QTree_Bool) : (memOut_QTree_Bool,MemOut_QTree_Bool) > (memOut_QTree_Bool_rbuf,MemOut_QTree_Bool) */
  MemOut_QTree_Bool_t memOut_QTree_Bool_buf;
  assign memOut_QTree_Bool_r = (! memOut_QTree_Bool_buf[0]);
  assign memOut_QTree_Bool_rbuf_d = (memOut_QTree_Bool_buf[0] ? memOut_QTree_Bool_buf :
                                     memOut_QTree_Bool_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memOut_QTree_Bool_buf <= {67'd0, 1'd0};
    else
      if ((memOut_QTree_Bool_rbuf_r && memOut_QTree_Bool_buf[0]))
        memOut_QTree_Bool_buf <= {67'd0, 1'd0};
      else if (((! memOut_QTree_Bool_rbuf_r) && (! memOut_QTree_Bool_buf[0])))
        memOut_QTree_Bool_buf <= memOut_QTree_Bool_d;
  
  /* mergectrl (Ty C5,
           Ty Pointer_QTree_Bool) : [(m1a84_1_argbuf,Pointer_QTree_Bool),
                                     (m2a85_1_argbuf,Pointer_QTree_Bool),
                                     (m3a86_1_argbuf,Pointer_QTree_Bool),
                                     (q4a90_1_argbuf,Pointer_QTree_Bool),
                                     (t4a91_1_argbuf,Pointer_QTree_Bool)] > (readMerge_choice_QTree_Bool,C5) (readMerge_data_QTree_Bool,Pointer_QTree_Bool) */
  logic [4:0] m1a84_1_argbuf_select_d;
  assign m1a84_1_argbuf_select_d = ((| m1a84_1_argbuf_select_q) ? m1a84_1_argbuf_select_q :
                                    (m1a84_1_argbuf_d[0] ? 5'd1 :
                                     (m2a85_1_argbuf_d[0] ? 5'd2 :
                                      (m3a86_1_argbuf_d[0] ? 5'd4 :
                                       (q4a90_1_argbuf_d[0] ? 5'd8 :
                                        (t4a91_1_argbuf_d[0] ? 5'd16 :
                                         5'd0))))));
  logic [4:0] m1a84_1_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m1a84_1_argbuf_select_q <= 5'd0;
    else
      m1a84_1_argbuf_select_q <= (m1a84_1_argbuf_done ? 5'd0 :
                                  m1a84_1_argbuf_select_d);
  logic [1:0] m1a84_1_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m1a84_1_argbuf_emit_q <= 2'd0;
    else
      m1a84_1_argbuf_emit_q <= (m1a84_1_argbuf_done ? 2'd0 :
                                m1a84_1_argbuf_emit_d);
  logic [1:0] m1a84_1_argbuf_emit_d;
  assign m1a84_1_argbuf_emit_d = (m1a84_1_argbuf_emit_q | ({readMerge_choice_QTree_Bool_d[0],
                                                            readMerge_data_QTree_Bool_d[0]} & {readMerge_choice_QTree_Bool_r,
                                                                                               readMerge_data_QTree_Bool_r}));
  logic m1a84_1_argbuf_done;
  assign m1a84_1_argbuf_done = (& m1a84_1_argbuf_emit_d);
  assign {t4a91_1_argbuf_r,
          q4a90_1_argbuf_r,
          m3a86_1_argbuf_r,
          m2a85_1_argbuf_r,
          m1a84_1_argbuf_r} = (m1a84_1_argbuf_done ? m1a84_1_argbuf_select_d :
                               5'd0);
  assign readMerge_data_QTree_Bool_d = ((m1a84_1_argbuf_select_d[0] && (! m1a84_1_argbuf_emit_q[0])) ? m1a84_1_argbuf_d :
                                        ((m1a84_1_argbuf_select_d[1] && (! m1a84_1_argbuf_emit_q[0])) ? m2a85_1_argbuf_d :
                                         ((m1a84_1_argbuf_select_d[2] && (! m1a84_1_argbuf_emit_q[0])) ? m3a86_1_argbuf_d :
                                          ((m1a84_1_argbuf_select_d[3] && (! m1a84_1_argbuf_emit_q[0])) ? q4a90_1_argbuf_d :
                                           ((m1a84_1_argbuf_select_d[4] && (! m1a84_1_argbuf_emit_q[0])) ? t4a91_1_argbuf_d :
                                            {16'd0, 1'd0})))));
  assign readMerge_choice_QTree_Bool_d = ((m1a84_1_argbuf_select_d[0] && (! m1a84_1_argbuf_emit_q[1])) ? C1_5_dc(1'd1) :
                                          ((m1a84_1_argbuf_select_d[1] && (! m1a84_1_argbuf_emit_q[1])) ? C2_5_dc(1'd1) :
                                           ((m1a84_1_argbuf_select_d[2] && (! m1a84_1_argbuf_emit_q[1])) ? C3_5_dc(1'd1) :
                                            ((m1a84_1_argbuf_select_d[3] && (! m1a84_1_argbuf_emit_q[1])) ? C4_5_dc(1'd1) :
                                             ((m1a84_1_argbuf_select_d[4] && (! m1a84_1_argbuf_emit_q[1])) ? C5_5_dc(1'd1) :
                                              {3'd0, 1'd0})))));
  
  /* demux (Ty C5,
       Ty QTree_Bool) : (readMerge_choice_QTree_Bool,C5) (destructReadOut_QTree_Bool,QTree_Bool) > [(readPointer_QTree_Boolm1a84_1_argbuf,QTree_Bool),
                                                                                                    (readPointer_QTree_Boolm2a85_1_argbuf,QTree_Bool),
                                                                                                    (readPointer_QTree_Boolm3a86_1_argbuf,QTree_Bool),
                                                                                                    (readPointer_QTree_Boolq4a90_1_argbuf,QTree_Bool),
                                                                                                    (readPointer_QTree_Boolt4a91_1_argbuf,QTree_Bool)] */
  logic [4:0] destructReadOut_QTree_Bool_onehotd;
  always_comb
    if ((readMerge_choice_QTree_Bool_d[0] && destructReadOut_QTree_Bool_d[0]))
      unique case (readMerge_choice_QTree_Bool_d[3:1])
        3'd0: destructReadOut_QTree_Bool_onehotd = 5'd1;
        3'd1: destructReadOut_QTree_Bool_onehotd = 5'd2;
        3'd2: destructReadOut_QTree_Bool_onehotd = 5'd4;
        3'd3: destructReadOut_QTree_Bool_onehotd = 5'd8;
        3'd4: destructReadOut_QTree_Bool_onehotd = 5'd16;
        default: destructReadOut_QTree_Bool_onehotd = 5'd0;
      endcase
    else destructReadOut_QTree_Bool_onehotd = 5'd0;
  assign readPointer_QTree_Boolm1a84_1_argbuf_d = {destructReadOut_QTree_Bool_d[66:1],
                                                   destructReadOut_QTree_Bool_onehotd[0]};
  assign readPointer_QTree_Boolm2a85_1_argbuf_d = {destructReadOut_QTree_Bool_d[66:1],
                                                   destructReadOut_QTree_Bool_onehotd[1]};
  assign readPointer_QTree_Boolm3a86_1_argbuf_d = {destructReadOut_QTree_Bool_d[66:1],
                                                   destructReadOut_QTree_Bool_onehotd[2]};
  assign readPointer_QTree_Boolq4a90_1_argbuf_d = {destructReadOut_QTree_Bool_d[66:1],
                                                   destructReadOut_QTree_Bool_onehotd[3]};
  assign readPointer_QTree_Boolt4a91_1_argbuf_d = {destructReadOut_QTree_Bool_d[66:1],
                                                   destructReadOut_QTree_Bool_onehotd[4]};
  assign destructReadOut_QTree_Bool_r = (| (destructReadOut_QTree_Bool_onehotd & {readPointer_QTree_Boolt4a91_1_argbuf_r,
                                                                                  readPointer_QTree_Boolq4a90_1_argbuf_r,
                                                                                  readPointer_QTree_Boolm3a86_1_argbuf_r,
                                                                                  readPointer_QTree_Boolm2a85_1_argbuf_r,
                                                                                  readPointer_QTree_Boolm1a84_1_argbuf_r}));
  assign readMerge_choice_QTree_Bool_r = destructReadOut_QTree_Bool_r;
  
  /* destruct (Ty Pointer_QTree_Bool,
          Dcon Pointer_QTree_Bool) : (readMerge_data_QTree_Bool,Pointer_QTree_Bool) > [(destructReadIn_QTree_Bool,Word16#)] */
  assign destructReadIn_QTree_Bool_d = {readMerge_data_QTree_Bool_d[16:1],
                                        readMerge_data_QTree_Bool_d[0]};
  assign readMerge_data_QTree_Bool_r = destructReadIn_QTree_Bool_r;
  
  /* dcon (Ty MemIn_QTree_Bool,
      Dcon ReadIn_QTree_Bool) : [(destructReadIn_QTree_Bool,Word16#)] > (dconReadIn_QTree_Bool,MemIn_QTree_Bool) */
  assign dconReadIn_QTree_Bool_d = ReadIn_QTree_Bool_dc((& {destructReadIn_QTree_Bool_d[0]}), destructReadIn_QTree_Bool_d);
  assign {destructReadIn_QTree_Bool_r} = {1 {(dconReadIn_QTree_Bool_r && dconReadIn_QTree_Bool_d[0])}};
  
  /* destruct (Ty MemOut_QTree_Bool,
          Dcon ReadOut_QTree_Bool) : (memReadOut_QTree_Bool,MemOut_QTree_Bool) > [(destructReadOut_QTree_Bool,QTree_Bool)] */
  assign destructReadOut_QTree_Bool_d = {memReadOut_QTree_Bool_d[67:2],
                                         memReadOut_QTree_Bool_d[0]};
  assign memReadOut_QTree_Bool_r = destructReadOut_QTree_Bool_r;
  
  /* mergectrl (Ty C35,
           Ty QTree_Bool) : [(lizzieLet10_1_1_argbuf,QTree_Bool),
                             (lizzieLet11_1_1_argbuf,QTree_Bool),
                             (lizzieLet12_1_1_argbuf,QTree_Bool),
                             (lizzieLet15_1_1_argbuf,QTree_Bool),
                             (lizzieLet18_1_argbuf,QTree_Bool),
                             (lizzieLet19_1_argbuf,QTree_Bool),
                             (lizzieLet23_1_argbuf,QTree_Bool),
                             (lizzieLet24_1_argbuf,QTree_Bool),
                             (lizzieLet28_1_argbuf,QTree_Bool),
                             (lizzieLet29_1_argbuf,QTree_Bool),
                             (lizzieLet30_1_argbuf,QTree_Bool),
                             (lizzieLet31_1_argbuf,QTree_Bool),
                             (lizzieLet34_1_argbuf,QTree_Bool),
                             (lizzieLet35_1_argbuf,QTree_Bool),
                             (lizzieLet36_1_argbuf,QTree_Bool),
                             (lizzieLet37_1_argbuf,QTree_Bool),
                             (lizzieLet39_1_argbuf,QTree_Bool),
                             (lizzieLet3_1_argbuf,QTree_Bool),
                             (lizzieLet40_1_argbuf,QTree_Bool),
                             (lizzieLet42_1_argbuf,QTree_Bool),
                             (lizzieLet43_1_argbuf,QTree_Bool),
                             (lizzieLet44_1_argbuf,QTree_Bool),
                             (lizzieLet47_1_argbuf,QTree_Bool),
                             (lizzieLet50_1_argbuf,QTree_Bool),
                             (lizzieLet51_1_argbuf,QTree_Bool),
                             (lizzieLet53_1_argbuf,QTree_Bool),
                             (lizzieLet55_1_argbuf,QTree_Bool),
                             (lizzieLet56_1_argbuf,QTree_Bool),
                             (lizzieLet59_1_argbuf,QTree_Bool),
                             (lizzieLet64_1_argbuf,QTree_Bool),
                             (lizzieLet69_1_argbuf,QTree_Bool),
                             (lizzieLet6_1_argbuf,QTree_Bool),
                             (lizzieLet7_1_argbuf,QTree_Bool),
                             (lizzieLet9_1_1_argbuf,QTree_Bool),
                             (dummy_write_QTree_Bool,QTree_Bool)] > (writeMerge_choice_QTree_Bool,C35) (writeMerge_data_QTree_Bool,QTree_Bool) */
  logic [34:0] lizzieLet10_1_1_argbuf_select_d;
  assign lizzieLet10_1_1_argbuf_select_d = ((| lizzieLet10_1_1_argbuf_select_q) ? lizzieLet10_1_1_argbuf_select_q :
                                            (lizzieLet10_1_1_argbuf_d[0] ? 35'd1 :
                                             (lizzieLet11_1_1_argbuf_d[0] ? 35'd2 :
                                              (lizzieLet12_1_1_argbuf_d[0] ? 35'd4 :
                                               (lizzieLet15_1_1_argbuf_d[0] ? 35'd8 :
                                                (lizzieLet18_1_argbuf_d[0] ? 35'd16 :
                                                 (lizzieLet19_1_argbuf_d[0] ? 35'd32 :
                                                  (lizzieLet23_1_argbuf_d[0] ? 35'd64 :
                                                   (lizzieLet24_1_argbuf_d[0] ? 35'd128 :
                                                    (lizzieLet28_1_argbuf_d[0] ? 35'd256 :
                                                     (lizzieLet29_1_argbuf_d[0] ? 35'd512 :
                                                      (lizzieLet30_1_argbuf_d[0] ? 35'd1024 :
                                                       (lizzieLet31_1_argbuf_d[0] ? 35'd2048 :
                                                        (lizzieLet34_1_argbuf_d[0] ? 35'd4096 :
                                                         (lizzieLet35_1_argbuf_d[0] ? 35'd8192 :
                                                          (lizzieLet36_1_argbuf_d[0] ? 35'd16384 :
                                                           (lizzieLet37_1_argbuf_d[0] ? 35'd32768 :
                                                            (lizzieLet39_1_argbuf_d[0] ? 35'd65536 :
                                                             (lizzieLet3_1_argbuf_d[0] ? 35'd131072 :
                                                              (lizzieLet40_1_argbuf_d[0] ? 35'd262144 :
                                                               (lizzieLet42_1_argbuf_d[0] ? 35'd524288 :
                                                                (lizzieLet43_1_argbuf_d[0] ? 35'd1048576 :
                                                                 (lizzieLet44_1_argbuf_d[0] ? 35'd2097152 :
                                                                  (lizzieLet47_1_argbuf_d[0] ? 35'd4194304 :
                                                                   (lizzieLet50_1_argbuf_d[0] ? 35'd8388608 :
                                                                    (lizzieLet51_1_argbuf_d[0] ? 35'd16777216 :
                                                                     (lizzieLet53_1_argbuf_d[0] ? 35'd33554432 :
                                                                      (lizzieLet55_1_argbuf_d[0] ? 35'd67108864 :
                                                                       (lizzieLet56_1_argbuf_d[0] ? 35'd134217728 :
                                                                        (lizzieLet59_1_argbuf_d[0] ? 35'd268435456 :
                                                                         (lizzieLet64_1_argbuf_d[0] ? 35'd536870912 :
                                                                          (lizzieLet69_1_argbuf_d[0] ? 35'd1073741824 :
                                                                           (lizzieLet6_1_argbuf_d[0] ? 35'd2147483648 :
                                                                            (lizzieLet7_1_argbuf_d[0] ? 35'd4294967296 :
                                                                             (lizzieLet9_1_1_argbuf_d[0] ? 35'd8589934592 :
                                                                              (dummy_write_QTree_Bool_d[0] ? 35'd17179869184 :
                                                                               35'd0))))))))))))))))))))))))))))))))))));
  logic [34:0] lizzieLet10_1_1_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet10_1_1_argbuf_select_q <= 35'd0;
    else
      lizzieLet10_1_1_argbuf_select_q <= (lizzieLet10_1_1_argbuf_done ? 35'd0 :
                                          lizzieLet10_1_1_argbuf_select_d);
  logic [1:0] lizzieLet10_1_1_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet10_1_1_argbuf_emit_q <= 2'd0;
    else
      lizzieLet10_1_1_argbuf_emit_q <= (lizzieLet10_1_1_argbuf_done ? 2'd0 :
                                        lizzieLet10_1_1_argbuf_emit_d);
  logic [1:0] lizzieLet10_1_1_argbuf_emit_d;
  assign lizzieLet10_1_1_argbuf_emit_d = (lizzieLet10_1_1_argbuf_emit_q | ({writeMerge_choice_QTree_Bool_d[0],
                                                                            writeMerge_data_QTree_Bool_d[0]} & {writeMerge_choice_QTree_Bool_r,
                                                                                                                writeMerge_data_QTree_Bool_r}));
  logic lizzieLet10_1_1_argbuf_done;
  assign lizzieLet10_1_1_argbuf_done = (& lizzieLet10_1_1_argbuf_emit_d);
  assign {dummy_write_QTree_Bool_r,
          lizzieLet9_1_1_argbuf_r,
          lizzieLet7_1_argbuf_r,
          lizzieLet6_1_argbuf_r,
          lizzieLet69_1_argbuf_r,
          lizzieLet64_1_argbuf_r,
          lizzieLet59_1_argbuf_r,
          lizzieLet56_1_argbuf_r,
          lizzieLet55_1_argbuf_r,
          lizzieLet53_1_argbuf_r,
          lizzieLet51_1_argbuf_r,
          lizzieLet50_1_argbuf_r,
          lizzieLet47_1_argbuf_r,
          lizzieLet44_1_argbuf_r,
          lizzieLet43_1_argbuf_r,
          lizzieLet42_1_argbuf_r,
          lizzieLet40_1_argbuf_r,
          lizzieLet3_1_argbuf_r,
          lizzieLet39_1_argbuf_r,
          lizzieLet37_1_argbuf_r,
          lizzieLet36_1_argbuf_r,
          lizzieLet35_1_argbuf_r,
          lizzieLet34_1_argbuf_r,
          lizzieLet31_1_argbuf_r,
          lizzieLet30_1_argbuf_r,
          lizzieLet29_1_argbuf_r,
          lizzieLet28_1_argbuf_r,
          lizzieLet24_1_argbuf_r,
          lizzieLet23_1_argbuf_r,
          lizzieLet19_1_argbuf_r,
          lizzieLet18_1_argbuf_r,
          lizzieLet15_1_1_argbuf_r,
          lizzieLet12_1_1_argbuf_r,
          lizzieLet11_1_1_argbuf_r,
          lizzieLet10_1_1_argbuf_r} = (lizzieLet10_1_1_argbuf_done ? lizzieLet10_1_1_argbuf_select_d :
                                       35'd0);
  assign writeMerge_data_QTree_Bool_d = ((lizzieLet10_1_1_argbuf_select_d[0] && (! lizzieLet10_1_1_argbuf_emit_q[0])) ? lizzieLet10_1_1_argbuf_d :
                                         ((lizzieLet10_1_1_argbuf_select_d[1] && (! lizzieLet10_1_1_argbuf_emit_q[0])) ? lizzieLet11_1_1_argbuf_d :
                                          ((lizzieLet10_1_1_argbuf_select_d[2] && (! lizzieLet10_1_1_argbuf_emit_q[0])) ? lizzieLet12_1_1_argbuf_d :
                                           ((lizzieLet10_1_1_argbuf_select_d[3] && (! lizzieLet10_1_1_argbuf_emit_q[0])) ? lizzieLet15_1_1_argbuf_d :
                                            ((lizzieLet10_1_1_argbuf_select_d[4] && (! lizzieLet10_1_1_argbuf_emit_q[0])) ? lizzieLet18_1_argbuf_d :
                                             ((lizzieLet10_1_1_argbuf_select_d[5] && (! lizzieLet10_1_1_argbuf_emit_q[0])) ? lizzieLet19_1_argbuf_d :
                                              ((lizzieLet10_1_1_argbuf_select_d[6] && (! lizzieLet10_1_1_argbuf_emit_q[0])) ? lizzieLet23_1_argbuf_d :
                                               ((lizzieLet10_1_1_argbuf_select_d[7] && (! lizzieLet10_1_1_argbuf_emit_q[0])) ? lizzieLet24_1_argbuf_d :
                                                ((lizzieLet10_1_1_argbuf_select_d[8] && (! lizzieLet10_1_1_argbuf_emit_q[0])) ? lizzieLet28_1_argbuf_d :
                                                 ((lizzieLet10_1_1_argbuf_select_d[9] && (! lizzieLet10_1_1_argbuf_emit_q[0])) ? lizzieLet29_1_argbuf_d :
                                                  ((lizzieLet10_1_1_argbuf_select_d[10] && (! lizzieLet10_1_1_argbuf_emit_q[0])) ? lizzieLet30_1_argbuf_d :
                                                   ((lizzieLet10_1_1_argbuf_select_d[11] && (! lizzieLet10_1_1_argbuf_emit_q[0])) ? lizzieLet31_1_argbuf_d :
                                                    ((lizzieLet10_1_1_argbuf_select_d[12] && (! lizzieLet10_1_1_argbuf_emit_q[0])) ? lizzieLet34_1_argbuf_d :
                                                     ((lizzieLet10_1_1_argbuf_select_d[13] && (! lizzieLet10_1_1_argbuf_emit_q[0])) ? lizzieLet35_1_argbuf_d :
                                                      ((lizzieLet10_1_1_argbuf_select_d[14] && (! lizzieLet10_1_1_argbuf_emit_q[0])) ? lizzieLet36_1_argbuf_d :
                                                       ((lizzieLet10_1_1_argbuf_select_d[15] && (! lizzieLet10_1_1_argbuf_emit_q[0])) ? lizzieLet37_1_argbuf_d :
                                                        ((lizzieLet10_1_1_argbuf_select_d[16] && (! lizzieLet10_1_1_argbuf_emit_q[0])) ? lizzieLet39_1_argbuf_d :
                                                         ((lizzieLet10_1_1_argbuf_select_d[17] && (! lizzieLet10_1_1_argbuf_emit_q[0])) ? lizzieLet3_1_argbuf_d :
                                                          ((lizzieLet10_1_1_argbuf_select_d[18] && (! lizzieLet10_1_1_argbuf_emit_q[0])) ? lizzieLet40_1_argbuf_d :
                                                           ((lizzieLet10_1_1_argbuf_select_d[19] && (! lizzieLet10_1_1_argbuf_emit_q[0])) ? lizzieLet42_1_argbuf_d :
                                                            ((lizzieLet10_1_1_argbuf_select_d[20] && (! lizzieLet10_1_1_argbuf_emit_q[0])) ? lizzieLet43_1_argbuf_d :
                                                             ((lizzieLet10_1_1_argbuf_select_d[21] && (! lizzieLet10_1_1_argbuf_emit_q[0])) ? lizzieLet44_1_argbuf_d :
                                                              ((lizzieLet10_1_1_argbuf_select_d[22] && (! lizzieLet10_1_1_argbuf_emit_q[0])) ? lizzieLet47_1_argbuf_d :
                                                               ((lizzieLet10_1_1_argbuf_select_d[23] && (! lizzieLet10_1_1_argbuf_emit_q[0])) ? lizzieLet50_1_argbuf_d :
                                                                ((lizzieLet10_1_1_argbuf_select_d[24] && (! lizzieLet10_1_1_argbuf_emit_q[0])) ? lizzieLet51_1_argbuf_d :
                                                                 ((lizzieLet10_1_1_argbuf_select_d[25] && (! lizzieLet10_1_1_argbuf_emit_q[0])) ? lizzieLet53_1_argbuf_d :
                                                                  ((lizzieLet10_1_1_argbuf_select_d[26] && (! lizzieLet10_1_1_argbuf_emit_q[0])) ? lizzieLet55_1_argbuf_d :
                                                                   ((lizzieLet10_1_1_argbuf_select_d[27] && (! lizzieLet10_1_1_argbuf_emit_q[0])) ? lizzieLet56_1_argbuf_d :
                                                                    ((lizzieLet10_1_1_argbuf_select_d[28] && (! lizzieLet10_1_1_argbuf_emit_q[0])) ? lizzieLet59_1_argbuf_d :
                                                                     ((lizzieLet10_1_1_argbuf_select_d[29] && (! lizzieLet10_1_1_argbuf_emit_q[0])) ? lizzieLet64_1_argbuf_d :
                                                                      ((lizzieLet10_1_1_argbuf_select_d[30] && (! lizzieLet10_1_1_argbuf_emit_q[0])) ? lizzieLet69_1_argbuf_d :
                                                                       ((lizzieLet10_1_1_argbuf_select_d[31] && (! lizzieLet10_1_1_argbuf_emit_q[0])) ? lizzieLet6_1_argbuf_d :
                                                                        ((lizzieLet10_1_1_argbuf_select_d[32] && (! lizzieLet10_1_1_argbuf_emit_q[0])) ? lizzieLet7_1_argbuf_d :
                                                                         ((lizzieLet10_1_1_argbuf_select_d[33] && (! lizzieLet10_1_1_argbuf_emit_q[0])) ? lizzieLet9_1_1_argbuf_d :
                                                                          ((lizzieLet10_1_1_argbuf_select_d[34] && (! lizzieLet10_1_1_argbuf_emit_q[0])) ? dummy_write_QTree_Bool_d :
                                                                           {66'd0,
                                                                            1'd0})))))))))))))))))))))))))))))))))));
  assign writeMerge_choice_QTree_Bool_d = ((lizzieLet10_1_1_argbuf_select_d[0] && (! lizzieLet10_1_1_argbuf_emit_q[1])) ? C1_35_dc(1'd1) :
                                           ((lizzieLet10_1_1_argbuf_select_d[1] && (! lizzieLet10_1_1_argbuf_emit_q[1])) ? C2_35_dc(1'd1) :
                                            ((lizzieLet10_1_1_argbuf_select_d[2] && (! lizzieLet10_1_1_argbuf_emit_q[1])) ? C3_35_dc(1'd1) :
                                             ((lizzieLet10_1_1_argbuf_select_d[3] && (! lizzieLet10_1_1_argbuf_emit_q[1])) ? C4_35_dc(1'd1) :
                                              ((lizzieLet10_1_1_argbuf_select_d[4] && (! lizzieLet10_1_1_argbuf_emit_q[1])) ? C5_35_dc(1'd1) :
                                               ((lizzieLet10_1_1_argbuf_select_d[5] && (! lizzieLet10_1_1_argbuf_emit_q[1])) ? C6_35_dc(1'd1) :
                                                ((lizzieLet10_1_1_argbuf_select_d[6] && (! lizzieLet10_1_1_argbuf_emit_q[1])) ? C7_35_dc(1'd1) :
                                                 ((lizzieLet10_1_1_argbuf_select_d[7] && (! lizzieLet10_1_1_argbuf_emit_q[1])) ? C8_35_dc(1'd1) :
                                                  ((lizzieLet10_1_1_argbuf_select_d[8] && (! lizzieLet10_1_1_argbuf_emit_q[1])) ? C9_35_dc(1'd1) :
                                                   ((lizzieLet10_1_1_argbuf_select_d[9] && (! lizzieLet10_1_1_argbuf_emit_q[1])) ? C10_35_dc(1'd1) :
                                                    ((lizzieLet10_1_1_argbuf_select_d[10] && (! lizzieLet10_1_1_argbuf_emit_q[1])) ? C11_35_dc(1'd1) :
                                                     ((lizzieLet10_1_1_argbuf_select_d[11] && (! lizzieLet10_1_1_argbuf_emit_q[1])) ? C12_35_dc(1'd1) :
                                                      ((lizzieLet10_1_1_argbuf_select_d[12] && (! lizzieLet10_1_1_argbuf_emit_q[1])) ? C13_35_dc(1'd1) :
                                                       ((lizzieLet10_1_1_argbuf_select_d[13] && (! lizzieLet10_1_1_argbuf_emit_q[1])) ? C14_35_dc(1'd1) :
                                                        ((lizzieLet10_1_1_argbuf_select_d[14] && (! lizzieLet10_1_1_argbuf_emit_q[1])) ? C15_35_dc(1'd1) :
                                                         ((lizzieLet10_1_1_argbuf_select_d[15] && (! lizzieLet10_1_1_argbuf_emit_q[1])) ? C16_35_dc(1'd1) :
                                                          ((lizzieLet10_1_1_argbuf_select_d[16] && (! lizzieLet10_1_1_argbuf_emit_q[1])) ? C17_35_dc(1'd1) :
                                                           ((lizzieLet10_1_1_argbuf_select_d[17] && (! lizzieLet10_1_1_argbuf_emit_q[1])) ? C18_35_dc(1'd1) :
                                                            ((lizzieLet10_1_1_argbuf_select_d[18] && (! lizzieLet10_1_1_argbuf_emit_q[1])) ? C19_35_dc(1'd1) :
                                                             ((lizzieLet10_1_1_argbuf_select_d[19] && (! lizzieLet10_1_1_argbuf_emit_q[1])) ? C20_35_dc(1'd1) :
                                                              ((lizzieLet10_1_1_argbuf_select_d[20] && (! lizzieLet10_1_1_argbuf_emit_q[1])) ? C21_35_dc(1'd1) :
                                                               ((lizzieLet10_1_1_argbuf_select_d[21] && (! lizzieLet10_1_1_argbuf_emit_q[1])) ? C22_35_dc(1'd1) :
                                                                ((lizzieLet10_1_1_argbuf_select_d[22] && (! lizzieLet10_1_1_argbuf_emit_q[1])) ? C23_35_dc(1'd1) :
                                                                 ((lizzieLet10_1_1_argbuf_select_d[23] && (! lizzieLet10_1_1_argbuf_emit_q[1])) ? C24_35_dc(1'd1) :
                                                                  ((lizzieLet10_1_1_argbuf_select_d[24] && (! lizzieLet10_1_1_argbuf_emit_q[1])) ? C25_35_dc(1'd1) :
                                                                   ((lizzieLet10_1_1_argbuf_select_d[25] && (! lizzieLet10_1_1_argbuf_emit_q[1])) ? C26_35_dc(1'd1) :
                                                                    ((lizzieLet10_1_1_argbuf_select_d[26] && (! lizzieLet10_1_1_argbuf_emit_q[1])) ? C27_35_dc(1'd1) :
                                                                     ((lizzieLet10_1_1_argbuf_select_d[27] && (! lizzieLet10_1_1_argbuf_emit_q[1])) ? C28_35_dc(1'd1) :
                                                                      ((lizzieLet10_1_1_argbuf_select_d[28] && (! lizzieLet10_1_1_argbuf_emit_q[1])) ? C29_35_dc(1'd1) :
                                                                       ((lizzieLet10_1_1_argbuf_select_d[29] && (! lizzieLet10_1_1_argbuf_emit_q[1])) ? C30_35_dc(1'd1) :
                                                                        ((lizzieLet10_1_1_argbuf_select_d[30] && (! lizzieLet10_1_1_argbuf_emit_q[1])) ? C31_35_dc(1'd1) :
                                                                         ((lizzieLet10_1_1_argbuf_select_d[31] && (! lizzieLet10_1_1_argbuf_emit_q[1])) ? C32_35_dc(1'd1) :
                                                                          ((lizzieLet10_1_1_argbuf_select_d[32] && (! lizzieLet10_1_1_argbuf_emit_q[1])) ? C33_35_dc(1'd1) :
                                                                           ((lizzieLet10_1_1_argbuf_select_d[33] && (! lizzieLet10_1_1_argbuf_emit_q[1])) ? C34_35_dc(1'd1) :
                                                                            ((lizzieLet10_1_1_argbuf_select_d[34] && (! lizzieLet10_1_1_argbuf_emit_q[1])) ? C35_35_dc(1'd1) :
                                                                             {6'd0,
                                                                              1'd0})))))))))))))))))))))))))))))))))));
  
  /* demux (Ty C35,
       Ty Pointer_QTree_Bool) : (writeMerge_choice_QTree_Bool,C35) (demuxWriteResult_QTree_Bool,Pointer_QTree_Bool) > [(writeQTree_BoollizzieLet10_1_1_argbuf,Pointer_QTree_Bool),
                                                                                                                       (writeQTree_BoollizzieLet11_1_1_argbuf,Pointer_QTree_Bool),
                                                                                                                       (writeQTree_BoollizzieLet12_1_1_argbuf,Pointer_QTree_Bool),
                                                                                                                       (writeQTree_BoollizzieLet15_1_1_argbuf,Pointer_QTree_Bool),
                                                                                                                       (writeQTree_BoollizzieLet18_1_argbuf,Pointer_QTree_Bool),
                                                                                                                       (writeQTree_BoollizzieLet19_1_argbuf,Pointer_QTree_Bool),
                                                                                                                       (writeQTree_BoollizzieLet23_1_argbuf,Pointer_QTree_Bool),
                                                                                                                       (writeQTree_BoollizzieLet24_1_argbuf,Pointer_QTree_Bool),
                                                                                                                       (writeQTree_BoollizzieLet28_1_argbuf,Pointer_QTree_Bool),
                                                                                                                       (writeQTree_BoollizzieLet29_1_argbuf,Pointer_QTree_Bool),
                                                                                                                       (writeQTree_BoollizzieLet30_1_argbuf,Pointer_QTree_Bool),
                                                                                                                       (writeQTree_BoollizzieLet31_1_argbuf,Pointer_QTree_Bool),
                                                                                                                       (writeQTree_BoollizzieLet34_1_argbuf,Pointer_QTree_Bool),
                                                                                                                       (writeQTree_BoollizzieLet35_1_argbuf,Pointer_QTree_Bool),
                                                                                                                       (writeQTree_BoollizzieLet36_1_argbuf,Pointer_QTree_Bool),
                                                                                                                       (writeQTree_BoollizzieLet37_1_argbuf,Pointer_QTree_Bool),
                                                                                                                       (writeQTree_BoollizzieLet39_1_argbuf,Pointer_QTree_Bool),
                                                                                                                       (writeQTree_BoollizzieLet3_1_argbuf,Pointer_QTree_Bool),
                                                                                                                       (writeQTree_BoollizzieLet40_1_argbuf,Pointer_QTree_Bool),
                                                                                                                       (writeQTree_BoollizzieLet42_1_argbuf,Pointer_QTree_Bool),
                                                                                                                       (writeQTree_BoollizzieLet43_1_argbuf,Pointer_QTree_Bool),
                                                                                                                       (writeQTree_BoollizzieLet44_1_argbuf,Pointer_QTree_Bool),
                                                                                                                       (writeQTree_BoollizzieLet47_1_argbuf,Pointer_QTree_Bool),
                                                                                                                       (writeQTree_BoollizzieLet50_1_argbuf,Pointer_QTree_Bool),
                                                                                                                       (writeQTree_BoollizzieLet51_1_argbuf,Pointer_QTree_Bool),
                                                                                                                       (writeQTree_BoollizzieLet53_1_argbuf,Pointer_QTree_Bool),
                                                                                                                       (writeQTree_BoollizzieLet55_1_argbuf,Pointer_QTree_Bool),
                                                                                                                       (writeQTree_BoollizzieLet56_1_argbuf,Pointer_QTree_Bool),
                                                                                                                       (writeQTree_BoollizzieLet59_1_argbuf,Pointer_QTree_Bool),
                                                                                                                       (writeQTree_BoollizzieLet64_1_argbuf,Pointer_QTree_Bool),
                                                                                                                       (writeQTree_BoollizzieLet69_1_argbuf,Pointer_QTree_Bool),
                                                                                                                       (writeQTree_BoollizzieLet6_1_argbuf,Pointer_QTree_Bool),
                                                                                                                       (writeQTree_BoollizzieLet7_1_argbuf,Pointer_QTree_Bool),
                                                                                                                       (writeQTree_BoollizzieLet9_1_1_argbuf,Pointer_QTree_Bool),
                                                                                                                       (dummy_write_QTree_Bool_sink,Pointer_QTree_Bool)] */
  logic [34:0] demuxWriteResult_QTree_Bool_onehotd;
  always_comb
    if ((writeMerge_choice_QTree_Bool_d[0] && demuxWriteResult_QTree_Bool_d[0]))
      unique case (writeMerge_choice_QTree_Bool_d[6:1])
        6'd0: demuxWriteResult_QTree_Bool_onehotd = 35'd1;
        6'd1: demuxWriteResult_QTree_Bool_onehotd = 35'd2;
        6'd2: demuxWriteResult_QTree_Bool_onehotd = 35'd4;
        6'd3: demuxWriteResult_QTree_Bool_onehotd = 35'd8;
        6'd4: demuxWriteResult_QTree_Bool_onehotd = 35'd16;
        6'd5: demuxWriteResult_QTree_Bool_onehotd = 35'd32;
        6'd6: demuxWriteResult_QTree_Bool_onehotd = 35'd64;
        6'd7: demuxWriteResult_QTree_Bool_onehotd = 35'd128;
        6'd8: demuxWriteResult_QTree_Bool_onehotd = 35'd256;
        6'd9: demuxWriteResult_QTree_Bool_onehotd = 35'd512;
        6'd10: demuxWriteResult_QTree_Bool_onehotd = 35'd1024;
        6'd11: demuxWriteResult_QTree_Bool_onehotd = 35'd2048;
        6'd12: demuxWriteResult_QTree_Bool_onehotd = 35'd4096;
        6'd13: demuxWriteResult_QTree_Bool_onehotd = 35'd8192;
        6'd14: demuxWriteResult_QTree_Bool_onehotd = 35'd16384;
        6'd15: demuxWriteResult_QTree_Bool_onehotd = 35'd32768;
        6'd16: demuxWriteResult_QTree_Bool_onehotd = 35'd65536;
        6'd17: demuxWriteResult_QTree_Bool_onehotd = 35'd131072;
        6'd18: demuxWriteResult_QTree_Bool_onehotd = 35'd262144;
        6'd19: demuxWriteResult_QTree_Bool_onehotd = 35'd524288;
        6'd20: demuxWriteResult_QTree_Bool_onehotd = 35'd1048576;
        6'd21: demuxWriteResult_QTree_Bool_onehotd = 35'd2097152;
        6'd22: demuxWriteResult_QTree_Bool_onehotd = 35'd4194304;
        6'd23: demuxWriteResult_QTree_Bool_onehotd = 35'd8388608;
        6'd24: demuxWriteResult_QTree_Bool_onehotd = 35'd16777216;
        6'd25: demuxWriteResult_QTree_Bool_onehotd = 35'd33554432;
        6'd26: demuxWriteResult_QTree_Bool_onehotd = 35'd67108864;
        6'd27: demuxWriteResult_QTree_Bool_onehotd = 35'd134217728;
        6'd28: demuxWriteResult_QTree_Bool_onehotd = 35'd268435456;
        6'd29: demuxWriteResult_QTree_Bool_onehotd = 35'd536870912;
        6'd30: demuxWriteResult_QTree_Bool_onehotd = 35'd1073741824;
        6'd31: demuxWriteResult_QTree_Bool_onehotd = 35'd2147483648;
        6'd32: demuxWriteResult_QTree_Bool_onehotd = 35'd4294967296;
        6'd33: demuxWriteResult_QTree_Bool_onehotd = 35'd8589934592;
        6'd34: demuxWriteResult_QTree_Bool_onehotd = 35'd17179869184;
        default: demuxWriteResult_QTree_Bool_onehotd = 35'd0;
      endcase
    else demuxWriteResult_QTree_Bool_onehotd = 35'd0;
  assign writeQTree_BoollizzieLet10_1_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                    demuxWriteResult_QTree_Bool_onehotd[0]};
  assign writeQTree_BoollizzieLet11_1_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                    demuxWriteResult_QTree_Bool_onehotd[1]};
  assign writeQTree_BoollizzieLet12_1_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                    demuxWriteResult_QTree_Bool_onehotd[2]};
  assign writeQTree_BoollizzieLet15_1_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                    demuxWriteResult_QTree_Bool_onehotd[3]};
  assign writeQTree_BoollizzieLet18_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                  demuxWriteResult_QTree_Bool_onehotd[4]};
  assign writeQTree_BoollizzieLet19_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                  demuxWriteResult_QTree_Bool_onehotd[5]};
  assign writeQTree_BoollizzieLet23_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                  demuxWriteResult_QTree_Bool_onehotd[6]};
  assign writeQTree_BoollizzieLet24_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                  demuxWriteResult_QTree_Bool_onehotd[7]};
  assign writeQTree_BoollizzieLet28_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                  demuxWriteResult_QTree_Bool_onehotd[8]};
  assign writeQTree_BoollizzieLet29_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                  demuxWriteResult_QTree_Bool_onehotd[9]};
  assign writeQTree_BoollizzieLet30_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                  demuxWriteResult_QTree_Bool_onehotd[10]};
  assign writeQTree_BoollizzieLet31_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                  demuxWriteResult_QTree_Bool_onehotd[11]};
  assign writeQTree_BoollizzieLet34_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                  demuxWriteResult_QTree_Bool_onehotd[12]};
  assign writeQTree_BoollizzieLet35_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                  demuxWriteResult_QTree_Bool_onehotd[13]};
  assign writeQTree_BoollizzieLet36_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                  demuxWriteResult_QTree_Bool_onehotd[14]};
  assign writeQTree_BoollizzieLet37_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                  demuxWriteResult_QTree_Bool_onehotd[15]};
  assign writeQTree_BoollizzieLet39_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                  demuxWriteResult_QTree_Bool_onehotd[16]};
  assign writeQTree_BoollizzieLet3_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                 demuxWriteResult_QTree_Bool_onehotd[17]};
  assign writeQTree_BoollizzieLet40_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                  demuxWriteResult_QTree_Bool_onehotd[18]};
  assign writeQTree_BoollizzieLet42_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                  demuxWriteResult_QTree_Bool_onehotd[19]};
  assign writeQTree_BoollizzieLet43_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                  demuxWriteResult_QTree_Bool_onehotd[20]};
  assign writeQTree_BoollizzieLet44_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                  demuxWriteResult_QTree_Bool_onehotd[21]};
  assign writeQTree_BoollizzieLet47_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                  demuxWriteResult_QTree_Bool_onehotd[22]};
  assign writeQTree_BoollizzieLet50_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                  demuxWriteResult_QTree_Bool_onehotd[23]};
  assign writeQTree_BoollizzieLet51_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                  demuxWriteResult_QTree_Bool_onehotd[24]};
  assign writeQTree_BoollizzieLet53_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                  demuxWriteResult_QTree_Bool_onehotd[25]};
  assign writeQTree_BoollizzieLet55_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                  demuxWriteResult_QTree_Bool_onehotd[26]};
  assign writeQTree_BoollizzieLet56_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                  demuxWriteResult_QTree_Bool_onehotd[27]};
  assign writeQTree_BoollizzieLet59_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                  demuxWriteResult_QTree_Bool_onehotd[28]};
  assign writeQTree_BoollizzieLet64_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                  demuxWriteResult_QTree_Bool_onehotd[29]};
  assign writeQTree_BoollizzieLet69_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                  demuxWriteResult_QTree_Bool_onehotd[30]};
  assign writeQTree_BoollizzieLet6_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                 demuxWriteResult_QTree_Bool_onehotd[31]};
  assign writeQTree_BoollizzieLet7_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                 demuxWriteResult_QTree_Bool_onehotd[32]};
  assign writeQTree_BoollizzieLet9_1_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                   demuxWriteResult_QTree_Bool_onehotd[33]};
  assign dummy_write_QTree_Bool_sink_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                          demuxWriteResult_QTree_Bool_onehotd[34]};
  assign demuxWriteResult_QTree_Bool_r = (| (demuxWriteResult_QTree_Bool_onehotd & {dummy_write_QTree_Bool_sink_r,
                                                                                    writeQTree_BoollizzieLet9_1_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet7_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet6_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet69_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet64_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet59_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet56_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet55_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet53_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet51_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet50_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet47_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet44_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet43_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet42_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet40_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet3_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet39_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet37_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet36_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet35_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet34_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet31_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet30_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet29_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet28_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet24_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet23_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet19_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet18_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet15_1_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet12_1_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet11_1_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet10_1_1_argbuf_r}));
  assign writeMerge_choice_QTree_Bool_r = demuxWriteResult_QTree_Bool_r;
  
  /* dcon (Ty MemIn_QTree_Bool,
      Dcon WriteIn_QTree_Bool) : [(forkHP1_QTree_Boo3,Word16#),
                                  (writeMerge_data_QTree_Bool,QTree_Bool)] > (dconWriteIn_QTree_Bool,MemIn_QTree_Bool) */
  assign dconWriteIn_QTree_Bool_d = WriteIn_QTree_Bool_dc((& {forkHP1_QTree_Boo3_d[0],
                                                              writeMerge_data_QTree_Bool_d[0]}), forkHP1_QTree_Boo3_d, writeMerge_data_QTree_Bool_d);
  assign {forkHP1_QTree_Boo3_r,
          writeMerge_data_QTree_Bool_r} = {2 {(dconWriteIn_QTree_Bool_r && dconWriteIn_QTree_Bool_d[0])}};
  
  /* dcon (Ty Pointer_QTree_Bool,
      Dcon Pointer_QTree_Bool) : [(forkHP1_QTree_Boo4,Word16#)] > (dconPtr_QTree_Bool,Pointer_QTree_Bool) */
  assign dconPtr_QTree_Bool_d = Pointer_QTree_Bool_dc((& {forkHP1_QTree_Boo4_d[0]}), forkHP1_QTree_Boo4_d);
  assign {forkHP1_QTree_Boo4_r} = {1 {(dconPtr_QTree_Bool_r && dconPtr_QTree_Bool_d[0])}};
  
  /* demux (Ty MemOut_QTree_Bool,
       Ty Pointer_QTree_Bool) : (memWriteOut_QTree_Bool,MemOut_QTree_Bool) (dconPtr_QTree_Bool,Pointer_QTree_Bool) > [(_171,Pointer_QTree_Bool),
                                                                                                                      (demuxWriteResult_QTree_Bool,Pointer_QTree_Bool)] */
  logic [1:0] dconPtr_QTree_Bool_onehotd;
  always_comb
    if ((memWriteOut_QTree_Bool_d[0] && dconPtr_QTree_Bool_d[0]))
      unique case (memWriteOut_QTree_Bool_d[1:1])
        1'd0: dconPtr_QTree_Bool_onehotd = 2'd1;
        1'd1: dconPtr_QTree_Bool_onehotd = 2'd2;
        default: dconPtr_QTree_Bool_onehotd = 2'd0;
      endcase
    else dconPtr_QTree_Bool_onehotd = 2'd0;
  assign _171_d = {dconPtr_QTree_Bool_d[16:1],
                   dconPtr_QTree_Bool_onehotd[0]};
  assign demuxWriteResult_QTree_Bool_d = {dconPtr_QTree_Bool_d[16:1],
                                          dconPtr_QTree_Bool_onehotd[1]};
  assign dconPtr_QTree_Bool_r = (| (dconPtr_QTree_Bool_onehotd & {demuxWriteResult_QTree_Bool_r,
                                                                  _171_r}));
  assign memWriteOut_QTree_Bool_r = dconPtr_QTree_Bool_r;
  
  /* const (Ty Word16#,Lit 0) : (goFor_2,Go) > (initHP_CTf,Word16#) */
  assign initHP_CTf_d = {16'd0, goFor_2_d[0]};
  assign goFor_2_r = initHP_CTf_r;
  
  /* const (Ty Word16#,Lit 1) : (incrHP_CTf1,Go) > (incrHP_CTf,Word16#) */
  assign incrHP_CTf_d = {16'd1, incrHP_CTf1_d[0]};
  assign incrHP_CTf1_r = incrHP_CTf_r;
  
  /* merge (Ty Go) : [(goFor_3,Go),
                 (incrHP_CTf2,Go)] > (incrHP_mergeCTf,Go) */
  logic [1:0] incrHP_mergeCTf_selected;
  logic [1:0] incrHP_mergeCTf_select;
  always_comb
    begin
      incrHP_mergeCTf_selected = 2'd0;
      if ((| incrHP_mergeCTf_select))
        incrHP_mergeCTf_selected = incrHP_mergeCTf_select;
      else
        if (goFor_3_d[0]) incrHP_mergeCTf_selected[0] = 1'd1;
        else if (incrHP_CTf2_d[0]) incrHP_mergeCTf_selected[1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeCTf_select <= 2'd0;
    else
      incrHP_mergeCTf_select <= (incrHP_mergeCTf_r ? 2'd0 :
                                 incrHP_mergeCTf_selected);
  always_comb
    if (incrHP_mergeCTf_selected[0]) incrHP_mergeCTf_d = goFor_3_d;
    else if (incrHP_mergeCTf_selected[1])
      incrHP_mergeCTf_d = incrHP_CTf2_d;
    else incrHP_mergeCTf_d = 1'd0;
  assign {incrHP_CTf2_r,
          goFor_3_r} = (incrHP_mergeCTf_r ? incrHP_mergeCTf_selected :
                        2'd0);
  
  /* fork (Ty Go) : (incrHP_mergeCTf_buf,Go) > [(incrHP_CTf1,Go),
                                           (incrHP_CTf2,Go)] */
  logic [1:0] incrHP_mergeCTf_buf_emitted;
  logic [1:0] incrHP_mergeCTf_buf_done;
  assign incrHP_CTf1_d = (incrHP_mergeCTf_buf_d[0] && (! incrHP_mergeCTf_buf_emitted[0]));
  assign incrHP_CTf2_d = (incrHP_mergeCTf_buf_d[0] && (! incrHP_mergeCTf_buf_emitted[1]));
  assign incrHP_mergeCTf_buf_done = (incrHP_mergeCTf_buf_emitted | ({incrHP_CTf2_d[0],
                                                                     incrHP_CTf1_d[0]} & {incrHP_CTf2_r,
                                                                                          incrHP_CTf1_r}));
  assign incrHP_mergeCTf_buf_r = (& incrHP_mergeCTf_buf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeCTf_buf_emitted <= 2'd0;
    else
      incrHP_mergeCTf_buf_emitted <= (incrHP_mergeCTf_buf_r ? 2'd0 :
                                      incrHP_mergeCTf_buf_done);
  
  /* op_add (Ty Word16#) : (incrHP_CTf,Word16#) (forkHP1_CTf,Word16#) > (addHP_CTf,Word16#) */
  assign addHP_CTf_d = {(incrHP_CTf_d[16:1] + forkHP1_CTf_d[16:1]),
                        (incrHP_CTf_d[0] && forkHP1_CTf_d[0])};
  assign {incrHP_CTf_r,
          forkHP1_CTf_r} = {2 {(addHP_CTf_r && addHP_CTf_d[0])}};
  
  /* merge (Ty Word16#) : [(initHP_CTf,Word16#),
                      (addHP_CTf,Word16#)] > (mergeHP_CTf,Word16#) */
  logic [1:0] mergeHP_CTf_selected;
  logic [1:0] mergeHP_CTf_select;
  always_comb
    begin
      mergeHP_CTf_selected = 2'd0;
      if ((| mergeHP_CTf_select))
        mergeHP_CTf_selected = mergeHP_CTf_select;
      else
        if (initHP_CTf_d[0]) mergeHP_CTf_selected[0] = 1'd1;
        else if (addHP_CTf_d[0]) mergeHP_CTf_selected[1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_CTf_select <= 2'd0;
    else
      mergeHP_CTf_select <= (mergeHP_CTf_r ? 2'd0 :
                             mergeHP_CTf_selected);
  always_comb
    if (mergeHP_CTf_selected[0]) mergeHP_CTf_d = initHP_CTf_d;
    else if (mergeHP_CTf_selected[1]) mergeHP_CTf_d = addHP_CTf_d;
    else mergeHP_CTf_d = {16'd0, 1'd0};
  assign {addHP_CTf_r,
          initHP_CTf_r} = (mergeHP_CTf_r ? mergeHP_CTf_selected :
                           2'd0);
  
  /* buf (Ty Go) : (incrHP_mergeCTf,Go) > (incrHP_mergeCTf_buf,Go) */
  Go_t incrHP_mergeCTf_bufchan_d;
  logic incrHP_mergeCTf_bufchan_r;
  assign incrHP_mergeCTf_r = ((! incrHP_mergeCTf_bufchan_d[0]) || incrHP_mergeCTf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeCTf_bufchan_d <= 1'd0;
    else
      if (incrHP_mergeCTf_r)
        incrHP_mergeCTf_bufchan_d <= incrHP_mergeCTf_d;
  Go_t incrHP_mergeCTf_bufchan_buf;
  assign incrHP_mergeCTf_bufchan_r = (! incrHP_mergeCTf_bufchan_buf[0]);
  assign incrHP_mergeCTf_buf_d = (incrHP_mergeCTf_bufchan_buf[0] ? incrHP_mergeCTf_bufchan_buf :
                                  incrHP_mergeCTf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeCTf_bufchan_buf <= 1'd0;
    else
      if ((incrHP_mergeCTf_buf_r && incrHP_mergeCTf_bufchan_buf[0]))
        incrHP_mergeCTf_bufchan_buf <= 1'd0;
      else if (((! incrHP_mergeCTf_buf_r) && (! incrHP_mergeCTf_bufchan_buf[0])))
        incrHP_mergeCTf_bufchan_buf <= incrHP_mergeCTf_bufchan_d;
  
  /* buf (Ty Word16#) : (mergeHP_CTf,Word16#) > (mergeHP_CTf_buf,Word16#) */
  \Word16#_t  mergeHP_CTf_bufchan_d;
  logic mergeHP_CTf_bufchan_r;
  assign mergeHP_CTf_r = ((! mergeHP_CTf_bufchan_d[0]) || mergeHP_CTf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_CTf_bufchan_d <= {16'd0, 1'd0};
    else if (mergeHP_CTf_r) mergeHP_CTf_bufchan_d <= mergeHP_CTf_d;
  \Word16#_t  mergeHP_CTf_bufchan_buf;
  assign mergeHP_CTf_bufchan_r = (! mergeHP_CTf_bufchan_buf[0]);
  assign mergeHP_CTf_buf_d = (mergeHP_CTf_bufchan_buf[0] ? mergeHP_CTf_bufchan_buf :
                              mergeHP_CTf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_CTf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((mergeHP_CTf_buf_r && mergeHP_CTf_bufchan_buf[0]))
        mergeHP_CTf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! mergeHP_CTf_buf_r) && (! mergeHP_CTf_bufchan_buf[0])))
        mergeHP_CTf_bufchan_buf <= mergeHP_CTf_bufchan_d;
  
  /* fork (Ty Word16#) : (mergeHP_CTf_buf,Word16#) > [(forkHP1_CTf,Word16#),
                                                 (forkHP1_CT2,Word16#),
                                                 (forkHP1_CT3,Word16#)] */
  logic [2:0] mergeHP_CTf_buf_emitted;
  logic [2:0] mergeHP_CTf_buf_done;
  assign forkHP1_CTf_d = {mergeHP_CTf_buf_d[16:1],
                          (mergeHP_CTf_buf_d[0] && (! mergeHP_CTf_buf_emitted[0]))};
  assign forkHP1_CT2_d = {mergeHP_CTf_buf_d[16:1],
                          (mergeHP_CTf_buf_d[0] && (! mergeHP_CTf_buf_emitted[1]))};
  assign forkHP1_CT3_d = {mergeHP_CTf_buf_d[16:1],
                          (mergeHP_CTf_buf_d[0] && (! mergeHP_CTf_buf_emitted[2]))};
  assign mergeHP_CTf_buf_done = (mergeHP_CTf_buf_emitted | ({forkHP1_CT3_d[0],
                                                             forkHP1_CT2_d[0],
                                                             forkHP1_CTf_d[0]} & {forkHP1_CT3_r,
                                                                                  forkHP1_CT2_r,
                                                                                  forkHP1_CTf_r}));
  assign mergeHP_CTf_buf_r = (& mergeHP_CTf_buf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_CTf_buf_emitted <= 3'd0;
    else
      mergeHP_CTf_buf_emitted <= (mergeHP_CTf_buf_r ? 3'd0 :
                                  mergeHP_CTf_buf_done);
  
  /* mergectrl (Ty C2,Ty MemIn_CTf) : [(dconReadIn_CTf,MemIn_CTf),
                                  (dconWriteIn_CTf,MemIn_CTf)] > (memMergeChoice_CTf,C2) (memMergeIn_CTf,MemIn_CTf) */
  logic [1:0] dconReadIn_CTf_select_d;
  assign dconReadIn_CTf_select_d = ((| dconReadIn_CTf_select_q) ? dconReadIn_CTf_select_q :
                                    (dconReadIn_CTf_d[0] ? 2'd1 :
                                     (dconWriteIn_CTf_d[0] ? 2'd2 :
                                      2'd0)));
  logic [1:0] dconReadIn_CTf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) dconReadIn_CTf_select_q <= 2'd0;
    else
      dconReadIn_CTf_select_q <= (dconReadIn_CTf_done ? 2'd0 :
                                  dconReadIn_CTf_select_d);
  logic [1:0] dconReadIn_CTf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) dconReadIn_CTf_emit_q <= 2'd0;
    else
      dconReadIn_CTf_emit_q <= (dconReadIn_CTf_done ? 2'd0 :
                                dconReadIn_CTf_emit_d);
  logic [1:0] dconReadIn_CTf_emit_d;
  assign dconReadIn_CTf_emit_d = (dconReadIn_CTf_emit_q | ({memMergeChoice_CTf_d[0],
                                                            memMergeIn_CTf_d[0]} & {memMergeChoice_CTf_r,
                                                                                    memMergeIn_CTf_r}));
  logic dconReadIn_CTf_done;
  assign dconReadIn_CTf_done = (& dconReadIn_CTf_emit_d);
  assign {dconWriteIn_CTf_r,
          dconReadIn_CTf_r} = (dconReadIn_CTf_done ? dconReadIn_CTf_select_d :
                               2'd0);
  assign memMergeIn_CTf_d = ((dconReadIn_CTf_select_d[0] && (! dconReadIn_CTf_emit_q[0])) ? dconReadIn_CTf_d :
                             ((dconReadIn_CTf_select_d[1] && (! dconReadIn_CTf_emit_q[0])) ? dconWriteIn_CTf_d :
                              {180'd0, 1'd0}));
  assign memMergeChoice_CTf_d = ((dconReadIn_CTf_select_d[0] && (! dconReadIn_CTf_emit_q[1])) ? C1_2_dc(1'd1) :
                                 ((dconReadIn_CTf_select_d[1] && (! dconReadIn_CTf_emit_q[1])) ? C2_2_dc(1'd1) :
                                  {1'd0, 1'd0}));
  
  /* bram (Ty MemIn_CTf,
      Ty MemOut_CTf) : (memMergeIn_CTf_dbuf,MemIn_CTf) > (memOut_CTf,MemOut_CTf) */
  logic [162:0] memMergeIn_CTf_dbuf_mem[65535:0];
  logic [15:0] memMergeIn_CTf_dbuf_address;
  logic [162:0] memMergeIn_CTf_dbuf_din;
  logic [162:0] memOut_CTf_q;
  logic memOut_CTf_valid;
  logic memMergeIn_CTf_dbuf_we;
  logic memOut_CTf_we;
  assign memMergeIn_CTf_dbuf_din = memMergeIn_CTf_dbuf_d[180:18];
  assign memMergeIn_CTf_dbuf_address = memMergeIn_CTf_dbuf_d[17:2];
  assign memMergeIn_CTf_dbuf_we = (memMergeIn_CTf_dbuf_d[1:1] && memMergeIn_CTf_dbuf_d[0]);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        memOut_CTf_we <= 1'd0;
        memOut_CTf_valid <= 1'd0;
      end
    else
      begin
        memOut_CTf_we <= memMergeIn_CTf_dbuf_we;
        memOut_CTf_valid <= memMergeIn_CTf_dbuf_d[0];
        if (memMergeIn_CTf_dbuf_we)
          begin
            memMergeIn_CTf_dbuf_mem[memMergeIn_CTf_dbuf_address] <= memMergeIn_CTf_dbuf_din;
            memOut_CTf_q <= memMergeIn_CTf_dbuf_din;
          end
        else
          memOut_CTf_q <= memMergeIn_CTf_dbuf_mem[memMergeIn_CTf_dbuf_address];
      end
  assign memOut_CTf_d = {memOut_CTf_q,
                         memOut_CTf_we,
                         memOut_CTf_valid};
  assign memMergeIn_CTf_dbuf_r = ((! memOut_CTf_valid) || memOut_CTf_r);
  logic [31:0] profiling_MemIn_CTf_read;
  logic [31:0] profiling_MemIn_CTf_write;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        profiling_MemIn_CTf_write <= 0;
        profiling_MemIn_CTf_read <= 0;
      end
    else
      if ((memMergeIn_CTf_dbuf_we == 1'd1))
        profiling_MemIn_CTf_write <= (profiling_MemIn_CTf_write + 1);
      else
        if ((memOut_CTf_valid == 1'd1))
          profiling_MemIn_CTf_read <= (profiling_MemIn_CTf_read + 1);
  
  /* demux (Ty C2,
       Ty MemOut_CTf) : (memMergeChoice_CTf,C2) (memOut_CTf_dbuf,MemOut_CTf) > [(memReadOut_CTf,MemOut_CTf),
                                                                                (memWriteOut_CTf,MemOut_CTf)] */
  logic [1:0] memOut_CTf_dbuf_onehotd;
  always_comb
    if ((memMergeChoice_CTf_d[0] && memOut_CTf_dbuf_d[0]))
      unique case (memMergeChoice_CTf_d[1:1])
        1'd0: memOut_CTf_dbuf_onehotd = 2'd1;
        1'd1: memOut_CTf_dbuf_onehotd = 2'd2;
        default: memOut_CTf_dbuf_onehotd = 2'd0;
      endcase
    else memOut_CTf_dbuf_onehotd = 2'd0;
  assign memReadOut_CTf_d = {memOut_CTf_dbuf_d[164:1],
                             memOut_CTf_dbuf_onehotd[0]};
  assign memWriteOut_CTf_d = {memOut_CTf_dbuf_d[164:1],
                              memOut_CTf_dbuf_onehotd[1]};
  assign memOut_CTf_dbuf_r = (| (memOut_CTf_dbuf_onehotd & {memWriteOut_CTf_r,
                                                            memReadOut_CTf_r}));
  assign memMergeChoice_CTf_r = memOut_CTf_dbuf_r;
  
  /* dbuf (Ty MemIn_CTf) : (memMergeIn_CTf_rbuf,MemIn_CTf) > (memMergeIn_CTf_dbuf,MemIn_CTf) */
  assign memMergeIn_CTf_rbuf_r = ((! memMergeIn_CTf_dbuf_d[0]) || memMergeIn_CTf_dbuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memMergeIn_CTf_dbuf_d <= {180'd0, 1'd0};
    else
      if (memMergeIn_CTf_rbuf_r)
        memMergeIn_CTf_dbuf_d <= memMergeIn_CTf_rbuf_d;
  
  /* rbuf (Ty MemIn_CTf) : (memMergeIn_CTf,MemIn_CTf) > (memMergeIn_CTf_rbuf,MemIn_CTf) */
  MemIn_CTf_t memMergeIn_CTf_buf;
  assign memMergeIn_CTf_r = (! memMergeIn_CTf_buf[0]);
  assign memMergeIn_CTf_rbuf_d = (memMergeIn_CTf_buf[0] ? memMergeIn_CTf_buf :
                                  memMergeIn_CTf_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memMergeIn_CTf_buf <= {180'd0, 1'd0};
    else
      if ((memMergeIn_CTf_rbuf_r && memMergeIn_CTf_buf[0]))
        memMergeIn_CTf_buf <= {180'd0, 1'd0};
      else if (((! memMergeIn_CTf_rbuf_r) && (! memMergeIn_CTf_buf[0])))
        memMergeIn_CTf_buf <= memMergeIn_CTf_d;
  
  /* dbuf (Ty MemOut_CTf) : (memOut_CTf_rbuf,MemOut_CTf) > (memOut_CTf_dbuf,MemOut_CTf) */
  assign memOut_CTf_rbuf_r = ((! memOut_CTf_dbuf_d[0]) || memOut_CTf_dbuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memOut_CTf_dbuf_d <= {164'd0, 1'd0};
    else if (memOut_CTf_rbuf_r) memOut_CTf_dbuf_d <= memOut_CTf_rbuf_d;
  
  /* rbuf (Ty MemOut_CTf) : (memOut_CTf,MemOut_CTf) > (memOut_CTf_rbuf,MemOut_CTf) */
  MemOut_CTf_t memOut_CTf_buf;
  assign memOut_CTf_r = (! memOut_CTf_buf[0]);
  assign memOut_CTf_rbuf_d = (memOut_CTf_buf[0] ? memOut_CTf_buf :
                              memOut_CTf_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memOut_CTf_buf <= {164'd0, 1'd0};
    else
      if ((memOut_CTf_rbuf_r && memOut_CTf_buf[0]))
        memOut_CTf_buf <= {164'd0, 1'd0};
      else if (((! memOut_CTf_rbuf_r) && (! memOut_CTf_buf[0])))
        memOut_CTf_buf <= memOut_CTf_d;
  
  /* destruct (Ty Pointer_CTf,
          Dcon Pointer_CTf) : (scfarg_0_1_argbuf,Pointer_CTf) > [(destructReadIn_CTf,Word16#)] */
  assign destructReadIn_CTf_d = {scfarg_0_1_argbuf_d[16:1],
                                 scfarg_0_1_argbuf_d[0]};
  assign scfarg_0_1_argbuf_r = destructReadIn_CTf_r;
  
  /* dcon (Ty MemIn_CTf,
      Dcon ReadIn_CTf) : [(destructReadIn_CTf,Word16#)] > (dconReadIn_CTf,MemIn_CTf) */
  assign dconReadIn_CTf_d = ReadIn_CTf_dc((& {destructReadIn_CTf_d[0]}), destructReadIn_CTf_d);
  assign {destructReadIn_CTf_r} = {1 {(dconReadIn_CTf_r && dconReadIn_CTf_d[0])}};
  
  /* destruct (Ty MemOut_CTf,
          Dcon ReadOut_CTf) : (memReadOut_CTf,MemOut_CTf) > [(readPointer_CTfscfarg_0_1_argbuf,CTf)] */
  assign readPointer_CTfscfarg_0_1_argbuf_d = {memReadOut_CTf_d[164:2],
                                               memReadOut_CTf_d[0]};
  assign memReadOut_CTf_r = readPointer_CTfscfarg_0_1_argbuf_r;
  
  /* mergectrl (Ty C5,Ty CTf) : [(lizzieLet41_1_argbuf,CTf),
                            (lizzieLet57_1_argbuf,CTf),
                            (lizzieLet61_1_argbuf,CTf),
                            (lizzieLet62_1_argbuf,CTf),
                            (lizzieLet63_1_argbuf,CTf)] > (writeMerge_choice_CTf,C5) (writeMerge_data_CTf,CTf) */
  logic [4:0] lizzieLet41_1_argbuf_select_d;
  assign lizzieLet41_1_argbuf_select_d = ((| lizzieLet41_1_argbuf_select_q) ? lizzieLet41_1_argbuf_select_q :
                                          (lizzieLet41_1_argbuf_d[0] ? 5'd1 :
                                           (lizzieLet57_1_argbuf_d[0] ? 5'd2 :
                                            (lizzieLet61_1_argbuf_d[0] ? 5'd4 :
                                             (lizzieLet62_1_argbuf_d[0] ? 5'd8 :
                                              (lizzieLet63_1_argbuf_d[0] ? 5'd16 :
                                               5'd0))))));
  logic [4:0] lizzieLet41_1_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet41_1_argbuf_select_q <= 5'd0;
    else
      lizzieLet41_1_argbuf_select_q <= (lizzieLet41_1_argbuf_done ? 5'd0 :
                                        lizzieLet41_1_argbuf_select_d);
  logic [1:0] lizzieLet41_1_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet41_1_argbuf_emit_q <= 2'd0;
    else
      lizzieLet41_1_argbuf_emit_q <= (lizzieLet41_1_argbuf_done ? 2'd0 :
                                      lizzieLet41_1_argbuf_emit_d);
  logic [1:0] lizzieLet41_1_argbuf_emit_d;
  assign lizzieLet41_1_argbuf_emit_d = (lizzieLet41_1_argbuf_emit_q | ({writeMerge_choice_CTf_d[0],
                                                                        writeMerge_data_CTf_d[0]} & {writeMerge_choice_CTf_r,
                                                                                                     writeMerge_data_CTf_r}));
  logic lizzieLet41_1_argbuf_done;
  assign lizzieLet41_1_argbuf_done = (& lizzieLet41_1_argbuf_emit_d);
  assign {lizzieLet63_1_argbuf_r,
          lizzieLet62_1_argbuf_r,
          lizzieLet61_1_argbuf_r,
          lizzieLet57_1_argbuf_r,
          lizzieLet41_1_argbuf_r} = (lizzieLet41_1_argbuf_done ? lizzieLet41_1_argbuf_select_d :
                                     5'd0);
  assign writeMerge_data_CTf_d = ((lizzieLet41_1_argbuf_select_d[0] && (! lizzieLet41_1_argbuf_emit_q[0])) ? lizzieLet41_1_argbuf_d :
                                  ((lizzieLet41_1_argbuf_select_d[1] && (! lizzieLet41_1_argbuf_emit_q[0])) ? lizzieLet57_1_argbuf_d :
                                   ((lizzieLet41_1_argbuf_select_d[2] && (! lizzieLet41_1_argbuf_emit_q[0])) ? lizzieLet61_1_argbuf_d :
                                    ((lizzieLet41_1_argbuf_select_d[3] && (! lizzieLet41_1_argbuf_emit_q[0])) ? lizzieLet62_1_argbuf_d :
                                     ((lizzieLet41_1_argbuf_select_d[4] && (! lizzieLet41_1_argbuf_emit_q[0])) ? lizzieLet63_1_argbuf_d :
                                      {163'd0, 1'd0})))));
  assign writeMerge_choice_CTf_d = ((lizzieLet41_1_argbuf_select_d[0] && (! lizzieLet41_1_argbuf_emit_q[1])) ? C1_5_dc(1'd1) :
                                    ((lizzieLet41_1_argbuf_select_d[1] && (! lizzieLet41_1_argbuf_emit_q[1])) ? C2_5_dc(1'd1) :
                                     ((lizzieLet41_1_argbuf_select_d[2] && (! lizzieLet41_1_argbuf_emit_q[1])) ? C3_5_dc(1'd1) :
                                      ((lizzieLet41_1_argbuf_select_d[3] && (! lizzieLet41_1_argbuf_emit_q[1])) ? C4_5_dc(1'd1) :
                                       ((lizzieLet41_1_argbuf_select_d[4] && (! lizzieLet41_1_argbuf_emit_q[1])) ? C5_5_dc(1'd1) :
                                        {3'd0, 1'd0})))));
  
  /* demux (Ty C5,
       Ty Pointer_CTf) : (writeMerge_choice_CTf,C5) (demuxWriteResult_CTf,Pointer_CTf) > [(writeCTflizzieLet41_1_argbuf,Pointer_CTf),
                                                                                          (writeCTflizzieLet57_1_argbuf,Pointer_CTf),
                                                                                          (writeCTflizzieLet61_1_argbuf,Pointer_CTf),
                                                                                          (writeCTflizzieLet62_1_argbuf,Pointer_CTf),
                                                                                          (writeCTflizzieLet63_1_argbuf,Pointer_CTf)] */
  logic [4:0] demuxWriteResult_CTf_onehotd;
  always_comb
    if ((writeMerge_choice_CTf_d[0] && demuxWriteResult_CTf_d[0]))
      unique case (writeMerge_choice_CTf_d[3:1])
        3'd0: demuxWriteResult_CTf_onehotd = 5'd1;
        3'd1: demuxWriteResult_CTf_onehotd = 5'd2;
        3'd2: demuxWriteResult_CTf_onehotd = 5'd4;
        3'd3: demuxWriteResult_CTf_onehotd = 5'd8;
        3'd4: demuxWriteResult_CTf_onehotd = 5'd16;
        default: demuxWriteResult_CTf_onehotd = 5'd0;
      endcase
    else demuxWriteResult_CTf_onehotd = 5'd0;
  assign writeCTflizzieLet41_1_argbuf_d = {demuxWriteResult_CTf_d[16:1],
                                           demuxWriteResult_CTf_onehotd[0]};
  assign writeCTflizzieLet57_1_argbuf_d = {demuxWriteResult_CTf_d[16:1],
                                           demuxWriteResult_CTf_onehotd[1]};
  assign writeCTflizzieLet61_1_argbuf_d = {demuxWriteResult_CTf_d[16:1],
                                           demuxWriteResult_CTf_onehotd[2]};
  assign writeCTflizzieLet62_1_argbuf_d = {demuxWriteResult_CTf_d[16:1],
                                           demuxWriteResult_CTf_onehotd[3]};
  assign writeCTflizzieLet63_1_argbuf_d = {demuxWriteResult_CTf_d[16:1],
                                           demuxWriteResult_CTf_onehotd[4]};
  assign demuxWriteResult_CTf_r = (| (demuxWriteResult_CTf_onehotd & {writeCTflizzieLet63_1_argbuf_r,
                                                                      writeCTflizzieLet62_1_argbuf_r,
                                                                      writeCTflizzieLet61_1_argbuf_r,
                                                                      writeCTflizzieLet57_1_argbuf_r,
                                                                      writeCTflizzieLet41_1_argbuf_r}));
  assign writeMerge_choice_CTf_r = demuxWriteResult_CTf_r;
  
  /* dcon (Ty MemIn_CTf,Dcon WriteIn_CTf) : [(forkHP1_CT2,Word16#),
                                        (writeMerge_data_CTf,CTf)] > (dconWriteIn_CTf,MemIn_CTf) */
  assign dconWriteIn_CTf_d = WriteIn_CTf_dc((& {forkHP1_CT2_d[0],
                                                writeMerge_data_CTf_d[0]}), forkHP1_CT2_d, writeMerge_data_CTf_d);
  assign {forkHP1_CT2_r,
          writeMerge_data_CTf_r} = {2 {(dconWriteIn_CTf_r && dconWriteIn_CTf_d[0])}};
  
  /* dcon (Ty Pointer_CTf,
      Dcon Pointer_CTf) : [(forkHP1_CT3,Word16#)] > (dconPtr_CTf,Pointer_CTf) */
  assign dconPtr_CTf_d = Pointer_CTf_dc((& {forkHP1_CT3_d[0]}), forkHP1_CT3_d);
  assign {forkHP1_CT3_r} = {1 {(dconPtr_CTf_r && dconPtr_CTf_d[0])}};
  
  /* demux (Ty MemOut_CTf,
       Ty Pointer_CTf) : (memWriteOut_CTf,MemOut_CTf) (dconPtr_CTf,Pointer_CTf) > [(_170,Pointer_CTf),
                                                                                   (demuxWriteResult_CTf,Pointer_CTf)] */
  logic [1:0] dconPtr_CTf_onehotd;
  always_comb
    if ((memWriteOut_CTf_d[0] && dconPtr_CTf_d[0]))
      unique case (memWriteOut_CTf_d[1:1])
        1'd0: dconPtr_CTf_onehotd = 2'd1;
        1'd1: dconPtr_CTf_onehotd = 2'd2;
        default: dconPtr_CTf_onehotd = 2'd0;
      endcase
    else dconPtr_CTf_onehotd = 2'd0;
  assign _170_d = {dconPtr_CTf_d[16:1], dconPtr_CTf_onehotd[0]};
  assign demuxWriteResult_CTf_d = {dconPtr_CTf_d[16:1],
                                   dconPtr_CTf_onehotd[1]};
  assign dconPtr_CTf_r = (| (dconPtr_CTf_onehotd & {demuxWriteResult_CTf_r,
                                                    _170_r}));
  assign memWriteOut_CTf_r = dconPtr_CTf_r;
  
  /* const (Ty Word16#,
       Lit 0) : (goFor_4,Go) > (initHP_CTf'''''''''''',Word16#) */
  assign \initHP_CTf''''''''''''_d  = {16'd0, goFor_4_d[0]};
  assign goFor_4_r = \initHP_CTf''''''''''''_r ;
  
  /* const (Ty Word16#,
       Lit 1) : (incrHP_CTf''''''''''''1,Go) > (incrHP_CTf'''''''''''',Word16#) */
  assign \incrHP_CTf''''''''''''_d  = {16'd1,
                                       \incrHP_CTf''''''''''''1_d [0]};
  assign \incrHP_CTf''''''''''''1_r  = \incrHP_CTf''''''''''''_r ;
  
  /* merge (Ty Go) : [(goFor_5,Go),
                 (incrHP_CTf''''''''''''2,Go)] > (incrHP_mergeCTf'''''''''''',Go) */
  logic [1:0] \incrHP_mergeCTf''''''''''''_selected ;
  logic [1:0] \incrHP_mergeCTf''''''''''''_select ;
  always_comb
    begin
      \incrHP_mergeCTf''''''''''''_selected  = 2'd0;
      if ((| \incrHP_mergeCTf''''''''''''_select ))
        \incrHP_mergeCTf''''''''''''_selected  = \incrHP_mergeCTf''''''''''''_select ;
      else
        if (goFor_5_d[0]) \incrHP_mergeCTf''''''''''''_selected [0] = 1'd1;
        else if (\incrHP_CTf''''''''''''2_d [0])
          \incrHP_mergeCTf''''''''''''_selected [1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \incrHP_mergeCTf''''''''''''_select  <= 2'd0;
    else
      \incrHP_mergeCTf''''''''''''_select  <= (\incrHP_mergeCTf''''''''''''_r  ? 2'd0 :
                                               \incrHP_mergeCTf''''''''''''_selected );
  always_comb
    if (\incrHP_mergeCTf''''''''''''_selected [0])
      \incrHP_mergeCTf''''''''''''_d  = goFor_5_d;
    else if (\incrHP_mergeCTf''''''''''''_selected [1])
      \incrHP_mergeCTf''''''''''''_d  = \incrHP_CTf''''''''''''2_d ;
    else \incrHP_mergeCTf''''''''''''_d  = 1'd0;
  assign {\incrHP_CTf''''''''''''2_r ,
          goFor_5_r} = (\incrHP_mergeCTf''''''''''''_r  ? \incrHP_mergeCTf''''''''''''_selected  :
                        2'd0);
  
  /* fork (Ty Go) : (incrHP_mergeCTf''''''''''''_buf,Go) > [(incrHP_CTf''''''''''''1,Go),
                                                       (incrHP_CTf''''''''''''2,Go)] */
  logic [1:0] \incrHP_mergeCTf''''''''''''_buf_emitted ;
  logic [1:0] \incrHP_mergeCTf''''''''''''_buf_done ;
  assign \incrHP_CTf''''''''''''1_d  = (\incrHP_mergeCTf''''''''''''_buf_d [0] && (! \incrHP_mergeCTf''''''''''''_buf_emitted [0]));
  assign \incrHP_CTf''''''''''''2_d  = (\incrHP_mergeCTf''''''''''''_buf_d [0] && (! \incrHP_mergeCTf''''''''''''_buf_emitted [1]));
  assign \incrHP_mergeCTf''''''''''''_buf_done  = (\incrHP_mergeCTf''''''''''''_buf_emitted  | ({\incrHP_CTf''''''''''''2_d [0],
                                                                                                 \incrHP_CTf''''''''''''1_d [0]} & {\incrHP_CTf''''''''''''2_r ,
                                                                                                                                    \incrHP_CTf''''''''''''1_r }));
  assign \incrHP_mergeCTf''''''''''''_buf_r  = (& \incrHP_mergeCTf''''''''''''_buf_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \incrHP_mergeCTf''''''''''''_buf_emitted  <= 2'd0;
    else
      \incrHP_mergeCTf''''''''''''_buf_emitted  <= (\incrHP_mergeCTf''''''''''''_buf_r  ? 2'd0 :
                                                    \incrHP_mergeCTf''''''''''''_buf_done );
  
  /* op_add (Ty Word16#) : (incrHP_CTf'''''''''''',Word16#) (forkHP1_CTf'''''''''''',Word16#) > (addHP_CTf'''''''''''',Word16#) */
  assign \addHP_CTf''''''''''''_d  = {(\incrHP_CTf''''''''''''_d [16:1] + \forkHP1_CTf''''''''''''_d [16:1]),
                                      (\incrHP_CTf''''''''''''_d [0] && \forkHP1_CTf''''''''''''_d [0])};
  assign {\incrHP_CTf''''''''''''_r ,
          \forkHP1_CTf''''''''''''_r } = {2 {(\addHP_CTf''''''''''''_r  && \addHP_CTf''''''''''''_d [0])}};
  
  /* merge (Ty Word16#) : [(initHP_CTf'''''''''''',Word16#),
                      (addHP_CTf'''''''''''',Word16#)] > (mergeHP_CTf'''''''''''',Word16#) */
  logic [1:0] \mergeHP_CTf''''''''''''_selected ;
  logic [1:0] \mergeHP_CTf''''''''''''_select ;
  always_comb
    begin
      \mergeHP_CTf''''''''''''_selected  = 2'd0;
      if ((| \mergeHP_CTf''''''''''''_select ))
        \mergeHP_CTf''''''''''''_selected  = \mergeHP_CTf''''''''''''_select ;
      else
        if (\initHP_CTf''''''''''''_d [0])
          \mergeHP_CTf''''''''''''_selected [0] = 1'd1;
        else if (\addHP_CTf''''''''''''_d [0])
          \mergeHP_CTf''''''''''''_selected [1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \mergeHP_CTf''''''''''''_select  <= 2'd0;
    else
      \mergeHP_CTf''''''''''''_select  <= (\mergeHP_CTf''''''''''''_r  ? 2'd0 :
                                           \mergeHP_CTf''''''''''''_selected );
  always_comb
    if (\mergeHP_CTf''''''''''''_selected [0])
      \mergeHP_CTf''''''''''''_d  = \initHP_CTf''''''''''''_d ;
    else if (\mergeHP_CTf''''''''''''_selected [1])
      \mergeHP_CTf''''''''''''_d  = \addHP_CTf''''''''''''_d ;
    else \mergeHP_CTf''''''''''''_d  = {16'd0, 1'd0};
  assign {\addHP_CTf''''''''''''_r ,
          \initHP_CTf''''''''''''_r } = (\mergeHP_CTf''''''''''''_r  ? \mergeHP_CTf''''''''''''_selected  :
                                         2'd0);
  
  /* buf (Ty Go) : (incrHP_mergeCTf'''''''''''',Go) > (incrHP_mergeCTf''''''''''''_buf,Go) */
  Go_t \incrHP_mergeCTf''''''''''''_bufchan_d ;
  logic \incrHP_mergeCTf''''''''''''_bufchan_r ;
  assign \incrHP_mergeCTf''''''''''''_r  = ((! \incrHP_mergeCTf''''''''''''_bufchan_d [0]) || \incrHP_mergeCTf''''''''''''_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \incrHP_mergeCTf''''''''''''_bufchan_d  <= 1'd0;
    else
      if (\incrHP_mergeCTf''''''''''''_r )
        \incrHP_mergeCTf''''''''''''_bufchan_d  <= \incrHP_mergeCTf''''''''''''_d ;
  Go_t \incrHP_mergeCTf''''''''''''_bufchan_buf ;
  assign \incrHP_mergeCTf''''''''''''_bufchan_r  = (! \incrHP_mergeCTf''''''''''''_bufchan_buf [0]);
  assign \incrHP_mergeCTf''''''''''''_buf_d  = (\incrHP_mergeCTf''''''''''''_bufchan_buf [0] ? \incrHP_mergeCTf''''''''''''_bufchan_buf  :
                                                \incrHP_mergeCTf''''''''''''_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \incrHP_mergeCTf''''''''''''_bufchan_buf  <= 1'd0;
    else
      if ((\incrHP_mergeCTf''''''''''''_buf_r  && \incrHP_mergeCTf''''''''''''_bufchan_buf [0]))
        \incrHP_mergeCTf''''''''''''_bufchan_buf  <= 1'd0;
      else if (((! \incrHP_mergeCTf''''''''''''_buf_r ) && (! \incrHP_mergeCTf''''''''''''_bufchan_buf [0])))
        \incrHP_mergeCTf''''''''''''_bufchan_buf  <= \incrHP_mergeCTf''''''''''''_bufchan_d ;
  
  /* buf (Ty Word16#) : (mergeHP_CTf'''''''''''',Word16#) > (mergeHP_CTf''''''''''''_buf,Word16#) */
  \Word16#_t  \mergeHP_CTf''''''''''''_bufchan_d ;
  logic \mergeHP_CTf''''''''''''_bufchan_r ;
  assign \mergeHP_CTf''''''''''''_r  = ((! \mergeHP_CTf''''''''''''_bufchan_d [0]) || \mergeHP_CTf''''''''''''_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \mergeHP_CTf''''''''''''_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\mergeHP_CTf''''''''''''_r )
        \mergeHP_CTf''''''''''''_bufchan_d  <= \mergeHP_CTf''''''''''''_d ;
  \Word16#_t  \mergeHP_CTf''''''''''''_bufchan_buf ;
  assign \mergeHP_CTf''''''''''''_bufchan_r  = (! \mergeHP_CTf''''''''''''_bufchan_buf [0]);
  assign \mergeHP_CTf''''''''''''_buf_d  = (\mergeHP_CTf''''''''''''_bufchan_buf [0] ? \mergeHP_CTf''''''''''''_bufchan_buf  :
                                            \mergeHP_CTf''''''''''''_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \mergeHP_CTf''''''''''''_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((\mergeHP_CTf''''''''''''_buf_r  && \mergeHP_CTf''''''''''''_bufchan_buf [0]))
        \mergeHP_CTf''''''''''''_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! \mergeHP_CTf''''''''''''_buf_r ) && (! \mergeHP_CTf''''''''''''_bufchan_buf [0])))
        \mergeHP_CTf''''''''''''_bufchan_buf  <= \mergeHP_CTf''''''''''''_bufchan_d ;
  
  /* fork (Ty Word16#) : (mergeHP_CTf''''''''''''_buf,Word16#) > [(forkHP1_CTf'''''''''''',Word16#),
                                                             (forkHP1_CTf'''''''''''2,Word16#),
                                                             (forkHP1_CTf'''''''''''3,Word16#)] */
  logic [2:0] \mergeHP_CTf''''''''''''_buf_emitted ;
  logic [2:0] \mergeHP_CTf''''''''''''_buf_done ;
  assign \forkHP1_CTf''''''''''''_d  = {\mergeHP_CTf''''''''''''_buf_d [16:1],
                                        (\mergeHP_CTf''''''''''''_buf_d [0] && (! \mergeHP_CTf''''''''''''_buf_emitted [0]))};
  assign \forkHP1_CTf'''''''''''2_d  = {\mergeHP_CTf''''''''''''_buf_d [16:1],
                                        (\mergeHP_CTf''''''''''''_buf_d [0] && (! \mergeHP_CTf''''''''''''_buf_emitted [1]))};
  assign \forkHP1_CTf'''''''''''3_d  = {\mergeHP_CTf''''''''''''_buf_d [16:1],
                                        (\mergeHP_CTf''''''''''''_buf_d [0] && (! \mergeHP_CTf''''''''''''_buf_emitted [2]))};
  assign \mergeHP_CTf''''''''''''_buf_done  = (\mergeHP_CTf''''''''''''_buf_emitted  | ({\forkHP1_CTf'''''''''''3_d [0],
                                                                                         \forkHP1_CTf'''''''''''2_d [0],
                                                                                         \forkHP1_CTf''''''''''''_d [0]} & {\forkHP1_CTf'''''''''''3_r ,
                                                                                                                            \forkHP1_CTf'''''''''''2_r ,
                                                                                                                            \forkHP1_CTf''''''''''''_r }));
  assign \mergeHP_CTf''''''''''''_buf_r  = (& \mergeHP_CTf''''''''''''_buf_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \mergeHP_CTf''''''''''''_buf_emitted  <= 3'd0;
    else
      \mergeHP_CTf''''''''''''_buf_emitted  <= (\mergeHP_CTf''''''''''''_buf_r  ? 3'd0 :
                                                \mergeHP_CTf''''''''''''_buf_done );
  
  /* mergectrl (Ty C2,
           Ty MemIn_CTf'''''''''''') : [(dconReadIn_CTf'''''''''''',MemIn_CTf''''''''''''),
                                        (dconWriteIn_CTf'''''''''''',MemIn_CTf'''''''''''')] > (memMergeChoice_CTf'''''''''''',C2) (memMergeIn_CTf'''''''''''',MemIn_CTf'''''''''''') */
  logic [1:0] \dconReadIn_CTf''''''''''''_select_d ;
  assign \dconReadIn_CTf''''''''''''_select_d  = ((| \dconReadIn_CTf''''''''''''_select_q ) ? \dconReadIn_CTf''''''''''''_select_q  :
                                                  (\dconReadIn_CTf''''''''''''_d [0] ? 2'd1 :
                                                   (\dconWriteIn_CTf''''''''''''_d [0] ? 2'd2 :
                                                    2'd0)));
  logic [1:0] \dconReadIn_CTf''''''''''''_select_q ;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \dconReadIn_CTf''''''''''''_select_q  <= 2'd0;
    else
      \dconReadIn_CTf''''''''''''_select_q  <= (\dconReadIn_CTf''''''''''''_done  ? 2'd0 :
                                                \dconReadIn_CTf''''''''''''_select_d );
  logic [1:0] \dconReadIn_CTf''''''''''''_emit_q ;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \dconReadIn_CTf''''''''''''_emit_q  <= 2'd0;
    else
      \dconReadIn_CTf''''''''''''_emit_q  <= (\dconReadIn_CTf''''''''''''_done  ? 2'd0 :
                                              \dconReadIn_CTf''''''''''''_emit_d );
  logic [1:0] \dconReadIn_CTf''''''''''''_emit_d ;
  assign \dconReadIn_CTf''''''''''''_emit_d  = (\dconReadIn_CTf''''''''''''_emit_q  | ({\memMergeChoice_CTf''''''''''''_d [0],
                                                                                        \memMergeIn_CTf''''''''''''_d [0]} & {\memMergeChoice_CTf''''''''''''_r ,
                                                                                                                              \memMergeIn_CTf''''''''''''_r }));
  logic \dconReadIn_CTf''''''''''''_done ;
  assign \dconReadIn_CTf''''''''''''_done  = (& \dconReadIn_CTf''''''''''''_emit_d );
  assign {\dconWriteIn_CTf''''''''''''_r ,
          \dconReadIn_CTf''''''''''''_r } = (\dconReadIn_CTf''''''''''''_done  ? \dconReadIn_CTf''''''''''''_select_d  :
                                             2'd0);
  assign \memMergeIn_CTf''''''''''''_d  = ((\dconReadIn_CTf''''''''''''_select_d [0] && (! \dconReadIn_CTf''''''''''''_emit_q [0])) ? \dconReadIn_CTf''''''''''''_d  :
                                           ((\dconReadIn_CTf''''''''''''_select_d [1] && (! \dconReadIn_CTf''''''''''''_emit_q [0])) ? \dconWriteIn_CTf''''''''''''_d  :
                                            {132'd0, 1'd0}));
  assign \memMergeChoice_CTf''''''''''''_d  = ((\dconReadIn_CTf''''''''''''_select_d [0] && (! \dconReadIn_CTf''''''''''''_emit_q [1])) ? C1_2_dc(1'd1) :
                                               ((\dconReadIn_CTf''''''''''''_select_d [1] && (! \dconReadIn_CTf''''''''''''_emit_q [1])) ? C2_2_dc(1'd1) :
                                                {1'd0, 1'd0}));
  
  /* bram (Ty MemIn_CTf'''''''''''',
      Ty MemOut_CTf'''''''''''') : (memMergeIn_CTf''''''''''''_dbuf,MemIn_CTf'''''''''''') > (memOut_CTf'''''''''''',MemOut_CTf'''''''''''') */
  logic [114:0] \memMergeIn_CTf''''''''''''_dbuf_mem [65535:0];
  logic [15:0] \memMergeIn_CTf''''''''''''_dbuf_address ;
  logic [114:0] \memMergeIn_CTf''''''''''''_dbuf_din ;
  logic [114:0] \memOut_CTf''''''''''''_q ;
  logic \memOut_CTf''''''''''''_valid ;
  logic \memMergeIn_CTf''''''''''''_dbuf_we ;
  logic \memOut_CTf''''''''''''_we ;
  assign \memMergeIn_CTf''''''''''''_dbuf_din  = \memMergeIn_CTf''''''''''''_dbuf_d [132:18];
  assign \memMergeIn_CTf''''''''''''_dbuf_address  = \memMergeIn_CTf''''''''''''_dbuf_d [17:2];
  assign \memMergeIn_CTf''''''''''''_dbuf_we  = (\memMergeIn_CTf''''''''''''_dbuf_d [1:1] && \memMergeIn_CTf''''''''''''_dbuf_d [0]);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        \memOut_CTf''''''''''''_we  <= 1'd0;
        \memOut_CTf''''''''''''_valid  <= 1'd0;
      end
    else
      begin
        \memOut_CTf''''''''''''_we  <= \memMergeIn_CTf''''''''''''_dbuf_we ;
        \memOut_CTf''''''''''''_valid  <= \memMergeIn_CTf''''''''''''_dbuf_d [0];
        if (\memMergeIn_CTf''''''''''''_dbuf_we )
          begin
            \memMergeIn_CTf''''''''''''_dbuf_mem [\memMergeIn_CTf''''''''''''_dbuf_address ] <= \memMergeIn_CTf''''''''''''_dbuf_din ;
            \memOut_CTf''''''''''''_q  <= \memMergeIn_CTf''''''''''''_dbuf_din ;
          end
        else
          \memOut_CTf''''''''''''_q  <= \memMergeIn_CTf''''''''''''_dbuf_mem [\memMergeIn_CTf''''''''''''_dbuf_address ];
      end
  assign \memOut_CTf''''''''''''_d  = {\memOut_CTf''''''''''''_q ,
                                       \memOut_CTf''''''''''''_we ,
                                       \memOut_CTf''''''''''''_valid };
  assign \memMergeIn_CTf''''''''''''_dbuf_r  = ((! \memOut_CTf''''''''''''_valid ) || \memOut_CTf''''''''''''_r );
  logic [31:0] \profiling_MemIn_CTf''''''''''''_read ;
  logic [31:0] \profiling_MemIn_CTf''''''''''''_write ;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        \profiling_MemIn_CTf''''''''''''_write  <= 0;
        \profiling_MemIn_CTf''''''''''''_read  <= 0;
      end
    else
      if ((\memMergeIn_CTf''''''''''''_dbuf_we  == 1'd1))
        \profiling_MemIn_CTf''''''''''''_write  <= (\profiling_MemIn_CTf''''''''''''_write  + 1);
      else
        if ((\memOut_CTf''''''''''''_valid  == 1'd1))
          \profiling_MemIn_CTf''''''''''''_read  <= (\profiling_MemIn_CTf''''''''''''_read  + 1);
  
  /* demux (Ty C2,
       Ty MemOut_CTf'''''''''''') : (memMergeChoice_CTf'''''''''''',C2) (memOut_CTf''''''''''''_dbuf,MemOut_CTf'''''''''''') > [(memReadOut_CTf'''''''''''',MemOut_CTf''''''''''''),
                                                                                                                                (memWriteOut_CTf'''''''''''',MemOut_CTf'''''''''''')] */
  logic [1:0] \memOut_CTf''''''''''''_dbuf_onehotd ;
  always_comb
    if ((\memMergeChoice_CTf''''''''''''_d [0] && \memOut_CTf''''''''''''_dbuf_d [0]))
      unique case (\memMergeChoice_CTf''''''''''''_d [1:1])
        1'd0: \memOut_CTf''''''''''''_dbuf_onehotd  = 2'd1;
        1'd1: \memOut_CTf''''''''''''_dbuf_onehotd  = 2'd2;
        default: \memOut_CTf''''''''''''_dbuf_onehotd  = 2'd0;
      endcase
    else \memOut_CTf''''''''''''_dbuf_onehotd  = 2'd0;
  assign \memReadOut_CTf''''''''''''_d  = {\memOut_CTf''''''''''''_dbuf_d [116:1],
                                           \memOut_CTf''''''''''''_dbuf_onehotd [0]};
  assign \memWriteOut_CTf''''''''''''_d  = {\memOut_CTf''''''''''''_dbuf_d [116:1],
                                            \memOut_CTf''''''''''''_dbuf_onehotd [1]};
  assign \memOut_CTf''''''''''''_dbuf_r  = (| (\memOut_CTf''''''''''''_dbuf_onehotd  & {\memWriteOut_CTf''''''''''''_r ,
                                                                                        \memReadOut_CTf''''''''''''_r }));
  assign \memMergeChoice_CTf''''''''''''_r  = \memOut_CTf''''''''''''_dbuf_r ;
  
  /* dbuf (Ty MemIn_CTf'''''''''''') : (memMergeIn_CTf''''''''''''_rbuf,MemIn_CTf'''''''''''') > (memMergeIn_CTf''''''''''''_dbuf,MemIn_CTf'''''''''''') */
  assign \memMergeIn_CTf''''''''''''_rbuf_r  = ((! \memMergeIn_CTf''''''''''''_dbuf_d [0]) || \memMergeIn_CTf''''''''''''_dbuf_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \memMergeIn_CTf''''''''''''_dbuf_d  <= {132'd0, 1'd0};
    else
      if (\memMergeIn_CTf''''''''''''_rbuf_r )
        \memMergeIn_CTf''''''''''''_dbuf_d  <= \memMergeIn_CTf''''''''''''_rbuf_d ;
  
  /* rbuf (Ty MemIn_CTf'''''''''''') : (memMergeIn_CTf'''''''''''',MemIn_CTf'''''''''''') > (memMergeIn_CTf''''''''''''_rbuf,MemIn_CTf'''''''''''') */
  \MemIn_CTf''''''''''''_t  \memMergeIn_CTf''''''''''''_buf ;
  assign \memMergeIn_CTf''''''''''''_r  = (! \memMergeIn_CTf''''''''''''_buf [0]);
  assign \memMergeIn_CTf''''''''''''_rbuf_d  = (\memMergeIn_CTf''''''''''''_buf [0] ? \memMergeIn_CTf''''''''''''_buf  :
                                                \memMergeIn_CTf''''''''''''_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \memMergeIn_CTf''''''''''''_buf  <= {132'd0, 1'd0};
    else
      if ((\memMergeIn_CTf''''''''''''_rbuf_r  && \memMergeIn_CTf''''''''''''_buf [0]))
        \memMergeIn_CTf''''''''''''_buf  <= {132'd0, 1'd0};
      else if (((! \memMergeIn_CTf''''''''''''_rbuf_r ) && (! \memMergeIn_CTf''''''''''''_buf [0])))
        \memMergeIn_CTf''''''''''''_buf  <= \memMergeIn_CTf''''''''''''_d ;
  
  /* dbuf (Ty MemOut_CTf'''''''''''') : (memOut_CTf''''''''''''_rbuf,MemOut_CTf'''''''''''') > (memOut_CTf''''''''''''_dbuf,MemOut_CTf'''''''''''') */
  assign \memOut_CTf''''''''''''_rbuf_r  = ((! \memOut_CTf''''''''''''_dbuf_d [0]) || \memOut_CTf''''''''''''_dbuf_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \memOut_CTf''''''''''''_dbuf_d  <= {116'd0, 1'd0};
    else
      if (\memOut_CTf''''''''''''_rbuf_r )
        \memOut_CTf''''''''''''_dbuf_d  <= \memOut_CTf''''''''''''_rbuf_d ;
  
  /* rbuf (Ty MemOut_CTf'''''''''''') : (memOut_CTf'''''''''''',MemOut_CTf'''''''''''') > (memOut_CTf''''''''''''_rbuf,MemOut_CTf'''''''''''') */
  \MemOut_CTf''''''''''''_t  \memOut_CTf''''''''''''_buf ;
  assign \memOut_CTf''''''''''''_r  = (! \memOut_CTf''''''''''''_buf [0]);
  assign \memOut_CTf''''''''''''_rbuf_d  = (\memOut_CTf''''''''''''_buf [0] ? \memOut_CTf''''''''''''_buf  :
                                            \memOut_CTf''''''''''''_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \memOut_CTf''''''''''''_buf  <= {116'd0, 1'd0};
    else
      if ((\memOut_CTf''''''''''''_rbuf_r  && \memOut_CTf''''''''''''_buf [0]))
        \memOut_CTf''''''''''''_buf  <= {116'd0, 1'd0};
      else if (((! \memOut_CTf''''''''''''_rbuf_r ) && (! \memOut_CTf''''''''''''_buf [0])))
        \memOut_CTf''''''''''''_buf  <= \memOut_CTf''''''''''''_d ;
  
  /* destruct (Ty Pointer_CTf'''''''''''',
          Dcon Pointer_CTf'''''''''''') : (scfarg_0_1_1_argbuf,Pointer_CTf'''''''''''') > [(destructReadIn_CTf'''''''''''',Word16#)] */
  assign \destructReadIn_CTf''''''''''''_d  = {scfarg_0_1_1_argbuf_d[16:1],
                                               scfarg_0_1_1_argbuf_d[0]};
  assign scfarg_0_1_1_argbuf_r = \destructReadIn_CTf''''''''''''_r ;
  
  /* dcon (Ty MemIn_CTf'''''''''''',
      Dcon ReadIn_CTf'''''''''''') : [(destructReadIn_CTf'''''''''''',Word16#)] > (dconReadIn_CTf'''''''''''',MemIn_CTf'''''''''''') */
  assign \dconReadIn_CTf''''''''''''_d  = \ReadIn_CTf''''''''''''_dc ((& {\destructReadIn_CTf''''''''''''_d [0]}), \destructReadIn_CTf''''''''''''_d );
  assign {\destructReadIn_CTf''''''''''''_r } = {1 {(\dconReadIn_CTf''''''''''''_r  && \dconReadIn_CTf''''''''''''_d [0])}};
  
  /* destruct (Ty MemOut_CTf'''''''''''',
          Dcon ReadOut_CTf'''''''''''') : (memReadOut_CTf'''''''''''',MemOut_CTf'''''''''''') > [(readPointer_CTf''''''''''''scfarg_0_1_1_argbuf,CTf'''''''''''')] */
  assign \readPointer_CTf''''''''''''scfarg_0_1_1_argbuf_d  = {\memReadOut_CTf''''''''''''_d [116:2],
                                                               \memReadOut_CTf''''''''''''_d [0]};
  assign \memReadOut_CTf''''''''''''_r  = \readPointer_CTf''''''''''''scfarg_0_1_1_argbuf_r ;
  
  /* mergectrl (Ty C5,
           Ty CTf'''''''''''') : [(lizzieLet54_1_argbuf,CTf''''''''''''),
                                  (lizzieLet58_1_argbuf,CTf''''''''''''),
                                  (lizzieLet66_1_argbuf,CTf''''''''''''),
                                  (lizzieLet67_1_argbuf,CTf''''''''''''),
                                  (lizzieLet68_1_argbuf,CTf'''''''''''')] > (writeMerge_choice_CTf'''''''''''',C5) (writeMerge_data_CTf'''''''''''',CTf'''''''''''') */
  logic [4:0] lizzieLet54_1_argbuf_select_d;
  assign lizzieLet54_1_argbuf_select_d = ((| lizzieLet54_1_argbuf_select_q) ? lizzieLet54_1_argbuf_select_q :
                                          (lizzieLet54_1_argbuf_d[0] ? 5'd1 :
                                           (lizzieLet58_1_argbuf_d[0] ? 5'd2 :
                                            (lizzieLet66_1_argbuf_d[0] ? 5'd4 :
                                             (lizzieLet67_1_argbuf_d[0] ? 5'd8 :
                                              (lizzieLet68_1_argbuf_d[0] ? 5'd16 :
                                               5'd0))))));
  logic [4:0] lizzieLet54_1_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet54_1_argbuf_select_q <= 5'd0;
    else
      lizzieLet54_1_argbuf_select_q <= (lizzieLet54_1_argbuf_done ? 5'd0 :
                                        lizzieLet54_1_argbuf_select_d);
  logic [1:0] lizzieLet54_1_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet54_1_argbuf_emit_q <= 2'd0;
    else
      lizzieLet54_1_argbuf_emit_q <= (lizzieLet54_1_argbuf_done ? 2'd0 :
                                      lizzieLet54_1_argbuf_emit_d);
  logic [1:0] lizzieLet54_1_argbuf_emit_d;
  assign lizzieLet54_1_argbuf_emit_d = (lizzieLet54_1_argbuf_emit_q | ({\writeMerge_choice_CTf''''''''''''_d [0],
                                                                        \writeMerge_data_CTf''''''''''''_d [0]} & {\writeMerge_choice_CTf''''''''''''_r ,
                                                                                                                   \writeMerge_data_CTf''''''''''''_r }));
  logic lizzieLet54_1_argbuf_done;
  assign lizzieLet54_1_argbuf_done = (& lizzieLet54_1_argbuf_emit_d);
  assign {lizzieLet68_1_argbuf_r,
          lizzieLet67_1_argbuf_r,
          lizzieLet66_1_argbuf_r,
          lizzieLet58_1_argbuf_r,
          lizzieLet54_1_argbuf_r} = (lizzieLet54_1_argbuf_done ? lizzieLet54_1_argbuf_select_d :
                                     5'd0);
  assign \writeMerge_data_CTf''''''''''''_d  = ((lizzieLet54_1_argbuf_select_d[0] && (! lizzieLet54_1_argbuf_emit_q[0])) ? lizzieLet54_1_argbuf_d :
                                                ((lizzieLet54_1_argbuf_select_d[1] && (! lizzieLet54_1_argbuf_emit_q[0])) ? lizzieLet58_1_argbuf_d :
                                                 ((lizzieLet54_1_argbuf_select_d[2] && (! lizzieLet54_1_argbuf_emit_q[0])) ? lizzieLet66_1_argbuf_d :
                                                  ((lizzieLet54_1_argbuf_select_d[3] && (! lizzieLet54_1_argbuf_emit_q[0])) ? lizzieLet67_1_argbuf_d :
                                                   ((lizzieLet54_1_argbuf_select_d[4] && (! lizzieLet54_1_argbuf_emit_q[0])) ? lizzieLet68_1_argbuf_d :
                                                    {115'd0, 1'd0})))));
  assign \writeMerge_choice_CTf''''''''''''_d  = ((lizzieLet54_1_argbuf_select_d[0] && (! lizzieLet54_1_argbuf_emit_q[1])) ? C1_5_dc(1'd1) :
                                                  ((lizzieLet54_1_argbuf_select_d[1] && (! lizzieLet54_1_argbuf_emit_q[1])) ? C2_5_dc(1'd1) :
                                                   ((lizzieLet54_1_argbuf_select_d[2] && (! lizzieLet54_1_argbuf_emit_q[1])) ? C3_5_dc(1'd1) :
                                                    ((lizzieLet54_1_argbuf_select_d[3] && (! lizzieLet54_1_argbuf_emit_q[1])) ? C4_5_dc(1'd1) :
                                                     ((lizzieLet54_1_argbuf_select_d[4] && (! lizzieLet54_1_argbuf_emit_q[1])) ? C5_5_dc(1'd1) :
                                                      {3'd0, 1'd0})))));
  
  /* demux (Ty C5,
       Ty Pointer_CTf'''''''''''') : (writeMerge_choice_CTf'''''''''''',C5) (demuxWriteResult_CTf'''''''''''',Pointer_CTf'''''''''''') > [(writeCTf''''''''''''lizzieLet54_1_argbuf,Pointer_CTf''''''''''''),
                                                                                                                                          (writeCTf''''''''''''lizzieLet58_1_argbuf,Pointer_CTf''''''''''''),
                                                                                                                                          (writeCTf''''''''''''lizzieLet66_1_argbuf,Pointer_CTf''''''''''''),
                                                                                                                                          (writeCTf''''''''''''lizzieLet67_1_argbuf,Pointer_CTf''''''''''''),
                                                                                                                                          (writeCTf''''''''''''lizzieLet68_1_argbuf,Pointer_CTf'''''''''''')] */
  logic [4:0] \demuxWriteResult_CTf''''''''''''_onehotd ;
  always_comb
    if ((\writeMerge_choice_CTf''''''''''''_d [0] && \demuxWriteResult_CTf''''''''''''_d [0]))
      unique case (\writeMerge_choice_CTf''''''''''''_d [3:1])
        3'd0: \demuxWriteResult_CTf''''''''''''_onehotd  = 5'd1;
        3'd1: \demuxWriteResult_CTf''''''''''''_onehotd  = 5'd2;
        3'd2: \demuxWriteResult_CTf''''''''''''_onehotd  = 5'd4;
        3'd3: \demuxWriteResult_CTf''''''''''''_onehotd  = 5'd8;
        3'd4: \demuxWriteResult_CTf''''''''''''_onehotd  = 5'd16;
        default: \demuxWriteResult_CTf''''''''''''_onehotd  = 5'd0;
      endcase
    else \demuxWriteResult_CTf''''''''''''_onehotd  = 5'd0;
  assign \writeCTf''''''''''''lizzieLet54_1_argbuf_d  = {\demuxWriteResult_CTf''''''''''''_d [16:1],
                                                         \demuxWriteResult_CTf''''''''''''_onehotd [0]};
  assign \writeCTf''''''''''''lizzieLet58_1_argbuf_d  = {\demuxWriteResult_CTf''''''''''''_d [16:1],
                                                         \demuxWriteResult_CTf''''''''''''_onehotd [1]};
  assign \writeCTf''''''''''''lizzieLet66_1_argbuf_d  = {\demuxWriteResult_CTf''''''''''''_d [16:1],
                                                         \demuxWriteResult_CTf''''''''''''_onehotd [2]};
  assign \writeCTf''''''''''''lizzieLet67_1_argbuf_d  = {\demuxWriteResult_CTf''''''''''''_d [16:1],
                                                         \demuxWriteResult_CTf''''''''''''_onehotd [3]};
  assign \writeCTf''''''''''''lizzieLet68_1_argbuf_d  = {\demuxWriteResult_CTf''''''''''''_d [16:1],
                                                         \demuxWriteResult_CTf''''''''''''_onehotd [4]};
  assign \demuxWriteResult_CTf''''''''''''_r  = (| (\demuxWriteResult_CTf''''''''''''_onehotd  & {\writeCTf''''''''''''lizzieLet68_1_argbuf_r ,
                                                                                                  \writeCTf''''''''''''lizzieLet67_1_argbuf_r ,
                                                                                                  \writeCTf''''''''''''lizzieLet66_1_argbuf_r ,
                                                                                                  \writeCTf''''''''''''lizzieLet58_1_argbuf_r ,
                                                                                                  \writeCTf''''''''''''lizzieLet54_1_argbuf_r }));
  assign \writeMerge_choice_CTf''''''''''''_r  = \demuxWriteResult_CTf''''''''''''_r ;
  
  /* dcon (Ty MemIn_CTf'''''''''''',
      Dcon WriteIn_CTf'''''''''''') : [(forkHP1_CTf'''''''''''2,Word16#),
                                       (writeMerge_data_CTf'''''''''''',CTf'''''''''''')] > (dconWriteIn_CTf'''''''''''',MemIn_CTf'''''''''''') */
  assign \dconWriteIn_CTf''''''''''''_d  = \WriteIn_CTf''''''''''''_dc ((& {\forkHP1_CTf'''''''''''2_d [0],
                                                                            \writeMerge_data_CTf''''''''''''_d [0]}), \forkHP1_CTf'''''''''''2_d , \writeMerge_data_CTf''''''''''''_d );
  assign {\forkHP1_CTf'''''''''''2_r ,
          \writeMerge_data_CTf''''''''''''_r } = {2 {(\dconWriteIn_CTf''''''''''''_r  && \dconWriteIn_CTf''''''''''''_d [0])}};
  
  /* dcon (Ty Pointer_CTf'''''''''''',
      Dcon Pointer_CTf'''''''''''') : [(forkHP1_CTf'''''''''''3,Word16#)] > (dconPtr_CTf'''''''''''',Pointer_CTf'''''''''''') */
  assign \dconPtr_CTf''''''''''''_d  = \Pointer_CTf''''''''''''_dc ((& {\forkHP1_CTf'''''''''''3_d [0]}), \forkHP1_CTf'''''''''''3_d );
  assign {\forkHP1_CTf'''''''''''3_r } = {1 {(\dconPtr_CTf''''''''''''_r  && \dconPtr_CTf''''''''''''_d [0])}};
  
  /* demux (Ty MemOut_CTf'''''''''''',
       Ty Pointer_CTf'''''''''''') : (memWriteOut_CTf'''''''''''',MemOut_CTf'''''''''''') (dconPtr_CTf'''''''''''',Pointer_CTf'''''''''''') > [(_169,Pointer_CTf''''''''''''),
                                                                                                                                               (demuxWriteResult_CTf'''''''''''',Pointer_CTf'''''''''''')] */
  logic [1:0] \dconPtr_CTf''''''''''''_onehotd ;
  always_comb
    if ((\memWriteOut_CTf''''''''''''_d [0] && \dconPtr_CTf''''''''''''_d [0]))
      unique case (\memWriteOut_CTf''''''''''''_d [1:1])
        1'd0: \dconPtr_CTf''''''''''''_onehotd  = 2'd1;
        1'd1: \dconPtr_CTf''''''''''''_onehotd  = 2'd2;
        default: \dconPtr_CTf''''''''''''_onehotd  = 2'd0;
      endcase
    else \dconPtr_CTf''''''''''''_onehotd  = 2'd0;
  assign _169_d = {\dconPtr_CTf''''''''''''_d [16:1],
                   \dconPtr_CTf''''''''''''_onehotd [0]};
  assign \demuxWriteResult_CTf''''''''''''_d  = {\dconPtr_CTf''''''''''''_d [16:1],
                                                 \dconPtr_CTf''''''''''''_onehotd [1]};
  assign \dconPtr_CTf''''''''''''_r  = (| (\dconPtr_CTf''''''''''''_onehotd  & {\demuxWriteResult_CTf''''''''''''_r ,
                                                                                _169_r}));
  assign \memWriteOut_CTf''''''''''''_r  = \dconPtr_CTf''''''''''''_r ;
  
  /* buf (Ty Go) : (goFork,Go) > (go_1_argbuf,Go) */
  Go_t goFork_bufchan_d;
  logic goFork_bufchan_r;
  assign goFork_r = ((! goFork_bufchan_d[0]) || goFork_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) goFork_bufchan_d <= 1'd0;
    else if (goFork_r) goFork_bufchan_d <= goFork_d;
  Go_t goFork_bufchan_buf;
  assign goFork_bufchan_r = (! goFork_bufchan_buf[0]);
  assign go_1_argbuf_d = (goFork_bufchan_buf[0] ? goFork_bufchan_buf :
                          goFork_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) goFork_bufchan_buf <= 1'd0;
    else
      if ((go_1_argbuf_r && goFork_bufchan_buf[0]))
        goFork_bufchan_buf <= 1'd0;
      else if (((! go_1_argbuf_r) && (! goFork_bufchan_buf[0])))
        goFork_bufchan_buf <= goFork_bufchan_d;
  
  /* source (Ty Go) : > (sourceGo,Go) */
  
  /* source (Ty Pointer_QTree_Bool) : > (m1a81_0,Pointer_QTree_Bool) */
  
  /* source (Ty Pointer_QTree_Bool) : > (m2a82_1,Pointer_QTree_Bool) */
  
  /* source (Ty Pointer_QTree_Bool) : > (m3a83_2,Pointer_QTree_Bool) */
  
  /* destruct (Ty TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf'''''''''''',
          Dcon TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf'''''''''''') : (call_f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf''''''''''''_1,TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf'''''''''''') > [(call_f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf''''''''''''go_3,Go),
                                                                                                                                                                                                                                                                         (call_f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf''''''''''''q4a90,Pointer_QTree_Bool),
                                                                                                                                                                                                                                                                         (call_f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf''''''''''''t4a91,Pointer_QTree_Bool),
                                                                                                                                                                                                                                                                         (call_f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf''''''''''''sc_0_1,Pointer_CTf'''''''''''')] */
  logic [3:0] \call_f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf''''''''''''_1_emitted ;
  logic [3:0] \call_f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf''''''''''''_1_done ;
  assign \call_f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf''''''''''''go_3_d  = (\call_f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf''''''''''''_1_d [0] && (! \call_f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf''''''''''''_1_emitted [0]));
  assign \call_f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf''''''''''''q4a90_d  = {\call_f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf''''''''''''_1_d [16:1],
                                                                                                                 (\call_f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf''''''''''''_1_d [0] && (! \call_f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf''''''''''''_1_emitted [1]))};
  assign \call_f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf''''''''''''t4a91_d  = {\call_f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf''''''''''''_1_d [32:17],
                                                                                                                 (\call_f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf''''''''''''_1_d [0] && (! \call_f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf''''''''''''_1_emitted [2]))};
  assign \call_f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf''''''''''''sc_0_1_d  = {\call_f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf''''''''''''_1_d [48:33],
                                                                                                                  (\call_f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf''''''''''''_1_d [0] && (! \call_f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf''''''''''''_1_emitted [3]))};
  assign \call_f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf''''''''''''_1_done  = (\call_f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf''''''''''''_1_emitted  | ({\call_f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf''''''''''''sc_0_1_d [0],
                                                                                                                                                                                                                             \call_f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf''''''''''''t4a91_d [0],
                                                                                                                                                                                                                             \call_f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf''''''''''''q4a90_d [0],
                                                                                                                                                                                                                             \call_f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf''''''''''''go_3_d [0]} & {\call_f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf''''''''''''sc_0_1_r ,
                                                                                                                                                                                                                                                                                                                                        \call_f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf''''''''''''t4a91_r ,
                                                                                                                                                                                                                                                                                                                                        \call_f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf''''''''''''q4a90_r ,
                                                                                                                                                                                                                                                                                                                                        \call_f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf''''''''''''go_3_r }));
  assign \call_f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf''''''''''''_1_r  = (& \call_f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf''''''''''''_1_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \call_f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf''''''''''''_1_emitted  <= 4'd0;
    else
      \call_f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf''''''''''''_1_emitted  <= (\call_f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf''''''''''''_1_r  ? 4'd0 :
                                                                                                                  \call_f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf''''''''''''_1_done );
  
  /* rbuf (Ty Go) : (call_f''''''''''''_goConst,Go) > (call_f''''''''''''_initBufi,Go) */
  Go_t \call_f''''''''''''_goConst_buf ;
  assign \call_f''''''''''''_goConst_r  = (! \call_f''''''''''''_goConst_buf [0]);
  assign \call_f''''''''''''_initBufi_d  = (\call_f''''''''''''_goConst_buf [0] ? \call_f''''''''''''_goConst_buf  :
                                            \call_f''''''''''''_goConst_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \call_f''''''''''''_goConst_buf  <= 1'd0;
    else
      if ((\call_f''''''''''''_initBufi_r  && \call_f''''''''''''_goConst_buf [0]))
        \call_f''''''''''''_goConst_buf  <= 1'd0;
      else if (((! \call_f''''''''''''_initBufi_r ) && (! \call_f''''''''''''_goConst_buf [0])))
        \call_f''''''''''''_goConst_buf  <= \call_f''''''''''''_goConst_d ;
  
  /* mergectrl (Ty C5,Ty Go) : [(call_f''''''''''''_goMux1,Go),
                           (lizzieLet65_3Lcall_f''''''''''''3_1_argbuf,Go),
                           (lizzieLet65_3Lcall_f''''''''''''2_1_argbuf,Go),
                           (lizzieLet65_3Lcall_f''''''''''''1_1_argbuf,Go),
                           (lizzieLet45_4QNode_Bool_3QNode_Bool_1_argbuf,Go)] > (go_3_goMux_choice,C5) (go_3_goMux_data,Go) */
  logic [4:0] \call_f''''''''''''_goMux1_select_d ;
  assign \call_f''''''''''''_goMux1_select_d  = ((| \call_f''''''''''''_goMux1_select_q ) ? \call_f''''''''''''_goMux1_select_q  :
                                                 (\call_f''''''''''''_goMux1_d [0] ? 5'd1 :
                                                  (\lizzieLet65_3Lcall_f''''''''''''3_1_argbuf_d [0] ? 5'd2 :
                                                   (\lizzieLet65_3Lcall_f''''''''''''2_1_argbuf_d [0] ? 5'd4 :
                                                    (\lizzieLet65_3Lcall_f''''''''''''1_1_argbuf_d [0] ? 5'd8 :
                                                     (lizzieLet45_4QNode_Bool_3QNode_Bool_1_argbuf_d[0] ? 5'd16 :
                                                      5'd0))))));
  logic [4:0] \call_f''''''''''''_goMux1_select_q ;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \call_f''''''''''''_goMux1_select_q  <= 5'd0;
    else
      \call_f''''''''''''_goMux1_select_q  <= (\call_f''''''''''''_goMux1_done  ? 5'd0 :
                                               \call_f''''''''''''_goMux1_select_d );
  logic [1:0] \call_f''''''''''''_goMux1_emit_q ;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \call_f''''''''''''_goMux1_emit_q  <= 2'd0;
    else
      \call_f''''''''''''_goMux1_emit_q  <= (\call_f''''''''''''_goMux1_done  ? 2'd0 :
                                             \call_f''''''''''''_goMux1_emit_d );
  logic [1:0] \call_f''''''''''''_goMux1_emit_d ;
  assign \call_f''''''''''''_goMux1_emit_d  = (\call_f''''''''''''_goMux1_emit_q  | ({go_3_goMux_choice_d[0],
                                                                                      go_3_goMux_data_d[0]} & {go_3_goMux_choice_r,
                                                                                                               go_3_goMux_data_r}));
  logic \call_f''''''''''''_goMux1_done ;
  assign \call_f''''''''''''_goMux1_done  = (& \call_f''''''''''''_goMux1_emit_d );
  assign {lizzieLet45_4QNode_Bool_3QNode_Bool_1_argbuf_r,
          \lizzieLet65_3Lcall_f''''''''''''1_1_argbuf_r ,
          \lizzieLet65_3Lcall_f''''''''''''2_1_argbuf_r ,
          \lizzieLet65_3Lcall_f''''''''''''3_1_argbuf_r ,
          \call_f''''''''''''_goMux1_r } = (\call_f''''''''''''_goMux1_done  ? \call_f''''''''''''_goMux1_select_d  :
                                            5'd0);
  assign go_3_goMux_data_d = ((\call_f''''''''''''_goMux1_select_d [0] && (! \call_f''''''''''''_goMux1_emit_q [0])) ? \call_f''''''''''''_goMux1_d  :
                              ((\call_f''''''''''''_goMux1_select_d [1] && (! \call_f''''''''''''_goMux1_emit_q [0])) ? \lizzieLet65_3Lcall_f''''''''''''3_1_argbuf_d  :
                               ((\call_f''''''''''''_goMux1_select_d [2] && (! \call_f''''''''''''_goMux1_emit_q [0])) ? \lizzieLet65_3Lcall_f''''''''''''2_1_argbuf_d  :
                                ((\call_f''''''''''''_goMux1_select_d [3] && (! \call_f''''''''''''_goMux1_emit_q [0])) ? \lizzieLet65_3Lcall_f''''''''''''1_1_argbuf_d  :
                                 ((\call_f''''''''''''_goMux1_select_d [4] && (! \call_f''''''''''''_goMux1_emit_q [0])) ? lizzieLet45_4QNode_Bool_3QNode_Bool_1_argbuf_d :
                                  1'd0)))));
  assign go_3_goMux_choice_d = ((\call_f''''''''''''_goMux1_select_d [0] && (! \call_f''''''''''''_goMux1_emit_q [1])) ? C1_5_dc(1'd1) :
                                ((\call_f''''''''''''_goMux1_select_d [1] && (! \call_f''''''''''''_goMux1_emit_q [1])) ? C2_5_dc(1'd1) :
                                 ((\call_f''''''''''''_goMux1_select_d [2] && (! \call_f''''''''''''_goMux1_emit_q [1])) ? C3_5_dc(1'd1) :
                                  ((\call_f''''''''''''_goMux1_select_d [3] && (! \call_f''''''''''''_goMux1_emit_q [1])) ? C4_5_dc(1'd1) :
                                   ((\call_f''''''''''''_goMux1_select_d [4] && (! \call_f''''''''''''_goMux1_emit_q [1])) ? C5_5_dc(1'd1) :
                                    {3'd0, 1'd0})))));
  
  /* fork (Ty Go) : (call_f''''''''''''_initBuf,Go) > [(call_f''''''''''''_unlockFork1,Go),
                                                  (call_f''''''''''''_unlockFork2,Go),
                                                  (call_f''''''''''''_unlockFork3,Go),
                                                  (call_f''''''''''''_unlockFork4,Go)] */
  logic [3:0] \call_f''''''''''''_initBuf_emitted ;
  logic [3:0] \call_f''''''''''''_initBuf_done ;
  assign \call_f''''''''''''_unlockFork1_d  = (\call_f''''''''''''_initBuf_d [0] && (! \call_f''''''''''''_initBuf_emitted [0]));
  assign \call_f''''''''''''_unlockFork2_d  = (\call_f''''''''''''_initBuf_d [0] && (! \call_f''''''''''''_initBuf_emitted [1]));
  assign \call_f''''''''''''_unlockFork3_d  = (\call_f''''''''''''_initBuf_d [0] && (! \call_f''''''''''''_initBuf_emitted [2]));
  assign \call_f''''''''''''_unlockFork4_d  = (\call_f''''''''''''_initBuf_d [0] && (! \call_f''''''''''''_initBuf_emitted [3]));
  assign \call_f''''''''''''_initBuf_done  = (\call_f''''''''''''_initBuf_emitted  | ({\call_f''''''''''''_unlockFork4_d [0],
                                                                                       \call_f''''''''''''_unlockFork3_d [0],
                                                                                       \call_f''''''''''''_unlockFork2_d [0],
                                                                                       \call_f''''''''''''_unlockFork1_d [0]} & {\call_f''''''''''''_unlockFork4_r ,
                                                                                                                                 \call_f''''''''''''_unlockFork3_r ,
                                                                                                                                 \call_f''''''''''''_unlockFork2_r ,
                                                                                                                                 \call_f''''''''''''_unlockFork1_r }));
  assign \call_f''''''''''''_initBuf_r  = (& \call_f''''''''''''_initBuf_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \call_f''''''''''''_initBuf_emitted  <= 4'd0;
    else
      \call_f''''''''''''_initBuf_emitted  <= (\call_f''''''''''''_initBuf_r  ? 4'd0 :
                                               \call_f''''''''''''_initBuf_done );
  
  /* initbuf (Ty Go,
         Dcon Go) : (call_f''''''''''''_initBufi,Go) > (call_f''''''''''''_initBuf,Go) */
  assign \call_f''''''''''''_initBufi_r  = ((! \call_f''''''''''''_initBuf_d [0]) || \call_f''''''''''''_initBuf_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \call_f''''''''''''_initBuf_d  <= Go_dc(1'd1);
    else
      if (\call_f''''''''''''_initBufi_r )
        \call_f''''''''''''_initBuf_d  <= \call_f''''''''''''_initBufi_d ;
  
  /* mux (Ty Go,
     Ty Go) : (call_f''''''''''''_unlockFork1,Go) [(call_f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf''''''''''''go_3,Go)] > (call_f''''''''''''_goMux1,Go) */
  assign \call_f''''''''''''_goMux1_d  = (\call_f''''''''''''_unlockFork1_d [0] && \call_f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf''''''''''''go_3_d [0]);
  assign \call_f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf''''''''''''go_3_r  = (\call_f''''''''''''_goMux1_r  && (\call_f''''''''''''_unlockFork1_d [0] && \call_f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf''''''''''''go_3_d [0]));
  assign \call_f''''''''''''_unlockFork1_r  = (\call_f''''''''''''_goMux1_r  && (\call_f''''''''''''_unlockFork1_d [0] && \call_f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf''''''''''''go_3_d [0]));
  
  /* mux (Ty Go,
     Ty Pointer_QTree_Bool) : (call_f''''''''''''_unlockFork2,Go) [(call_f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf''''''''''''q4a90,Pointer_QTree_Bool)] > (call_f''''''''''''_goMux2,Pointer_QTree_Bool) */
  assign \call_f''''''''''''_goMux2_d  = {\call_f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf''''''''''''q4a90_d [16:1],
                                          (\call_f''''''''''''_unlockFork2_d [0] && \call_f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf''''''''''''q4a90_d [0])};
  assign \call_f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf''''''''''''q4a90_r  = (\call_f''''''''''''_goMux2_r  && (\call_f''''''''''''_unlockFork2_d [0] && \call_f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf''''''''''''q4a90_d [0]));
  assign \call_f''''''''''''_unlockFork2_r  = (\call_f''''''''''''_goMux2_r  && (\call_f''''''''''''_unlockFork2_d [0] && \call_f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf''''''''''''q4a90_d [0]));
  
  /* mux (Ty Go,
     Ty Pointer_QTree_Bool) : (call_f''''''''''''_unlockFork3,Go) [(call_f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf''''''''''''t4a91,Pointer_QTree_Bool)] > (call_f''''''''''''_goMux3,Pointer_QTree_Bool) */
  assign \call_f''''''''''''_goMux3_d  = {\call_f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf''''''''''''t4a91_d [16:1],
                                          (\call_f''''''''''''_unlockFork3_d [0] && \call_f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf''''''''''''t4a91_d [0])};
  assign \call_f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf''''''''''''t4a91_r  = (\call_f''''''''''''_goMux3_r  && (\call_f''''''''''''_unlockFork3_d [0] && \call_f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf''''''''''''t4a91_d [0]));
  assign \call_f''''''''''''_unlockFork3_r  = (\call_f''''''''''''_goMux3_r  && (\call_f''''''''''''_unlockFork3_d [0] && \call_f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf''''''''''''t4a91_d [0]));
  
  /* mux (Ty Go,
     Ty Pointer_CTf'''''''''''') : (call_f''''''''''''_unlockFork4,Go) [(call_f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf''''''''''''sc_0_1,Pointer_CTf'''''''''''')] > (call_f''''''''''''_goMux4,Pointer_CTf'''''''''''') */
  assign \call_f''''''''''''_goMux4_d  = {\call_f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf''''''''''''sc_0_1_d [16:1],
                                          (\call_f''''''''''''_unlockFork4_d [0] && \call_f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf''''''''''''sc_0_1_d [0])};
  assign \call_f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf''''''''''''sc_0_1_r  = (\call_f''''''''''''_goMux4_r  && (\call_f''''''''''''_unlockFork4_d [0] && \call_f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf''''''''''''sc_0_1_d [0]));
  assign \call_f''''''''''''_unlockFork4_r  = (\call_f''''''''''''_goMux4_r  && (\call_f''''''''''''_unlockFork4_d [0] && \call_f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf''''''''''''sc_0_1_d [0]));
  
  /* destruct (Ty TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf,
          Dcon TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf) : (call_fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf_1,TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf) > [(call_fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfgo_2,Go),
                                                                                                                                                                                                                                                                                        (call_fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfm1a84,Pointer_QTree_Bool),
                                                                                                                                                                                                                                                                                        (call_fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfm2a85,Pointer_QTree_Bool),
                                                                                                                                                                                                                                                                                        (call_fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfm3a86,Pointer_QTree_Bool),
                                                                                                                                                                                                                                                                                        (call_fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfsc_0,Pointer_CTf)] */
  logic [4:0] call_fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf_1_emitted;
  logic [4:0] call_fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf_1_done;
  assign call_fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfgo_2_d = (call_fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf_1_d[0] && (! call_fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf_1_emitted[0]));
  assign call_fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfm1a84_d = {call_fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf_1_d[16:1],
                                                                                                            (call_fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf_1_d[0] && (! call_fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf_1_emitted[1]))};
  assign call_fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfm2a85_d = {call_fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf_1_d[32:17],
                                                                                                            (call_fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf_1_d[0] && (! call_fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf_1_emitted[2]))};
  assign call_fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfm3a86_d = {call_fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf_1_d[48:33],
                                                                                                            (call_fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf_1_d[0] && (! call_fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf_1_emitted[3]))};
  assign call_fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfsc_0_d = {call_fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf_1_d[64:49],
                                                                                                           (call_fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf_1_d[0] && (! call_fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf_1_emitted[4]))};
  assign call_fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf_1_done = (call_fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf_1_emitted | ({call_fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfsc_0_d[0],
                                                                                                                                                                                                                   call_fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfm3a86_d[0],
                                                                                                                                                                                                                   call_fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfm2a85_d[0],
                                                                                                                                                                                                                   call_fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfm1a84_d[0],
                                                                                                                                                                                                                   call_fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfgo_2_d[0]} & {call_fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfsc_0_r,
                                                                                                                                                                                                                                                                                                                         call_fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfm3a86_r,
                                                                                                                                                                                                                                                                                                                         call_fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfm2a85_r,
                                                                                                                                                                                                                                                                                                                         call_fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfm1a84_r,
                                                                                                                                                                                                                                                                                                                         call_fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfgo_2_r}));
  assign call_fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf_1_r = (& call_fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf_1_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      call_fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf_1_emitted <= 5'd0;
    else
      call_fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf_1_emitted <= (call_fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf_1_r ? 5'd0 :
                                                                                                             call_fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf_1_done);
  
  /* rbuf (Ty Go) : (call_f_goConst,Go) > (call_f_initBufi,Go) */
  Go_t call_f_goConst_buf;
  assign call_f_goConst_r = (! call_f_goConst_buf[0]);
  assign call_f_initBufi_d = (call_f_goConst_buf[0] ? call_f_goConst_buf :
                              call_f_goConst_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_f_goConst_buf <= 1'd0;
    else
      if ((call_f_initBufi_r && call_f_goConst_buf[0]))
        call_f_goConst_buf <= 1'd0;
      else if (((! call_f_initBufi_r) && (! call_f_goConst_buf[0])))
        call_f_goConst_buf <= call_f_goConst_d;
  
  /* mergectrl (Ty C5,Ty Go) : [(call_f_goMux1,Go),
                           (lizzieLet60_3Lcall_f3_1_argbuf,Go),
                           (lizzieLet60_3Lcall_f2_1_argbuf,Go),
                           (lizzieLet60_3Lcall_f1_1_argbuf,Go),
                           (lizzieLet0_4QNode_Bool_4QNode_Bool_4QNode_Bool_1_argbuf,Go)] > (go_2_goMux_choice,C5) (go_2_goMux_data,Go) */
  logic [4:0] call_f_goMux1_select_d;
  assign call_f_goMux1_select_d = ((| call_f_goMux1_select_q) ? call_f_goMux1_select_q :
                                   (call_f_goMux1_d[0] ? 5'd1 :
                                    (lizzieLet60_3Lcall_f3_1_argbuf_d[0] ? 5'd2 :
                                     (lizzieLet60_3Lcall_f2_1_argbuf_d[0] ? 5'd4 :
                                      (lizzieLet60_3Lcall_f1_1_argbuf_d[0] ? 5'd8 :
                                       (lizzieLet0_4QNode_Bool_4QNode_Bool_4QNode_Bool_1_argbuf_d[0] ? 5'd16 :
                                        5'd0))))));
  logic [4:0] call_f_goMux1_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_f_goMux1_select_q <= 5'd0;
    else
      call_f_goMux1_select_q <= (call_f_goMux1_done ? 5'd0 :
                                 call_f_goMux1_select_d);
  logic [1:0] call_f_goMux1_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_f_goMux1_emit_q <= 2'd0;
    else
      call_f_goMux1_emit_q <= (call_f_goMux1_done ? 2'd0 :
                               call_f_goMux1_emit_d);
  logic [1:0] call_f_goMux1_emit_d;
  assign call_f_goMux1_emit_d = (call_f_goMux1_emit_q | ({go_2_goMux_choice_d[0],
                                                          go_2_goMux_data_d[0]} & {go_2_goMux_choice_r,
                                                                                   go_2_goMux_data_r}));
  logic call_f_goMux1_done;
  assign call_f_goMux1_done = (& call_f_goMux1_emit_d);
  assign {lizzieLet0_4QNode_Bool_4QNode_Bool_4QNode_Bool_1_argbuf_r,
          lizzieLet60_3Lcall_f1_1_argbuf_r,
          lizzieLet60_3Lcall_f2_1_argbuf_r,
          lizzieLet60_3Lcall_f3_1_argbuf_r,
          call_f_goMux1_r} = (call_f_goMux1_done ? call_f_goMux1_select_d :
                              5'd0);
  assign go_2_goMux_data_d = ((call_f_goMux1_select_d[0] && (! call_f_goMux1_emit_q[0])) ? call_f_goMux1_d :
                              ((call_f_goMux1_select_d[1] && (! call_f_goMux1_emit_q[0])) ? lizzieLet60_3Lcall_f3_1_argbuf_d :
                               ((call_f_goMux1_select_d[2] && (! call_f_goMux1_emit_q[0])) ? lizzieLet60_3Lcall_f2_1_argbuf_d :
                                ((call_f_goMux1_select_d[3] && (! call_f_goMux1_emit_q[0])) ? lizzieLet60_3Lcall_f1_1_argbuf_d :
                                 ((call_f_goMux1_select_d[4] && (! call_f_goMux1_emit_q[0])) ? lizzieLet0_4QNode_Bool_4QNode_Bool_4QNode_Bool_1_argbuf_d :
                                  1'd0)))));
  assign go_2_goMux_choice_d = ((call_f_goMux1_select_d[0] && (! call_f_goMux1_emit_q[1])) ? C1_5_dc(1'd1) :
                                ((call_f_goMux1_select_d[1] && (! call_f_goMux1_emit_q[1])) ? C2_5_dc(1'd1) :
                                 ((call_f_goMux1_select_d[2] && (! call_f_goMux1_emit_q[1])) ? C3_5_dc(1'd1) :
                                  ((call_f_goMux1_select_d[3] && (! call_f_goMux1_emit_q[1])) ? C4_5_dc(1'd1) :
                                   ((call_f_goMux1_select_d[4] && (! call_f_goMux1_emit_q[1])) ? C5_5_dc(1'd1) :
                                    {3'd0, 1'd0})))));
  
  /* fork (Ty Go) : (call_f_initBuf,Go) > [(call_f_unlockFork1,Go),
                                      (call_f_unlockFork2,Go),
                                      (call_f_unlockFork3,Go),
                                      (call_f_unlockFork4,Go),
                                      (call_f_unlockFork5,Go)] */
  logic [4:0] call_f_initBuf_emitted;
  logic [4:0] call_f_initBuf_done;
  assign call_f_unlockFork1_d = (call_f_initBuf_d[0] && (! call_f_initBuf_emitted[0]));
  assign call_f_unlockFork2_d = (call_f_initBuf_d[0] && (! call_f_initBuf_emitted[1]));
  assign call_f_unlockFork3_d = (call_f_initBuf_d[0] && (! call_f_initBuf_emitted[2]));
  assign call_f_unlockFork4_d = (call_f_initBuf_d[0] && (! call_f_initBuf_emitted[3]));
  assign call_f_unlockFork5_d = (call_f_initBuf_d[0] && (! call_f_initBuf_emitted[4]));
  assign call_f_initBuf_done = (call_f_initBuf_emitted | ({call_f_unlockFork5_d[0],
                                                           call_f_unlockFork4_d[0],
                                                           call_f_unlockFork3_d[0],
                                                           call_f_unlockFork2_d[0],
                                                           call_f_unlockFork1_d[0]} & {call_f_unlockFork5_r,
                                                                                       call_f_unlockFork4_r,
                                                                                       call_f_unlockFork3_r,
                                                                                       call_f_unlockFork2_r,
                                                                                       call_f_unlockFork1_r}));
  assign call_f_initBuf_r = (& call_f_initBuf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_f_initBuf_emitted <= 5'd0;
    else
      call_f_initBuf_emitted <= (call_f_initBuf_r ? 5'd0 :
                                 call_f_initBuf_done);
  
  /* initbuf (Ty Go,
         Dcon Go) : (call_f_initBufi,Go) > (call_f_initBuf,Go) */
  assign call_f_initBufi_r = ((! call_f_initBuf_d[0]) || call_f_initBuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_f_initBuf_d <= Go_dc(1'd1);
    else if (call_f_initBufi_r) call_f_initBuf_d <= call_f_initBufi_d;
  
  /* mux (Ty Go,
     Ty Go) : (call_f_unlockFork1,Go) [(call_fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfgo_2,Go)] > (call_f_goMux1,Go) */
  assign call_f_goMux1_d = (call_f_unlockFork1_d[0] && call_fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfgo_2_d[0]);
  assign call_fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfgo_2_r = (call_f_goMux1_r && (call_f_unlockFork1_d[0] && call_fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfgo_2_d[0]));
  assign call_f_unlockFork1_r = (call_f_goMux1_r && (call_f_unlockFork1_d[0] && call_fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfgo_2_d[0]));
  
  /* mux (Ty Go,
     Ty Pointer_QTree_Bool) : (call_f_unlockFork2,Go) [(call_fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfm1a84,Pointer_QTree_Bool)] > (call_f_goMux2,Pointer_QTree_Bool) */
  assign call_f_goMux2_d = {call_fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfm1a84_d[16:1],
                            (call_f_unlockFork2_d[0] && call_fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfm1a84_d[0])};
  assign call_fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfm1a84_r = (call_f_goMux2_r && (call_f_unlockFork2_d[0] && call_fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfm1a84_d[0]));
  assign call_f_unlockFork2_r = (call_f_goMux2_r && (call_f_unlockFork2_d[0] && call_fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfm1a84_d[0]));
  
  /* mux (Ty Go,
     Ty Pointer_QTree_Bool) : (call_f_unlockFork3,Go) [(call_fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfm2a85,Pointer_QTree_Bool)] > (call_f_goMux3,Pointer_QTree_Bool) */
  assign call_f_goMux3_d = {call_fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfm2a85_d[16:1],
                            (call_f_unlockFork3_d[0] && call_fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfm2a85_d[0])};
  assign call_fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfm2a85_r = (call_f_goMux3_r && (call_f_unlockFork3_d[0] && call_fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfm2a85_d[0]));
  assign call_f_unlockFork3_r = (call_f_goMux3_r && (call_f_unlockFork3_d[0] && call_fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfm2a85_d[0]));
  
  /* mux (Ty Go,
     Ty Pointer_QTree_Bool) : (call_f_unlockFork4,Go) [(call_fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfm3a86,Pointer_QTree_Bool)] > (call_f_goMux4,Pointer_QTree_Bool) */
  assign call_f_goMux4_d = {call_fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfm3a86_d[16:1],
                            (call_f_unlockFork4_d[0] && call_fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfm3a86_d[0])};
  assign call_fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfm3a86_r = (call_f_goMux4_r && (call_f_unlockFork4_d[0] && call_fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfm3a86_d[0]));
  assign call_f_unlockFork4_r = (call_f_goMux4_r && (call_f_unlockFork4_d[0] && call_fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfm3a86_d[0]));
  
  /* mux (Ty Go,
     Ty Pointer_CTf) : (call_f_unlockFork5,Go) [(call_fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfsc_0,Pointer_CTf)] > (call_f_goMux5,Pointer_CTf) */
  assign call_f_goMux5_d = {call_fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfsc_0_d[16:1],
                            (call_f_unlockFork5_d[0] && call_fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfsc_0_d[0])};
  assign call_fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfsc_0_r = (call_f_goMux5_r && (call_f_unlockFork5_d[0] && call_fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfsc_0_d[0]));
  assign call_f_unlockFork5_r = (call_f_goMux5_r && (call_f_unlockFork5_d[0] && call_fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfsc_0_d[0]));
  
  /* buf (Ty QTree_Bool) : (es_0_1es_1_1es_2_1es_3_1QNode_Bool,QTree_Bool) > (lizzieLet10_1_1_argbuf,QTree_Bool) */
  QTree_Bool_t es_0_1es_1_1es_2_1es_3_1QNode_Bool_bufchan_d;
  logic es_0_1es_1_1es_2_1es_3_1QNode_Bool_bufchan_r;
  assign es_0_1es_1_1es_2_1es_3_1QNode_Bool_r = ((! es_0_1es_1_1es_2_1es_3_1QNode_Bool_bufchan_d[0]) || es_0_1es_1_1es_2_1es_3_1QNode_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_0_1es_1_1es_2_1es_3_1QNode_Bool_bufchan_d <= {66'd0, 1'd0};
    else
      if (es_0_1es_1_1es_2_1es_3_1QNode_Bool_r)
        es_0_1es_1_1es_2_1es_3_1QNode_Bool_bufchan_d <= es_0_1es_1_1es_2_1es_3_1QNode_Bool_d;
  QTree_Bool_t es_0_1es_1_1es_2_1es_3_1QNode_Bool_bufchan_buf;
  assign es_0_1es_1_1es_2_1es_3_1QNode_Bool_bufchan_r = (! es_0_1es_1_1es_2_1es_3_1QNode_Bool_bufchan_buf[0]);
  assign lizzieLet10_1_1_argbuf_d = (es_0_1es_1_1es_2_1es_3_1QNode_Bool_bufchan_buf[0] ? es_0_1es_1_1es_2_1es_3_1QNode_Bool_bufchan_buf :
                                     es_0_1es_1_1es_2_1es_3_1QNode_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_0_1es_1_1es_2_1es_3_1QNode_Bool_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((lizzieLet10_1_1_argbuf_r && es_0_1es_1_1es_2_1es_3_1QNode_Bool_bufchan_buf[0]))
        es_0_1es_1_1es_2_1es_3_1QNode_Bool_bufchan_buf <= {66'd0, 1'd0};
      else if (((! lizzieLet10_1_1_argbuf_r) && (! es_0_1es_1_1es_2_1es_3_1QNode_Bool_bufchan_buf[0])))
        es_0_1es_1_1es_2_1es_3_1QNode_Bool_bufchan_buf <= es_0_1es_1_1es_2_1es_3_1QNode_Bool_bufchan_d;
  
  /* buf (Ty QTree_Bool) : (es_4_1es_5_1es_6_1es_7_1QNode_Bool,QTree_Bool) > (lizzieLet35_1_argbuf,QTree_Bool) */
  QTree_Bool_t es_4_1es_5_1es_6_1es_7_1QNode_Bool_bufchan_d;
  logic es_4_1es_5_1es_6_1es_7_1QNode_Bool_bufchan_r;
  assign es_4_1es_5_1es_6_1es_7_1QNode_Bool_r = ((! es_4_1es_5_1es_6_1es_7_1QNode_Bool_bufchan_d[0]) || es_4_1es_5_1es_6_1es_7_1QNode_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_4_1es_5_1es_6_1es_7_1QNode_Bool_bufchan_d <= {66'd0, 1'd0};
    else
      if (es_4_1es_5_1es_6_1es_7_1QNode_Bool_r)
        es_4_1es_5_1es_6_1es_7_1QNode_Bool_bufchan_d <= es_4_1es_5_1es_6_1es_7_1QNode_Bool_d;
  QTree_Bool_t es_4_1es_5_1es_6_1es_7_1QNode_Bool_bufchan_buf;
  assign es_4_1es_5_1es_6_1es_7_1QNode_Bool_bufchan_r = (! es_4_1es_5_1es_6_1es_7_1QNode_Bool_bufchan_buf[0]);
  assign lizzieLet35_1_argbuf_d = (es_4_1es_5_1es_6_1es_7_1QNode_Bool_bufchan_buf[0] ? es_4_1es_5_1es_6_1es_7_1QNode_Bool_bufchan_buf :
                                   es_4_1es_5_1es_6_1es_7_1QNode_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_4_1es_5_1es_6_1es_7_1QNode_Bool_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((lizzieLet35_1_argbuf_r && es_4_1es_5_1es_6_1es_7_1QNode_Bool_bufchan_buf[0]))
        es_4_1es_5_1es_6_1es_7_1QNode_Bool_bufchan_buf <= {66'd0, 1'd0};
      else if (((! lizzieLet35_1_argbuf_r) && (! es_4_1es_5_1es_6_1es_7_1QNode_Bool_bufchan_buf[0])))
        es_4_1es_5_1es_6_1es_7_1QNode_Bool_bufchan_buf <= es_4_1es_5_1es_6_1es_7_1QNode_Bool_bufchan_d;
  
  /* buf (Ty QTree_Bool) : (es_8_1es_9_1es_10_1es_11_1QNode_Bool,QTree_Bool) > (lizzieLet39_1_argbuf,QTree_Bool) */
  QTree_Bool_t es_8_1es_9_1es_10_1es_11_1QNode_Bool_bufchan_d;
  logic es_8_1es_9_1es_10_1es_11_1QNode_Bool_bufchan_r;
  assign es_8_1es_9_1es_10_1es_11_1QNode_Bool_r = ((! es_8_1es_9_1es_10_1es_11_1QNode_Bool_bufchan_d[0]) || es_8_1es_9_1es_10_1es_11_1QNode_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_8_1es_9_1es_10_1es_11_1QNode_Bool_bufchan_d <= {66'd0, 1'd0};
    else
      if (es_8_1es_9_1es_10_1es_11_1QNode_Bool_r)
        es_8_1es_9_1es_10_1es_11_1QNode_Bool_bufchan_d <= es_8_1es_9_1es_10_1es_11_1QNode_Bool_d;
  QTree_Bool_t es_8_1es_9_1es_10_1es_11_1QNode_Bool_bufchan_buf;
  assign es_8_1es_9_1es_10_1es_11_1QNode_Bool_bufchan_r = (! es_8_1es_9_1es_10_1es_11_1QNode_Bool_bufchan_buf[0]);
  assign lizzieLet39_1_argbuf_d = (es_8_1es_9_1es_10_1es_11_1QNode_Bool_bufchan_buf[0] ? es_8_1es_9_1es_10_1es_11_1QNode_Bool_bufchan_buf :
                                   es_8_1es_9_1es_10_1es_11_1QNode_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_8_1es_9_1es_10_1es_11_1QNode_Bool_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((lizzieLet39_1_argbuf_r && es_8_1es_9_1es_10_1es_11_1QNode_Bool_bufchan_buf[0]))
        es_8_1es_9_1es_10_1es_11_1QNode_Bool_bufchan_buf <= {66'd0, 1'd0};
      else if (((! lizzieLet39_1_argbuf_r) && (! es_8_1es_9_1es_10_1es_11_1QNode_Bool_bufchan_buf[0])))
        es_8_1es_9_1es_10_1es_11_1QNode_Bool_bufchan_buf <= es_8_1es_9_1es_10_1es_11_1QNode_Bool_bufchan_d;
  
  /* mergectrl (Ty C12,
           Ty TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool) : [(f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_1,TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool),
                                                                  (f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool2,TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool),
                                                                  (f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool3,TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool),
                                                                  (f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool4,TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool),
                                                                  (f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool5,TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool),
                                                                  (f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool6,TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool),
                                                                  (f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool7,TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool),
                                                                  (f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool8,TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool),
                                                                  (f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool9,TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool),
                                                                  (f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool10,TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool),
                                                                  (f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool11,TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool),
                                                                  (f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool12,TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool)] > (f''''''''''''_choice,C12) (f''''''''''''_data,TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool) */
  logic [11:0] \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_1_select_d ;
  assign \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_1_select_d  = ((| \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_1_select_q ) ? \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_1_select_q  :
                                                                                      (\f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_1_d [0] ? 12'd1 :
                                                                                       (\f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool2_d [0] ? 12'd2 :
                                                                                        (\f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool3_d [0] ? 12'd4 :
                                                                                         (\f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool4_d [0] ? 12'd8 :
                                                                                          (\f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool5_d [0] ? 12'd16 :
                                                                                           (\f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool6_d [0] ? 12'd32 :
                                                                                            (\f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool7_d [0] ? 12'd64 :
                                                                                             (\f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool8_d [0] ? 12'd128 :
                                                                                              (\f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool9_d [0] ? 12'd256 :
                                                                                               (\f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool10_d [0] ? 12'd512 :
                                                                                                (\f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool11_d [0] ? 12'd1024 :
                                                                                                 (\f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool12_d [0] ? 12'd2048 :
                                                                                                  12'd0)))))))))))));
  logic [11:0] \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_1_select_q ;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_1_select_q  <= 12'd0;
    else
      \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_1_select_q  <= (\f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_1_done  ? 12'd0 :
                                                                                    \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_1_select_d );
  logic [1:0] \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_1_emit_q ;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_1_emit_q  <= 2'd0;
    else
      \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_1_emit_q  <= (\f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_1_done  ? 2'd0 :
                                                                                  \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_1_emit_d );
  logic [1:0] \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_1_emit_d ;
  assign \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_1_emit_d  = (\f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_1_emit_q  | ({\f''''''''''''_choice_d [0],
                                                                                                                                                                \f''''''''''''_data_d [0]} & {\f''''''''''''_choice_r ,
                                                                                                                                                                                              \f''''''''''''_data_r }));
  logic \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_1_done ;
  assign \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_1_done  = (& \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_1_emit_d );
  assign {\f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool12_r ,
          \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool11_r ,
          \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool10_r ,
          \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool9_r ,
          \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool8_r ,
          \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool7_r ,
          \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool6_r ,
          \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool5_r ,
          \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool4_r ,
          \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool3_r ,
          \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool2_r ,
          \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_1_r } = (\f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_1_done  ? \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_1_select_d  :
                                                                                 12'd0);
  assign \f''''''''''''_data_d  = ((\f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_1_select_d [0] && (! \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_1_emit_q [0])) ? \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_1_d  :
                                   ((\f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_1_select_d [1] && (! \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_1_emit_q [0])) ? \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool2_d  :
                                    ((\f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_1_select_d [2] && (! \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_1_emit_q [0])) ? \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool3_d  :
                                     ((\f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_1_select_d [3] && (! \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_1_emit_q [0])) ? \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool4_d  :
                                      ((\f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_1_select_d [4] && (! \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_1_emit_q [0])) ? \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool5_d  :
                                       ((\f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_1_select_d [5] && (! \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_1_emit_q [0])) ? \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool6_d  :
                                        ((\f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_1_select_d [6] && (! \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_1_emit_q [0])) ? \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool7_d  :
                                         ((\f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_1_select_d [7] && (! \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_1_emit_q [0])) ? \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool8_d  :
                                          ((\f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_1_select_d [8] && (! \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_1_emit_q [0])) ? \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool9_d  :
                                           ((\f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_1_select_d [9] && (! \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_1_emit_q [0])) ? \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool10_d  :
                                            ((\f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_1_select_d [10] && (! \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_1_emit_q [0])) ? \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool11_d  :
                                             ((\f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_1_select_d [11] && (! \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_1_emit_q [0])) ? \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool12_d  :
                                              {32'd0, 1'd0}))))))))))));
  assign \f''''''''''''_choice_d  = ((\f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_1_select_d [0] && (! \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_1_emit_q [1])) ? C1_12_dc(1'd1) :
                                     ((\f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_1_select_d [1] && (! \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_1_emit_q [1])) ? C2_12_dc(1'd1) :
                                      ((\f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_1_select_d [2] && (! \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_1_emit_q [1])) ? C3_12_dc(1'd1) :
                                       ((\f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_1_select_d [3] && (! \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_1_emit_q [1])) ? C4_12_dc(1'd1) :
                                        ((\f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_1_select_d [4] && (! \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_1_emit_q [1])) ? C5_12_dc(1'd1) :
                                         ((\f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_1_select_d [5] && (! \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_1_emit_q [1])) ? C6_12_dc(1'd1) :
                                          ((\f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_1_select_d [6] && (! \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_1_emit_q [1])) ? C7_12_dc(1'd1) :
                                           ((\f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_1_select_d [7] && (! \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_1_emit_q [1])) ? C8_12_dc(1'd1) :
                                            ((\f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_1_select_d [8] && (! \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_1_emit_q [1])) ? C9_12_dc(1'd1) :
                                             ((\f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_1_select_d [9] && (! \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_1_emit_q [1])) ? C10_12_dc(1'd1) :
                                              ((\f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_1_select_d [10] && (! \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_1_emit_q [1])) ? C11_12_dc(1'd1) :
                                               ((\f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_1_select_d [11] && (! \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_1_emit_q [1])) ? C12_12_dc(1'd1) :
                                                {4'd0, 1'd0}))))))))))));
  
  /* fork (Ty Go) : (f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolgo_5,Go) > [(go_5_1,Go),
                                                                                        (go_5_2,Go)] */
  logic [1:0] \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolgo_5_emitted ;
  logic [1:0] \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolgo_5_done ;
  assign go_5_1_d = (\f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolgo_5_d [0] && (! \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolgo_5_emitted [0]));
  assign go_5_2_d = (\f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolgo_5_d [0] && (! \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolgo_5_emitted [1]));
  assign \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolgo_5_done  = (\f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolgo_5_emitted  | ({go_5_2_d[0],
                                                                                                                                                                   go_5_1_d[0]} & {go_5_2_r,
                                                                                                                                                                                   go_5_1_r}));
  assign \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolgo_5_r  = (& \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolgo_5_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolgo_5_emitted  <= 2'd0;
    else
      \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolgo_5_emitted  <= (\f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolgo_5_r  ? 2'd0 :
                                                                                     \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolgo_5_done );
  
  /* buf (Ty Pointer_QTree_Bool) : (f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolq4a90_1,Pointer_QTree_Bool) > (q4a90_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolq4a90_1_bufchan_d ;
  logic \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolq4a90_1_bufchan_r ;
  assign \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolq4a90_1_r  = ((! \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolq4a90_1_bufchan_d [0]) || \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolq4a90_1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolq4a90_1_bufchan_d  <= {16'd0,
                                                                                          1'd0};
    else
      if (\f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolq4a90_1_r )
        \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolq4a90_1_bufchan_d  <= \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolq4a90_1_d ;
  Pointer_QTree_Bool_t \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolq4a90_1_bufchan_buf ;
  assign \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolq4a90_1_bufchan_r  = (! \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolq4a90_1_bufchan_buf [0]);
  assign q4a90_1_1_argbuf_d = (\f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolq4a90_1_bufchan_buf [0] ? \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolq4a90_1_bufchan_buf  :
                               \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolq4a90_1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolq4a90_1_bufchan_buf  <= {16'd0,
                                                                                            1'd0};
    else
      if ((q4a90_1_1_argbuf_r && \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolq4a90_1_bufchan_buf [0]))
        \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolq4a90_1_bufchan_buf  <= {16'd0,
                                                                                              1'd0};
      else if (((! q4a90_1_1_argbuf_r) && (! \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolq4a90_1_bufchan_buf [0])))
        \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolq4a90_1_bufchan_buf  <= \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolq4a90_1_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Bool) : (f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolt4a91_1,Pointer_QTree_Bool) > (t4a91_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolt4a91_1_bufchan_d ;
  logic \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolt4a91_1_bufchan_r ;
  assign \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolt4a91_1_r  = ((! \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolt4a91_1_bufchan_d [0]) || \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolt4a91_1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolt4a91_1_bufchan_d  <= {16'd0,
                                                                                          1'd0};
    else
      if (\f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolt4a91_1_r )
        \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolt4a91_1_bufchan_d  <= \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolt4a91_1_d ;
  Pointer_QTree_Bool_t \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolt4a91_1_bufchan_buf ;
  assign \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolt4a91_1_bufchan_r  = (! \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolt4a91_1_bufchan_buf [0]);
  assign t4a91_1_1_argbuf_d = (\f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolt4a91_1_bufchan_buf [0] ? \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolt4a91_1_bufchan_buf  :
                               \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolt4a91_1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolt4a91_1_bufchan_buf  <= {16'd0,
                                                                                            1'd0};
    else
      if ((t4a91_1_1_argbuf_r && \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolt4a91_1_bufchan_buf [0]))
        \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolt4a91_1_bufchan_buf  <= {16'd0,
                                                                                              1'd0};
      else if (((! t4a91_1_1_argbuf_r) && (! \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolt4a91_1_bufchan_buf [0])))
        \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolt4a91_1_bufchan_buf  <= \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolt4a91_1_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Bool) : (f''''''''''''_1,Pointer_QTree_Bool) > (f''''''''''''_resbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t \f''''''''''''_1_bufchan_d ;
  logic \f''''''''''''_1_bufchan_r ;
  assign \f''''''''''''_1_r  = ((! \f''''''''''''_1_bufchan_d [0]) || \f''''''''''''_1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \f''''''''''''_1_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\f''''''''''''_1_r )
        \f''''''''''''_1_bufchan_d  <= \f''''''''''''_1_d ;
  Pointer_QTree_Bool_t \f''''''''''''_1_bufchan_buf ;
  assign \f''''''''''''_1_bufchan_r  = (! \f''''''''''''_1_bufchan_buf [0]);
  assign \f''''''''''''_resbuf_d  = (\f''''''''''''_1_bufchan_buf [0] ? \f''''''''''''_1_bufchan_buf  :
                                     \f''''''''''''_1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''''''_1_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((\f''''''''''''_resbuf_r  && \f''''''''''''_1_bufchan_buf [0]))
        \f''''''''''''_1_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! \f''''''''''''_resbuf_r ) && (! \f''''''''''''_1_bufchan_buf [0])))
        \f''''''''''''_1_bufchan_buf  <= \f''''''''''''_1_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Bool) : (f''''''''''''_10,Pointer_QTree_Bool) > (f''''''''''''_10_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t \f''''''''''''_10_bufchan_d ;
  logic \f''''''''''''_10_bufchan_r ;
  assign \f''''''''''''_10_r  = ((! \f''''''''''''_10_bufchan_d [0]) || \f''''''''''''_10_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \f''''''''''''_10_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\f''''''''''''_10_r )
        \f''''''''''''_10_bufchan_d  <= \f''''''''''''_10_d ;
  Pointer_QTree_Bool_t \f''''''''''''_10_bufchan_buf ;
  assign \f''''''''''''_10_bufchan_r  = (! \f''''''''''''_10_bufchan_buf [0]);
  assign \f''''''''''''_10_argbuf_d  = (\f''''''''''''_10_bufchan_buf [0] ? \f''''''''''''_10_bufchan_buf  :
                                        \f''''''''''''_10_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''''''_10_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((\f''''''''''''_10_argbuf_r  && \f''''''''''''_10_bufchan_buf [0]))
        \f''''''''''''_10_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! \f''''''''''''_10_argbuf_r ) && (! \f''''''''''''_10_bufchan_buf [0])))
        \f''''''''''''_10_bufchan_buf  <= \f''''''''''''_10_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Bool) : (f''''''''''''_11,Pointer_QTree_Bool) > (f''''''''''''_11_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t \f''''''''''''_11_bufchan_d ;
  logic \f''''''''''''_11_bufchan_r ;
  assign \f''''''''''''_11_r  = ((! \f''''''''''''_11_bufchan_d [0]) || \f''''''''''''_11_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \f''''''''''''_11_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\f''''''''''''_11_r )
        \f''''''''''''_11_bufchan_d  <= \f''''''''''''_11_d ;
  Pointer_QTree_Bool_t \f''''''''''''_11_bufchan_buf ;
  assign \f''''''''''''_11_bufchan_r  = (! \f''''''''''''_11_bufchan_buf [0]);
  assign \f''''''''''''_11_argbuf_d  = (\f''''''''''''_11_bufchan_buf [0] ? \f''''''''''''_11_bufchan_buf  :
                                        \f''''''''''''_11_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''''''_11_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((\f''''''''''''_11_argbuf_r  && \f''''''''''''_11_bufchan_buf [0]))
        \f''''''''''''_11_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! \f''''''''''''_11_argbuf_r ) && (! \f''''''''''''_11_bufchan_buf [0])))
        \f''''''''''''_11_bufchan_buf  <= \f''''''''''''_11_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Bool) : (f''''''''''''_12,Pointer_QTree_Bool) > (f''''''''''''_12_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t \f''''''''''''_12_bufchan_d ;
  logic \f''''''''''''_12_bufchan_r ;
  assign \f''''''''''''_12_r  = ((! \f''''''''''''_12_bufchan_d [0]) || \f''''''''''''_12_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \f''''''''''''_12_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\f''''''''''''_12_r )
        \f''''''''''''_12_bufchan_d  <= \f''''''''''''_12_d ;
  Pointer_QTree_Bool_t \f''''''''''''_12_bufchan_buf ;
  assign \f''''''''''''_12_bufchan_r  = (! \f''''''''''''_12_bufchan_buf [0]);
  assign \f''''''''''''_12_argbuf_d  = (\f''''''''''''_12_bufchan_buf [0] ? \f''''''''''''_12_bufchan_buf  :
                                        \f''''''''''''_12_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''''''_12_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((\f''''''''''''_12_argbuf_r  && \f''''''''''''_12_bufchan_buf [0]))
        \f''''''''''''_12_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! \f''''''''''''_12_argbuf_r ) && (! \f''''''''''''_12_bufchan_buf [0])))
        \f''''''''''''_12_bufchan_buf  <= \f''''''''''''_12_bufchan_d ;
  
  /* dcon (Ty QTree_Bool,
      Dcon QNode_Bool) : [(f''''''''''''_12_argbuf,Pointer_QTree_Bool),
                          (f''''''''''''_11_argbuf,Pointer_QTree_Bool),
                          (f''''''''''''_10_argbuf,Pointer_QTree_Bool),
                          (f''''''''''''_9_argbuf,Pointer_QTree_Bool)] > (es_8_1es_9_1es_10_1es_11_1QNode_Bool,QTree_Bool) */
  assign es_8_1es_9_1es_10_1es_11_1QNode_Bool_d = QNode_Bool_dc((& {\f''''''''''''_12_argbuf_d [0],
                                                                    \f''''''''''''_11_argbuf_d [0],
                                                                    \f''''''''''''_10_argbuf_d [0],
                                                                    \f''''''''''''_9_argbuf_d [0]}), \f''''''''''''_12_argbuf_d , \f''''''''''''_11_argbuf_d , \f''''''''''''_10_argbuf_d , \f''''''''''''_9_argbuf_d );
  assign {\f''''''''''''_12_argbuf_r ,
          \f''''''''''''_11_argbuf_r ,
          \f''''''''''''_10_argbuf_r ,
          \f''''''''''''_9_argbuf_r } = {4 {(es_8_1es_9_1es_10_1es_11_1QNode_Bool_r && es_8_1es_9_1es_10_1es_11_1QNode_Bool_d[0])}};
  
  /* buf (Ty Pointer_QTree_Bool) : (f''''''''''''_2,Pointer_QTree_Bool) > (f''''''''''''_2_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t \f''''''''''''_2_bufchan_d ;
  logic \f''''''''''''_2_bufchan_r ;
  assign \f''''''''''''_2_r  = ((! \f''''''''''''_2_bufchan_d [0]) || \f''''''''''''_2_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \f''''''''''''_2_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\f''''''''''''_2_r )
        \f''''''''''''_2_bufchan_d  <= \f''''''''''''_2_d ;
  Pointer_QTree_Bool_t \f''''''''''''_2_bufchan_buf ;
  assign \f''''''''''''_2_bufchan_r  = (! \f''''''''''''_2_bufchan_buf [0]);
  assign \f''''''''''''_2_argbuf_d  = (\f''''''''''''_2_bufchan_buf [0] ? \f''''''''''''_2_bufchan_buf  :
                                       \f''''''''''''_2_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''''''_2_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((\f''''''''''''_2_argbuf_r  && \f''''''''''''_2_bufchan_buf [0]))
        \f''''''''''''_2_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! \f''''''''''''_2_argbuf_r ) && (! \f''''''''''''_2_bufchan_buf [0])))
        \f''''''''''''_2_bufchan_buf  <= \f''''''''''''_2_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Bool) : (f''''''''''''_3,Pointer_QTree_Bool) > (f''''''''''''_3_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t \f''''''''''''_3_bufchan_d ;
  logic \f''''''''''''_3_bufchan_r ;
  assign \f''''''''''''_3_r  = ((! \f''''''''''''_3_bufchan_d [0]) || \f''''''''''''_3_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \f''''''''''''_3_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\f''''''''''''_3_r )
        \f''''''''''''_3_bufchan_d  <= \f''''''''''''_3_d ;
  Pointer_QTree_Bool_t \f''''''''''''_3_bufchan_buf ;
  assign \f''''''''''''_3_bufchan_r  = (! \f''''''''''''_3_bufchan_buf [0]);
  assign \f''''''''''''_3_argbuf_d  = (\f''''''''''''_3_bufchan_buf [0] ? \f''''''''''''_3_bufchan_buf  :
                                       \f''''''''''''_3_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''''''_3_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((\f''''''''''''_3_argbuf_r  && \f''''''''''''_3_bufchan_buf [0]))
        \f''''''''''''_3_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! \f''''''''''''_3_argbuf_r ) && (! \f''''''''''''_3_bufchan_buf [0])))
        \f''''''''''''_3_bufchan_buf  <= \f''''''''''''_3_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Bool) : (f''''''''''''_4,Pointer_QTree_Bool) > (f''''''''''''_4_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t \f''''''''''''_4_bufchan_d ;
  logic \f''''''''''''_4_bufchan_r ;
  assign \f''''''''''''_4_r  = ((! \f''''''''''''_4_bufchan_d [0]) || \f''''''''''''_4_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \f''''''''''''_4_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\f''''''''''''_4_r )
        \f''''''''''''_4_bufchan_d  <= \f''''''''''''_4_d ;
  Pointer_QTree_Bool_t \f''''''''''''_4_bufchan_buf ;
  assign \f''''''''''''_4_bufchan_r  = (! \f''''''''''''_4_bufchan_buf [0]);
  assign \f''''''''''''_4_argbuf_d  = (\f''''''''''''_4_bufchan_buf [0] ? \f''''''''''''_4_bufchan_buf  :
                                       \f''''''''''''_4_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''''''_4_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((\f''''''''''''_4_argbuf_r  && \f''''''''''''_4_bufchan_buf [0]))
        \f''''''''''''_4_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! \f''''''''''''_4_argbuf_r ) && (! \f''''''''''''_4_bufchan_buf [0])))
        \f''''''''''''_4_bufchan_buf  <= \f''''''''''''_4_bufchan_d ;
  
  /* dcon (Ty QTree_Bool,
      Dcon QNode_Bool) : [(f''''''''''''_4_argbuf,Pointer_QTree_Bool),
                          (f''''''''''''_3_argbuf,Pointer_QTree_Bool),
                          (f''''''''''''_2_argbuf,Pointer_QTree_Bool),
                          (f''''''''''''_resbuf,Pointer_QTree_Bool)] > (es_0_1es_1_1es_2_1es_3_1QNode_Bool,QTree_Bool) */
  assign es_0_1es_1_1es_2_1es_3_1QNode_Bool_d = QNode_Bool_dc((& {\f''''''''''''_4_argbuf_d [0],
                                                                  \f''''''''''''_3_argbuf_d [0],
                                                                  \f''''''''''''_2_argbuf_d [0],
                                                                  \f''''''''''''_resbuf_d [0]}), \f''''''''''''_4_argbuf_d , \f''''''''''''_3_argbuf_d , \f''''''''''''_2_argbuf_d , \f''''''''''''_resbuf_d );
  assign {\f''''''''''''_4_argbuf_r ,
          \f''''''''''''_3_argbuf_r ,
          \f''''''''''''_2_argbuf_r ,
          \f''''''''''''_resbuf_r } = {4 {(es_0_1es_1_1es_2_1es_3_1QNode_Bool_r && es_0_1es_1_1es_2_1es_3_1QNode_Bool_d[0])}};
  
  /* buf (Ty Pointer_QTree_Bool) : (f''''''''''''_5,Pointer_QTree_Bool) > (f''''''''''''_5_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t \f''''''''''''_5_bufchan_d ;
  logic \f''''''''''''_5_bufchan_r ;
  assign \f''''''''''''_5_r  = ((! \f''''''''''''_5_bufchan_d [0]) || \f''''''''''''_5_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \f''''''''''''_5_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\f''''''''''''_5_r )
        \f''''''''''''_5_bufchan_d  <= \f''''''''''''_5_d ;
  Pointer_QTree_Bool_t \f''''''''''''_5_bufchan_buf ;
  assign \f''''''''''''_5_bufchan_r  = (! \f''''''''''''_5_bufchan_buf [0]);
  assign \f''''''''''''_5_argbuf_d  = (\f''''''''''''_5_bufchan_buf [0] ? \f''''''''''''_5_bufchan_buf  :
                                       \f''''''''''''_5_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''''''_5_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((\f''''''''''''_5_argbuf_r  && \f''''''''''''_5_bufchan_buf [0]))
        \f''''''''''''_5_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! \f''''''''''''_5_argbuf_r ) && (! \f''''''''''''_5_bufchan_buf [0])))
        \f''''''''''''_5_bufchan_buf  <= \f''''''''''''_5_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Bool) : (f''''''''''''_6,Pointer_QTree_Bool) > (f''''''''''''_6_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t \f''''''''''''_6_bufchan_d ;
  logic \f''''''''''''_6_bufchan_r ;
  assign \f''''''''''''_6_r  = ((! \f''''''''''''_6_bufchan_d [0]) || \f''''''''''''_6_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \f''''''''''''_6_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\f''''''''''''_6_r )
        \f''''''''''''_6_bufchan_d  <= \f''''''''''''_6_d ;
  Pointer_QTree_Bool_t \f''''''''''''_6_bufchan_buf ;
  assign \f''''''''''''_6_bufchan_r  = (! \f''''''''''''_6_bufchan_buf [0]);
  assign \f''''''''''''_6_argbuf_d  = (\f''''''''''''_6_bufchan_buf [0] ? \f''''''''''''_6_bufchan_buf  :
                                       \f''''''''''''_6_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''''''_6_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((\f''''''''''''_6_argbuf_r  && \f''''''''''''_6_bufchan_buf [0]))
        \f''''''''''''_6_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! \f''''''''''''_6_argbuf_r ) && (! \f''''''''''''_6_bufchan_buf [0])))
        \f''''''''''''_6_bufchan_buf  <= \f''''''''''''_6_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Bool) : (f''''''''''''_7,Pointer_QTree_Bool) > (f''''''''''''_7_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t \f''''''''''''_7_bufchan_d ;
  logic \f''''''''''''_7_bufchan_r ;
  assign \f''''''''''''_7_r  = ((! \f''''''''''''_7_bufchan_d [0]) || \f''''''''''''_7_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \f''''''''''''_7_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\f''''''''''''_7_r )
        \f''''''''''''_7_bufchan_d  <= \f''''''''''''_7_d ;
  Pointer_QTree_Bool_t \f''''''''''''_7_bufchan_buf ;
  assign \f''''''''''''_7_bufchan_r  = (! \f''''''''''''_7_bufchan_buf [0]);
  assign \f''''''''''''_7_argbuf_d  = (\f''''''''''''_7_bufchan_buf [0] ? \f''''''''''''_7_bufchan_buf  :
                                       \f''''''''''''_7_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''''''_7_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((\f''''''''''''_7_argbuf_r  && \f''''''''''''_7_bufchan_buf [0]))
        \f''''''''''''_7_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! \f''''''''''''_7_argbuf_r ) && (! \f''''''''''''_7_bufchan_buf [0])))
        \f''''''''''''_7_bufchan_buf  <= \f''''''''''''_7_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Bool) : (f''''''''''''_8,Pointer_QTree_Bool) > (f''''''''''''_8_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t \f''''''''''''_8_bufchan_d ;
  logic \f''''''''''''_8_bufchan_r ;
  assign \f''''''''''''_8_r  = ((! \f''''''''''''_8_bufchan_d [0]) || \f''''''''''''_8_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \f''''''''''''_8_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\f''''''''''''_8_r )
        \f''''''''''''_8_bufchan_d  <= \f''''''''''''_8_d ;
  Pointer_QTree_Bool_t \f''''''''''''_8_bufchan_buf ;
  assign \f''''''''''''_8_bufchan_r  = (! \f''''''''''''_8_bufchan_buf [0]);
  assign \f''''''''''''_8_argbuf_d  = (\f''''''''''''_8_bufchan_buf [0] ? \f''''''''''''_8_bufchan_buf  :
                                       \f''''''''''''_8_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''''''_8_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((\f''''''''''''_8_argbuf_r  && \f''''''''''''_8_bufchan_buf [0]))
        \f''''''''''''_8_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! \f''''''''''''_8_argbuf_r ) && (! \f''''''''''''_8_bufchan_buf [0])))
        \f''''''''''''_8_bufchan_buf  <= \f''''''''''''_8_bufchan_d ;
  
  /* dcon (Ty QTree_Bool,
      Dcon QNode_Bool) : [(f''''''''''''_8_argbuf,Pointer_QTree_Bool),
                          (f''''''''''''_7_argbuf,Pointer_QTree_Bool),
                          (f''''''''''''_6_argbuf,Pointer_QTree_Bool),
                          (f''''''''''''_5_argbuf,Pointer_QTree_Bool)] > (es_4_1es_5_1es_6_1es_7_1QNode_Bool,QTree_Bool) */
  assign es_4_1es_5_1es_6_1es_7_1QNode_Bool_d = QNode_Bool_dc((& {\f''''''''''''_8_argbuf_d [0],
                                                                  \f''''''''''''_7_argbuf_d [0],
                                                                  \f''''''''''''_6_argbuf_d [0],
                                                                  \f''''''''''''_5_argbuf_d [0]}), \f''''''''''''_8_argbuf_d , \f''''''''''''_7_argbuf_d , \f''''''''''''_6_argbuf_d , \f''''''''''''_5_argbuf_d );
  assign {\f''''''''''''_8_argbuf_r ,
          \f''''''''''''_7_argbuf_r ,
          \f''''''''''''_6_argbuf_r ,
          \f''''''''''''_5_argbuf_r } = {4 {(es_4_1es_5_1es_6_1es_7_1QNode_Bool_r && es_4_1es_5_1es_6_1es_7_1QNode_Bool_d[0])}};
  
  /* buf (Ty Pointer_QTree_Bool) : (f''''''''''''_9,Pointer_QTree_Bool) > (f''''''''''''_9_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t \f''''''''''''_9_bufchan_d ;
  logic \f''''''''''''_9_bufchan_r ;
  assign \f''''''''''''_9_r  = ((! \f''''''''''''_9_bufchan_d [0]) || \f''''''''''''_9_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \f''''''''''''_9_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\f''''''''''''_9_r )
        \f''''''''''''_9_bufchan_d  <= \f''''''''''''_9_d ;
  Pointer_QTree_Bool_t \f''''''''''''_9_bufchan_buf ;
  assign \f''''''''''''_9_bufchan_r  = (! \f''''''''''''_9_bufchan_buf [0]);
  assign \f''''''''''''_9_argbuf_d  = (\f''''''''''''_9_bufchan_buf [0] ? \f''''''''''''_9_bufchan_buf  :
                                       \f''''''''''''_9_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''''''_9_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((\f''''''''''''_9_argbuf_r  && \f''''''''''''_9_bufchan_buf [0]))
        \f''''''''''''_9_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! \f''''''''''''_9_argbuf_r ) && (! \f''''''''''''_9_bufchan_buf [0])))
        \f''''''''''''_9_bufchan_buf  <= \f''''''''''''_9_bufchan_d ;
  
  /* demux (Ty C12,
       Ty Pointer_QTree_Bool) : (f''''''''''''_choice,C12) (lizzieLet65_4Lf''''''''''''sbos_1_merge_merge_fork_2,Pointer_QTree_Bool) > [(f''''''''''''_1,Pointer_QTree_Bool),
                                                                                                                                        (f''''''''''''_2,Pointer_QTree_Bool),
                                                                                                                                        (f''''''''''''_3,Pointer_QTree_Bool),
                                                                                                                                        (f''''''''''''_4,Pointer_QTree_Bool),
                                                                                                                                        (f''''''''''''_5,Pointer_QTree_Bool),
                                                                                                                                        (f''''''''''''_6,Pointer_QTree_Bool),
                                                                                                                                        (f''''''''''''_7,Pointer_QTree_Bool),
                                                                                                                                        (f''''''''''''_8,Pointer_QTree_Bool),
                                                                                                                                        (f''''''''''''_9,Pointer_QTree_Bool),
                                                                                                                                        (f''''''''''''_10,Pointer_QTree_Bool),
                                                                                                                                        (f''''''''''''_11,Pointer_QTree_Bool),
                                                                                                                                        (f''''''''''''_12,Pointer_QTree_Bool)] */
  logic [11:0] \lizzieLet65_4Lf''''''''''''sbos_1_merge_merge_fork_2_onehotd ;
  always_comb
    if ((\f''''''''''''_choice_d [0] && \lizzieLet65_4Lf''''''''''''sbos_1_merge_merge_fork_2_d [0]))
      unique case (\f''''''''''''_choice_d [4:1])
        4'd0:
          \lizzieLet65_4Lf''''''''''''sbos_1_merge_merge_fork_2_onehotd  = 12'd1;
        4'd1:
          \lizzieLet65_4Lf''''''''''''sbos_1_merge_merge_fork_2_onehotd  = 12'd2;
        4'd2:
          \lizzieLet65_4Lf''''''''''''sbos_1_merge_merge_fork_2_onehotd  = 12'd4;
        4'd3:
          \lizzieLet65_4Lf''''''''''''sbos_1_merge_merge_fork_2_onehotd  = 12'd8;
        4'd4:
          \lizzieLet65_4Lf''''''''''''sbos_1_merge_merge_fork_2_onehotd  = 12'd16;
        4'd5:
          \lizzieLet65_4Lf''''''''''''sbos_1_merge_merge_fork_2_onehotd  = 12'd32;
        4'd6:
          \lizzieLet65_4Lf''''''''''''sbos_1_merge_merge_fork_2_onehotd  = 12'd64;
        4'd7:
          \lizzieLet65_4Lf''''''''''''sbos_1_merge_merge_fork_2_onehotd  = 12'd128;
        4'd8:
          \lizzieLet65_4Lf''''''''''''sbos_1_merge_merge_fork_2_onehotd  = 12'd256;
        4'd9:
          \lizzieLet65_4Lf''''''''''''sbos_1_merge_merge_fork_2_onehotd  = 12'd512;
        4'd10:
          \lizzieLet65_4Lf''''''''''''sbos_1_merge_merge_fork_2_onehotd  = 12'd1024;
        4'd11:
          \lizzieLet65_4Lf''''''''''''sbos_1_merge_merge_fork_2_onehotd  = 12'd2048;
        default:
          \lizzieLet65_4Lf''''''''''''sbos_1_merge_merge_fork_2_onehotd  = 12'd0;
      endcase
    else
      \lizzieLet65_4Lf''''''''''''sbos_1_merge_merge_fork_2_onehotd  = 12'd0;
  assign \f''''''''''''_1_d  = {\lizzieLet65_4Lf''''''''''''sbos_1_merge_merge_fork_2_d [16:1],
                                \lizzieLet65_4Lf''''''''''''sbos_1_merge_merge_fork_2_onehotd [0]};
  assign \f''''''''''''_2_d  = {\lizzieLet65_4Lf''''''''''''sbos_1_merge_merge_fork_2_d [16:1],
                                \lizzieLet65_4Lf''''''''''''sbos_1_merge_merge_fork_2_onehotd [1]};
  assign \f''''''''''''_3_d  = {\lizzieLet65_4Lf''''''''''''sbos_1_merge_merge_fork_2_d [16:1],
                                \lizzieLet65_4Lf''''''''''''sbos_1_merge_merge_fork_2_onehotd [2]};
  assign \f''''''''''''_4_d  = {\lizzieLet65_4Lf''''''''''''sbos_1_merge_merge_fork_2_d [16:1],
                                \lizzieLet65_4Lf''''''''''''sbos_1_merge_merge_fork_2_onehotd [3]};
  assign \f''''''''''''_5_d  = {\lizzieLet65_4Lf''''''''''''sbos_1_merge_merge_fork_2_d [16:1],
                                \lizzieLet65_4Lf''''''''''''sbos_1_merge_merge_fork_2_onehotd [4]};
  assign \f''''''''''''_6_d  = {\lizzieLet65_4Lf''''''''''''sbos_1_merge_merge_fork_2_d [16:1],
                                \lizzieLet65_4Lf''''''''''''sbos_1_merge_merge_fork_2_onehotd [5]};
  assign \f''''''''''''_7_d  = {\lizzieLet65_4Lf''''''''''''sbos_1_merge_merge_fork_2_d [16:1],
                                \lizzieLet65_4Lf''''''''''''sbos_1_merge_merge_fork_2_onehotd [6]};
  assign \f''''''''''''_8_d  = {\lizzieLet65_4Lf''''''''''''sbos_1_merge_merge_fork_2_d [16:1],
                                \lizzieLet65_4Lf''''''''''''sbos_1_merge_merge_fork_2_onehotd [7]};
  assign \f''''''''''''_9_d  = {\lizzieLet65_4Lf''''''''''''sbos_1_merge_merge_fork_2_d [16:1],
                                \lizzieLet65_4Lf''''''''''''sbos_1_merge_merge_fork_2_onehotd [8]};
  assign \f''''''''''''_10_d  = {\lizzieLet65_4Lf''''''''''''sbos_1_merge_merge_fork_2_d [16:1],
                                 \lizzieLet65_4Lf''''''''''''sbos_1_merge_merge_fork_2_onehotd [9]};
  assign \f''''''''''''_11_d  = {\lizzieLet65_4Lf''''''''''''sbos_1_merge_merge_fork_2_d [16:1],
                                 \lizzieLet65_4Lf''''''''''''sbos_1_merge_merge_fork_2_onehotd [10]};
  assign \f''''''''''''_12_d  = {\lizzieLet65_4Lf''''''''''''sbos_1_merge_merge_fork_2_d [16:1],
                                 \lizzieLet65_4Lf''''''''''''sbos_1_merge_merge_fork_2_onehotd [11]};
  assign \lizzieLet65_4Lf''''''''''''sbos_1_merge_merge_fork_2_r  = (| (\lizzieLet65_4Lf''''''''''''sbos_1_merge_merge_fork_2_onehotd  & {\f''''''''''''_12_r ,
                                                                                                                                          \f''''''''''''_11_r ,
                                                                                                                                          \f''''''''''''_10_r ,
                                                                                                                                          \f''''''''''''_9_r ,
                                                                                                                                          \f''''''''''''_8_r ,
                                                                                                                                          \f''''''''''''_7_r ,
                                                                                                                                          \f''''''''''''_6_r ,
                                                                                                                                          \f''''''''''''_5_r ,
                                                                                                                                          \f''''''''''''_4_r ,
                                                                                                                                          \f''''''''''''_3_r ,
                                                                                                                                          \f''''''''''''_2_r ,
                                                                                                                                          \f''''''''''''_1_r }));
  assign \f''''''''''''_choice_r  = \lizzieLet65_4Lf''''''''''''sbos_1_merge_merge_fork_2_r ;
  
  /* destruct (Ty TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool,
          Dcon TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool) : (f''''''''''''_data,TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool) > [(f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolgo_5,Go),
                                                                                                                                          (f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolq4a90_1,Pointer_QTree_Bool),
                                                                                                                                          (f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolt4a91_1,Pointer_QTree_Bool)] */
  logic [2:0] \f''''''''''''_data_emitted ;
  logic [2:0] \f''''''''''''_data_done ;
  assign \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolgo_5_d  = (\f''''''''''''_data_d [0] && (! \f''''''''''''_data_emitted [0]));
  assign \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolq4a90_1_d  = {\f''''''''''''_data_d [16:1],
                                                                                    (\f''''''''''''_data_d [0] && (! \f''''''''''''_data_emitted [1]))};
  assign \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolt4a91_1_d  = {\f''''''''''''_data_d [32:17],
                                                                                    (\f''''''''''''_data_d [0] && (! \f''''''''''''_data_emitted [2]))};
  assign \f''''''''''''_data_done  = (\f''''''''''''_data_emitted  | ({\f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolt4a91_1_d [0],
                                                                       \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolq4a90_1_d [0],
                                                                       \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolgo_5_d [0]} & {\f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolt4a91_1_r ,
                                                                                                                                                   \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolq4a90_1_r ,
                                                                                                                                                   \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolgo_5_r }));
  assign \f''''''''''''_data_r  = (& \f''''''''''''_data_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \f''''''''''''_data_emitted  <= 3'd0;
    else
      \f''''''''''''_data_emitted  <= (\f''''''''''''_data_r  ? 3'd0 :
                                       \f''''''''''''_data_done );
  
  /* destruct (Ty TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool,
          Dcon TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool) : (fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1,TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool) > [(fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgo_4,Go),
                                                                                                                                                                                                                                         (fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm1a84_1,Pointer_QTree_Bool),
                                                                                                                                                                                                                                         (fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm2a85_1,Pointer_QTree_Bool),
                                                                                                                                                                                                                                         (fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm3a86_1,Pointer_QTree_Bool)] */
  logic [3:0] fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1_emitted;
  logic [3:0] fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1_done;
  assign fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgo_4_d = (fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1_d[0] && (! fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1_emitted[0]));
  assign fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm1a84_1_d = {fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1_d[16:1],
                                                                                           (fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1_d[0] && (! fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1_emitted[1]))};
  assign fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm2a85_1_d = {fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1_d[32:17],
                                                                                           (fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1_d[0] && (! fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1_emitted[2]))};
  assign fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm3a86_1_d = {fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1_d[48:33],
                                                                                           (fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1_d[0] && (! fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1_emitted[3]))};
  assign fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1_done = (fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1_emitted | ({fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm3a86_1_d[0],
                                                                                                                                                                             fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm2a85_1_d[0],
                                                                                                                                                                             fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm1a84_1_d[0],
                                                                                                                                                                             fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgo_4_d[0]} & {fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm3a86_1_r,
                                                                                                                                                                                                                                                                fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm2a85_1_r,
                                                                                                                                                                                                                                                                fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm1a84_1_r,
                                                                                                                                                                                                                                                                fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgo_4_r}));
  assign fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1_r = (& fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1_emitted <= 4'd0;
    else
      fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1_emitted <= (fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1_r ? 4'd0 :
                                                                                          fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1_done);
  
  /* fork (Ty Go) : (fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgo_4,Go) > [(go_4_1,Go),
                                                                                                 (go_4_2,Go)] */
  logic [1:0] fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgo_4_emitted;
  logic [1:0] fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgo_4_done;
  assign go_4_1_d = (fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgo_4_d[0] && (! fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgo_4_emitted[0]));
  assign go_4_2_d = (fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgo_4_d[0] && (! fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgo_4_emitted[1]));
  assign fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgo_4_done = (fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgo_4_emitted | ({go_4_2_d[0],
                                                                                                                                                                                 go_4_1_d[0]} & {go_4_2_r,
                                                                                                                                                                                                 go_4_1_r}));
  assign fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgo_4_r = (& fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgo_4_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgo_4_emitted <= 2'd0;
    else
      fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgo_4_emitted <= (fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgo_4_r ? 2'd0 :
                                                                                            fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgo_4_done);
  
  /* buf (Ty Pointer_QTree_Bool) : (fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm1a84_1,Pointer_QTree_Bool) > (m1a84_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm1a84_1_bufchan_d;
  logic fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm1a84_1_bufchan_r;
  assign fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm1a84_1_r = ((! fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm1a84_1_bufchan_d[0]) || fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm1a84_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm1a84_1_bufchan_d <= {16'd0,
                                                                                                 1'd0};
    else
      if (fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm1a84_1_r)
        fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm1a84_1_bufchan_d <= fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm1a84_1_d;
  Pointer_QTree_Bool_t fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm1a84_1_bufchan_buf;
  assign fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm1a84_1_bufchan_r = (! fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm1a84_1_bufchan_buf[0]);
  assign m1a84_1_1_argbuf_d = (fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm1a84_1_bufchan_buf[0] ? fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm1a84_1_bufchan_buf :
                               fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm1a84_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm1a84_1_bufchan_buf <= {16'd0,
                                                                                                   1'd0};
    else
      if ((m1a84_1_1_argbuf_r && fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm1a84_1_bufchan_buf[0]))
        fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm1a84_1_bufchan_buf <= {16'd0,
                                                                                                     1'd0};
      else if (((! m1a84_1_1_argbuf_r) && (! fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm1a84_1_bufchan_buf[0])))
        fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm1a84_1_bufchan_buf <= fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm1a84_1_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm2a85_1,Pointer_QTree_Bool) > (m2a85_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm2a85_1_bufchan_d;
  logic fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm2a85_1_bufchan_r;
  assign fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm2a85_1_r = ((! fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm2a85_1_bufchan_d[0]) || fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm2a85_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm2a85_1_bufchan_d <= {16'd0,
                                                                                                 1'd0};
    else
      if (fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm2a85_1_r)
        fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm2a85_1_bufchan_d <= fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm2a85_1_d;
  Pointer_QTree_Bool_t fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm2a85_1_bufchan_buf;
  assign fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm2a85_1_bufchan_r = (! fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm2a85_1_bufchan_buf[0]);
  assign m2a85_1_1_argbuf_d = (fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm2a85_1_bufchan_buf[0] ? fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm2a85_1_bufchan_buf :
                               fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm2a85_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm2a85_1_bufchan_buf <= {16'd0,
                                                                                                   1'd0};
    else
      if ((m2a85_1_1_argbuf_r && fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm2a85_1_bufchan_buf[0]))
        fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm2a85_1_bufchan_buf <= {16'd0,
                                                                                                     1'd0};
      else if (((! m2a85_1_1_argbuf_r) && (! fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm2a85_1_bufchan_buf[0])))
        fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm2a85_1_bufchan_buf <= fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm2a85_1_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm3a86_1,Pointer_QTree_Bool) > (m3a86_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm3a86_1_bufchan_d;
  logic fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm3a86_1_bufchan_r;
  assign fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm3a86_1_r = ((! fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm3a86_1_bufchan_d[0]) || fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm3a86_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm3a86_1_bufchan_d <= {16'd0,
                                                                                                 1'd0};
    else
      if (fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm3a86_1_r)
        fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm3a86_1_bufchan_d <= fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm3a86_1_d;
  Pointer_QTree_Bool_t fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm3a86_1_bufchan_buf;
  assign fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm3a86_1_bufchan_r = (! fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm3a86_1_bufchan_buf[0]);
  assign m3a86_1_1_argbuf_d = (fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm3a86_1_bufchan_buf[0] ? fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm3a86_1_bufchan_buf :
                               fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm3a86_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm3a86_1_bufchan_buf <= {16'd0,
                                                                                                   1'd0};
    else
      if ((m3a86_1_1_argbuf_r && fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm3a86_1_bufchan_buf[0]))
        fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm3a86_1_bufchan_buf <= {16'd0,
                                                                                                     1'd0};
      else if (((! m3a86_1_1_argbuf_r) && (! fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm3a86_1_bufchan_buf[0])))
        fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm3a86_1_bufchan_buf <= fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm3a86_1_bufchan_d;
  
  /* sink (Ty Pointer_QTree_Bool) : (f_resbuf,Pointer_QTree_Bool) > */
  assign {f_resbuf_r, f_resbuf_dout} = {f_resbuf_rout, f_resbuf_d};
  
  /* dcon (Ty TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool,
      Dcon TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool) : [(go_1_argbuf,Go),
                                                                                    (m1a81_0,Pointer_QTree_Bool),
                                                                                    (m2a82_1,Pointer_QTree_Bool),
                                                                                    (m3a83_2,Pointer_QTree_Bool)] > (fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1,TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool) */
  assign fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1_d = TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_dc((& {go_1_argbuf_d[0],
                                                                                                                                                                 m1a81_0_d[0],
                                                                                                                                                                 m2a82_1_d[0],
                                                                                                                                                                 m3a83_2_d[0]}), go_1_argbuf_d, m1a81_0_d, m2a82_1_d, m3a83_2_d);
  assign {go_1_argbuf_r,
          m1a81_0_r,
          m2a82_1_r,
          m3a83_2_r} = {4 {(fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1_r && fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1_d[0])}};
  
  /* fork (Ty C5) : (go_2_goMux_choice,C5) > [(go_2_goMux_choice_1,C5),
                                         (go_2_goMux_choice_2,C5),
                                         (go_2_goMux_choice_3,C5),
                                         (go_2_goMux_choice_4,C5)] */
  logic [3:0] go_2_goMux_choice_emitted;
  logic [3:0] go_2_goMux_choice_done;
  assign go_2_goMux_choice_1_d = {go_2_goMux_choice_d[3:1],
                                  (go_2_goMux_choice_d[0] && (! go_2_goMux_choice_emitted[0]))};
  assign go_2_goMux_choice_2_d = {go_2_goMux_choice_d[3:1],
                                  (go_2_goMux_choice_d[0] && (! go_2_goMux_choice_emitted[1]))};
  assign go_2_goMux_choice_3_d = {go_2_goMux_choice_d[3:1],
                                  (go_2_goMux_choice_d[0] && (! go_2_goMux_choice_emitted[2]))};
  assign go_2_goMux_choice_4_d = {go_2_goMux_choice_d[3:1],
                                  (go_2_goMux_choice_d[0] && (! go_2_goMux_choice_emitted[3]))};
  assign go_2_goMux_choice_done = (go_2_goMux_choice_emitted | ({go_2_goMux_choice_4_d[0],
                                                                 go_2_goMux_choice_3_d[0],
                                                                 go_2_goMux_choice_2_d[0],
                                                                 go_2_goMux_choice_1_d[0]} & {go_2_goMux_choice_4_r,
                                                                                              go_2_goMux_choice_3_r,
                                                                                              go_2_goMux_choice_2_r,
                                                                                              go_2_goMux_choice_1_r}));
  assign go_2_goMux_choice_r = (& go_2_goMux_choice_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_2_goMux_choice_emitted <= 4'd0;
    else
      go_2_goMux_choice_emitted <= (go_2_goMux_choice_r ? 4'd0 :
                                    go_2_goMux_choice_done);
  
  /* mux (Ty C5,
     Ty Pointer_QTree_Bool) : (go_2_goMux_choice_1,C5) [(call_f_goMux2,Pointer_QTree_Bool),
                                                        (q3a8J_1_1_argbuf,Pointer_QTree_Bool),
                                                        (q2a8I_2_1_argbuf,Pointer_QTree_Bool),
                                                        (q1a8H_3_1_argbuf,Pointer_QTree_Bool),
                                                        (lizzieLet0_4QNode_Bool_4QNode_Bool_3QNode_Bool_1_argbuf,Pointer_QTree_Bool)] > (m1a84_goMux_mux,Pointer_QTree_Bool) */
  logic [16:0] m1a84_goMux_mux_mux;
  logic [4:0] m1a84_goMux_mux_onehot;
  always_comb
    unique case (go_2_goMux_choice_1_d[3:1])
      3'd0:
        {m1a84_goMux_mux_onehot, m1a84_goMux_mux_mux} = {5'd1,
                                                         call_f_goMux2_d};
      3'd1:
        {m1a84_goMux_mux_onehot, m1a84_goMux_mux_mux} = {5'd2,
                                                         q3a8J_1_1_argbuf_d};
      3'd2:
        {m1a84_goMux_mux_onehot, m1a84_goMux_mux_mux} = {5'd4,
                                                         q2a8I_2_1_argbuf_d};
      3'd3:
        {m1a84_goMux_mux_onehot, m1a84_goMux_mux_mux} = {5'd8,
                                                         q1a8H_3_1_argbuf_d};
      3'd4:
        {m1a84_goMux_mux_onehot, m1a84_goMux_mux_mux} = {5'd16,
                                                         lizzieLet0_4QNode_Bool_4QNode_Bool_3QNode_Bool_1_argbuf_d};
      default:
        {m1a84_goMux_mux_onehot, m1a84_goMux_mux_mux} = {5'd0,
                                                         {16'd0, 1'd0}};
    endcase
  assign m1a84_goMux_mux_d = {m1a84_goMux_mux_mux[16:1],
                              (m1a84_goMux_mux_mux[0] && go_2_goMux_choice_1_d[0])};
  assign go_2_goMux_choice_1_r = (m1a84_goMux_mux_d[0] && m1a84_goMux_mux_r);
  assign {lizzieLet0_4QNode_Bool_4QNode_Bool_3QNode_Bool_1_argbuf_r,
          q1a8H_3_1_argbuf_r,
          q2a8I_2_1_argbuf_r,
          q3a8J_1_1_argbuf_r,
          call_f_goMux2_r} = (go_2_goMux_choice_1_r ? m1a84_goMux_mux_onehot :
                              5'd0);
  
  /* mux (Ty C5,
     Ty Pointer_QTree_Bool) : (go_2_goMux_choice_2,C5) [(call_f_goMux3,Pointer_QTree_Bool),
                                                        (t3a8T_1_1_argbuf,Pointer_QTree_Bool),
                                                        (t2a8S_2_1_argbuf,Pointer_QTree_Bool),
                                                        (t1a8R_3_1_argbuf,Pointer_QTree_Bool),
                                                        (lizzieLet0_4QNode_Bool_4QNode_Bool_12QNode_Bool_1_argbuf,Pointer_QTree_Bool)] > (m2a85_goMux_mux,Pointer_QTree_Bool) */
  logic [16:0] m2a85_goMux_mux_mux;
  logic [4:0] m2a85_goMux_mux_onehot;
  always_comb
    unique case (go_2_goMux_choice_2_d[3:1])
      3'd0:
        {m2a85_goMux_mux_onehot, m2a85_goMux_mux_mux} = {5'd1,
                                                         call_f_goMux3_d};
      3'd1:
        {m2a85_goMux_mux_onehot, m2a85_goMux_mux_mux} = {5'd2,
                                                         t3a8T_1_1_argbuf_d};
      3'd2:
        {m2a85_goMux_mux_onehot, m2a85_goMux_mux_mux} = {5'd4,
                                                         t2a8S_2_1_argbuf_d};
      3'd3:
        {m2a85_goMux_mux_onehot, m2a85_goMux_mux_mux} = {5'd8,
                                                         t1a8R_3_1_argbuf_d};
      3'd4:
        {m2a85_goMux_mux_onehot, m2a85_goMux_mux_mux} = {5'd16,
                                                         lizzieLet0_4QNode_Bool_4QNode_Bool_12QNode_Bool_1_argbuf_d};
      default:
        {m2a85_goMux_mux_onehot, m2a85_goMux_mux_mux} = {5'd0,
                                                         {16'd0, 1'd0}};
    endcase
  assign m2a85_goMux_mux_d = {m2a85_goMux_mux_mux[16:1],
                              (m2a85_goMux_mux_mux[0] && go_2_goMux_choice_2_d[0])};
  assign go_2_goMux_choice_2_r = (m2a85_goMux_mux_d[0] && m2a85_goMux_mux_r);
  assign {lizzieLet0_4QNode_Bool_4QNode_Bool_12QNode_Bool_1_argbuf_r,
          t1a8R_3_1_argbuf_r,
          t2a8S_2_1_argbuf_r,
          t3a8T_1_1_argbuf_r,
          call_f_goMux3_r} = (go_2_goMux_choice_2_r ? m2a85_goMux_mux_onehot :
                              5'd0);
  
  /* mux (Ty C5,
     Ty Pointer_QTree_Bool) : (go_2_goMux_choice_3,C5) [(call_f_goMux4,Pointer_QTree_Bool),
                                                        (t3'a8Y_1_1_argbuf,Pointer_QTree_Bool),
                                                        (t2'a8X_2_1_argbuf,Pointer_QTree_Bool),
                                                        (t1'a8W_3_1_argbuf,Pointer_QTree_Bool),
                                                        (t4'a8Z_1_argbuf,Pointer_QTree_Bool)] > (m3a86_goMux_mux,Pointer_QTree_Bool) */
  logic [16:0] m3a86_goMux_mux_mux;
  logic [4:0] m3a86_goMux_mux_onehot;
  always_comb
    unique case (go_2_goMux_choice_3_d[3:1])
      3'd0:
        {m3a86_goMux_mux_onehot, m3a86_goMux_mux_mux} = {5'd1,
                                                         call_f_goMux4_d};
      3'd1:
        {m3a86_goMux_mux_onehot, m3a86_goMux_mux_mux} = {5'd2,
                                                         \t3'a8Y_1_1_argbuf_d };
      3'd2:
        {m3a86_goMux_mux_onehot, m3a86_goMux_mux_mux} = {5'd4,
                                                         \t2'a8X_2_1_argbuf_d };
      3'd3:
        {m3a86_goMux_mux_onehot, m3a86_goMux_mux_mux} = {5'd8,
                                                         \t1'a8W_3_1_argbuf_d };
      3'd4:
        {m3a86_goMux_mux_onehot, m3a86_goMux_mux_mux} = {5'd16,
                                                         \t4'a8Z_1_argbuf_d };
      default:
        {m3a86_goMux_mux_onehot, m3a86_goMux_mux_mux} = {5'd0,
                                                         {16'd0, 1'd0}};
    endcase
  assign m3a86_goMux_mux_d = {m3a86_goMux_mux_mux[16:1],
                              (m3a86_goMux_mux_mux[0] && go_2_goMux_choice_3_d[0])};
  assign go_2_goMux_choice_3_r = (m3a86_goMux_mux_d[0] && m3a86_goMux_mux_r);
  assign {\t4'a8Z_1_argbuf_r ,
          \t1'a8W_3_1_argbuf_r ,
          \t2'a8X_2_1_argbuf_r ,
          \t3'a8Y_1_1_argbuf_r ,
          call_f_goMux4_r} = (go_2_goMux_choice_3_r ? m3a86_goMux_mux_onehot :
                              5'd0);
  
  /* mux (Ty C5,
     Ty Pointer_CTf) : (go_2_goMux_choice_4,C5) [(call_f_goMux5,Pointer_CTf),
                                                 (sca2_1_argbuf,Pointer_CTf),
                                                 (sca1_1_argbuf,Pointer_CTf),
                                                 (sca0_1_argbuf,Pointer_CTf),
                                                 (sca3_1_argbuf,Pointer_CTf)] > (sc_0_goMux_mux,Pointer_CTf) */
  logic [16:0] sc_0_goMux_mux_mux;
  logic [4:0] sc_0_goMux_mux_onehot;
  always_comb
    unique case (go_2_goMux_choice_4_d[3:1])
      3'd0:
        {sc_0_goMux_mux_onehot, sc_0_goMux_mux_mux} = {5'd1,
                                                       call_f_goMux5_d};
      3'd1:
        {sc_0_goMux_mux_onehot, sc_0_goMux_mux_mux} = {5'd2,
                                                       sca2_1_argbuf_d};
      3'd2:
        {sc_0_goMux_mux_onehot, sc_0_goMux_mux_mux} = {5'd4,
                                                       sca1_1_argbuf_d};
      3'd3:
        {sc_0_goMux_mux_onehot, sc_0_goMux_mux_mux} = {5'd8,
                                                       sca0_1_argbuf_d};
      3'd4:
        {sc_0_goMux_mux_onehot, sc_0_goMux_mux_mux} = {5'd16,
                                                       sca3_1_argbuf_d};
      default:
        {sc_0_goMux_mux_onehot, sc_0_goMux_mux_mux} = {5'd0,
                                                       {16'd0, 1'd0}};
    endcase
  assign sc_0_goMux_mux_d = {sc_0_goMux_mux_mux[16:1],
                             (sc_0_goMux_mux_mux[0] && go_2_goMux_choice_4_d[0])};
  assign go_2_goMux_choice_4_r = (sc_0_goMux_mux_d[0] && sc_0_goMux_mux_r);
  assign {sca3_1_argbuf_r,
          sca0_1_argbuf_r,
          sca1_1_argbuf_r,
          sca2_1_argbuf_r,
          call_f_goMux5_r} = (go_2_goMux_choice_4_r ? sc_0_goMux_mux_onehot :
                              5'd0);
  
  /* fork (Ty C5) : (go_3_goMux_choice,C5) > [(go_3_goMux_choice_1,C5),
                                         (go_3_goMux_choice_2,C5),
                                         (go_3_goMux_choice_3,C5)] */
  logic [2:0] go_3_goMux_choice_emitted;
  logic [2:0] go_3_goMux_choice_done;
  assign go_3_goMux_choice_1_d = {go_3_goMux_choice_d[3:1],
                                  (go_3_goMux_choice_d[0] && (! go_3_goMux_choice_emitted[0]))};
  assign go_3_goMux_choice_2_d = {go_3_goMux_choice_d[3:1],
                                  (go_3_goMux_choice_d[0] && (! go_3_goMux_choice_emitted[1]))};
  assign go_3_goMux_choice_3_d = {go_3_goMux_choice_d[3:1],
                                  (go_3_goMux_choice_d[0] && (! go_3_goMux_choice_emitted[2]))};
  assign go_3_goMux_choice_done = (go_3_goMux_choice_emitted | ({go_3_goMux_choice_3_d[0],
                                                                 go_3_goMux_choice_2_d[0],
                                                                 go_3_goMux_choice_1_d[0]} & {go_3_goMux_choice_3_r,
                                                                                              go_3_goMux_choice_2_r,
                                                                                              go_3_goMux_choice_1_r}));
  assign go_3_goMux_choice_r = (& go_3_goMux_choice_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_3_goMux_choice_emitted <= 3'd0;
    else
      go_3_goMux_choice_emitted <= (go_3_goMux_choice_r ? 3'd0 :
                                    go_3_goMux_choice_done);
  
  /* mux (Ty C5,
     Ty Pointer_QTree_Bool) : (go_3_goMux_choice_1,C5) [(call_f''''''''''''_goMux2,Pointer_QTree_Bool),
                                                        (q3a9a_1_1_argbuf,Pointer_QTree_Bool),
                                                        (q2a99_2_1_argbuf,Pointer_QTree_Bool),
                                                        (q1a98_3_1_argbuf,Pointer_QTree_Bool),
                                                        (lizzieLet45_4QNode_Bool_9QNode_Bool_1_argbuf,Pointer_QTree_Bool)] > (q4a90_goMux_mux,Pointer_QTree_Bool) */
  logic [16:0] q4a90_goMux_mux_mux;
  logic [4:0] q4a90_goMux_mux_onehot;
  always_comb
    unique case (go_3_goMux_choice_1_d[3:1])
      3'd0:
        {q4a90_goMux_mux_onehot, q4a90_goMux_mux_mux} = {5'd1,
                                                         \call_f''''''''''''_goMux2_d };
      3'd1:
        {q4a90_goMux_mux_onehot, q4a90_goMux_mux_mux} = {5'd2,
                                                         q3a9a_1_1_argbuf_d};
      3'd2:
        {q4a90_goMux_mux_onehot, q4a90_goMux_mux_mux} = {5'd4,
                                                         q2a99_2_1_argbuf_d};
      3'd3:
        {q4a90_goMux_mux_onehot, q4a90_goMux_mux_mux} = {5'd8,
                                                         q1a98_3_1_argbuf_d};
      3'd4:
        {q4a90_goMux_mux_onehot, q4a90_goMux_mux_mux} = {5'd16,
                                                         lizzieLet45_4QNode_Bool_9QNode_Bool_1_argbuf_d};
      default:
        {q4a90_goMux_mux_onehot, q4a90_goMux_mux_mux} = {5'd0,
                                                         {16'd0, 1'd0}};
    endcase
  assign q4a90_goMux_mux_d = {q4a90_goMux_mux_mux[16:1],
                              (q4a90_goMux_mux_mux[0] && go_3_goMux_choice_1_d[0])};
  assign go_3_goMux_choice_1_r = (q4a90_goMux_mux_d[0] && q4a90_goMux_mux_r);
  assign {lizzieLet45_4QNode_Bool_9QNode_Bool_1_argbuf_r,
          q1a98_3_1_argbuf_r,
          q2a99_2_1_argbuf_r,
          q3a9a_1_1_argbuf_r,
          \call_f''''''''''''_goMux2_r } = (go_3_goMux_choice_1_r ? q4a90_goMux_mux_onehot :
                                            5'd0);
  
  /* mux (Ty C5,
     Ty Pointer_QTree_Bool) : (go_3_goMux_choice_2,C5) [(call_f''''''''''''_goMux3,Pointer_QTree_Bool),
                                                        (t3a9f_1_1_argbuf,Pointer_QTree_Bool),
                                                        (t2a9e_2_1_argbuf,Pointer_QTree_Bool),
                                                        (t1a9d_3_1_argbuf,Pointer_QTree_Bool),
                                                        (t5a9g_1_argbuf,Pointer_QTree_Bool)] > (t4a91_goMux_mux,Pointer_QTree_Bool) */
  logic [16:0] t4a91_goMux_mux_mux;
  logic [4:0] t4a91_goMux_mux_onehot;
  always_comb
    unique case (go_3_goMux_choice_2_d[3:1])
      3'd0:
        {t4a91_goMux_mux_onehot, t4a91_goMux_mux_mux} = {5'd1,
                                                         \call_f''''''''''''_goMux3_d };
      3'd1:
        {t4a91_goMux_mux_onehot, t4a91_goMux_mux_mux} = {5'd2,
                                                         t3a9f_1_1_argbuf_d};
      3'd2:
        {t4a91_goMux_mux_onehot, t4a91_goMux_mux_mux} = {5'd4,
                                                         t2a9e_2_1_argbuf_d};
      3'd3:
        {t4a91_goMux_mux_onehot, t4a91_goMux_mux_mux} = {5'd8,
                                                         t1a9d_3_1_argbuf_d};
      3'd4:
        {t4a91_goMux_mux_onehot, t4a91_goMux_mux_mux} = {5'd16,
                                                         t5a9g_1_argbuf_d};
      default:
        {t4a91_goMux_mux_onehot, t4a91_goMux_mux_mux} = {5'd0,
                                                         {16'd0, 1'd0}};
    endcase
  assign t4a91_goMux_mux_d = {t4a91_goMux_mux_mux[16:1],
                              (t4a91_goMux_mux_mux[0] && go_3_goMux_choice_2_d[0])};
  assign go_3_goMux_choice_2_r = (t4a91_goMux_mux_d[0] && t4a91_goMux_mux_r);
  assign {t5a9g_1_argbuf_r,
          t1a9d_3_1_argbuf_r,
          t2a9e_2_1_argbuf_r,
          t3a9f_1_1_argbuf_r,
          \call_f''''''''''''_goMux3_r } = (go_3_goMux_choice_2_r ? t4a91_goMux_mux_onehot :
                                            5'd0);
  
  /* mux (Ty C5,
     Ty Pointer_CTf'''''''''''') : (go_3_goMux_choice_3,C5) [(call_f''''''''''''_goMux4,Pointer_CTf''''''''''''),
                                                             (sca2_1_1_argbuf,Pointer_CTf''''''''''''),
                                                             (sca1_1_1_argbuf,Pointer_CTf''''''''''''),
                                                             (sca0_1_1_argbuf,Pointer_CTf''''''''''''),
                                                             (sca3_1_1_argbuf,Pointer_CTf'''''''''''')] > (sc_0_1_goMux_mux,Pointer_CTf'''''''''''') */
  logic [16:0] sc_0_1_goMux_mux_mux;
  logic [4:0] sc_0_1_goMux_mux_onehot;
  always_comb
    unique case (go_3_goMux_choice_3_d[3:1])
      3'd0:
        {sc_0_1_goMux_mux_onehot, sc_0_1_goMux_mux_mux} = {5'd1,
                                                           \call_f''''''''''''_goMux4_d };
      3'd1:
        {sc_0_1_goMux_mux_onehot, sc_0_1_goMux_mux_mux} = {5'd2,
                                                           sca2_1_1_argbuf_d};
      3'd2:
        {sc_0_1_goMux_mux_onehot, sc_0_1_goMux_mux_mux} = {5'd4,
                                                           sca1_1_1_argbuf_d};
      3'd3:
        {sc_0_1_goMux_mux_onehot, sc_0_1_goMux_mux_mux} = {5'd8,
                                                           sca0_1_1_argbuf_d};
      3'd4:
        {sc_0_1_goMux_mux_onehot, sc_0_1_goMux_mux_mux} = {5'd16,
                                                           sca3_1_1_argbuf_d};
      default:
        {sc_0_1_goMux_mux_onehot, sc_0_1_goMux_mux_mux} = {5'd0,
                                                           {16'd0, 1'd0}};
    endcase
  assign sc_0_1_goMux_mux_d = {sc_0_1_goMux_mux_mux[16:1],
                               (sc_0_1_goMux_mux_mux[0] && go_3_goMux_choice_3_d[0])};
  assign go_3_goMux_choice_3_r = (sc_0_1_goMux_mux_d[0] && sc_0_1_goMux_mux_r);
  assign {sca3_1_1_argbuf_r,
          sca0_1_1_argbuf_r,
          sca1_1_1_argbuf_r,
          sca2_1_1_argbuf_r,
          \call_f''''''''''''_goMux4_r } = (go_3_goMux_choice_3_r ? sc_0_1_goMux_mux_onehot :
                                            5'd0);
  
  /* dcon (Ty CTf,Dcon Lfsbos) : [(go_4_1,Go)] > (go_4_1Lfsbos,CTf) */
  assign go_4_1Lfsbos_d = Lfsbos_dc((& {go_4_1_d[0]}), go_4_1_d);
  assign {go_4_1_r} = {1 {(go_4_1Lfsbos_r && go_4_1Lfsbos_d[0])}};
  
  /* buf (Ty CTf) : (go_4_1Lfsbos,CTf) > (lizzieLet57_1_argbuf,CTf) */
  CTf_t go_4_1Lfsbos_bufchan_d;
  logic go_4_1Lfsbos_bufchan_r;
  assign go_4_1Lfsbos_r = ((! go_4_1Lfsbos_bufchan_d[0]) || go_4_1Lfsbos_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_4_1Lfsbos_bufchan_d <= {163'd0, 1'd0};
    else if (go_4_1Lfsbos_r) go_4_1Lfsbos_bufchan_d <= go_4_1Lfsbos_d;
  CTf_t go_4_1Lfsbos_bufchan_buf;
  assign go_4_1Lfsbos_bufchan_r = (! go_4_1Lfsbos_bufchan_buf[0]);
  assign lizzieLet57_1_argbuf_d = (go_4_1Lfsbos_bufchan_buf[0] ? go_4_1Lfsbos_bufchan_buf :
                                   go_4_1Lfsbos_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_4_1Lfsbos_bufchan_buf <= {163'd0, 1'd0};
    else
      if ((lizzieLet57_1_argbuf_r && go_4_1Lfsbos_bufchan_buf[0]))
        go_4_1Lfsbos_bufchan_buf <= {163'd0, 1'd0};
      else if (((! lizzieLet57_1_argbuf_r) && (! go_4_1Lfsbos_bufchan_buf[0])))
        go_4_1Lfsbos_bufchan_buf <= go_4_1Lfsbos_bufchan_d;
  
  /* buf (Ty Go) : (go_4_2,Go) > (go_4_2_argbuf,Go) */
  Go_t go_4_2_bufchan_d;
  logic go_4_2_bufchan_r;
  assign go_4_2_r = ((! go_4_2_bufchan_d[0]) || go_4_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_4_2_bufchan_d <= 1'd0;
    else if (go_4_2_r) go_4_2_bufchan_d <= go_4_2_d;
  Go_t go_4_2_bufchan_buf;
  assign go_4_2_bufchan_r = (! go_4_2_bufchan_buf[0]);
  assign go_4_2_argbuf_d = (go_4_2_bufchan_buf[0] ? go_4_2_bufchan_buf :
                            go_4_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_4_2_bufchan_buf <= 1'd0;
    else
      if ((go_4_2_argbuf_r && go_4_2_bufchan_buf[0]))
        go_4_2_bufchan_buf <= 1'd0;
      else if (((! go_4_2_argbuf_r) && (! go_4_2_bufchan_buf[0])))
        go_4_2_bufchan_buf <= go_4_2_bufchan_d;
  
  /* dcon (Ty TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf,
      Dcon TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf) : [(go_4_2_argbuf,Go),
                                                                                                  (m1a84_1_1_argbuf,Pointer_QTree_Bool),
                                                                                                  (m2a85_1_1_argbuf,Pointer_QTree_Bool),
                                                                                                  (m3a86_1_1_argbuf,Pointer_QTree_Bool),
                                                                                                  (lizzieLet33_1_argbuf,Pointer_CTf)] > (call_fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf_1,TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf) */
  assign call_fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf_1_d = TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf_dc((& {go_4_2_argbuf_d[0],
                                                                                                                                                                                                  m1a84_1_1_argbuf_d[0],
                                                                                                                                                                                                  m2a85_1_1_argbuf_d[0],
                                                                                                                                                                                                  m3a86_1_1_argbuf_d[0],
                                                                                                                                                                                                  lizzieLet33_1_argbuf_d[0]}), go_4_2_argbuf_d, m1a84_1_1_argbuf_d, m2a85_1_1_argbuf_d, m3a86_1_1_argbuf_d, lizzieLet33_1_argbuf_d);
  assign {go_4_2_argbuf_r,
          m1a84_1_1_argbuf_r,
          m2a85_1_1_argbuf_r,
          m3a86_1_1_argbuf_r,
          lizzieLet33_1_argbuf_r} = {5 {(call_fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf_1_r && call_fTupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf_1_d[0])}};
  
  /* dcon (Ty CTf'''''''''''',
      Dcon Lf''''''''''''sbos) : [(go_5_1,Go)] > (go_5_1Lf''''''''''''sbos,CTf'''''''''''') */
  assign \go_5_1Lf''''''''''''sbos_d  = \Lf''''''''''''sbos_dc ((& {go_5_1_d[0]}), go_5_1_d);
  assign {go_5_1_r} = {1 {(\go_5_1Lf''''''''''''sbos_r  && \go_5_1Lf''''''''''''sbos_d [0])}};
  
  /* buf (Ty CTf'''''''''''') : (go_5_1Lf''''''''''''sbos,CTf'''''''''''') > (lizzieLet58_1_argbuf,CTf'''''''''''') */
  \CTf''''''''''''_t  \go_5_1Lf''''''''''''sbos_bufchan_d ;
  logic \go_5_1Lf''''''''''''sbos_bufchan_r ;
  assign \go_5_1Lf''''''''''''sbos_r  = ((! \go_5_1Lf''''''''''''sbos_bufchan_d [0]) || \go_5_1Lf''''''''''''sbos_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \go_5_1Lf''''''''''''sbos_bufchan_d  <= {115'd0, 1'd0};
    else
      if (\go_5_1Lf''''''''''''sbos_r )
        \go_5_1Lf''''''''''''sbos_bufchan_d  <= \go_5_1Lf''''''''''''sbos_d ;
  \CTf''''''''''''_t  \go_5_1Lf''''''''''''sbos_bufchan_buf ;
  assign \go_5_1Lf''''''''''''sbos_bufchan_r  = (! \go_5_1Lf''''''''''''sbos_bufchan_buf [0]);
  assign lizzieLet58_1_argbuf_d = (\go_5_1Lf''''''''''''sbos_bufchan_buf [0] ? \go_5_1Lf''''''''''''sbos_bufchan_buf  :
                                   \go_5_1Lf''''''''''''sbos_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \go_5_1Lf''''''''''''sbos_bufchan_buf  <= {115'd0, 1'd0};
    else
      if ((lizzieLet58_1_argbuf_r && \go_5_1Lf''''''''''''sbos_bufchan_buf [0]))
        \go_5_1Lf''''''''''''sbos_bufchan_buf  <= {115'd0, 1'd0};
      else if (((! lizzieLet58_1_argbuf_r) && (! \go_5_1Lf''''''''''''sbos_bufchan_buf [0])))
        \go_5_1Lf''''''''''''sbos_bufchan_buf  <= \go_5_1Lf''''''''''''sbos_bufchan_d ;
  
  /* buf (Ty Go) : (go_5_2,Go) > (go_5_2_argbuf,Go) */
  Go_t go_5_2_bufchan_d;
  logic go_5_2_bufchan_r;
  assign go_5_2_r = ((! go_5_2_bufchan_d[0]) || go_5_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_5_2_bufchan_d <= 1'd0;
    else if (go_5_2_r) go_5_2_bufchan_d <= go_5_2_d;
  Go_t go_5_2_bufchan_buf;
  assign go_5_2_bufchan_r = (! go_5_2_bufchan_buf[0]);
  assign go_5_2_argbuf_d = (go_5_2_bufchan_buf[0] ? go_5_2_bufchan_buf :
                            go_5_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_5_2_bufchan_buf <= 1'd0;
    else
      if ((go_5_2_argbuf_r && go_5_2_bufchan_buf[0]))
        go_5_2_bufchan_buf <= 1'd0;
      else if (((! go_5_2_argbuf_r) && (! go_5_2_bufchan_buf[0])))
        go_5_2_bufchan_buf <= go_5_2_bufchan_d;
  
  /* dcon (Ty TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf'''''''''''',
      Dcon TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf'''''''''''') : [(go_5_2_argbuf,Go),
                                                                                         (q4a90_1_1_argbuf,Pointer_QTree_Bool),
                                                                                         (t4a91_1_1_argbuf,Pointer_QTree_Bool),
                                                                                         (lizzieLet7_1_1_argbuf,Pointer_CTf'''''''''''')] > (call_f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf''''''''''''_1,TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf'''''''''''') */
  assign \call_f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf''''''''''''_1_d  = \TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf''''''''''''_dc ((& {go_5_2_argbuf_d[0],
                                                                                                                                                                                                q4a90_1_1_argbuf_d[0],
                                                                                                                                                                                                t4a91_1_1_argbuf_d[0],
                                                                                                                                                                                                lizzieLet7_1_1_argbuf_d[0]}), go_5_2_argbuf_d, q4a90_1_1_argbuf_d, t4a91_1_1_argbuf_d, lizzieLet7_1_1_argbuf_d);
  assign {go_5_2_argbuf_r,
          q4a90_1_1_argbuf_r,
          t4a91_1_1_argbuf_r,
          lizzieLet7_1_1_argbuf_r} = {4 {(\call_f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf''''''''''''_1_r  && \call_f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf''''''''''''_1_d [0])}};
  
  /* dcon (Ty QTree_Bool,
      Dcon QVal_Bool) : [(go_6_1MyTrue,MyBool)] > (lizzieLet0_1_1QVal_Bool,QTree_Bool) */
  assign lizzieLet0_1_1QVal_Bool_d = QVal_Bool_dc((& {go_6_1MyTrue_d[0]}), go_6_1MyTrue_d);
  assign {go_6_1MyTrue_r} = {1 {(lizzieLet0_1_1QVal_Bool_r && lizzieLet0_1_1QVal_Bool_d[0])}};
  
  /* fork (Ty C40) : (go_7_goMux_choice,C40) > [(go_7_goMux_choice_1,C40),
                                           (go_7_goMux_choice_2,C40)] */
  logic [1:0] go_7_goMux_choice_emitted;
  logic [1:0] go_7_goMux_choice_done;
  assign go_7_goMux_choice_1_d = {go_7_goMux_choice_d[6:1],
                                  (go_7_goMux_choice_d[0] && (! go_7_goMux_choice_emitted[0]))};
  assign go_7_goMux_choice_2_d = {go_7_goMux_choice_d[6:1],
                                  (go_7_goMux_choice_d[0] && (! go_7_goMux_choice_emitted[1]))};
  assign go_7_goMux_choice_done = (go_7_goMux_choice_emitted | ({go_7_goMux_choice_2_d[0],
                                                                 go_7_goMux_choice_1_d[0]} & {go_7_goMux_choice_2_r,
                                                                                              go_7_goMux_choice_1_r}));
  assign go_7_goMux_choice_r = (& go_7_goMux_choice_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_7_goMux_choice_emitted <= 2'd0;
    else
      go_7_goMux_choice_emitted <= (go_7_goMux_choice_r ? 2'd0 :
                                    go_7_goMux_choice_done);
  
  /* mux (Ty C40,
     Ty Pointer_QTree_Bool) : (go_7_goMux_choice_1,C40) [(lizzieLet0_4QNone_Bool_6QNone_Bool_1_argbuf,Pointer_QTree_Bool),
                                                         (contRet_0_1_argbuf,Pointer_QTree_Bool),
                                                         (lizzieLet0_4QNone_Bool_4QVal_Bool_4QNone_Bool_1_argbuf,Pointer_QTree_Bool),
                                                         (lizzieLet8_1_argbuf,Pointer_QTree_Bool),
                                                         (lizzieLet4_1_argbuf,Pointer_QTree_Bool),
                                                         (lizzieLet5_1_argbuf,Pointer_QTree_Bool),
                                                         (lizzieLet9_1_argbuf,Pointer_QTree_Bool),
                                                         (lizzieLet10_1_argbuf,Pointer_QTree_Bool),
                                                         (lizzieLet0_4QNone_Bool_4QNode_Bool_4QNone_Bool_1_argbuf,Pointer_QTree_Bool),
                                                         (lizzieLet11_1_argbuf,Pointer_QTree_Bool),
                                                         (lizzieLet12_1_argbuf,Pointer_QTree_Bool),
                                                         (lizzieLet13_1_argbuf,Pointer_QTree_Bool),
                                                         (lizzieLet14_1_argbuf,Pointer_QTree_Bool),
                                                         (lizzieLet0_4QVal_Bool_4QNone_Bool_4QNone_Bool_1_argbuf,Pointer_QTree_Bool),
                                                         (lizzieLet15_1_argbuf,Pointer_QTree_Bool),
                                                         (lizzieLet16_1_argbuf,Pointer_QTree_Bool),
                                                         (lizzieLet17_1_argbuf,Pointer_QTree_Bool),
                                                         (lizzieLet16_1_1_argbuf,Pointer_QTree_Bool),
                                                         (lizzieLet17_1_1_argbuf,Pointer_QTree_Bool),
                                                         (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_3MyFalse_1_argbuf,Pointer_QTree_Bool),
                                                         (lizzieLet21_1_argbuf,Pointer_QTree_Bool),
                                                         (lizzieLet22_1_argbuf,Pointer_QTree_Bool),
                                                         (lizzieLet18_1_1_argbuf,Pointer_QTree_Bool),
                                                         (lizzieLet19_1_1_argbuf,Pointer_QTree_Bool),
                                                         (lizzieLet26_1_argbuf,Pointer_QTree_Bool),
                                                         (lizzieLet27_1_argbuf,Pointer_QTree_Bool),
                                                         (lizzieLet20_1_argbuf,Pointer_QTree_Bool),
                                                         (lizzieLet21_1_1_argbuf,Pointer_QTree_Bool),
                                                         (lizzieLet22_1_1_argbuf,Pointer_QTree_Bool),
                                                         (lizzieLet23_1_1_argbuf,Pointer_QTree_Bool),
                                                         (lizzieLet0_4QNode_Bool_4QNone_Bool_5QNone_Bool_1_argbuf,Pointer_QTree_Bool),
                                                         (lizzieLet24_1_1_argbuf,Pointer_QTree_Bool),
                                                         (lizzieLet25_1_argbuf,Pointer_QTree_Bool),
                                                         (lizzieLet26_1_1_argbuf,Pointer_QTree_Bool),
                                                         (lizzieLet27_1_1_argbuf,Pointer_QTree_Bool),
                                                         (lizzieLet28_1_1_argbuf,Pointer_QTree_Bool),
                                                         (lizzieLet29_1_1_argbuf,Pointer_QTree_Bool),
                                                         (lizzieLet30_1_1_argbuf,Pointer_QTree_Bool),
                                                         (lizzieLet31_1_1_argbuf,Pointer_QTree_Bool),
                                                         (lizzieLet32_1_argbuf,Pointer_QTree_Bool)] > (srtarg_0_goMux_mux,Pointer_QTree_Bool) */
  logic [16:0] srtarg_0_goMux_mux_mux;
  logic [39:0] srtarg_0_goMux_mux_onehot;
  always_comb
    unique case (go_7_goMux_choice_1_d[6:1])
      6'd0:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {40'd1,
                                                               lizzieLet0_4QNone_Bool_6QNone_Bool_1_argbuf_d};
      6'd1:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {40'd2,
                                                               contRet_0_1_argbuf_d};
      6'd2:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {40'd4,
                                                               lizzieLet0_4QNone_Bool_4QVal_Bool_4QNone_Bool_1_argbuf_d};
      6'd3:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {40'd8,
                                                               lizzieLet8_1_argbuf_d};
      6'd4:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {40'd16,
                                                               lizzieLet4_1_argbuf_d};
      6'd5:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {40'd32,
                                                               lizzieLet5_1_argbuf_d};
      6'd6:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {40'd64,
                                                               lizzieLet9_1_argbuf_d};
      6'd7:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {40'd128,
                                                               lizzieLet10_1_argbuf_d};
      6'd8:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {40'd256,
                                                               lizzieLet0_4QNone_Bool_4QNode_Bool_4QNone_Bool_1_argbuf_d};
      6'd9:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {40'd512,
                                                               lizzieLet11_1_argbuf_d};
      6'd10:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {40'd1024,
                                                               lizzieLet12_1_argbuf_d};
      6'd11:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {40'd2048,
                                                               lizzieLet13_1_argbuf_d};
      6'd12:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {40'd4096,
                                                               lizzieLet14_1_argbuf_d};
      6'd13:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {40'd8192,
                                                               lizzieLet0_4QVal_Bool_4QNone_Bool_4QNone_Bool_1_argbuf_d};
      6'd14:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {40'd16384,
                                                               lizzieLet15_1_argbuf_d};
      6'd15:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {40'd32768,
                                                               lizzieLet16_1_argbuf_d};
      6'd16:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {40'd65536,
                                                               lizzieLet17_1_argbuf_d};
      6'd17:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {40'd131072,
                                                               lizzieLet16_1_1_argbuf_d};
      6'd18:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {40'd262144,
                                                               lizzieLet17_1_1_argbuf_d};
      6'd19:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {40'd524288,
                                                               lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_3MyFalse_1_argbuf_d};
      6'd20:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {40'd1048576,
                                                               lizzieLet21_1_argbuf_d};
      6'd21:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {40'd2097152,
                                                               lizzieLet22_1_argbuf_d};
      6'd22:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {40'd4194304,
                                                               lizzieLet18_1_1_argbuf_d};
      6'd23:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {40'd8388608,
                                                               lizzieLet19_1_1_argbuf_d};
      6'd24:
        {srtarg_0_goMux_mux_onehot,
         srtarg_0_goMux_mux_mux} = {40'd16777216, lizzieLet26_1_argbuf_d};
      6'd25:
        {srtarg_0_goMux_mux_onehot,
         srtarg_0_goMux_mux_mux} = {40'd33554432, lizzieLet27_1_argbuf_d};
      6'd26:
        {srtarg_0_goMux_mux_onehot,
         srtarg_0_goMux_mux_mux} = {40'd67108864, lizzieLet20_1_argbuf_d};
      6'd27:
        {srtarg_0_goMux_mux_onehot,
         srtarg_0_goMux_mux_mux} = {40'd134217728,
                                    lizzieLet21_1_1_argbuf_d};
      6'd28:
        {srtarg_0_goMux_mux_onehot,
         srtarg_0_goMux_mux_mux} = {40'd268435456,
                                    lizzieLet22_1_1_argbuf_d};
      6'd29:
        {srtarg_0_goMux_mux_onehot,
         srtarg_0_goMux_mux_mux} = {40'd536870912,
                                    lizzieLet23_1_1_argbuf_d};
      6'd30:
        {srtarg_0_goMux_mux_onehot,
         srtarg_0_goMux_mux_mux} = {40'd1073741824,
                                    lizzieLet0_4QNode_Bool_4QNone_Bool_5QNone_Bool_1_argbuf_d};
      6'd31:
        {srtarg_0_goMux_mux_onehot,
         srtarg_0_goMux_mux_mux} = {40'd2147483648,
                                    lizzieLet24_1_1_argbuf_d};
      6'd32:
        {srtarg_0_goMux_mux_onehot,
         srtarg_0_goMux_mux_mux} = {40'd4294967296, lizzieLet25_1_argbuf_d};
      6'd33:
        {srtarg_0_goMux_mux_onehot,
         srtarg_0_goMux_mux_mux} = {40'd8589934592,
                                    lizzieLet26_1_1_argbuf_d};
      6'd34:
        {srtarg_0_goMux_mux_onehot,
         srtarg_0_goMux_mux_mux} = {40'd17179869184,
                                    lizzieLet27_1_1_argbuf_d};
      6'd35:
        {srtarg_0_goMux_mux_onehot,
         srtarg_0_goMux_mux_mux} = {40'd34359738368,
                                    lizzieLet28_1_1_argbuf_d};
      6'd36:
        {srtarg_0_goMux_mux_onehot,
         srtarg_0_goMux_mux_mux} = {40'd68719476736,
                                    lizzieLet29_1_1_argbuf_d};
      6'd37:
        {srtarg_0_goMux_mux_onehot,
         srtarg_0_goMux_mux_mux} = {40'd137438953472,
                                    lizzieLet30_1_1_argbuf_d};
      6'd38:
        {srtarg_0_goMux_mux_onehot,
         srtarg_0_goMux_mux_mux} = {40'd274877906944,
                                    lizzieLet31_1_1_argbuf_d};
      6'd39:
        {srtarg_0_goMux_mux_onehot,
         srtarg_0_goMux_mux_mux} = {40'd549755813888,
                                    lizzieLet32_1_argbuf_d};
      default:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {40'd0,
                                                               {16'd0, 1'd0}};
    endcase
  assign srtarg_0_goMux_mux_d = {srtarg_0_goMux_mux_mux[16:1],
                                 (srtarg_0_goMux_mux_mux[0] && go_7_goMux_choice_1_d[0])};
  assign go_7_goMux_choice_1_r = (srtarg_0_goMux_mux_d[0] && srtarg_0_goMux_mux_r);
  assign {lizzieLet32_1_argbuf_r,
          lizzieLet31_1_1_argbuf_r,
          lizzieLet30_1_1_argbuf_r,
          lizzieLet29_1_1_argbuf_r,
          lizzieLet28_1_1_argbuf_r,
          lizzieLet27_1_1_argbuf_r,
          lizzieLet26_1_1_argbuf_r,
          lizzieLet25_1_argbuf_r,
          lizzieLet24_1_1_argbuf_r,
          lizzieLet0_4QNode_Bool_4QNone_Bool_5QNone_Bool_1_argbuf_r,
          lizzieLet23_1_1_argbuf_r,
          lizzieLet22_1_1_argbuf_r,
          lizzieLet21_1_1_argbuf_r,
          lizzieLet20_1_argbuf_r,
          lizzieLet27_1_argbuf_r,
          lizzieLet26_1_argbuf_r,
          lizzieLet19_1_1_argbuf_r,
          lizzieLet18_1_1_argbuf_r,
          lizzieLet22_1_argbuf_r,
          lizzieLet21_1_argbuf_r,
          lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_3MyFalse_1_argbuf_r,
          lizzieLet17_1_1_argbuf_r,
          lizzieLet16_1_1_argbuf_r,
          lizzieLet17_1_argbuf_r,
          lizzieLet16_1_argbuf_r,
          lizzieLet15_1_argbuf_r,
          lizzieLet0_4QVal_Bool_4QNone_Bool_4QNone_Bool_1_argbuf_r,
          lizzieLet14_1_argbuf_r,
          lizzieLet13_1_argbuf_r,
          lizzieLet12_1_argbuf_r,
          lizzieLet11_1_argbuf_r,
          lizzieLet0_4QNone_Bool_4QNode_Bool_4QNone_Bool_1_argbuf_r,
          lizzieLet10_1_argbuf_r,
          lizzieLet9_1_argbuf_r,
          lizzieLet5_1_argbuf_r,
          lizzieLet4_1_argbuf_r,
          lizzieLet8_1_argbuf_r,
          lizzieLet0_4QNone_Bool_4QVal_Bool_4QNone_Bool_1_argbuf_r,
          contRet_0_1_argbuf_r,
          lizzieLet0_4QNone_Bool_6QNone_Bool_1_argbuf_r} = (go_7_goMux_choice_1_r ? srtarg_0_goMux_mux_onehot :
                                                            40'd0);
  
  /* mux (Ty C40,
     Ty Pointer_CTf) : (go_7_goMux_choice_2,C40) [(lizzieLet0_4QNone_Bool_7QNone_Bool_1_argbuf,Pointer_CTf),
                                                  (sc_0_5_1_argbuf,Pointer_CTf),
                                                  (lizzieLet0_4QNone_Bool_4QVal_Bool_5QNone_Bool_1_argbuf,Pointer_CTf),
                                                  (lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_2MyFalse_1_argbuf,Pointer_CTf),
                                                  (lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_2MyTrue_1_argbuf,Pointer_CTf),
                                                  (lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_2MyTrue_1_argbuf,Pointer_CTf),
                                                  (lizzieLet0_4QNone_Bool_4QVal_Bool_5QNode_Bool_1_argbuf,Pointer_CTf),
                                                  (lizzieLet0_4QNone_Bool_4QVal_Bool_5QError_Bool_1_argbuf,Pointer_CTf),
                                                  (lizzieLet0_4QNone_Bool_4QNode_Bool_5QNone_Bool_1_argbuf,Pointer_CTf),
                                                  (lizzieLet0_4QNone_Bool_4QNode_Bool_5QVal_Bool_1_argbuf,Pointer_CTf),
                                                  (lizzieLet0_4QNone_Bool_4QNode_Bool_5QNode_Bool_1_argbuf,Pointer_CTf),
                                                  (lizzieLet0_4QNone_Bool_4QNode_Bool_5QError_Bool_1_argbuf,Pointer_CTf),
                                                  (lizzieLet0_4QNone_Bool_7QError_Bool_1_argbuf,Pointer_CTf),
                                                  (lizzieLet0_4QVal_Bool_4QNone_Bool_5QNone_Bool_1_argbuf,Pointer_CTf),
                                                  (lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_2MyFalse_1_argbuf,Pointer_CTf),
                                                  (lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_2MyTrue_1_argbuf,Pointer_CTf),
                                                  (lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_2MyTrue_1_argbuf,Pointer_CTf),
                                                  (lizzieLet0_4QVal_Bool_4QNone_Bool_5QNode_Bool_1_argbuf,Pointer_CTf),
                                                  (lizzieLet0_4QVal_Bool_4QNone_Bool_5QError_Bool_1_argbuf,Pointer_CTf),
                                                  (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_4MyFalse_1_argbuf,Pointer_CTf),
                                                  (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QNone_Bool_1_argbuf,Pointer_CTf),
                                                  (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QVal_Bool_1_argbuf,Pointer_CTf),
                                                  (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QNode_Bool_1_argbuf,Pointer_CTf),
                                                  (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QError_Bool_1_argbuf,Pointer_CTf),
                                                  (lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QNone_Bool_1_argbuf,Pointer_CTf),
                                                  (lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QVal_Bool_1_argbuf,Pointer_CTf),
                                                  (lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QNode_Bool_1_argbuf,Pointer_CTf),
                                                  (lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QError_Bool_1_argbuf,Pointer_CTf),
                                                  (lizzieLet0_4QVal_Bool_7QNode_Bool_1_argbuf,Pointer_CTf),
                                                  (lizzieLet0_4QVal_Bool_7QError_Bool_1_argbuf,Pointer_CTf),
                                                  (lizzieLet0_4QNode_Bool_4QNone_Bool_6QNone_Bool_1_argbuf,Pointer_CTf),
                                                  (lizzieLet0_4QNode_Bool_4QNone_Bool_6QVal_Bool_1_argbuf,Pointer_CTf),
                                                  (lizzieLet0_4QNode_Bool_4QNone_Bool_6QNode_Bool_1_argbuf,Pointer_CTf),
                                                  (lizzieLet0_4QNode_Bool_4QNone_Bool_6QError_Bool_1_argbuf,Pointer_CTf),
                                                  (lizzieLet0_4QNode_Bool_6QVal_Bool_1_argbuf,Pointer_CTf),
                                                  (lizzieLet0_4QNode_Bool_4QNode_Bool_5QNone_Bool_1_argbuf,Pointer_CTf),
                                                  (lizzieLet0_4QNode_Bool_4QNode_Bool_5QVal_Bool_1_argbuf,Pointer_CTf),
                                                  (lizzieLet0_4QNode_Bool_4QNode_Bool_5QError_Bool_1_argbuf,Pointer_CTf),
                                                  (lizzieLet0_4QNode_Bool_6QError_Bool_1_argbuf,Pointer_CTf),
                                                  (lizzieLet0_9QError_Bool_1_argbuf,Pointer_CTf)] > (scfarg_0_goMux_mux,Pointer_CTf) */
  logic [16:0] scfarg_0_goMux_mux_mux;
  logic [39:0] scfarg_0_goMux_mux_onehot;
  always_comb
    unique case (go_7_goMux_choice_2_d[6:1])
      6'd0:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {40'd1,
                                                               lizzieLet0_4QNone_Bool_7QNone_Bool_1_argbuf_d};
      6'd1:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {40'd2,
                                                               sc_0_5_1_argbuf_d};
      6'd2:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {40'd4,
                                                               lizzieLet0_4QNone_Bool_4QVal_Bool_5QNone_Bool_1_argbuf_d};
      6'd3:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {40'd8,
                                                               lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_2MyFalse_1_argbuf_d};
      6'd4:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {40'd16,
                                                               lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_2MyTrue_1_argbuf_d};
      6'd5:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {40'd32,
                                                               lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_2MyTrue_1_argbuf_d};
      6'd6:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {40'd64,
                                                               lizzieLet0_4QNone_Bool_4QVal_Bool_5QNode_Bool_1_argbuf_d};
      6'd7:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {40'd128,
                                                               lizzieLet0_4QNone_Bool_4QVal_Bool_5QError_Bool_1_argbuf_d};
      6'd8:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {40'd256,
                                                               lizzieLet0_4QNone_Bool_4QNode_Bool_5QNone_Bool_1_argbuf_d};
      6'd9:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {40'd512,
                                                               lizzieLet0_4QNone_Bool_4QNode_Bool_5QVal_Bool_1_argbuf_d};
      6'd10:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {40'd1024,
                                                               lizzieLet0_4QNone_Bool_4QNode_Bool_5QNode_Bool_1_argbuf_d};
      6'd11:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {40'd2048,
                                                               lizzieLet0_4QNone_Bool_4QNode_Bool_5QError_Bool_1_argbuf_d};
      6'd12:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {40'd4096,
                                                               lizzieLet0_4QNone_Bool_7QError_Bool_1_argbuf_d};
      6'd13:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {40'd8192,
                                                               lizzieLet0_4QVal_Bool_4QNone_Bool_5QNone_Bool_1_argbuf_d};
      6'd14:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {40'd16384,
                                                               lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_2MyFalse_1_argbuf_d};
      6'd15:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {40'd32768,
                                                               lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_2MyTrue_1_argbuf_d};
      6'd16:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {40'd65536,
                                                               lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_2MyTrue_1_argbuf_d};
      6'd17:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {40'd131072,
                                                               lizzieLet0_4QVal_Bool_4QNone_Bool_5QNode_Bool_1_argbuf_d};
      6'd18:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {40'd262144,
                                                               lizzieLet0_4QVal_Bool_4QNone_Bool_5QError_Bool_1_argbuf_d};
      6'd19:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {40'd524288,
                                                               lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_4MyFalse_1_argbuf_d};
      6'd20:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {40'd1048576,
                                                               lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QNone_Bool_1_argbuf_d};
      6'd21:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {40'd2097152,
                                                               lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QVal_Bool_1_argbuf_d};
      6'd22:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {40'd4194304,
                                                               lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QNode_Bool_1_argbuf_d};
      6'd23:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {40'd8388608,
                                                               lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QError_Bool_1_argbuf_d};
      6'd24:
        {scfarg_0_goMux_mux_onehot,
         scfarg_0_goMux_mux_mux} = {40'd16777216,
                                    lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QNone_Bool_1_argbuf_d};
      6'd25:
        {scfarg_0_goMux_mux_onehot,
         scfarg_0_goMux_mux_mux} = {40'd33554432,
                                    lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QVal_Bool_1_argbuf_d};
      6'd26:
        {scfarg_0_goMux_mux_onehot,
         scfarg_0_goMux_mux_mux} = {40'd67108864,
                                    lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QNode_Bool_1_argbuf_d};
      6'd27:
        {scfarg_0_goMux_mux_onehot,
         scfarg_0_goMux_mux_mux} = {40'd134217728,
                                    lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QError_Bool_1_argbuf_d};
      6'd28:
        {scfarg_0_goMux_mux_onehot,
         scfarg_0_goMux_mux_mux} = {40'd268435456,
                                    lizzieLet0_4QVal_Bool_7QNode_Bool_1_argbuf_d};
      6'd29:
        {scfarg_0_goMux_mux_onehot,
         scfarg_0_goMux_mux_mux} = {40'd536870912,
                                    lizzieLet0_4QVal_Bool_7QError_Bool_1_argbuf_d};
      6'd30:
        {scfarg_0_goMux_mux_onehot,
         scfarg_0_goMux_mux_mux} = {40'd1073741824,
                                    lizzieLet0_4QNode_Bool_4QNone_Bool_6QNone_Bool_1_argbuf_d};
      6'd31:
        {scfarg_0_goMux_mux_onehot,
         scfarg_0_goMux_mux_mux} = {40'd2147483648,
                                    lizzieLet0_4QNode_Bool_4QNone_Bool_6QVal_Bool_1_argbuf_d};
      6'd32:
        {scfarg_0_goMux_mux_onehot,
         scfarg_0_goMux_mux_mux} = {40'd4294967296,
                                    lizzieLet0_4QNode_Bool_4QNone_Bool_6QNode_Bool_1_argbuf_d};
      6'd33:
        {scfarg_0_goMux_mux_onehot,
         scfarg_0_goMux_mux_mux} = {40'd8589934592,
                                    lizzieLet0_4QNode_Bool_4QNone_Bool_6QError_Bool_1_argbuf_d};
      6'd34:
        {scfarg_0_goMux_mux_onehot,
         scfarg_0_goMux_mux_mux} = {40'd17179869184,
                                    lizzieLet0_4QNode_Bool_6QVal_Bool_1_argbuf_d};
      6'd35:
        {scfarg_0_goMux_mux_onehot,
         scfarg_0_goMux_mux_mux} = {40'd34359738368,
                                    lizzieLet0_4QNode_Bool_4QNode_Bool_5QNone_Bool_1_argbuf_d};
      6'd36:
        {scfarg_0_goMux_mux_onehot,
         scfarg_0_goMux_mux_mux} = {40'd68719476736,
                                    lizzieLet0_4QNode_Bool_4QNode_Bool_5QVal_Bool_1_argbuf_d};
      6'd37:
        {scfarg_0_goMux_mux_onehot,
         scfarg_0_goMux_mux_mux} = {40'd137438953472,
                                    lizzieLet0_4QNode_Bool_4QNode_Bool_5QError_Bool_1_argbuf_d};
      6'd38:
        {scfarg_0_goMux_mux_onehot,
         scfarg_0_goMux_mux_mux} = {40'd274877906944,
                                    lizzieLet0_4QNode_Bool_6QError_Bool_1_argbuf_d};
      6'd39:
        {scfarg_0_goMux_mux_onehot,
         scfarg_0_goMux_mux_mux} = {40'd549755813888,
                                    lizzieLet0_9QError_Bool_1_argbuf_d};
      default:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {40'd0,
                                                               {16'd0, 1'd0}};
    endcase
  assign scfarg_0_goMux_mux_d = {scfarg_0_goMux_mux_mux[16:1],
                                 (scfarg_0_goMux_mux_mux[0] && go_7_goMux_choice_2_d[0])};
  assign go_7_goMux_choice_2_r = (scfarg_0_goMux_mux_d[0] && scfarg_0_goMux_mux_r);
  assign {lizzieLet0_9QError_Bool_1_argbuf_r,
          lizzieLet0_4QNode_Bool_6QError_Bool_1_argbuf_r,
          lizzieLet0_4QNode_Bool_4QNode_Bool_5QError_Bool_1_argbuf_r,
          lizzieLet0_4QNode_Bool_4QNode_Bool_5QVal_Bool_1_argbuf_r,
          lizzieLet0_4QNode_Bool_4QNode_Bool_5QNone_Bool_1_argbuf_r,
          lizzieLet0_4QNode_Bool_6QVal_Bool_1_argbuf_r,
          lizzieLet0_4QNode_Bool_4QNone_Bool_6QError_Bool_1_argbuf_r,
          lizzieLet0_4QNode_Bool_4QNone_Bool_6QNode_Bool_1_argbuf_r,
          lizzieLet0_4QNode_Bool_4QNone_Bool_6QVal_Bool_1_argbuf_r,
          lizzieLet0_4QNode_Bool_4QNone_Bool_6QNone_Bool_1_argbuf_r,
          lizzieLet0_4QVal_Bool_7QError_Bool_1_argbuf_r,
          lizzieLet0_4QVal_Bool_7QNode_Bool_1_argbuf_r,
          lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QError_Bool_1_argbuf_r,
          lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QNode_Bool_1_argbuf_r,
          lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QVal_Bool_1_argbuf_r,
          lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QNone_Bool_1_argbuf_r,
          lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QError_Bool_1_argbuf_r,
          lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QNode_Bool_1_argbuf_r,
          lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QVal_Bool_1_argbuf_r,
          lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QNone_Bool_1_argbuf_r,
          lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_4MyFalse_1_argbuf_r,
          lizzieLet0_4QVal_Bool_4QNone_Bool_5QError_Bool_1_argbuf_r,
          lizzieLet0_4QVal_Bool_4QNone_Bool_5QNode_Bool_1_argbuf_r,
          lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_2MyTrue_1_argbuf_r,
          lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_2MyTrue_1_argbuf_r,
          lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_2MyFalse_1_argbuf_r,
          lizzieLet0_4QVal_Bool_4QNone_Bool_5QNone_Bool_1_argbuf_r,
          lizzieLet0_4QNone_Bool_7QError_Bool_1_argbuf_r,
          lizzieLet0_4QNone_Bool_4QNode_Bool_5QError_Bool_1_argbuf_r,
          lizzieLet0_4QNone_Bool_4QNode_Bool_5QNode_Bool_1_argbuf_r,
          lizzieLet0_4QNone_Bool_4QNode_Bool_5QVal_Bool_1_argbuf_r,
          lizzieLet0_4QNone_Bool_4QNode_Bool_5QNone_Bool_1_argbuf_r,
          lizzieLet0_4QNone_Bool_4QVal_Bool_5QError_Bool_1_argbuf_r,
          lizzieLet0_4QNone_Bool_4QVal_Bool_5QNode_Bool_1_argbuf_r,
          lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_2MyTrue_1_argbuf_r,
          lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_2MyTrue_1_argbuf_r,
          lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_2MyFalse_1_argbuf_r,
          lizzieLet0_4QNone_Bool_4QVal_Bool_5QNone_Bool_1_argbuf_r,
          sc_0_5_1_argbuf_r,
          lizzieLet0_4QNone_Bool_7QNone_Bool_1_argbuf_r} = (go_7_goMux_choice_2_r ? scfarg_0_goMux_mux_onehot :
                                                            40'd0);
  
  /* fork (Ty C12) : (go_8_goMux_choice,C12) > [(go_8_goMux_choice_1,C12),
                                           (go_8_goMux_choice_2,C12)] */
  logic [1:0] go_8_goMux_choice_emitted;
  logic [1:0] go_8_goMux_choice_done;
  assign go_8_goMux_choice_1_d = {go_8_goMux_choice_d[4:1],
                                  (go_8_goMux_choice_d[0] && (! go_8_goMux_choice_emitted[0]))};
  assign go_8_goMux_choice_2_d = {go_8_goMux_choice_d[4:1],
                                  (go_8_goMux_choice_d[0] && (! go_8_goMux_choice_emitted[1]))};
  assign go_8_goMux_choice_done = (go_8_goMux_choice_emitted | ({go_8_goMux_choice_2_d[0],
                                                                 go_8_goMux_choice_1_d[0]} & {go_8_goMux_choice_2_r,
                                                                                              go_8_goMux_choice_1_r}));
  assign go_8_goMux_choice_r = (& go_8_goMux_choice_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_8_goMux_choice_emitted <= 2'd0;
    else
      go_8_goMux_choice_emitted <= (go_8_goMux_choice_r ? 2'd0 :
                                    go_8_goMux_choice_done);
  
  /* mux (Ty C12,
     Ty Pointer_QTree_Bool) : (go_8_goMux_choice_1,C12) [(lizzieLet45_7QNone_Bool_1_argbuf,Pointer_QTree_Bool),
                                                         (contRet_0_1_1_argbuf,Pointer_QTree_Bool),
                                                         (lizzieLet45_4QVal_Bool_4QNone_Bool_1_argbuf,Pointer_QTree_Bool),
                                                         (lizzieLet1_1_1_argbuf,Pointer_QTree_Bool),
                                                         (lizzieLet48_1_argbuf,Pointer_QTree_Bool),
                                                         (lizzieLet49_1_argbuf,Pointer_QTree_Bool),
                                                         (lizzieLet2_1_1_argbuf,Pointer_QTree_Bool),
                                                         (lizzieLet3_1_1_argbuf,Pointer_QTree_Bool),
                                                         (lizzieLet45_4QNode_Bool_4QNone_Bool_1_argbuf,Pointer_QTree_Bool),
                                                         (lizzieLet4_1_1_argbuf,Pointer_QTree_Bool),
                                                         (lizzieLet5_1_1_argbuf,Pointer_QTree_Bool),
                                                         (lizzieLet6_1_1_argbuf,Pointer_QTree_Bool)] > (srtarg_0_1_goMux_mux,Pointer_QTree_Bool) */
  logic [16:0] srtarg_0_1_goMux_mux_mux;
  logic [11:0] srtarg_0_1_goMux_mux_onehot;
  always_comb
    unique case (go_8_goMux_choice_1_d[4:1])
      4'd0:
        {srtarg_0_1_goMux_mux_onehot, srtarg_0_1_goMux_mux_mux} = {12'd1,
                                                                   lizzieLet45_7QNone_Bool_1_argbuf_d};
      4'd1:
        {srtarg_0_1_goMux_mux_onehot, srtarg_0_1_goMux_mux_mux} = {12'd2,
                                                                   contRet_0_1_1_argbuf_d};
      4'd2:
        {srtarg_0_1_goMux_mux_onehot, srtarg_0_1_goMux_mux_mux} = {12'd4,
                                                                   lizzieLet45_4QVal_Bool_4QNone_Bool_1_argbuf_d};
      4'd3:
        {srtarg_0_1_goMux_mux_onehot, srtarg_0_1_goMux_mux_mux} = {12'd8,
                                                                   lizzieLet1_1_1_argbuf_d};
      4'd4:
        {srtarg_0_1_goMux_mux_onehot, srtarg_0_1_goMux_mux_mux} = {12'd16,
                                                                   lizzieLet48_1_argbuf_d};
      4'd5:
        {srtarg_0_1_goMux_mux_onehot, srtarg_0_1_goMux_mux_mux} = {12'd32,
                                                                   lizzieLet49_1_argbuf_d};
      4'd6:
        {srtarg_0_1_goMux_mux_onehot, srtarg_0_1_goMux_mux_mux} = {12'd64,
                                                                   lizzieLet2_1_1_argbuf_d};
      4'd7:
        {srtarg_0_1_goMux_mux_onehot, srtarg_0_1_goMux_mux_mux} = {12'd128,
                                                                   lizzieLet3_1_1_argbuf_d};
      4'd8:
        {srtarg_0_1_goMux_mux_onehot, srtarg_0_1_goMux_mux_mux} = {12'd256,
                                                                   lizzieLet45_4QNode_Bool_4QNone_Bool_1_argbuf_d};
      4'd9:
        {srtarg_0_1_goMux_mux_onehot, srtarg_0_1_goMux_mux_mux} = {12'd512,
                                                                   lizzieLet4_1_1_argbuf_d};
      4'd10:
        {srtarg_0_1_goMux_mux_onehot,
         srtarg_0_1_goMux_mux_mux} = {12'd1024, lizzieLet5_1_1_argbuf_d};
      4'd11:
        {srtarg_0_1_goMux_mux_onehot,
         srtarg_0_1_goMux_mux_mux} = {12'd2048, lizzieLet6_1_1_argbuf_d};
      default:
        {srtarg_0_1_goMux_mux_onehot, srtarg_0_1_goMux_mux_mux} = {12'd0,
                                                                   {16'd0, 1'd0}};
    endcase
  assign srtarg_0_1_goMux_mux_d = {srtarg_0_1_goMux_mux_mux[16:1],
                                   (srtarg_0_1_goMux_mux_mux[0] && go_8_goMux_choice_1_d[0])};
  assign go_8_goMux_choice_1_r = (srtarg_0_1_goMux_mux_d[0] && srtarg_0_1_goMux_mux_r);
  assign {lizzieLet6_1_1_argbuf_r,
          lizzieLet5_1_1_argbuf_r,
          lizzieLet4_1_1_argbuf_r,
          lizzieLet45_4QNode_Bool_4QNone_Bool_1_argbuf_r,
          lizzieLet3_1_1_argbuf_r,
          lizzieLet2_1_1_argbuf_r,
          lizzieLet49_1_argbuf_r,
          lizzieLet48_1_argbuf_r,
          lizzieLet1_1_1_argbuf_r,
          lizzieLet45_4QVal_Bool_4QNone_Bool_1_argbuf_r,
          contRet_0_1_1_argbuf_r,
          lizzieLet45_7QNone_Bool_1_argbuf_r} = (go_8_goMux_choice_1_r ? srtarg_0_1_goMux_mux_onehot :
                                                 12'd0);
  
  /* mux (Ty C12,
     Ty Pointer_CTf'''''''''''') : (go_8_goMux_choice_2,C12) [(lizzieLet45_6QNone_Bool_1_argbuf,Pointer_CTf''''''''''''),
                                                              (sc_0_9_1_argbuf,Pointer_CTf''''''''''''),
                                                              (lizzieLet45_4QVal_Bool_5QNone_Bool_1_argbuf,Pointer_CTf''''''''''''),
                                                              (lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_2MyFalse_1_argbuf,Pointer_CTf''''''''''''),
                                                              (lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_2MyTrue_1_argbuf,Pointer_CTf''''''''''''),
                                                              (lizzieLet45_4QVal_Bool_6QVal_Bool_2MyTrue_1_argbuf,Pointer_CTf''''''''''''),
                                                              (lizzieLet45_4QVal_Bool_5QNode_Bool_1_argbuf,Pointer_CTf''''''''''''),
                                                              (lizzieLet45_4QVal_Bool_5QError_Bool_1_argbuf,Pointer_CTf''''''''''''),
                                                              (lizzieLet45_4QNode_Bool_5QNone_Bool_1_argbuf,Pointer_CTf''''''''''''),
                                                              (lizzieLet45_4QNode_Bool_5QVal_Bool_1_argbuf,Pointer_CTf''''''''''''),
                                                              (lizzieLet45_4QNode_Bool_5QError_Bool_1_argbuf,Pointer_CTf''''''''''''),
                                                              (lizzieLet45_6QError_Bool_1_argbuf,Pointer_CTf'''''''''''')] > (scfarg_0_1_goMux_mux,Pointer_CTf'''''''''''') */
  logic [16:0] scfarg_0_1_goMux_mux_mux;
  logic [11:0] scfarg_0_1_goMux_mux_onehot;
  always_comb
    unique case (go_8_goMux_choice_2_d[4:1])
      4'd0:
        {scfarg_0_1_goMux_mux_onehot, scfarg_0_1_goMux_mux_mux} = {12'd1,
                                                                   lizzieLet45_6QNone_Bool_1_argbuf_d};
      4'd1:
        {scfarg_0_1_goMux_mux_onehot, scfarg_0_1_goMux_mux_mux} = {12'd2,
                                                                   sc_0_9_1_argbuf_d};
      4'd2:
        {scfarg_0_1_goMux_mux_onehot, scfarg_0_1_goMux_mux_mux} = {12'd4,
                                                                   lizzieLet45_4QVal_Bool_5QNone_Bool_1_argbuf_d};
      4'd3:
        {scfarg_0_1_goMux_mux_onehot, scfarg_0_1_goMux_mux_mux} = {12'd8,
                                                                   lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_2MyFalse_1_argbuf_d};
      4'd4:
        {scfarg_0_1_goMux_mux_onehot, scfarg_0_1_goMux_mux_mux} = {12'd16,
                                                                   lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_2MyTrue_1_argbuf_d};
      4'd5:
        {scfarg_0_1_goMux_mux_onehot, scfarg_0_1_goMux_mux_mux} = {12'd32,
                                                                   lizzieLet45_4QVal_Bool_6QVal_Bool_2MyTrue_1_argbuf_d};
      4'd6:
        {scfarg_0_1_goMux_mux_onehot, scfarg_0_1_goMux_mux_mux} = {12'd64,
                                                                   lizzieLet45_4QVal_Bool_5QNode_Bool_1_argbuf_d};
      4'd7:
        {scfarg_0_1_goMux_mux_onehot, scfarg_0_1_goMux_mux_mux} = {12'd128,
                                                                   lizzieLet45_4QVal_Bool_5QError_Bool_1_argbuf_d};
      4'd8:
        {scfarg_0_1_goMux_mux_onehot, scfarg_0_1_goMux_mux_mux} = {12'd256,
                                                                   lizzieLet45_4QNode_Bool_5QNone_Bool_1_argbuf_d};
      4'd9:
        {scfarg_0_1_goMux_mux_onehot, scfarg_0_1_goMux_mux_mux} = {12'd512,
                                                                   lizzieLet45_4QNode_Bool_5QVal_Bool_1_argbuf_d};
      4'd10:
        {scfarg_0_1_goMux_mux_onehot,
         scfarg_0_1_goMux_mux_mux} = {12'd1024,
                                      lizzieLet45_4QNode_Bool_5QError_Bool_1_argbuf_d};
      4'd11:
        {scfarg_0_1_goMux_mux_onehot,
         scfarg_0_1_goMux_mux_mux} = {12'd2048,
                                      lizzieLet45_6QError_Bool_1_argbuf_d};
      default:
        {scfarg_0_1_goMux_mux_onehot, scfarg_0_1_goMux_mux_mux} = {12'd0,
                                                                   {16'd0, 1'd0}};
    endcase
  assign scfarg_0_1_goMux_mux_d = {scfarg_0_1_goMux_mux_mux[16:1],
                                   (scfarg_0_1_goMux_mux_mux[0] && go_8_goMux_choice_2_d[0])};
  assign go_8_goMux_choice_2_r = (scfarg_0_1_goMux_mux_d[0] && scfarg_0_1_goMux_mux_r);
  assign {lizzieLet45_6QError_Bool_1_argbuf_r,
          lizzieLet45_4QNode_Bool_5QError_Bool_1_argbuf_r,
          lizzieLet45_4QNode_Bool_5QVal_Bool_1_argbuf_r,
          lizzieLet45_4QNode_Bool_5QNone_Bool_1_argbuf_r,
          lizzieLet45_4QVal_Bool_5QError_Bool_1_argbuf_r,
          lizzieLet45_4QVal_Bool_5QNode_Bool_1_argbuf_r,
          lizzieLet45_4QVal_Bool_6QVal_Bool_2MyTrue_1_argbuf_r,
          lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_2MyTrue_1_argbuf_r,
          lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_2MyFalse_1_argbuf_r,
          lizzieLet45_4QVal_Bool_5QNone_Bool_1_argbuf_r,
          sc_0_9_1_argbuf_r,
          lizzieLet45_6QNone_Bool_1_argbuf_r} = (go_8_goMux_choice_2_r ? scfarg_0_1_goMux_mux_onehot :
                                                 12'd0);
  
  /* destruct (Ty QTree_Bool,
          Dcon QNode_Bool) : (lizzieLet0_1QNode_Bool,QTree_Bool) > [(q1a8H_destruct,Pointer_QTree_Bool),
                                                                    (q2a8I_destruct,Pointer_QTree_Bool),
                                                                    (q3a8J_destruct,Pointer_QTree_Bool),
                                                                    (q4a8K_destruct,Pointer_QTree_Bool)] */
  logic [3:0] lizzieLet0_1QNode_Bool_emitted;
  logic [3:0] lizzieLet0_1QNode_Bool_done;
  assign q1a8H_destruct_d = {lizzieLet0_1QNode_Bool_d[18:3],
                             (lizzieLet0_1QNode_Bool_d[0] && (! lizzieLet0_1QNode_Bool_emitted[0]))};
  assign q2a8I_destruct_d = {lizzieLet0_1QNode_Bool_d[34:19],
                             (lizzieLet0_1QNode_Bool_d[0] && (! lizzieLet0_1QNode_Bool_emitted[1]))};
  assign q3a8J_destruct_d = {lizzieLet0_1QNode_Bool_d[50:35],
                             (lizzieLet0_1QNode_Bool_d[0] && (! lizzieLet0_1QNode_Bool_emitted[2]))};
  assign q4a8K_destruct_d = {lizzieLet0_1QNode_Bool_d[66:51],
                             (lizzieLet0_1QNode_Bool_d[0] && (! lizzieLet0_1QNode_Bool_emitted[3]))};
  assign lizzieLet0_1QNode_Bool_done = (lizzieLet0_1QNode_Bool_emitted | ({q4a8K_destruct_d[0],
                                                                           q3a8J_destruct_d[0],
                                                                           q2a8I_destruct_d[0],
                                                                           q1a8H_destruct_d[0]} & {q4a8K_destruct_r,
                                                                                                   q3a8J_destruct_r,
                                                                                                   q2a8I_destruct_r,
                                                                                                   q1a8H_destruct_r}));
  assign lizzieLet0_1QNode_Bool_r = (& lizzieLet0_1QNode_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet0_1QNode_Bool_emitted <= 4'd0;
    else
      lizzieLet0_1QNode_Bool_emitted <= (lizzieLet0_1QNode_Bool_r ? 4'd0 :
                                         lizzieLet0_1QNode_Bool_done);
  
  /* destruct (Ty QTree_Bool,
          Dcon QVal_Bool) : (lizzieLet0_1QVal_Bool,QTree_Bool) > [(v1a8m_destruct,MyBool)] */
  assign v1a8m_destruct_d = {lizzieLet0_1QVal_Bool_d[3:3],
                             lizzieLet0_1QVal_Bool_d[0]};
  assign lizzieLet0_1QVal_Bool_r = v1a8m_destruct_r;
  
  /* buf (Ty QTree_Bool) : (lizzieLet0_1_1QVal_Bool,QTree_Bool) > (lizzieLet59_1_argbuf,QTree_Bool) */
  QTree_Bool_t lizzieLet0_1_1QVal_Bool_bufchan_d;
  logic lizzieLet0_1_1QVal_Bool_bufchan_r;
  assign lizzieLet0_1_1QVal_Bool_r = ((! lizzieLet0_1_1QVal_Bool_bufchan_d[0]) || lizzieLet0_1_1QVal_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_1_1QVal_Bool_bufchan_d <= {66'd0, 1'd0};
    else
      if (lizzieLet0_1_1QVal_Bool_r)
        lizzieLet0_1_1QVal_Bool_bufchan_d <= lizzieLet0_1_1QVal_Bool_d;
  QTree_Bool_t lizzieLet0_1_1QVal_Bool_bufchan_buf;
  assign lizzieLet0_1_1QVal_Bool_bufchan_r = (! lizzieLet0_1_1QVal_Bool_bufchan_buf[0]);
  assign lizzieLet59_1_argbuf_d = (lizzieLet0_1_1QVal_Bool_bufchan_buf[0] ? lizzieLet0_1_1QVal_Bool_bufchan_buf :
                                   lizzieLet0_1_1QVal_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_1_1QVal_Bool_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((lizzieLet59_1_argbuf_r && lizzieLet0_1_1QVal_Bool_bufchan_buf[0]))
        lizzieLet0_1_1QVal_Bool_bufchan_buf <= {66'd0, 1'd0};
      else if (((! lizzieLet59_1_argbuf_r) && (! lizzieLet0_1_1QVal_Bool_bufchan_buf[0])))
        lizzieLet0_1_1QVal_Bool_bufchan_buf <= lizzieLet0_1_1QVal_Bool_bufchan_d;
  
  /* demux (Ty QTree_Bool,
       Ty QTree_Bool) : (lizzieLet0_2,QTree_Bool) (lizzieLet0_1,QTree_Bool) > [(_168,QTree_Bool),
                                                                               (lizzieLet0_1QVal_Bool,QTree_Bool),
                                                                               (lizzieLet0_1QNode_Bool,QTree_Bool),
                                                                               (_167,QTree_Bool)] */
  logic [3:0] lizzieLet0_1_onehotd;
  always_comb
    if ((lizzieLet0_2_d[0] && lizzieLet0_1_d[0]))
      unique case (lizzieLet0_2_d[2:1])
        2'd0: lizzieLet0_1_onehotd = 4'd1;
        2'd1: lizzieLet0_1_onehotd = 4'd2;
        2'd2: lizzieLet0_1_onehotd = 4'd4;
        2'd3: lizzieLet0_1_onehotd = 4'd8;
        default: lizzieLet0_1_onehotd = 4'd0;
      endcase
    else lizzieLet0_1_onehotd = 4'd0;
  assign _168_d = {lizzieLet0_1_d[66:1], lizzieLet0_1_onehotd[0]};
  assign lizzieLet0_1QVal_Bool_d = {lizzieLet0_1_d[66:1],
                                    lizzieLet0_1_onehotd[1]};
  assign lizzieLet0_1QNode_Bool_d = {lizzieLet0_1_d[66:1],
                                     lizzieLet0_1_onehotd[2]};
  assign _167_d = {lizzieLet0_1_d[66:1], lizzieLet0_1_onehotd[3]};
  assign lizzieLet0_1_r = (| (lizzieLet0_1_onehotd & {_167_r,
                                                      lizzieLet0_1QNode_Bool_r,
                                                      lizzieLet0_1QVal_Bool_r,
                                                      _168_r}));
  assign lizzieLet0_2_r = lizzieLet0_1_r;
  
  /* demux (Ty QTree_Bool,
       Ty Go) : (lizzieLet0_3,QTree_Bool) (go_2_goMux_data,Go) > [(lizzieLet0_3QNone_Bool,Go),
                                                                  (lizzieLet0_3QVal_Bool,Go),
                                                                  (lizzieLet0_3QNode_Bool,Go),
                                                                  (lizzieLet0_3QError_Bool,Go)] */
  logic [3:0] go_2_goMux_data_onehotd;
  always_comb
    if ((lizzieLet0_3_d[0] && go_2_goMux_data_d[0]))
      unique case (lizzieLet0_3_d[2:1])
        2'd0: go_2_goMux_data_onehotd = 4'd1;
        2'd1: go_2_goMux_data_onehotd = 4'd2;
        2'd2: go_2_goMux_data_onehotd = 4'd4;
        2'd3: go_2_goMux_data_onehotd = 4'd8;
        default: go_2_goMux_data_onehotd = 4'd0;
      endcase
    else go_2_goMux_data_onehotd = 4'd0;
  assign lizzieLet0_3QNone_Bool_d = go_2_goMux_data_onehotd[0];
  assign lizzieLet0_3QVal_Bool_d = go_2_goMux_data_onehotd[1];
  assign lizzieLet0_3QNode_Bool_d = go_2_goMux_data_onehotd[2];
  assign lizzieLet0_3QError_Bool_d = go_2_goMux_data_onehotd[3];
  assign go_2_goMux_data_r = (| (go_2_goMux_data_onehotd & {lizzieLet0_3QError_Bool_r,
                                                            lizzieLet0_3QNode_Bool_r,
                                                            lizzieLet0_3QVal_Bool_r,
                                                            lizzieLet0_3QNone_Bool_r}));
  assign lizzieLet0_3_r = go_2_goMux_data_r;
  
  /* fork (Ty Go) : (lizzieLet0_3QError_Bool,Go) > [(lizzieLet0_3QError_Bool_1,Go),
                                               (lizzieLet0_3QError_Bool_2,Go)] */
  logic [1:0] lizzieLet0_3QError_Bool_emitted;
  logic [1:0] lizzieLet0_3QError_Bool_done;
  assign lizzieLet0_3QError_Bool_1_d = (lizzieLet0_3QError_Bool_d[0] && (! lizzieLet0_3QError_Bool_emitted[0]));
  assign lizzieLet0_3QError_Bool_2_d = (lizzieLet0_3QError_Bool_d[0] && (! lizzieLet0_3QError_Bool_emitted[1]));
  assign lizzieLet0_3QError_Bool_done = (lizzieLet0_3QError_Bool_emitted | ({lizzieLet0_3QError_Bool_2_d[0],
                                                                             lizzieLet0_3QError_Bool_1_d[0]} & {lizzieLet0_3QError_Bool_2_r,
                                                                                                                lizzieLet0_3QError_Bool_1_r}));
  assign lizzieLet0_3QError_Bool_r = (& lizzieLet0_3QError_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet0_3QError_Bool_emitted <= 2'd0;
    else
      lizzieLet0_3QError_Bool_emitted <= (lizzieLet0_3QError_Bool_r ? 2'd0 :
                                          lizzieLet0_3QError_Bool_done);
  
  /* dcon (Ty QTree_Bool,
      Dcon QError_Bool) : [(lizzieLet0_3QError_Bool_1,Go)] > (lizzieLet0_3QError_Bool_1QError_Bool,QTree_Bool) */
  assign lizzieLet0_3QError_Bool_1QError_Bool_d = QError_Bool_dc((& {lizzieLet0_3QError_Bool_1_d[0]}), lizzieLet0_3QError_Bool_1_d);
  assign {lizzieLet0_3QError_Bool_1_r} = {1 {(lizzieLet0_3QError_Bool_1QError_Bool_r && lizzieLet0_3QError_Bool_1QError_Bool_d[0])}};
  
  /* buf (Ty QTree_Bool) : (lizzieLet0_3QError_Bool_1QError_Bool,QTree_Bool) > (lizzieLet44_1_argbuf,QTree_Bool) */
  QTree_Bool_t lizzieLet0_3QError_Bool_1QError_Bool_bufchan_d;
  logic lizzieLet0_3QError_Bool_1QError_Bool_bufchan_r;
  assign lizzieLet0_3QError_Bool_1QError_Bool_r = ((! lizzieLet0_3QError_Bool_1QError_Bool_bufchan_d[0]) || lizzieLet0_3QError_Bool_1QError_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_3QError_Bool_1QError_Bool_bufchan_d <= {66'd0, 1'd0};
    else
      if (lizzieLet0_3QError_Bool_1QError_Bool_r)
        lizzieLet0_3QError_Bool_1QError_Bool_bufchan_d <= lizzieLet0_3QError_Bool_1QError_Bool_d;
  QTree_Bool_t lizzieLet0_3QError_Bool_1QError_Bool_bufchan_buf;
  assign lizzieLet0_3QError_Bool_1QError_Bool_bufchan_r = (! lizzieLet0_3QError_Bool_1QError_Bool_bufchan_buf[0]);
  assign lizzieLet44_1_argbuf_d = (lizzieLet0_3QError_Bool_1QError_Bool_bufchan_buf[0] ? lizzieLet0_3QError_Bool_1QError_Bool_bufchan_buf :
                                   lizzieLet0_3QError_Bool_1QError_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_3QError_Bool_1QError_Bool_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((lizzieLet44_1_argbuf_r && lizzieLet0_3QError_Bool_1QError_Bool_bufchan_buf[0]))
        lizzieLet0_3QError_Bool_1QError_Bool_bufchan_buf <= {66'd0, 1'd0};
      else if (((! lizzieLet44_1_argbuf_r) && (! lizzieLet0_3QError_Bool_1QError_Bool_bufchan_buf[0])))
        lizzieLet0_3QError_Bool_1QError_Bool_bufchan_buf <= lizzieLet0_3QError_Bool_1QError_Bool_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet0_3QError_Bool_2,Go) > (lizzieLet0_3QError_Bool_2_argbuf,Go) */
  Go_t lizzieLet0_3QError_Bool_2_bufchan_d;
  logic lizzieLet0_3QError_Bool_2_bufchan_r;
  assign lizzieLet0_3QError_Bool_2_r = ((! lizzieLet0_3QError_Bool_2_bufchan_d[0]) || lizzieLet0_3QError_Bool_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet0_3QError_Bool_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet0_3QError_Bool_2_r)
        lizzieLet0_3QError_Bool_2_bufchan_d <= lizzieLet0_3QError_Bool_2_d;
  Go_t lizzieLet0_3QError_Bool_2_bufchan_buf;
  assign lizzieLet0_3QError_Bool_2_bufchan_r = (! lizzieLet0_3QError_Bool_2_bufchan_buf[0]);
  assign lizzieLet0_3QError_Bool_2_argbuf_d = (lizzieLet0_3QError_Bool_2_bufchan_buf[0] ? lizzieLet0_3QError_Bool_2_bufchan_buf :
                                               lizzieLet0_3QError_Bool_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet0_3QError_Bool_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet0_3QError_Bool_2_argbuf_r && lizzieLet0_3QError_Bool_2_bufchan_buf[0]))
        lizzieLet0_3QError_Bool_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet0_3QError_Bool_2_argbuf_r) && (! lizzieLet0_3QError_Bool_2_bufchan_buf[0])))
        lizzieLet0_3QError_Bool_2_bufchan_buf <= lizzieLet0_3QError_Bool_2_bufchan_d;
  
  /* demux (Ty QTree_Bool,
       Ty QTree_Bool) : (lizzieLet0_4,QTree_Bool) (readPointer_QTree_Boolm2a85_1_argbuf_rwb,QTree_Bool) > [(lizzieLet0_4QNone_Bool,QTree_Bool),
                                                                                                           (lizzieLet0_4QVal_Bool,QTree_Bool),
                                                                                                           (lizzieLet0_4QNode_Bool,QTree_Bool),
                                                                                                           (_166,QTree_Bool)] */
  logic [3:0] readPointer_QTree_Boolm2a85_1_argbuf_rwb_onehotd;
  always_comb
    if ((lizzieLet0_4_d[0] && readPointer_QTree_Boolm2a85_1_argbuf_rwb_d[0]))
      unique case (lizzieLet0_4_d[2:1])
        2'd0: readPointer_QTree_Boolm2a85_1_argbuf_rwb_onehotd = 4'd1;
        2'd1: readPointer_QTree_Boolm2a85_1_argbuf_rwb_onehotd = 4'd2;
        2'd2: readPointer_QTree_Boolm2a85_1_argbuf_rwb_onehotd = 4'd4;
        2'd3: readPointer_QTree_Boolm2a85_1_argbuf_rwb_onehotd = 4'd8;
        default: readPointer_QTree_Boolm2a85_1_argbuf_rwb_onehotd = 4'd0;
      endcase
    else readPointer_QTree_Boolm2a85_1_argbuf_rwb_onehotd = 4'd0;
  assign lizzieLet0_4QNone_Bool_d = {readPointer_QTree_Boolm2a85_1_argbuf_rwb_d[66:1],
                                     readPointer_QTree_Boolm2a85_1_argbuf_rwb_onehotd[0]};
  assign lizzieLet0_4QVal_Bool_d = {readPointer_QTree_Boolm2a85_1_argbuf_rwb_d[66:1],
                                    readPointer_QTree_Boolm2a85_1_argbuf_rwb_onehotd[1]};
  assign lizzieLet0_4QNode_Bool_d = {readPointer_QTree_Boolm2a85_1_argbuf_rwb_d[66:1],
                                     readPointer_QTree_Boolm2a85_1_argbuf_rwb_onehotd[2]};
  assign _166_d = {readPointer_QTree_Boolm2a85_1_argbuf_rwb_d[66:1],
                   readPointer_QTree_Boolm2a85_1_argbuf_rwb_onehotd[3]};
  assign readPointer_QTree_Boolm2a85_1_argbuf_rwb_r = (| (readPointer_QTree_Boolm2a85_1_argbuf_rwb_onehotd & {_166_r,
                                                                                                              lizzieLet0_4QNode_Bool_r,
                                                                                                              lizzieLet0_4QVal_Bool_r,
                                                                                                              lizzieLet0_4QNone_Bool_r}));
  assign lizzieLet0_4_r = readPointer_QTree_Boolm2a85_1_argbuf_rwb_r;
  
  /* fork (Ty QTree_Bool) : (lizzieLet0_4QNode_Bool,QTree_Bool) > [(lizzieLet0_4QNode_Bool_1,QTree_Bool),
                                                              (lizzieLet0_4QNode_Bool_2,QTree_Bool),
                                                              (lizzieLet0_4QNode_Bool_3,QTree_Bool),
                                                              (lizzieLet0_4QNode_Bool_4,QTree_Bool),
                                                              (lizzieLet0_4QNode_Bool_5,QTree_Bool),
                                                              (lizzieLet0_4QNode_Bool_6,QTree_Bool),
                                                              (lizzieLet0_4QNode_Bool_7,QTree_Bool),
                                                              (lizzieLet0_4QNode_Bool_8,QTree_Bool),
                                                              (lizzieLet0_4QNode_Bool_9,QTree_Bool),
                                                              (lizzieLet0_4QNode_Bool_10,QTree_Bool)] */
  logic [9:0] lizzieLet0_4QNode_Bool_emitted;
  logic [9:0] lizzieLet0_4QNode_Bool_done;
  assign lizzieLet0_4QNode_Bool_1_d = {lizzieLet0_4QNode_Bool_d[66:1],
                                       (lizzieLet0_4QNode_Bool_d[0] && (! lizzieLet0_4QNode_Bool_emitted[0]))};
  assign lizzieLet0_4QNode_Bool_2_d = {lizzieLet0_4QNode_Bool_d[66:1],
                                       (lizzieLet0_4QNode_Bool_d[0] && (! lizzieLet0_4QNode_Bool_emitted[1]))};
  assign lizzieLet0_4QNode_Bool_3_d = {lizzieLet0_4QNode_Bool_d[66:1],
                                       (lizzieLet0_4QNode_Bool_d[0] && (! lizzieLet0_4QNode_Bool_emitted[2]))};
  assign lizzieLet0_4QNode_Bool_4_d = {lizzieLet0_4QNode_Bool_d[66:1],
                                       (lizzieLet0_4QNode_Bool_d[0] && (! lizzieLet0_4QNode_Bool_emitted[3]))};
  assign lizzieLet0_4QNode_Bool_5_d = {lizzieLet0_4QNode_Bool_d[66:1],
                                       (lizzieLet0_4QNode_Bool_d[0] && (! lizzieLet0_4QNode_Bool_emitted[4]))};
  assign lizzieLet0_4QNode_Bool_6_d = {lizzieLet0_4QNode_Bool_d[66:1],
                                       (lizzieLet0_4QNode_Bool_d[0] && (! lizzieLet0_4QNode_Bool_emitted[5]))};
  assign lizzieLet0_4QNode_Bool_7_d = {lizzieLet0_4QNode_Bool_d[66:1],
                                       (lizzieLet0_4QNode_Bool_d[0] && (! lizzieLet0_4QNode_Bool_emitted[6]))};
  assign lizzieLet0_4QNode_Bool_8_d = {lizzieLet0_4QNode_Bool_d[66:1],
                                       (lizzieLet0_4QNode_Bool_d[0] && (! lizzieLet0_4QNode_Bool_emitted[7]))};
  assign lizzieLet0_4QNode_Bool_9_d = {lizzieLet0_4QNode_Bool_d[66:1],
                                       (lizzieLet0_4QNode_Bool_d[0] && (! lizzieLet0_4QNode_Bool_emitted[8]))};
  assign lizzieLet0_4QNode_Bool_10_d = {lizzieLet0_4QNode_Bool_d[66:1],
                                        (lizzieLet0_4QNode_Bool_d[0] && (! lizzieLet0_4QNode_Bool_emitted[9]))};
  assign lizzieLet0_4QNode_Bool_done = (lizzieLet0_4QNode_Bool_emitted | ({lizzieLet0_4QNode_Bool_10_d[0],
                                                                           lizzieLet0_4QNode_Bool_9_d[0],
                                                                           lizzieLet0_4QNode_Bool_8_d[0],
                                                                           lizzieLet0_4QNode_Bool_7_d[0],
                                                                           lizzieLet0_4QNode_Bool_6_d[0],
                                                                           lizzieLet0_4QNode_Bool_5_d[0],
                                                                           lizzieLet0_4QNode_Bool_4_d[0],
                                                                           lizzieLet0_4QNode_Bool_3_d[0],
                                                                           lizzieLet0_4QNode_Bool_2_d[0],
                                                                           lizzieLet0_4QNode_Bool_1_d[0]} & {lizzieLet0_4QNode_Bool_10_r,
                                                                                                             lizzieLet0_4QNode_Bool_9_r,
                                                                                                             lizzieLet0_4QNode_Bool_8_r,
                                                                                                             lizzieLet0_4QNode_Bool_7_r,
                                                                                                             lizzieLet0_4QNode_Bool_6_r,
                                                                                                             lizzieLet0_4QNode_Bool_5_r,
                                                                                                             lizzieLet0_4QNode_Bool_4_r,
                                                                                                             lizzieLet0_4QNode_Bool_3_r,
                                                                                                             lizzieLet0_4QNode_Bool_2_r,
                                                                                                             lizzieLet0_4QNode_Bool_1_r}));
  assign lizzieLet0_4QNode_Bool_r = (& lizzieLet0_4QNode_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet0_4QNode_Bool_emitted <= 10'd0;
    else
      lizzieLet0_4QNode_Bool_emitted <= (lizzieLet0_4QNode_Bool_r ? 10'd0 :
                                         lizzieLet0_4QNode_Bool_done);
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_QTree_Bool) : (lizzieLet0_4QNode_Bool_10,QTree_Bool) (q4a8K_destruct,Pointer_QTree_Bool) > [(lizzieLet0_4QNode_Bool_10QNone_Bool,Pointer_QTree_Bool),
                                                                                                              (_165,Pointer_QTree_Bool),
                                                                                                              (lizzieLet0_4QNode_Bool_10QNode_Bool,Pointer_QTree_Bool),
                                                                                                              (_164,Pointer_QTree_Bool)] */
  logic [3:0] q4a8K_destruct_onehotd;
  always_comb
    if ((lizzieLet0_4QNode_Bool_10_d[0] && q4a8K_destruct_d[0]))
      unique case (lizzieLet0_4QNode_Bool_10_d[2:1])
        2'd0: q4a8K_destruct_onehotd = 4'd1;
        2'd1: q4a8K_destruct_onehotd = 4'd2;
        2'd2: q4a8K_destruct_onehotd = 4'd4;
        2'd3: q4a8K_destruct_onehotd = 4'd8;
        default: q4a8K_destruct_onehotd = 4'd0;
      endcase
    else q4a8K_destruct_onehotd = 4'd0;
  assign lizzieLet0_4QNode_Bool_10QNone_Bool_d = {q4a8K_destruct_d[16:1],
                                                  q4a8K_destruct_onehotd[0]};
  assign _165_d = {q4a8K_destruct_d[16:1],
                   q4a8K_destruct_onehotd[1]};
  assign lizzieLet0_4QNode_Bool_10QNode_Bool_d = {q4a8K_destruct_d[16:1],
                                                  q4a8K_destruct_onehotd[2]};
  assign _164_d = {q4a8K_destruct_d[16:1],
                   q4a8K_destruct_onehotd[3]};
  assign q4a8K_destruct_r = (| (q4a8K_destruct_onehotd & {_164_r,
                                                          lizzieLet0_4QNode_Bool_10QNode_Bool_r,
                                                          _165_r,
                                                          lizzieLet0_4QNode_Bool_10QNone_Bool_r}));
  assign lizzieLet0_4QNode_Bool_10_r = q4a8K_destruct_r;
  
  /* destruct (Ty QTree_Bool,
          Dcon QNode_Bool) : (lizzieLet0_4QNode_Bool_1QNode_Bool,QTree_Bool) > [(t1a8R_destruct,Pointer_QTree_Bool),
                                                                                (t2a8S_destruct,Pointer_QTree_Bool),
                                                                                (t3a8T_destruct,Pointer_QTree_Bool),
                                                                                (t4a8U_destruct,Pointer_QTree_Bool)] */
  logic [3:0] lizzieLet0_4QNode_Bool_1QNode_Bool_emitted;
  logic [3:0] lizzieLet0_4QNode_Bool_1QNode_Bool_done;
  assign t1a8R_destruct_d = {lizzieLet0_4QNode_Bool_1QNode_Bool_d[18:3],
                             (lizzieLet0_4QNode_Bool_1QNode_Bool_d[0] && (! lizzieLet0_4QNode_Bool_1QNode_Bool_emitted[0]))};
  assign t2a8S_destruct_d = {lizzieLet0_4QNode_Bool_1QNode_Bool_d[34:19],
                             (lizzieLet0_4QNode_Bool_1QNode_Bool_d[0] && (! lizzieLet0_4QNode_Bool_1QNode_Bool_emitted[1]))};
  assign t3a8T_destruct_d = {lizzieLet0_4QNode_Bool_1QNode_Bool_d[50:35],
                             (lizzieLet0_4QNode_Bool_1QNode_Bool_d[0] && (! lizzieLet0_4QNode_Bool_1QNode_Bool_emitted[2]))};
  assign t4a8U_destruct_d = {lizzieLet0_4QNode_Bool_1QNode_Bool_d[66:51],
                             (lizzieLet0_4QNode_Bool_1QNode_Bool_d[0] && (! lizzieLet0_4QNode_Bool_1QNode_Bool_emitted[3]))};
  assign lizzieLet0_4QNode_Bool_1QNode_Bool_done = (lizzieLet0_4QNode_Bool_1QNode_Bool_emitted | ({t4a8U_destruct_d[0],
                                                                                                   t3a8T_destruct_d[0],
                                                                                                   t2a8S_destruct_d[0],
                                                                                                   t1a8R_destruct_d[0]} & {t4a8U_destruct_r,
                                                                                                                           t3a8T_destruct_r,
                                                                                                                           t2a8S_destruct_r,
                                                                                                                           t1a8R_destruct_r}));
  assign lizzieLet0_4QNode_Bool_1QNode_Bool_r = (& lizzieLet0_4QNode_Bool_1QNode_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNode_Bool_1QNode_Bool_emitted <= 4'd0;
    else
      lizzieLet0_4QNode_Bool_1QNode_Bool_emitted <= (lizzieLet0_4QNode_Bool_1QNode_Bool_r ? 4'd0 :
                                                     lizzieLet0_4QNode_Bool_1QNode_Bool_done);
  
  /* demux (Ty QTree_Bool,
       Ty QTree_Bool) : (lizzieLet0_4QNode_Bool_2,QTree_Bool) (lizzieLet0_4QNode_Bool_1,QTree_Bool) > [(_163,QTree_Bool),
                                                                                                       (_162,QTree_Bool),
                                                                                                       (lizzieLet0_4QNode_Bool_1QNode_Bool,QTree_Bool),
                                                                                                       (_161,QTree_Bool)] */
  logic [3:0] lizzieLet0_4QNode_Bool_1_onehotd;
  always_comb
    if ((lizzieLet0_4QNode_Bool_2_d[0] && lizzieLet0_4QNode_Bool_1_d[0]))
      unique case (lizzieLet0_4QNode_Bool_2_d[2:1])
        2'd0: lizzieLet0_4QNode_Bool_1_onehotd = 4'd1;
        2'd1: lizzieLet0_4QNode_Bool_1_onehotd = 4'd2;
        2'd2: lizzieLet0_4QNode_Bool_1_onehotd = 4'd4;
        2'd3: lizzieLet0_4QNode_Bool_1_onehotd = 4'd8;
        default: lizzieLet0_4QNode_Bool_1_onehotd = 4'd0;
      endcase
    else lizzieLet0_4QNode_Bool_1_onehotd = 4'd0;
  assign _163_d = {lizzieLet0_4QNode_Bool_1_d[66:1],
                   lizzieLet0_4QNode_Bool_1_onehotd[0]};
  assign _162_d = {lizzieLet0_4QNode_Bool_1_d[66:1],
                   lizzieLet0_4QNode_Bool_1_onehotd[1]};
  assign lizzieLet0_4QNode_Bool_1QNode_Bool_d = {lizzieLet0_4QNode_Bool_1_d[66:1],
                                                 lizzieLet0_4QNode_Bool_1_onehotd[2]};
  assign _161_d = {lizzieLet0_4QNode_Bool_1_d[66:1],
                   lizzieLet0_4QNode_Bool_1_onehotd[3]};
  assign lizzieLet0_4QNode_Bool_1_r = (| (lizzieLet0_4QNode_Bool_1_onehotd & {_161_r,
                                                                              lizzieLet0_4QNode_Bool_1QNode_Bool_r,
                                                                              _162_r,
                                                                              _163_r}));
  assign lizzieLet0_4QNode_Bool_2_r = lizzieLet0_4QNode_Bool_1_r;
  
  /* demux (Ty QTree_Bool,
       Ty Go) : (lizzieLet0_4QNode_Bool_3,QTree_Bool) (lizzieLet0_3QNode_Bool,Go) > [(lizzieLet0_4QNode_Bool_3QNone_Bool,Go),
                                                                                     (lizzieLet0_4QNode_Bool_3QVal_Bool,Go),
                                                                                     (lizzieLet0_4QNode_Bool_3QNode_Bool,Go),
                                                                                     (lizzieLet0_4QNode_Bool_3QError_Bool,Go)] */
  logic [3:0] lizzieLet0_3QNode_Bool_onehotd;
  always_comb
    if ((lizzieLet0_4QNode_Bool_3_d[0] && lizzieLet0_3QNode_Bool_d[0]))
      unique case (lizzieLet0_4QNode_Bool_3_d[2:1])
        2'd0: lizzieLet0_3QNode_Bool_onehotd = 4'd1;
        2'd1: lizzieLet0_3QNode_Bool_onehotd = 4'd2;
        2'd2: lizzieLet0_3QNode_Bool_onehotd = 4'd4;
        2'd3: lizzieLet0_3QNode_Bool_onehotd = 4'd8;
        default: lizzieLet0_3QNode_Bool_onehotd = 4'd0;
      endcase
    else lizzieLet0_3QNode_Bool_onehotd = 4'd0;
  assign lizzieLet0_4QNode_Bool_3QNone_Bool_d = lizzieLet0_3QNode_Bool_onehotd[0];
  assign lizzieLet0_4QNode_Bool_3QVal_Bool_d = lizzieLet0_3QNode_Bool_onehotd[1];
  assign lizzieLet0_4QNode_Bool_3QNode_Bool_d = lizzieLet0_3QNode_Bool_onehotd[2];
  assign lizzieLet0_4QNode_Bool_3QError_Bool_d = lizzieLet0_3QNode_Bool_onehotd[3];
  assign lizzieLet0_3QNode_Bool_r = (| (lizzieLet0_3QNode_Bool_onehotd & {lizzieLet0_4QNode_Bool_3QError_Bool_r,
                                                                          lizzieLet0_4QNode_Bool_3QNode_Bool_r,
                                                                          lizzieLet0_4QNode_Bool_3QVal_Bool_r,
                                                                          lizzieLet0_4QNode_Bool_3QNone_Bool_r}));
  assign lizzieLet0_4QNode_Bool_3_r = lizzieLet0_3QNode_Bool_r;
  
  /* fork (Ty Go) : (lizzieLet0_4QNode_Bool_3QError_Bool,Go) > [(lizzieLet0_4QNode_Bool_3QError_Bool_1,Go),
                                                           (lizzieLet0_4QNode_Bool_3QError_Bool_2,Go)] */
  logic [1:0] lizzieLet0_4QNode_Bool_3QError_Bool_emitted;
  logic [1:0] lizzieLet0_4QNode_Bool_3QError_Bool_done;
  assign lizzieLet0_4QNode_Bool_3QError_Bool_1_d = (lizzieLet0_4QNode_Bool_3QError_Bool_d[0] && (! lizzieLet0_4QNode_Bool_3QError_Bool_emitted[0]));
  assign lizzieLet0_4QNode_Bool_3QError_Bool_2_d = (lizzieLet0_4QNode_Bool_3QError_Bool_d[0] && (! lizzieLet0_4QNode_Bool_3QError_Bool_emitted[1]));
  assign lizzieLet0_4QNode_Bool_3QError_Bool_done = (lizzieLet0_4QNode_Bool_3QError_Bool_emitted | ({lizzieLet0_4QNode_Bool_3QError_Bool_2_d[0],
                                                                                                     lizzieLet0_4QNode_Bool_3QError_Bool_1_d[0]} & {lizzieLet0_4QNode_Bool_3QError_Bool_2_r,
                                                                                                                                                    lizzieLet0_4QNode_Bool_3QError_Bool_1_r}));
  assign lizzieLet0_4QNode_Bool_3QError_Bool_r = (& lizzieLet0_4QNode_Bool_3QError_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNode_Bool_3QError_Bool_emitted <= 2'd0;
    else
      lizzieLet0_4QNode_Bool_3QError_Bool_emitted <= (lizzieLet0_4QNode_Bool_3QError_Bool_r ? 2'd0 :
                                                      lizzieLet0_4QNode_Bool_3QError_Bool_done);
  
  /* dcon (Ty QTree_Bool,
      Dcon QError_Bool) : [(lizzieLet0_4QNode_Bool_3QError_Bool_1,Go)] > (lizzieLet0_4QNode_Bool_3QError_Bool_1QError_Bool,QTree_Bool) */
  assign lizzieLet0_4QNode_Bool_3QError_Bool_1QError_Bool_d = QError_Bool_dc((& {lizzieLet0_4QNode_Bool_3QError_Bool_1_d[0]}), lizzieLet0_4QNode_Bool_3QError_Bool_1_d);
  assign {lizzieLet0_4QNode_Bool_3QError_Bool_1_r} = {1 {(lizzieLet0_4QNode_Bool_3QError_Bool_1QError_Bool_r && lizzieLet0_4QNode_Bool_3QError_Bool_1QError_Bool_d[0])}};
  
  /* buf (Ty QTree_Bool) : (lizzieLet0_4QNode_Bool_3QError_Bool_1QError_Bool,QTree_Bool) > (lizzieLet43_1_argbuf,QTree_Bool) */
  QTree_Bool_t lizzieLet0_4QNode_Bool_3QError_Bool_1QError_Bool_bufchan_d;
  logic lizzieLet0_4QNode_Bool_3QError_Bool_1QError_Bool_bufchan_r;
  assign lizzieLet0_4QNode_Bool_3QError_Bool_1QError_Bool_r = ((! lizzieLet0_4QNode_Bool_3QError_Bool_1QError_Bool_bufchan_d[0]) || lizzieLet0_4QNode_Bool_3QError_Bool_1QError_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNode_Bool_3QError_Bool_1QError_Bool_bufchan_d <= {66'd0,
                                                                     1'd0};
    else
      if (lizzieLet0_4QNode_Bool_3QError_Bool_1QError_Bool_r)
        lizzieLet0_4QNode_Bool_3QError_Bool_1QError_Bool_bufchan_d <= lizzieLet0_4QNode_Bool_3QError_Bool_1QError_Bool_d;
  QTree_Bool_t lizzieLet0_4QNode_Bool_3QError_Bool_1QError_Bool_bufchan_buf;
  assign lizzieLet0_4QNode_Bool_3QError_Bool_1QError_Bool_bufchan_r = (! lizzieLet0_4QNode_Bool_3QError_Bool_1QError_Bool_bufchan_buf[0]);
  assign lizzieLet43_1_argbuf_d = (lizzieLet0_4QNode_Bool_3QError_Bool_1QError_Bool_bufchan_buf[0] ? lizzieLet0_4QNode_Bool_3QError_Bool_1QError_Bool_bufchan_buf :
                                   lizzieLet0_4QNode_Bool_3QError_Bool_1QError_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNode_Bool_3QError_Bool_1QError_Bool_bufchan_buf <= {66'd0,
                                                                       1'd0};
    else
      if ((lizzieLet43_1_argbuf_r && lizzieLet0_4QNode_Bool_3QError_Bool_1QError_Bool_bufchan_buf[0]))
        lizzieLet0_4QNode_Bool_3QError_Bool_1QError_Bool_bufchan_buf <= {66'd0,
                                                                         1'd0};
      else if (((! lizzieLet43_1_argbuf_r) && (! lizzieLet0_4QNode_Bool_3QError_Bool_1QError_Bool_bufchan_buf[0])))
        lizzieLet0_4QNode_Bool_3QError_Bool_1QError_Bool_bufchan_buf <= lizzieLet0_4QNode_Bool_3QError_Bool_1QError_Bool_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet0_4QNode_Bool_3QError_Bool_2,Go) > (lizzieLet0_4QNode_Bool_3QError_Bool_2_argbuf,Go) */
  Go_t lizzieLet0_4QNode_Bool_3QError_Bool_2_bufchan_d;
  logic lizzieLet0_4QNode_Bool_3QError_Bool_2_bufchan_r;
  assign lizzieLet0_4QNode_Bool_3QError_Bool_2_r = ((! lizzieLet0_4QNode_Bool_3QError_Bool_2_bufchan_d[0]) || lizzieLet0_4QNode_Bool_3QError_Bool_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNode_Bool_3QError_Bool_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet0_4QNode_Bool_3QError_Bool_2_r)
        lizzieLet0_4QNode_Bool_3QError_Bool_2_bufchan_d <= lizzieLet0_4QNode_Bool_3QError_Bool_2_d;
  Go_t lizzieLet0_4QNode_Bool_3QError_Bool_2_bufchan_buf;
  assign lizzieLet0_4QNode_Bool_3QError_Bool_2_bufchan_r = (! lizzieLet0_4QNode_Bool_3QError_Bool_2_bufchan_buf[0]);
  assign lizzieLet0_4QNode_Bool_3QError_Bool_2_argbuf_d = (lizzieLet0_4QNode_Bool_3QError_Bool_2_bufchan_buf[0] ? lizzieLet0_4QNode_Bool_3QError_Bool_2_bufchan_buf :
                                                           lizzieLet0_4QNode_Bool_3QError_Bool_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNode_Bool_3QError_Bool_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet0_4QNode_Bool_3QError_Bool_2_argbuf_r && lizzieLet0_4QNode_Bool_3QError_Bool_2_bufchan_buf[0]))
        lizzieLet0_4QNode_Bool_3QError_Bool_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet0_4QNode_Bool_3QError_Bool_2_argbuf_r) && (! lizzieLet0_4QNode_Bool_3QError_Bool_2_bufchan_buf[0])))
        lizzieLet0_4QNode_Bool_3QError_Bool_2_bufchan_buf <= lizzieLet0_4QNode_Bool_3QError_Bool_2_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet0_4QNode_Bool_3QVal_Bool,Go) > [(lizzieLet0_4QNode_Bool_3QVal_Bool_1,Go),
                                                         (lizzieLet0_4QNode_Bool_3QVal_Bool_2,Go)] */
  logic [1:0] lizzieLet0_4QNode_Bool_3QVal_Bool_emitted;
  logic [1:0] lizzieLet0_4QNode_Bool_3QVal_Bool_done;
  assign lizzieLet0_4QNode_Bool_3QVal_Bool_1_d = (lizzieLet0_4QNode_Bool_3QVal_Bool_d[0] && (! lizzieLet0_4QNode_Bool_3QVal_Bool_emitted[0]));
  assign lizzieLet0_4QNode_Bool_3QVal_Bool_2_d = (lizzieLet0_4QNode_Bool_3QVal_Bool_d[0] && (! lizzieLet0_4QNode_Bool_3QVal_Bool_emitted[1]));
  assign lizzieLet0_4QNode_Bool_3QVal_Bool_done = (lizzieLet0_4QNode_Bool_3QVal_Bool_emitted | ({lizzieLet0_4QNode_Bool_3QVal_Bool_2_d[0],
                                                                                                 lizzieLet0_4QNode_Bool_3QVal_Bool_1_d[0]} & {lizzieLet0_4QNode_Bool_3QVal_Bool_2_r,
                                                                                                                                              lizzieLet0_4QNode_Bool_3QVal_Bool_1_r}));
  assign lizzieLet0_4QNode_Bool_3QVal_Bool_r = (& lizzieLet0_4QNode_Bool_3QVal_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNode_Bool_3QVal_Bool_emitted <= 2'd0;
    else
      lizzieLet0_4QNode_Bool_3QVal_Bool_emitted <= (lizzieLet0_4QNode_Bool_3QVal_Bool_r ? 2'd0 :
                                                    lizzieLet0_4QNode_Bool_3QVal_Bool_done);
  
  /* dcon (Ty QTree_Bool,
      Dcon QError_Bool) : [(lizzieLet0_4QNode_Bool_3QVal_Bool_1,Go)] > (lizzieLet0_4QNode_Bool_3QVal_Bool_1QError_Bool,QTree_Bool) */
  assign lizzieLet0_4QNode_Bool_3QVal_Bool_1QError_Bool_d = QError_Bool_dc((& {lizzieLet0_4QNode_Bool_3QVal_Bool_1_d[0]}), lizzieLet0_4QNode_Bool_3QVal_Bool_1_d);
  assign {lizzieLet0_4QNode_Bool_3QVal_Bool_1_r} = {1 {(lizzieLet0_4QNode_Bool_3QVal_Bool_1QError_Bool_r && lizzieLet0_4QNode_Bool_3QVal_Bool_1QError_Bool_d[0])}};
  
  /* buf (Ty QTree_Bool) : (lizzieLet0_4QNode_Bool_3QVal_Bool_1QError_Bool,QTree_Bool) > (lizzieLet37_1_argbuf,QTree_Bool) */
  QTree_Bool_t lizzieLet0_4QNode_Bool_3QVal_Bool_1QError_Bool_bufchan_d;
  logic lizzieLet0_4QNode_Bool_3QVal_Bool_1QError_Bool_bufchan_r;
  assign lizzieLet0_4QNode_Bool_3QVal_Bool_1QError_Bool_r = ((! lizzieLet0_4QNode_Bool_3QVal_Bool_1QError_Bool_bufchan_d[0]) || lizzieLet0_4QNode_Bool_3QVal_Bool_1QError_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNode_Bool_3QVal_Bool_1QError_Bool_bufchan_d <= {66'd0,
                                                                   1'd0};
    else
      if (lizzieLet0_4QNode_Bool_3QVal_Bool_1QError_Bool_r)
        lizzieLet0_4QNode_Bool_3QVal_Bool_1QError_Bool_bufchan_d <= lizzieLet0_4QNode_Bool_3QVal_Bool_1QError_Bool_d;
  QTree_Bool_t lizzieLet0_4QNode_Bool_3QVal_Bool_1QError_Bool_bufchan_buf;
  assign lizzieLet0_4QNode_Bool_3QVal_Bool_1QError_Bool_bufchan_r = (! lizzieLet0_4QNode_Bool_3QVal_Bool_1QError_Bool_bufchan_buf[0]);
  assign lizzieLet37_1_argbuf_d = (lizzieLet0_4QNode_Bool_3QVal_Bool_1QError_Bool_bufchan_buf[0] ? lizzieLet0_4QNode_Bool_3QVal_Bool_1QError_Bool_bufchan_buf :
                                   lizzieLet0_4QNode_Bool_3QVal_Bool_1QError_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNode_Bool_3QVal_Bool_1QError_Bool_bufchan_buf <= {66'd0,
                                                                     1'd0};
    else
      if ((lizzieLet37_1_argbuf_r && lizzieLet0_4QNode_Bool_3QVal_Bool_1QError_Bool_bufchan_buf[0]))
        lizzieLet0_4QNode_Bool_3QVal_Bool_1QError_Bool_bufchan_buf <= {66'd0,
                                                                       1'd0};
      else if (((! lizzieLet37_1_argbuf_r) && (! lizzieLet0_4QNode_Bool_3QVal_Bool_1QError_Bool_bufchan_buf[0])))
        lizzieLet0_4QNode_Bool_3QVal_Bool_1QError_Bool_bufchan_buf <= lizzieLet0_4QNode_Bool_3QVal_Bool_1QError_Bool_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet0_4QNode_Bool_3QVal_Bool_2,Go) > (lizzieLet0_4QNode_Bool_3QVal_Bool_2_argbuf,Go) */
  Go_t lizzieLet0_4QNode_Bool_3QVal_Bool_2_bufchan_d;
  logic lizzieLet0_4QNode_Bool_3QVal_Bool_2_bufchan_r;
  assign lizzieLet0_4QNode_Bool_3QVal_Bool_2_r = ((! lizzieLet0_4QNode_Bool_3QVal_Bool_2_bufchan_d[0]) || lizzieLet0_4QNode_Bool_3QVal_Bool_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNode_Bool_3QVal_Bool_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet0_4QNode_Bool_3QVal_Bool_2_r)
        lizzieLet0_4QNode_Bool_3QVal_Bool_2_bufchan_d <= lizzieLet0_4QNode_Bool_3QVal_Bool_2_d;
  Go_t lizzieLet0_4QNode_Bool_3QVal_Bool_2_bufchan_buf;
  assign lizzieLet0_4QNode_Bool_3QVal_Bool_2_bufchan_r = (! lizzieLet0_4QNode_Bool_3QVal_Bool_2_bufchan_buf[0]);
  assign lizzieLet0_4QNode_Bool_3QVal_Bool_2_argbuf_d = (lizzieLet0_4QNode_Bool_3QVal_Bool_2_bufchan_buf[0] ? lizzieLet0_4QNode_Bool_3QVal_Bool_2_bufchan_buf :
                                                         lizzieLet0_4QNode_Bool_3QVal_Bool_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNode_Bool_3QVal_Bool_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet0_4QNode_Bool_3QVal_Bool_2_argbuf_r && lizzieLet0_4QNode_Bool_3QVal_Bool_2_bufchan_buf[0]))
        lizzieLet0_4QNode_Bool_3QVal_Bool_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet0_4QNode_Bool_3QVal_Bool_2_argbuf_r) && (! lizzieLet0_4QNode_Bool_3QVal_Bool_2_bufchan_buf[0])))
        lizzieLet0_4QNode_Bool_3QVal_Bool_2_bufchan_buf <= lizzieLet0_4QNode_Bool_3QVal_Bool_2_bufchan_d;
  
  /* demux (Ty QTree_Bool,
       Ty QTree_Bool) : (lizzieLet0_4QNode_Bool_4,QTree_Bool) (lizzieLet0_5QNode_Bool,QTree_Bool) > [(lizzieLet0_4QNode_Bool_4QNone_Bool,QTree_Bool),
                                                                                                     (_160,QTree_Bool),
                                                                                                     (lizzieLet0_4QNode_Bool_4QNode_Bool,QTree_Bool),
                                                                                                     (_159,QTree_Bool)] */
  logic [3:0] lizzieLet0_5QNode_Bool_onehotd;
  always_comb
    if ((lizzieLet0_4QNode_Bool_4_d[0] && lizzieLet0_5QNode_Bool_d[0]))
      unique case (lizzieLet0_4QNode_Bool_4_d[2:1])
        2'd0: lizzieLet0_5QNode_Bool_onehotd = 4'd1;
        2'd1: lizzieLet0_5QNode_Bool_onehotd = 4'd2;
        2'd2: lizzieLet0_5QNode_Bool_onehotd = 4'd4;
        2'd3: lizzieLet0_5QNode_Bool_onehotd = 4'd8;
        default: lizzieLet0_5QNode_Bool_onehotd = 4'd0;
      endcase
    else lizzieLet0_5QNode_Bool_onehotd = 4'd0;
  assign lizzieLet0_4QNode_Bool_4QNone_Bool_d = {lizzieLet0_5QNode_Bool_d[66:1],
                                                 lizzieLet0_5QNode_Bool_onehotd[0]};
  assign _160_d = {lizzieLet0_5QNode_Bool_d[66:1],
                   lizzieLet0_5QNode_Bool_onehotd[1]};
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_d = {lizzieLet0_5QNode_Bool_d[66:1],
                                                 lizzieLet0_5QNode_Bool_onehotd[2]};
  assign _159_d = {lizzieLet0_5QNode_Bool_d[66:1],
                   lizzieLet0_5QNode_Bool_onehotd[3]};
  assign lizzieLet0_5QNode_Bool_r = (| (lizzieLet0_5QNode_Bool_onehotd & {_159_r,
                                                                          lizzieLet0_4QNode_Bool_4QNode_Bool_r,
                                                                          _160_r,
                                                                          lizzieLet0_4QNode_Bool_4QNone_Bool_r}));
  assign lizzieLet0_4QNode_Bool_4_r = lizzieLet0_5QNode_Bool_r;
  
  /* fork (Ty QTree_Bool) : (lizzieLet0_4QNode_Bool_4QNode_Bool,QTree_Bool) > [(lizzieLet0_4QNode_Bool_4QNode_Bool_1,QTree_Bool),
                                                                          (lizzieLet0_4QNode_Bool_4QNode_Bool_2,QTree_Bool),
                                                                          (lizzieLet0_4QNode_Bool_4QNode_Bool_3,QTree_Bool),
                                                                          (lizzieLet0_4QNode_Bool_4QNode_Bool_4,QTree_Bool),
                                                                          (lizzieLet0_4QNode_Bool_4QNode_Bool_5,QTree_Bool),
                                                                          (lizzieLet0_4QNode_Bool_4QNode_Bool_6,QTree_Bool),
                                                                          (lizzieLet0_4QNode_Bool_4QNode_Bool_7,QTree_Bool),
                                                                          (lizzieLet0_4QNode_Bool_4QNode_Bool_8,QTree_Bool),
                                                                          (lizzieLet0_4QNode_Bool_4QNode_Bool_9,QTree_Bool),
                                                                          (lizzieLet0_4QNode_Bool_4QNode_Bool_10,QTree_Bool),
                                                                          (lizzieLet0_4QNode_Bool_4QNode_Bool_11,QTree_Bool),
                                                                          (lizzieLet0_4QNode_Bool_4QNode_Bool_12,QTree_Bool)] */
  logic [11:0] lizzieLet0_4QNode_Bool_4QNode_Bool_emitted;
  logic [11:0] lizzieLet0_4QNode_Bool_4QNode_Bool_done;
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_1_d = {lizzieLet0_4QNode_Bool_4QNode_Bool_d[66:1],
                                                   (lizzieLet0_4QNode_Bool_4QNode_Bool_d[0] && (! lizzieLet0_4QNode_Bool_4QNode_Bool_emitted[0]))};
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_2_d = {lizzieLet0_4QNode_Bool_4QNode_Bool_d[66:1],
                                                   (lizzieLet0_4QNode_Bool_4QNode_Bool_d[0] && (! lizzieLet0_4QNode_Bool_4QNode_Bool_emitted[1]))};
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_3_d = {lizzieLet0_4QNode_Bool_4QNode_Bool_d[66:1],
                                                   (lizzieLet0_4QNode_Bool_4QNode_Bool_d[0] && (! lizzieLet0_4QNode_Bool_4QNode_Bool_emitted[2]))};
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_4_d = {lizzieLet0_4QNode_Bool_4QNode_Bool_d[66:1],
                                                   (lizzieLet0_4QNode_Bool_4QNode_Bool_d[0] && (! lizzieLet0_4QNode_Bool_4QNode_Bool_emitted[3]))};
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_5_d = {lizzieLet0_4QNode_Bool_4QNode_Bool_d[66:1],
                                                   (lizzieLet0_4QNode_Bool_4QNode_Bool_d[0] && (! lizzieLet0_4QNode_Bool_4QNode_Bool_emitted[4]))};
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_6_d = {lizzieLet0_4QNode_Bool_4QNode_Bool_d[66:1],
                                                   (lizzieLet0_4QNode_Bool_4QNode_Bool_d[0] && (! lizzieLet0_4QNode_Bool_4QNode_Bool_emitted[5]))};
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_7_d = {lizzieLet0_4QNode_Bool_4QNode_Bool_d[66:1],
                                                   (lizzieLet0_4QNode_Bool_4QNode_Bool_d[0] && (! lizzieLet0_4QNode_Bool_4QNode_Bool_emitted[6]))};
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_8_d = {lizzieLet0_4QNode_Bool_4QNode_Bool_d[66:1],
                                                   (lizzieLet0_4QNode_Bool_4QNode_Bool_d[0] && (! lizzieLet0_4QNode_Bool_4QNode_Bool_emitted[7]))};
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_9_d = {lizzieLet0_4QNode_Bool_4QNode_Bool_d[66:1],
                                                   (lizzieLet0_4QNode_Bool_4QNode_Bool_d[0] && (! lizzieLet0_4QNode_Bool_4QNode_Bool_emitted[8]))};
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_10_d = {lizzieLet0_4QNode_Bool_4QNode_Bool_d[66:1],
                                                    (lizzieLet0_4QNode_Bool_4QNode_Bool_d[0] && (! lizzieLet0_4QNode_Bool_4QNode_Bool_emitted[9]))};
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_11_d = {lizzieLet0_4QNode_Bool_4QNode_Bool_d[66:1],
                                                    (lizzieLet0_4QNode_Bool_4QNode_Bool_d[0] && (! lizzieLet0_4QNode_Bool_4QNode_Bool_emitted[10]))};
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_12_d = {lizzieLet0_4QNode_Bool_4QNode_Bool_d[66:1],
                                                    (lizzieLet0_4QNode_Bool_4QNode_Bool_d[0] && (! lizzieLet0_4QNode_Bool_4QNode_Bool_emitted[11]))};
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_done = (lizzieLet0_4QNode_Bool_4QNode_Bool_emitted | ({lizzieLet0_4QNode_Bool_4QNode_Bool_12_d[0],
                                                                                                   lizzieLet0_4QNode_Bool_4QNode_Bool_11_d[0],
                                                                                                   lizzieLet0_4QNode_Bool_4QNode_Bool_10_d[0],
                                                                                                   lizzieLet0_4QNode_Bool_4QNode_Bool_9_d[0],
                                                                                                   lizzieLet0_4QNode_Bool_4QNode_Bool_8_d[0],
                                                                                                   lizzieLet0_4QNode_Bool_4QNode_Bool_7_d[0],
                                                                                                   lizzieLet0_4QNode_Bool_4QNode_Bool_6_d[0],
                                                                                                   lizzieLet0_4QNode_Bool_4QNode_Bool_5_d[0],
                                                                                                   lizzieLet0_4QNode_Bool_4QNode_Bool_4_d[0],
                                                                                                   lizzieLet0_4QNode_Bool_4QNode_Bool_3_d[0],
                                                                                                   lizzieLet0_4QNode_Bool_4QNode_Bool_2_d[0],
                                                                                                   lizzieLet0_4QNode_Bool_4QNode_Bool_1_d[0]} & {lizzieLet0_4QNode_Bool_4QNode_Bool_12_r,
                                                                                                                                                 lizzieLet0_4QNode_Bool_4QNode_Bool_11_r,
                                                                                                                                                 lizzieLet0_4QNode_Bool_4QNode_Bool_10_r,
                                                                                                                                                 lizzieLet0_4QNode_Bool_4QNode_Bool_9_r,
                                                                                                                                                 lizzieLet0_4QNode_Bool_4QNode_Bool_8_r,
                                                                                                                                                 lizzieLet0_4QNode_Bool_4QNode_Bool_7_r,
                                                                                                                                                 lizzieLet0_4QNode_Bool_4QNode_Bool_6_r,
                                                                                                                                                 lizzieLet0_4QNode_Bool_4QNode_Bool_5_r,
                                                                                                                                                 lizzieLet0_4QNode_Bool_4QNode_Bool_4_r,
                                                                                                                                                 lizzieLet0_4QNode_Bool_4QNode_Bool_3_r,
                                                                                                                                                 lizzieLet0_4QNode_Bool_4QNode_Bool_2_r,
                                                                                                                                                 lizzieLet0_4QNode_Bool_4QNode_Bool_1_r}));
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_r = (& lizzieLet0_4QNode_Bool_4QNode_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNode_Bool_4QNode_Bool_emitted <= 12'd0;
    else
      lizzieLet0_4QNode_Bool_4QNode_Bool_emitted <= (lizzieLet0_4QNode_Bool_4QNode_Bool_r ? 12'd0 :
                                                     lizzieLet0_4QNode_Bool_4QNode_Bool_done);
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_QTree_Bool) : (lizzieLet0_4QNode_Bool_4QNode_Bool_10,QTree_Bool) (t2a8S_destruct,Pointer_QTree_Bool) > [(lizzieLet0_4QNode_Bool_4QNode_Bool_10QNone_Bool,Pointer_QTree_Bool),
                                                                                                                          (_158,Pointer_QTree_Bool),
                                                                                                                          (lizzieLet0_4QNode_Bool_4QNode_Bool_10QNode_Bool,Pointer_QTree_Bool),
                                                                                                                          (_157,Pointer_QTree_Bool)] */
  logic [3:0] t2a8S_destruct_onehotd;
  always_comb
    if ((lizzieLet0_4QNode_Bool_4QNode_Bool_10_d[0] && t2a8S_destruct_d[0]))
      unique case (lizzieLet0_4QNode_Bool_4QNode_Bool_10_d[2:1])
        2'd0: t2a8S_destruct_onehotd = 4'd1;
        2'd1: t2a8S_destruct_onehotd = 4'd2;
        2'd2: t2a8S_destruct_onehotd = 4'd4;
        2'd3: t2a8S_destruct_onehotd = 4'd8;
        default: t2a8S_destruct_onehotd = 4'd0;
      endcase
    else t2a8S_destruct_onehotd = 4'd0;
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_10QNone_Bool_d = {t2a8S_destruct_d[16:1],
                                                              t2a8S_destruct_onehotd[0]};
  assign _158_d = {t2a8S_destruct_d[16:1],
                   t2a8S_destruct_onehotd[1]};
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_10QNode_Bool_d = {t2a8S_destruct_d[16:1],
                                                              t2a8S_destruct_onehotd[2]};
  assign _157_d = {t2a8S_destruct_d[16:1],
                   t2a8S_destruct_onehotd[3]};
  assign t2a8S_destruct_r = (| (t2a8S_destruct_onehotd & {_157_r,
                                                          lizzieLet0_4QNode_Bool_4QNode_Bool_10QNode_Bool_r,
                                                          _158_r,
                                                          lizzieLet0_4QNode_Bool_4QNode_Bool_10QNone_Bool_r}));
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_10_r = t2a8S_destruct_r;
  
  /* buf (Ty Pointer_QTree_Bool) : (lizzieLet0_4QNode_Bool_4QNode_Bool_10QNone_Bool,Pointer_QTree_Bool) > (lizzieLet0_4QNode_Bool_4QNode_Bool_10QNone_Bool_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t lizzieLet0_4QNode_Bool_4QNode_Bool_10QNone_Bool_bufchan_d;
  logic lizzieLet0_4QNode_Bool_4QNode_Bool_10QNone_Bool_bufchan_r;
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_10QNone_Bool_r = ((! lizzieLet0_4QNode_Bool_4QNode_Bool_10QNone_Bool_bufchan_d[0]) || lizzieLet0_4QNode_Bool_4QNode_Bool_10QNone_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNode_Bool_4QNode_Bool_10QNone_Bool_bufchan_d <= {16'd0,
                                                                    1'd0};
    else
      if (lizzieLet0_4QNode_Bool_4QNode_Bool_10QNone_Bool_r)
        lizzieLet0_4QNode_Bool_4QNode_Bool_10QNone_Bool_bufchan_d <= lizzieLet0_4QNode_Bool_4QNode_Bool_10QNone_Bool_d;
  Pointer_QTree_Bool_t lizzieLet0_4QNode_Bool_4QNode_Bool_10QNone_Bool_bufchan_buf;
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_10QNone_Bool_bufchan_r = (! lizzieLet0_4QNode_Bool_4QNode_Bool_10QNone_Bool_bufchan_buf[0]);
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_10QNone_Bool_1_argbuf_d = (lizzieLet0_4QNode_Bool_4QNode_Bool_10QNone_Bool_bufchan_buf[0] ? lizzieLet0_4QNode_Bool_4QNode_Bool_10QNone_Bool_bufchan_buf :
                                                                       lizzieLet0_4QNode_Bool_4QNode_Bool_10QNone_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNode_Bool_4QNode_Bool_10QNone_Bool_bufchan_buf <= {16'd0,
                                                                      1'd0};
    else
      if ((lizzieLet0_4QNode_Bool_4QNode_Bool_10QNone_Bool_1_argbuf_r && lizzieLet0_4QNode_Bool_4QNode_Bool_10QNone_Bool_bufchan_buf[0]))
        lizzieLet0_4QNode_Bool_4QNode_Bool_10QNone_Bool_bufchan_buf <= {16'd0,
                                                                        1'd0};
      else if (((! lizzieLet0_4QNode_Bool_4QNode_Bool_10QNone_Bool_1_argbuf_r) && (! lizzieLet0_4QNode_Bool_4QNode_Bool_10QNone_Bool_bufchan_buf[0])))
        lizzieLet0_4QNode_Bool_4QNode_Bool_10QNone_Bool_bufchan_buf <= lizzieLet0_4QNode_Bool_4QNode_Bool_10QNone_Bool_bufchan_d;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_QTree_Bool) : (lizzieLet0_4QNode_Bool_4QNode_Bool_11,QTree_Bool) (t3a8T_destruct,Pointer_QTree_Bool) > [(lizzieLet0_4QNode_Bool_4QNode_Bool_11QNone_Bool,Pointer_QTree_Bool),
                                                                                                                          (_156,Pointer_QTree_Bool),
                                                                                                                          (lizzieLet0_4QNode_Bool_4QNode_Bool_11QNode_Bool,Pointer_QTree_Bool),
                                                                                                                          (_155,Pointer_QTree_Bool)] */
  logic [3:0] t3a8T_destruct_onehotd;
  always_comb
    if ((lizzieLet0_4QNode_Bool_4QNode_Bool_11_d[0] && t3a8T_destruct_d[0]))
      unique case (lizzieLet0_4QNode_Bool_4QNode_Bool_11_d[2:1])
        2'd0: t3a8T_destruct_onehotd = 4'd1;
        2'd1: t3a8T_destruct_onehotd = 4'd2;
        2'd2: t3a8T_destruct_onehotd = 4'd4;
        2'd3: t3a8T_destruct_onehotd = 4'd8;
        default: t3a8T_destruct_onehotd = 4'd0;
      endcase
    else t3a8T_destruct_onehotd = 4'd0;
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_11QNone_Bool_d = {t3a8T_destruct_d[16:1],
                                                              t3a8T_destruct_onehotd[0]};
  assign _156_d = {t3a8T_destruct_d[16:1],
                   t3a8T_destruct_onehotd[1]};
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_11QNode_Bool_d = {t3a8T_destruct_d[16:1],
                                                              t3a8T_destruct_onehotd[2]};
  assign _155_d = {t3a8T_destruct_d[16:1],
                   t3a8T_destruct_onehotd[3]};
  assign t3a8T_destruct_r = (| (t3a8T_destruct_onehotd & {_155_r,
                                                          lizzieLet0_4QNode_Bool_4QNode_Bool_11QNode_Bool_r,
                                                          _156_r,
                                                          lizzieLet0_4QNode_Bool_4QNode_Bool_11QNone_Bool_r}));
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_11_r = t3a8T_destruct_r;
  
  /* buf (Ty Pointer_QTree_Bool) : (lizzieLet0_4QNode_Bool_4QNode_Bool_11QNone_Bool,Pointer_QTree_Bool) > (lizzieLet0_4QNode_Bool_4QNode_Bool_11QNone_Bool_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t lizzieLet0_4QNode_Bool_4QNode_Bool_11QNone_Bool_bufchan_d;
  logic lizzieLet0_4QNode_Bool_4QNode_Bool_11QNone_Bool_bufchan_r;
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_11QNone_Bool_r = ((! lizzieLet0_4QNode_Bool_4QNode_Bool_11QNone_Bool_bufchan_d[0]) || lizzieLet0_4QNode_Bool_4QNode_Bool_11QNone_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNode_Bool_4QNode_Bool_11QNone_Bool_bufchan_d <= {16'd0,
                                                                    1'd0};
    else
      if (lizzieLet0_4QNode_Bool_4QNode_Bool_11QNone_Bool_r)
        lizzieLet0_4QNode_Bool_4QNode_Bool_11QNone_Bool_bufchan_d <= lizzieLet0_4QNode_Bool_4QNode_Bool_11QNone_Bool_d;
  Pointer_QTree_Bool_t lizzieLet0_4QNode_Bool_4QNode_Bool_11QNone_Bool_bufchan_buf;
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_11QNone_Bool_bufchan_r = (! lizzieLet0_4QNode_Bool_4QNode_Bool_11QNone_Bool_bufchan_buf[0]);
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_11QNone_Bool_1_argbuf_d = (lizzieLet0_4QNode_Bool_4QNode_Bool_11QNone_Bool_bufchan_buf[0] ? lizzieLet0_4QNode_Bool_4QNode_Bool_11QNone_Bool_bufchan_buf :
                                                                       lizzieLet0_4QNode_Bool_4QNode_Bool_11QNone_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNode_Bool_4QNode_Bool_11QNone_Bool_bufchan_buf <= {16'd0,
                                                                      1'd0};
    else
      if ((lizzieLet0_4QNode_Bool_4QNode_Bool_11QNone_Bool_1_argbuf_r && lizzieLet0_4QNode_Bool_4QNode_Bool_11QNone_Bool_bufchan_buf[0]))
        lizzieLet0_4QNode_Bool_4QNode_Bool_11QNone_Bool_bufchan_buf <= {16'd0,
                                                                        1'd0};
      else if (((! lizzieLet0_4QNode_Bool_4QNode_Bool_11QNone_Bool_1_argbuf_r) && (! lizzieLet0_4QNode_Bool_4QNode_Bool_11QNone_Bool_bufchan_buf[0])))
        lizzieLet0_4QNode_Bool_4QNode_Bool_11QNone_Bool_bufchan_buf <= lizzieLet0_4QNode_Bool_4QNode_Bool_11QNone_Bool_bufchan_d;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_QTree_Bool) : (lizzieLet0_4QNode_Bool_4QNode_Bool_12,QTree_Bool) (t4a8U_destruct,Pointer_QTree_Bool) > [(lizzieLet0_4QNode_Bool_4QNode_Bool_12QNone_Bool,Pointer_QTree_Bool),
                                                                                                                          (_154,Pointer_QTree_Bool),
                                                                                                                          (lizzieLet0_4QNode_Bool_4QNode_Bool_12QNode_Bool,Pointer_QTree_Bool),
                                                                                                                          (_153,Pointer_QTree_Bool)] */
  logic [3:0] t4a8U_destruct_onehotd;
  always_comb
    if ((lizzieLet0_4QNode_Bool_4QNode_Bool_12_d[0] && t4a8U_destruct_d[0]))
      unique case (lizzieLet0_4QNode_Bool_4QNode_Bool_12_d[2:1])
        2'd0: t4a8U_destruct_onehotd = 4'd1;
        2'd1: t4a8U_destruct_onehotd = 4'd2;
        2'd2: t4a8U_destruct_onehotd = 4'd4;
        2'd3: t4a8U_destruct_onehotd = 4'd8;
        default: t4a8U_destruct_onehotd = 4'd0;
      endcase
    else t4a8U_destruct_onehotd = 4'd0;
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_12QNone_Bool_d = {t4a8U_destruct_d[16:1],
                                                              t4a8U_destruct_onehotd[0]};
  assign _154_d = {t4a8U_destruct_d[16:1],
                   t4a8U_destruct_onehotd[1]};
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_12QNode_Bool_d = {t4a8U_destruct_d[16:1],
                                                              t4a8U_destruct_onehotd[2]};
  assign _153_d = {t4a8U_destruct_d[16:1],
                   t4a8U_destruct_onehotd[3]};
  assign t4a8U_destruct_r = (| (t4a8U_destruct_onehotd & {_153_r,
                                                          lizzieLet0_4QNode_Bool_4QNode_Bool_12QNode_Bool_r,
                                                          _154_r,
                                                          lizzieLet0_4QNode_Bool_4QNode_Bool_12QNone_Bool_r}));
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_12_r = t4a8U_destruct_r;
  
  /* buf (Ty Pointer_QTree_Bool) : (lizzieLet0_4QNode_Bool_4QNode_Bool_12QNode_Bool,Pointer_QTree_Bool) > (lizzieLet0_4QNode_Bool_4QNode_Bool_12QNode_Bool_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t lizzieLet0_4QNode_Bool_4QNode_Bool_12QNode_Bool_bufchan_d;
  logic lizzieLet0_4QNode_Bool_4QNode_Bool_12QNode_Bool_bufchan_r;
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_12QNode_Bool_r = ((! lizzieLet0_4QNode_Bool_4QNode_Bool_12QNode_Bool_bufchan_d[0]) || lizzieLet0_4QNode_Bool_4QNode_Bool_12QNode_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNode_Bool_4QNode_Bool_12QNode_Bool_bufchan_d <= {16'd0,
                                                                    1'd0};
    else
      if (lizzieLet0_4QNode_Bool_4QNode_Bool_12QNode_Bool_r)
        lizzieLet0_4QNode_Bool_4QNode_Bool_12QNode_Bool_bufchan_d <= lizzieLet0_4QNode_Bool_4QNode_Bool_12QNode_Bool_d;
  Pointer_QTree_Bool_t lizzieLet0_4QNode_Bool_4QNode_Bool_12QNode_Bool_bufchan_buf;
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_12QNode_Bool_bufchan_r = (! lizzieLet0_4QNode_Bool_4QNode_Bool_12QNode_Bool_bufchan_buf[0]);
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_12QNode_Bool_1_argbuf_d = (lizzieLet0_4QNode_Bool_4QNode_Bool_12QNode_Bool_bufchan_buf[0] ? lizzieLet0_4QNode_Bool_4QNode_Bool_12QNode_Bool_bufchan_buf :
                                                                       lizzieLet0_4QNode_Bool_4QNode_Bool_12QNode_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNode_Bool_4QNode_Bool_12QNode_Bool_bufchan_buf <= {16'd0,
                                                                      1'd0};
    else
      if ((lizzieLet0_4QNode_Bool_4QNode_Bool_12QNode_Bool_1_argbuf_r && lizzieLet0_4QNode_Bool_4QNode_Bool_12QNode_Bool_bufchan_buf[0]))
        lizzieLet0_4QNode_Bool_4QNode_Bool_12QNode_Bool_bufchan_buf <= {16'd0,
                                                                        1'd0};
      else if (((! lizzieLet0_4QNode_Bool_4QNode_Bool_12QNode_Bool_1_argbuf_r) && (! lizzieLet0_4QNode_Bool_4QNode_Bool_12QNode_Bool_bufchan_buf[0])))
        lizzieLet0_4QNode_Bool_4QNode_Bool_12QNode_Bool_bufchan_buf <= lizzieLet0_4QNode_Bool_4QNode_Bool_12QNode_Bool_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (lizzieLet0_4QNode_Bool_4QNode_Bool_12QNone_Bool,Pointer_QTree_Bool) > (lizzieLet0_4QNode_Bool_4QNode_Bool_12QNone_Bool_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t lizzieLet0_4QNode_Bool_4QNode_Bool_12QNone_Bool_bufchan_d;
  logic lizzieLet0_4QNode_Bool_4QNode_Bool_12QNone_Bool_bufchan_r;
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_12QNone_Bool_r = ((! lizzieLet0_4QNode_Bool_4QNode_Bool_12QNone_Bool_bufchan_d[0]) || lizzieLet0_4QNode_Bool_4QNode_Bool_12QNone_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNode_Bool_4QNode_Bool_12QNone_Bool_bufchan_d <= {16'd0,
                                                                    1'd0};
    else
      if (lizzieLet0_4QNode_Bool_4QNode_Bool_12QNone_Bool_r)
        lizzieLet0_4QNode_Bool_4QNode_Bool_12QNone_Bool_bufchan_d <= lizzieLet0_4QNode_Bool_4QNode_Bool_12QNone_Bool_d;
  Pointer_QTree_Bool_t lizzieLet0_4QNode_Bool_4QNode_Bool_12QNone_Bool_bufchan_buf;
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_12QNone_Bool_bufchan_r = (! lizzieLet0_4QNode_Bool_4QNode_Bool_12QNone_Bool_bufchan_buf[0]);
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_12QNone_Bool_1_argbuf_d = (lizzieLet0_4QNode_Bool_4QNode_Bool_12QNone_Bool_bufchan_buf[0] ? lizzieLet0_4QNode_Bool_4QNode_Bool_12QNone_Bool_bufchan_buf :
                                                                       lizzieLet0_4QNode_Bool_4QNode_Bool_12QNone_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNode_Bool_4QNode_Bool_12QNone_Bool_bufchan_buf <= {16'd0,
                                                                      1'd0};
    else
      if ((lizzieLet0_4QNode_Bool_4QNode_Bool_12QNone_Bool_1_argbuf_r && lizzieLet0_4QNode_Bool_4QNode_Bool_12QNone_Bool_bufchan_buf[0]))
        lizzieLet0_4QNode_Bool_4QNode_Bool_12QNone_Bool_bufchan_buf <= {16'd0,
                                                                        1'd0};
      else if (((! lizzieLet0_4QNode_Bool_4QNode_Bool_12QNone_Bool_1_argbuf_r) && (! lizzieLet0_4QNode_Bool_4QNode_Bool_12QNone_Bool_bufchan_buf[0])))
        lizzieLet0_4QNode_Bool_4QNode_Bool_12QNone_Bool_bufchan_buf <= lizzieLet0_4QNode_Bool_4QNode_Bool_12QNone_Bool_bufchan_d;
  
  /* destruct (Ty QTree_Bool,
          Dcon QNode_Bool) : (lizzieLet0_4QNode_Bool_4QNode_Bool_1QNode_Bool,QTree_Bool) > [(t1'a8W_destruct,Pointer_QTree_Bool),
                                                                                            (t2'a8X_destruct,Pointer_QTree_Bool),
                                                                                            (t3'a8Y_destruct,Pointer_QTree_Bool),
                                                                                            (t4'a8Z_destruct,Pointer_QTree_Bool)] */
  logic [3:0] lizzieLet0_4QNode_Bool_4QNode_Bool_1QNode_Bool_emitted;
  logic [3:0] lizzieLet0_4QNode_Bool_4QNode_Bool_1QNode_Bool_done;
  assign \t1'a8W_destruct_d  = {lizzieLet0_4QNode_Bool_4QNode_Bool_1QNode_Bool_d[18:3],
                                (lizzieLet0_4QNode_Bool_4QNode_Bool_1QNode_Bool_d[0] && (! lizzieLet0_4QNode_Bool_4QNode_Bool_1QNode_Bool_emitted[0]))};
  assign \t2'a8X_destruct_d  = {lizzieLet0_4QNode_Bool_4QNode_Bool_1QNode_Bool_d[34:19],
                                (lizzieLet0_4QNode_Bool_4QNode_Bool_1QNode_Bool_d[0] && (! lizzieLet0_4QNode_Bool_4QNode_Bool_1QNode_Bool_emitted[1]))};
  assign \t3'a8Y_destruct_d  = {lizzieLet0_4QNode_Bool_4QNode_Bool_1QNode_Bool_d[50:35],
                                (lizzieLet0_4QNode_Bool_4QNode_Bool_1QNode_Bool_d[0] && (! lizzieLet0_4QNode_Bool_4QNode_Bool_1QNode_Bool_emitted[2]))};
  assign \t4'a8Z_destruct_d  = {lizzieLet0_4QNode_Bool_4QNode_Bool_1QNode_Bool_d[66:51],
                                (lizzieLet0_4QNode_Bool_4QNode_Bool_1QNode_Bool_d[0] && (! lizzieLet0_4QNode_Bool_4QNode_Bool_1QNode_Bool_emitted[3]))};
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_1QNode_Bool_done = (lizzieLet0_4QNode_Bool_4QNode_Bool_1QNode_Bool_emitted | ({\t4'a8Z_destruct_d [0],
                                                                                                                           \t3'a8Y_destruct_d [0],
                                                                                                                           \t2'a8X_destruct_d [0],
                                                                                                                           \t1'a8W_destruct_d [0]} & {\t4'a8Z_destruct_r ,
                                                                                                                                                      \t3'a8Y_destruct_r ,
                                                                                                                                                      \t2'a8X_destruct_r ,
                                                                                                                                                      \t1'a8W_destruct_r }));
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_1QNode_Bool_r = (& lizzieLet0_4QNode_Bool_4QNode_Bool_1QNode_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNode_Bool_4QNode_Bool_1QNode_Bool_emitted <= 4'd0;
    else
      lizzieLet0_4QNode_Bool_4QNode_Bool_1QNode_Bool_emitted <= (lizzieLet0_4QNode_Bool_4QNode_Bool_1QNode_Bool_r ? 4'd0 :
                                                                 lizzieLet0_4QNode_Bool_4QNode_Bool_1QNode_Bool_done);
  
  /* demux (Ty QTree_Bool,
       Ty QTree_Bool) : (lizzieLet0_4QNode_Bool_4QNode_Bool_2,QTree_Bool) (lizzieLet0_4QNode_Bool_4QNode_Bool_1,QTree_Bool) > [(_152,QTree_Bool),
                                                                                                                               (_151,QTree_Bool),
                                                                                                                               (lizzieLet0_4QNode_Bool_4QNode_Bool_1QNode_Bool,QTree_Bool),
                                                                                                                               (_150,QTree_Bool)] */
  logic [3:0] lizzieLet0_4QNode_Bool_4QNode_Bool_1_onehotd;
  always_comb
    if ((lizzieLet0_4QNode_Bool_4QNode_Bool_2_d[0] && lizzieLet0_4QNode_Bool_4QNode_Bool_1_d[0]))
      unique case (lizzieLet0_4QNode_Bool_4QNode_Bool_2_d[2:1])
        2'd0: lizzieLet0_4QNode_Bool_4QNode_Bool_1_onehotd = 4'd1;
        2'd1: lizzieLet0_4QNode_Bool_4QNode_Bool_1_onehotd = 4'd2;
        2'd2: lizzieLet0_4QNode_Bool_4QNode_Bool_1_onehotd = 4'd4;
        2'd3: lizzieLet0_4QNode_Bool_4QNode_Bool_1_onehotd = 4'd8;
        default: lizzieLet0_4QNode_Bool_4QNode_Bool_1_onehotd = 4'd0;
      endcase
    else lizzieLet0_4QNode_Bool_4QNode_Bool_1_onehotd = 4'd0;
  assign _152_d = {lizzieLet0_4QNode_Bool_4QNode_Bool_1_d[66:1],
                   lizzieLet0_4QNode_Bool_4QNode_Bool_1_onehotd[0]};
  assign _151_d = {lizzieLet0_4QNode_Bool_4QNode_Bool_1_d[66:1],
                   lizzieLet0_4QNode_Bool_4QNode_Bool_1_onehotd[1]};
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_1QNode_Bool_d = {lizzieLet0_4QNode_Bool_4QNode_Bool_1_d[66:1],
                                                             lizzieLet0_4QNode_Bool_4QNode_Bool_1_onehotd[2]};
  assign _150_d = {lizzieLet0_4QNode_Bool_4QNode_Bool_1_d[66:1],
                   lizzieLet0_4QNode_Bool_4QNode_Bool_1_onehotd[3]};
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_1_r = (| (lizzieLet0_4QNode_Bool_4QNode_Bool_1_onehotd & {_150_r,
                                                                                                      lizzieLet0_4QNode_Bool_4QNode_Bool_1QNode_Bool_r,
                                                                                                      _151_r,
                                                                                                      _152_r}));
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_2_r = lizzieLet0_4QNode_Bool_4QNode_Bool_1_r;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_QTree_Bool) : (lizzieLet0_4QNode_Bool_4QNode_Bool_3,QTree_Bool) (lizzieLet0_4QNode_Bool_10QNode_Bool,Pointer_QTree_Bool) > [(lizzieLet0_4QNode_Bool_4QNode_Bool_3QNone_Bool,Pointer_QTree_Bool),
                                                                                                                                              (_149,Pointer_QTree_Bool),
                                                                                                                                              (lizzieLet0_4QNode_Bool_4QNode_Bool_3QNode_Bool,Pointer_QTree_Bool),
                                                                                                                                              (_148,Pointer_QTree_Bool)] */
  logic [3:0] lizzieLet0_4QNode_Bool_10QNode_Bool_onehotd;
  always_comb
    if ((lizzieLet0_4QNode_Bool_4QNode_Bool_3_d[0] && lizzieLet0_4QNode_Bool_10QNode_Bool_d[0]))
      unique case (lizzieLet0_4QNode_Bool_4QNode_Bool_3_d[2:1])
        2'd0: lizzieLet0_4QNode_Bool_10QNode_Bool_onehotd = 4'd1;
        2'd1: lizzieLet0_4QNode_Bool_10QNode_Bool_onehotd = 4'd2;
        2'd2: lizzieLet0_4QNode_Bool_10QNode_Bool_onehotd = 4'd4;
        2'd3: lizzieLet0_4QNode_Bool_10QNode_Bool_onehotd = 4'd8;
        default: lizzieLet0_4QNode_Bool_10QNode_Bool_onehotd = 4'd0;
      endcase
    else lizzieLet0_4QNode_Bool_10QNode_Bool_onehotd = 4'd0;
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_3QNone_Bool_d = {lizzieLet0_4QNode_Bool_10QNode_Bool_d[16:1],
                                                             lizzieLet0_4QNode_Bool_10QNode_Bool_onehotd[0]};
  assign _149_d = {lizzieLet0_4QNode_Bool_10QNode_Bool_d[16:1],
                   lizzieLet0_4QNode_Bool_10QNode_Bool_onehotd[1]};
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_3QNode_Bool_d = {lizzieLet0_4QNode_Bool_10QNode_Bool_d[16:1],
                                                             lizzieLet0_4QNode_Bool_10QNode_Bool_onehotd[2]};
  assign _148_d = {lizzieLet0_4QNode_Bool_10QNode_Bool_d[16:1],
                   lizzieLet0_4QNode_Bool_10QNode_Bool_onehotd[3]};
  assign lizzieLet0_4QNode_Bool_10QNode_Bool_r = (| (lizzieLet0_4QNode_Bool_10QNode_Bool_onehotd & {_148_r,
                                                                                                    lizzieLet0_4QNode_Bool_4QNode_Bool_3QNode_Bool_r,
                                                                                                    _149_r,
                                                                                                    lizzieLet0_4QNode_Bool_4QNode_Bool_3QNone_Bool_r}));
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_3_r = lizzieLet0_4QNode_Bool_10QNode_Bool_r;
  
  /* buf (Ty Pointer_QTree_Bool) : (lizzieLet0_4QNode_Bool_4QNode_Bool_3QNode_Bool,Pointer_QTree_Bool) > (lizzieLet0_4QNode_Bool_4QNode_Bool_3QNode_Bool_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t lizzieLet0_4QNode_Bool_4QNode_Bool_3QNode_Bool_bufchan_d;
  logic lizzieLet0_4QNode_Bool_4QNode_Bool_3QNode_Bool_bufchan_r;
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_3QNode_Bool_r = ((! lizzieLet0_4QNode_Bool_4QNode_Bool_3QNode_Bool_bufchan_d[0]) || lizzieLet0_4QNode_Bool_4QNode_Bool_3QNode_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNode_Bool_4QNode_Bool_3QNode_Bool_bufchan_d <= {16'd0,
                                                                   1'd0};
    else
      if (lizzieLet0_4QNode_Bool_4QNode_Bool_3QNode_Bool_r)
        lizzieLet0_4QNode_Bool_4QNode_Bool_3QNode_Bool_bufchan_d <= lizzieLet0_4QNode_Bool_4QNode_Bool_3QNode_Bool_d;
  Pointer_QTree_Bool_t lizzieLet0_4QNode_Bool_4QNode_Bool_3QNode_Bool_bufchan_buf;
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_3QNode_Bool_bufchan_r = (! lizzieLet0_4QNode_Bool_4QNode_Bool_3QNode_Bool_bufchan_buf[0]);
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_3QNode_Bool_1_argbuf_d = (lizzieLet0_4QNode_Bool_4QNode_Bool_3QNode_Bool_bufchan_buf[0] ? lizzieLet0_4QNode_Bool_4QNode_Bool_3QNode_Bool_bufchan_buf :
                                                                      lizzieLet0_4QNode_Bool_4QNode_Bool_3QNode_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNode_Bool_4QNode_Bool_3QNode_Bool_bufchan_buf <= {16'd0,
                                                                     1'd0};
    else
      if ((lizzieLet0_4QNode_Bool_4QNode_Bool_3QNode_Bool_1_argbuf_r && lizzieLet0_4QNode_Bool_4QNode_Bool_3QNode_Bool_bufchan_buf[0]))
        lizzieLet0_4QNode_Bool_4QNode_Bool_3QNode_Bool_bufchan_buf <= {16'd0,
                                                                       1'd0};
      else if (((! lizzieLet0_4QNode_Bool_4QNode_Bool_3QNode_Bool_1_argbuf_r) && (! lizzieLet0_4QNode_Bool_4QNode_Bool_3QNode_Bool_bufchan_buf[0])))
        lizzieLet0_4QNode_Bool_4QNode_Bool_3QNode_Bool_bufchan_buf <= lizzieLet0_4QNode_Bool_4QNode_Bool_3QNode_Bool_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (lizzieLet0_4QNode_Bool_4QNode_Bool_3QNone_Bool,Pointer_QTree_Bool) > (lizzieLet0_4QNode_Bool_4QNode_Bool_3QNone_Bool_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t lizzieLet0_4QNode_Bool_4QNode_Bool_3QNone_Bool_bufchan_d;
  logic lizzieLet0_4QNode_Bool_4QNode_Bool_3QNone_Bool_bufchan_r;
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_3QNone_Bool_r = ((! lizzieLet0_4QNode_Bool_4QNode_Bool_3QNone_Bool_bufchan_d[0]) || lizzieLet0_4QNode_Bool_4QNode_Bool_3QNone_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNode_Bool_4QNode_Bool_3QNone_Bool_bufchan_d <= {16'd0,
                                                                   1'd0};
    else
      if (lizzieLet0_4QNode_Bool_4QNode_Bool_3QNone_Bool_r)
        lizzieLet0_4QNode_Bool_4QNode_Bool_3QNone_Bool_bufchan_d <= lizzieLet0_4QNode_Bool_4QNode_Bool_3QNone_Bool_d;
  Pointer_QTree_Bool_t lizzieLet0_4QNode_Bool_4QNode_Bool_3QNone_Bool_bufchan_buf;
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_3QNone_Bool_bufchan_r = (! lizzieLet0_4QNode_Bool_4QNode_Bool_3QNone_Bool_bufchan_buf[0]);
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_3QNone_Bool_1_argbuf_d = (lizzieLet0_4QNode_Bool_4QNode_Bool_3QNone_Bool_bufchan_buf[0] ? lizzieLet0_4QNode_Bool_4QNode_Bool_3QNone_Bool_bufchan_buf :
                                                                      lizzieLet0_4QNode_Bool_4QNode_Bool_3QNone_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNode_Bool_4QNode_Bool_3QNone_Bool_bufchan_buf <= {16'd0,
                                                                     1'd0};
    else
      if ((lizzieLet0_4QNode_Bool_4QNode_Bool_3QNone_Bool_1_argbuf_r && lizzieLet0_4QNode_Bool_4QNode_Bool_3QNone_Bool_bufchan_buf[0]))
        lizzieLet0_4QNode_Bool_4QNode_Bool_3QNone_Bool_bufchan_buf <= {16'd0,
                                                                       1'd0};
      else if (((! lizzieLet0_4QNode_Bool_4QNode_Bool_3QNone_Bool_1_argbuf_r) && (! lizzieLet0_4QNode_Bool_4QNode_Bool_3QNone_Bool_bufchan_buf[0])))
        lizzieLet0_4QNode_Bool_4QNode_Bool_3QNone_Bool_bufchan_buf <= lizzieLet0_4QNode_Bool_4QNode_Bool_3QNone_Bool_bufchan_d;
  
  /* demux (Ty QTree_Bool,
       Ty Go) : (lizzieLet0_4QNode_Bool_4QNode_Bool_4,QTree_Bool) (lizzieLet0_4QNode_Bool_3QNode_Bool,Go) > [(lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool,Go),
                                                                                                             (lizzieLet0_4QNode_Bool_4QNode_Bool_4QVal_Bool,Go),
                                                                                                             (lizzieLet0_4QNode_Bool_4QNode_Bool_4QNode_Bool,Go),
                                                                                                             (lizzieLet0_4QNode_Bool_4QNode_Bool_4QError_Bool,Go)] */
  logic [3:0] lizzieLet0_4QNode_Bool_3QNode_Bool_onehotd;
  always_comb
    if ((lizzieLet0_4QNode_Bool_4QNode_Bool_4_d[0] && lizzieLet0_4QNode_Bool_3QNode_Bool_d[0]))
      unique case (lizzieLet0_4QNode_Bool_4QNode_Bool_4_d[2:1])
        2'd0: lizzieLet0_4QNode_Bool_3QNode_Bool_onehotd = 4'd1;
        2'd1: lizzieLet0_4QNode_Bool_3QNode_Bool_onehotd = 4'd2;
        2'd2: lizzieLet0_4QNode_Bool_3QNode_Bool_onehotd = 4'd4;
        2'd3: lizzieLet0_4QNode_Bool_3QNode_Bool_onehotd = 4'd8;
        default: lizzieLet0_4QNode_Bool_3QNode_Bool_onehotd = 4'd0;
      endcase
    else lizzieLet0_4QNode_Bool_3QNode_Bool_onehotd = 4'd0;
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_d = lizzieLet0_4QNode_Bool_3QNode_Bool_onehotd[0];
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_4QVal_Bool_d = lizzieLet0_4QNode_Bool_3QNode_Bool_onehotd[1];
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_4QNode_Bool_d = lizzieLet0_4QNode_Bool_3QNode_Bool_onehotd[2];
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_4QError_Bool_d = lizzieLet0_4QNode_Bool_3QNode_Bool_onehotd[3];
  assign lizzieLet0_4QNode_Bool_3QNode_Bool_r = (| (lizzieLet0_4QNode_Bool_3QNode_Bool_onehotd & {lizzieLet0_4QNode_Bool_4QNode_Bool_4QError_Bool_r,
                                                                                                  lizzieLet0_4QNode_Bool_4QNode_Bool_4QNode_Bool_r,
                                                                                                  lizzieLet0_4QNode_Bool_4QNode_Bool_4QVal_Bool_r,
                                                                                                  lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_r}));
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_4_r = lizzieLet0_4QNode_Bool_3QNode_Bool_r;
  
  /* fork (Ty Go) : (lizzieLet0_4QNode_Bool_4QNode_Bool_4QError_Bool,Go) > [(lizzieLet0_4QNode_Bool_4QNode_Bool_4QError_Bool_1,Go),
                                                                       (lizzieLet0_4QNode_Bool_4QNode_Bool_4QError_Bool_2,Go)] */
  logic [1:0] lizzieLet0_4QNode_Bool_4QNode_Bool_4QError_Bool_emitted;
  logic [1:0] lizzieLet0_4QNode_Bool_4QNode_Bool_4QError_Bool_done;
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_4QError_Bool_1_d = (lizzieLet0_4QNode_Bool_4QNode_Bool_4QError_Bool_d[0] && (! lizzieLet0_4QNode_Bool_4QNode_Bool_4QError_Bool_emitted[0]));
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_4QError_Bool_2_d = (lizzieLet0_4QNode_Bool_4QNode_Bool_4QError_Bool_d[0] && (! lizzieLet0_4QNode_Bool_4QNode_Bool_4QError_Bool_emitted[1]));
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_4QError_Bool_done = (lizzieLet0_4QNode_Bool_4QNode_Bool_4QError_Bool_emitted | ({lizzieLet0_4QNode_Bool_4QNode_Bool_4QError_Bool_2_d[0],
                                                                                                                             lizzieLet0_4QNode_Bool_4QNode_Bool_4QError_Bool_1_d[0]} & {lizzieLet0_4QNode_Bool_4QNode_Bool_4QError_Bool_2_r,
                                                                                                                                                                                        lizzieLet0_4QNode_Bool_4QNode_Bool_4QError_Bool_1_r}));
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_4QError_Bool_r = (& lizzieLet0_4QNode_Bool_4QNode_Bool_4QError_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNode_Bool_4QNode_Bool_4QError_Bool_emitted <= 2'd0;
    else
      lizzieLet0_4QNode_Bool_4QNode_Bool_4QError_Bool_emitted <= (lizzieLet0_4QNode_Bool_4QNode_Bool_4QError_Bool_r ? 2'd0 :
                                                                  lizzieLet0_4QNode_Bool_4QNode_Bool_4QError_Bool_done);
  
  /* dcon (Ty QTree_Bool,
      Dcon QError_Bool) : [(lizzieLet0_4QNode_Bool_4QNode_Bool_4QError_Bool_1,Go)] > (lizzieLet0_4QNode_Bool_4QNode_Bool_4QError_Bool_1QError_Bool,QTree_Bool) */
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_4QError_Bool_1QError_Bool_d = QError_Bool_dc((& {lizzieLet0_4QNode_Bool_4QNode_Bool_4QError_Bool_1_d[0]}), lizzieLet0_4QNode_Bool_4QNode_Bool_4QError_Bool_1_d);
  assign {lizzieLet0_4QNode_Bool_4QNode_Bool_4QError_Bool_1_r} = {1 {(lizzieLet0_4QNode_Bool_4QNode_Bool_4QError_Bool_1QError_Bool_r && lizzieLet0_4QNode_Bool_4QNode_Bool_4QError_Bool_1QError_Bool_d[0])}};
  
  /* buf (Ty QTree_Bool) : (lizzieLet0_4QNode_Bool_4QNode_Bool_4QError_Bool_1QError_Bool,QTree_Bool) > (lizzieLet42_1_argbuf,QTree_Bool) */
  QTree_Bool_t lizzieLet0_4QNode_Bool_4QNode_Bool_4QError_Bool_1QError_Bool_bufchan_d;
  logic lizzieLet0_4QNode_Bool_4QNode_Bool_4QError_Bool_1QError_Bool_bufchan_r;
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_4QError_Bool_1QError_Bool_r = ((! lizzieLet0_4QNode_Bool_4QNode_Bool_4QError_Bool_1QError_Bool_bufchan_d[0]) || lizzieLet0_4QNode_Bool_4QNode_Bool_4QError_Bool_1QError_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNode_Bool_4QNode_Bool_4QError_Bool_1QError_Bool_bufchan_d <= {66'd0,
                                                                                 1'd0};
    else
      if (lizzieLet0_4QNode_Bool_4QNode_Bool_4QError_Bool_1QError_Bool_r)
        lizzieLet0_4QNode_Bool_4QNode_Bool_4QError_Bool_1QError_Bool_bufchan_d <= lizzieLet0_4QNode_Bool_4QNode_Bool_4QError_Bool_1QError_Bool_d;
  QTree_Bool_t lizzieLet0_4QNode_Bool_4QNode_Bool_4QError_Bool_1QError_Bool_bufchan_buf;
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_4QError_Bool_1QError_Bool_bufchan_r = (! lizzieLet0_4QNode_Bool_4QNode_Bool_4QError_Bool_1QError_Bool_bufchan_buf[0]);
  assign lizzieLet42_1_argbuf_d = (lizzieLet0_4QNode_Bool_4QNode_Bool_4QError_Bool_1QError_Bool_bufchan_buf[0] ? lizzieLet0_4QNode_Bool_4QNode_Bool_4QError_Bool_1QError_Bool_bufchan_buf :
                                   lizzieLet0_4QNode_Bool_4QNode_Bool_4QError_Bool_1QError_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNode_Bool_4QNode_Bool_4QError_Bool_1QError_Bool_bufchan_buf <= {66'd0,
                                                                                   1'd0};
    else
      if ((lizzieLet42_1_argbuf_r && lizzieLet0_4QNode_Bool_4QNode_Bool_4QError_Bool_1QError_Bool_bufchan_buf[0]))
        lizzieLet0_4QNode_Bool_4QNode_Bool_4QError_Bool_1QError_Bool_bufchan_buf <= {66'd0,
                                                                                     1'd0};
      else if (((! lizzieLet42_1_argbuf_r) && (! lizzieLet0_4QNode_Bool_4QNode_Bool_4QError_Bool_1QError_Bool_bufchan_buf[0])))
        lizzieLet0_4QNode_Bool_4QNode_Bool_4QError_Bool_1QError_Bool_bufchan_buf <= lizzieLet0_4QNode_Bool_4QNode_Bool_4QError_Bool_1QError_Bool_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet0_4QNode_Bool_4QNode_Bool_4QError_Bool_2,Go) > (lizzieLet0_4QNode_Bool_4QNode_Bool_4QError_Bool_2_argbuf,Go) */
  Go_t lizzieLet0_4QNode_Bool_4QNode_Bool_4QError_Bool_2_bufchan_d;
  logic lizzieLet0_4QNode_Bool_4QNode_Bool_4QError_Bool_2_bufchan_r;
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_4QError_Bool_2_r = ((! lizzieLet0_4QNode_Bool_4QNode_Bool_4QError_Bool_2_bufchan_d[0]) || lizzieLet0_4QNode_Bool_4QNode_Bool_4QError_Bool_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNode_Bool_4QNode_Bool_4QError_Bool_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet0_4QNode_Bool_4QNode_Bool_4QError_Bool_2_r)
        lizzieLet0_4QNode_Bool_4QNode_Bool_4QError_Bool_2_bufchan_d <= lizzieLet0_4QNode_Bool_4QNode_Bool_4QError_Bool_2_d;
  Go_t lizzieLet0_4QNode_Bool_4QNode_Bool_4QError_Bool_2_bufchan_buf;
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_4QError_Bool_2_bufchan_r = (! lizzieLet0_4QNode_Bool_4QNode_Bool_4QError_Bool_2_bufchan_buf[0]);
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_4QError_Bool_2_argbuf_d = (lizzieLet0_4QNode_Bool_4QNode_Bool_4QError_Bool_2_bufchan_buf[0] ? lizzieLet0_4QNode_Bool_4QNode_Bool_4QError_Bool_2_bufchan_buf :
                                                                       lizzieLet0_4QNode_Bool_4QNode_Bool_4QError_Bool_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNode_Bool_4QNode_Bool_4QError_Bool_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet0_4QNode_Bool_4QNode_Bool_4QError_Bool_2_argbuf_r && lizzieLet0_4QNode_Bool_4QNode_Bool_4QError_Bool_2_bufchan_buf[0]))
        lizzieLet0_4QNode_Bool_4QNode_Bool_4QError_Bool_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet0_4QNode_Bool_4QNode_Bool_4QError_Bool_2_argbuf_r) && (! lizzieLet0_4QNode_Bool_4QNode_Bool_4QError_Bool_2_bufchan_buf[0])))
        lizzieLet0_4QNode_Bool_4QNode_Bool_4QError_Bool_2_bufchan_buf <= lizzieLet0_4QNode_Bool_4QNode_Bool_4QError_Bool_2_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet0_4QNode_Bool_4QNode_Bool_4QNode_Bool,Go) > (lizzieLet0_4QNode_Bool_4QNode_Bool_4QNode_Bool_1_argbuf,Go) */
  Go_t lizzieLet0_4QNode_Bool_4QNode_Bool_4QNode_Bool_bufchan_d;
  logic lizzieLet0_4QNode_Bool_4QNode_Bool_4QNode_Bool_bufchan_r;
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_4QNode_Bool_r = ((! lizzieLet0_4QNode_Bool_4QNode_Bool_4QNode_Bool_bufchan_d[0]) || lizzieLet0_4QNode_Bool_4QNode_Bool_4QNode_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNode_Bool_4QNode_Bool_4QNode_Bool_bufchan_d <= 1'd0;
    else
      if (lizzieLet0_4QNode_Bool_4QNode_Bool_4QNode_Bool_r)
        lizzieLet0_4QNode_Bool_4QNode_Bool_4QNode_Bool_bufchan_d <= lizzieLet0_4QNode_Bool_4QNode_Bool_4QNode_Bool_d;
  Go_t lizzieLet0_4QNode_Bool_4QNode_Bool_4QNode_Bool_bufchan_buf;
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_4QNode_Bool_bufchan_r = (! lizzieLet0_4QNode_Bool_4QNode_Bool_4QNode_Bool_bufchan_buf[0]);
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_4QNode_Bool_1_argbuf_d = (lizzieLet0_4QNode_Bool_4QNode_Bool_4QNode_Bool_bufchan_buf[0] ? lizzieLet0_4QNode_Bool_4QNode_Bool_4QNode_Bool_bufchan_buf :
                                                                      lizzieLet0_4QNode_Bool_4QNode_Bool_4QNode_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNode_Bool_4QNode_Bool_4QNode_Bool_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet0_4QNode_Bool_4QNode_Bool_4QNode_Bool_1_argbuf_r && lizzieLet0_4QNode_Bool_4QNode_Bool_4QNode_Bool_bufchan_buf[0]))
        lizzieLet0_4QNode_Bool_4QNode_Bool_4QNode_Bool_bufchan_buf <= 1'd0;
      else if (((! lizzieLet0_4QNode_Bool_4QNode_Bool_4QNode_Bool_1_argbuf_r) && (! lizzieLet0_4QNode_Bool_4QNode_Bool_4QNode_Bool_bufchan_buf[0])))
        lizzieLet0_4QNode_Bool_4QNode_Bool_4QNode_Bool_bufchan_buf <= lizzieLet0_4QNode_Bool_4QNode_Bool_4QNode_Bool_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool,Go) > [(lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_1,Go),
                                                                      (lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_2,Go),
                                                                      (lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_3,Go),
                                                                      (lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_4,Go),
                                                                      (lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_5,Go)] */
  logic [4:0] lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_emitted;
  logic [4:0] lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_done;
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_1_d = (lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_d[0] && (! lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_emitted[0]));
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_2_d = (lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_d[0] && (! lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_emitted[1]));
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_3_d = (lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_d[0] && (! lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_emitted[2]));
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_4_d = (lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_d[0] && (! lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_emitted[3]));
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_5_d = (lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_d[0] && (! lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_emitted[4]));
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_done = (lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_emitted | ({lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_5_d[0],
                                                                                                                           lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_4_d[0],
                                                                                                                           lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_3_d[0],
                                                                                                                           lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_2_d[0],
                                                                                                                           lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_1_d[0]} & {lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_5_r,
                                                                                                                                                                                     lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_4_r,
                                                                                                                                                                                     lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_3_r,
                                                                                                                                                                                     lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_2_r,
                                                                                                                                                                                     lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_1_r}));
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_r = (& lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_emitted <= 5'd0;
    else
      lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_emitted <= (lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_r ? 5'd0 :
                                                                 lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_done);
  
  /* buf (Ty Go) : (lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_1,Go) > (lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_1_argbuf,Go) */
  Go_t lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_1_bufchan_d;
  logic lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_1_bufchan_r;
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_1_r = ((! lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_1_bufchan_d[0]) || lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_1_bufchan_d <= 1'd0;
    else
      if (lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_1_r)
        lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_1_bufchan_d <= lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_1_d;
  Go_t lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_1_bufchan_buf;
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_1_bufchan_r = (! lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_1_bufchan_buf[0]);
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_1_argbuf_d = (lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_1_bufchan_buf[0] ? lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_1_bufchan_buf :
                                                                      lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_1_argbuf_r && lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_1_bufchan_buf[0]))
        lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_1_argbuf_r) && (! lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_1_bufchan_buf[0])))
        lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_1_bufchan_buf <= lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_1_bufchan_d;
  
  /* dcon (Ty TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool,
      Dcon TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool) : [(lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_1_argbuf,Go),
                                                               (lizzieLet0_4QNode_Bool_4QNode_Bool_3QNone_Bool_1_argbuf,Pointer_QTree_Bool),
                                                               (lizzieLet0_4QNode_Bool_4QNode_Bool_12QNone_Bool_1_argbuf,Pointer_QTree_Bool)] > (f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool9,TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool) */
  assign \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool9_d  = TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_dc((& {lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_1_argbuf_d[0],
                                                                                                                                    lizzieLet0_4QNode_Bool_4QNode_Bool_3QNone_Bool_1_argbuf_d[0],
                                                                                                                                    lizzieLet0_4QNode_Bool_4QNode_Bool_12QNone_Bool_1_argbuf_d[0]}), lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_1_argbuf_d, lizzieLet0_4QNode_Bool_4QNode_Bool_3QNone_Bool_1_argbuf_d, lizzieLet0_4QNode_Bool_4QNode_Bool_12QNone_Bool_1_argbuf_d);
  assign {lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_1_argbuf_r,
          lizzieLet0_4QNode_Bool_4QNode_Bool_3QNone_Bool_1_argbuf_r,
          lizzieLet0_4QNode_Bool_4QNode_Bool_12QNone_Bool_1_argbuf_r} = {3 {(\f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool9_r  && \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool9_d [0])}};
  
  /* buf (Ty Go) : (lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_2,Go) > (lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_2_argbuf,Go) */
  Go_t lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_2_bufchan_d;
  logic lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_2_bufchan_r;
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_2_r = ((! lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_2_bufchan_d[0]) || lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_2_r)
        lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_2_bufchan_d <= lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_2_d;
  Go_t lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_2_bufchan_buf;
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_2_bufchan_r = (! lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_2_bufchan_buf[0]);
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_2_argbuf_d = (lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_2_bufchan_buf[0] ? lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_2_bufchan_buf :
                                                                      lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_2_argbuf_r && lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_2_bufchan_buf[0]))
        lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_2_argbuf_r) && (! lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_2_bufchan_buf[0])))
        lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_2_bufchan_buf <= lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_2_bufchan_d;
  
  /* dcon (Ty TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool,
      Dcon TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool) : [(lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_2_argbuf,Go),
                                                               (lizzieLet0_4QNode_Bool_4QNode_Bool_8QNone_Bool_1_argbuf,Pointer_QTree_Bool),
                                                               (lizzieLet0_4QNode_Bool_4QNode_Bool_11QNone_Bool_1_argbuf,Pointer_QTree_Bool)] > (f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool10,TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool) */
  assign \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool10_d  = TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_dc((& {lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_2_argbuf_d[0],
                                                                                                                                     lizzieLet0_4QNode_Bool_4QNode_Bool_8QNone_Bool_1_argbuf_d[0],
                                                                                                                                     lizzieLet0_4QNode_Bool_4QNode_Bool_11QNone_Bool_1_argbuf_d[0]}), lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_2_argbuf_d, lizzieLet0_4QNode_Bool_4QNode_Bool_8QNone_Bool_1_argbuf_d, lizzieLet0_4QNode_Bool_4QNode_Bool_11QNone_Bool_1_argbuf_d);
  assign {lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_2_argbuf_r,
          lizzieLet0_4QNode_Bool_4QNode_Bool_8QNone_Bool_1_argbuf_r,
          lizzieLet0_4QNode_Bool_4QNode_Bool_11QNone_Bool_1_argbuf_r} = {3 {(\f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool10_r  && \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool10_d [0])}};
  
  /* buf (Ty Go) : (lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_3,Go) > (lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_3_argbuf,Go) */
  Go_t lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_3_bufchan_d;
  logic lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_3_bufchan_r;
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_3_r = ((! lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_3_bufchan_d[0]) || lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_3_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_3_bufchan_d <= 1'd0;
    else
      if (lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_3_r)
        lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_3_bufchan_d <= lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_3_d;
  Go_t lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_3_bufchan_buf;
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_3_bufchan_r = (! lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_3_bufchan_buf[0]);
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_3_argbuf_d = (lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_3_bufchan_buf[0] ? lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_3_bufchan_buf :
                                                                      lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_3_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_3_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_3_argbuf_r && lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_3_bufchan_buf[0]))
        lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_3_bufchan_buf <= 1'd0;
      else if (((! lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_3_argbuf_r) && (! lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_3_bufchan_buf[0])))
        lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_3_bufchan_buf <= lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_3_bufchan_d;
  
  /* dcon (Ty TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool,
      Dcon TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool) : [(lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_3_argbuf,Go),
                                                               (lizzieLet0_4QNode_Bool_4QNode_Bool_7QNone_Bool_1_argbuf,Pointer_QTree_Bool),
                                                               (lizzieLet0_4QNode_Bool_4QNode_Bool_10QNone_Bool_1_argbuf,Pointer_QTree_Bool)] > (f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool11,TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool) */
  assign \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool11_d  = TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_dc((& {lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_3_argbuf_d[0],
                                                                                                                                     lizzieLet0_4QNode_Bool_4QNode_Bool_7QNone_Bool_1_argbuf_d[0],
                                                                                                                                     lizzieLet0_4QNode_Bool_4QNode_Bool_10QNone_Bool_1_argbuf_d[0]}), lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_3_argbuf_d, lizzieLet0_4QNode_Bool_4QNode_Bool_7QNone_Bool_1_argbuf_d, lizzieLet0_4QNode_Bool_4QNode_Bool_10QNone_Bool_1_argbuf_d);
  assign {lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_3_argbuf_r,
          lizzieLet0_4QNode_Bool_4QNode_Bool_7QNone_Bool_1_argbuf_r,
          lizzieLet0_4QNode_Bool_4QNode_Bool_10QNone_Bool_1_argbuf_r} = {3 {(\f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool11_r  && \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool11_d [0])}};
  
  /* buf (Ty Go) : (lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_4,Go) > (lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_4_argbuf,Go) */
  Go_t lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_4_bufchan_d;
  logic lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_4_bufchan_r;
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_4_r = ((! lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_4_bufchan_d[0]) || lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_4_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_4_bufchan_d <= 1'd0;
    else
      if (lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_4_r)
        lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_4_bufchan_d <= lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_4_d;
  Go_t lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_4_bufchan_buf;
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_4_bufchan_r = (! lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_4_bufchan_buf[0]);
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_4_argbuf_d = (lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_4_bufchan_buf[0] ? lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_4_bufchan_buf :
                                                                      lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_4_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_4_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_4_argbuf_r && lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_4_bufchan_buf[0]))
        lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_4_bufchan_buf <= 1'd0;
      else if (((! lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_4_argbuf_r) && (! lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_4_bufchan_buf[0])))
        lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_4_bufchan_buf <= lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_4_bufchan_d;
  
  /* dcon (Ty TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool,
      Dcon TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool) : [(lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_4_argbuf,Go),
                                                               (lizzieLet0_4QNode_Bool_4QNode_Bool_6QNone_Bool_1_argbuf,Pointer_QTree_Bool),
                                                               (lizzieLet0_4QNode_Bool_4QNode_Bool_9QNone_Bool_1_argbuf,Pointer_QTree_Bool)] > (f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool12,TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool) */
  assign \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool12_d  = TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_dc((& {lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_4_argbuf_d[0],
                                                                                                                                     lizzieLet0_4QNode_Bool_4QNode_Bool_6QNone_Bool_1_argbuf_d[0],
                                                                                                                                     lizzieLet0_4QNode_Bool_4QNode_Bool_9QNone_Bool_1_argbuf_d[0]}), lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_4_argbuf_d, lizzieLet0_4QNode_Bool_4QNode_Bool_6QNone_Bool_1_argbuf_d, lizzieLet0_4QNode_Bool_4QNode_Bool_9QNone_Bool_1_argbuf_d);
  assign {lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_4_argbuf_r,
          lizzieLet0_4QNode_Bool_4QNode_Bool_6QNone_Bool_1_argbuf_r,
          lizzieLet0_4QNode_Bool_4QNode_Bool_9QNone_Bool_1_argbuf_r} = {3 {(\f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool12_r  && \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool12_d [0])}};
  
  /* buf (Ty Go) : (lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_5,Go) > (lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_5_argbuf,Go) */
  Go_t lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_5_bufchan_d;
  logic lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_5_bufchan_r;
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_5_r = ((! lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_5_bufchan_d[0]) || lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_5_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_5_bufchan_d <= 1'd0;
    else
      if (lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_5_r)
        lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_5_bufchan_d <= lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_5_d;
  Go_t lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_5_bufchan_buf;
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_5_bufchan_r = (! lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_5_bufchan_buf[0]);
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_5_argbuf_d = (lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_5_bufchan_buf[0] ? lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_5_bufchan_buf :
                                                                      lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_5_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_5_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_5_argbuf_r && lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_5_bufchan_buf[0]))
        lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_5_bufchan_buf <= 1'd0;
      else if (((! lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_5_argbuf_r) && (! lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_5_bufchan_buf[0])))
        lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_5_bufchan_buf <= lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_5_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet0_4QNode_Bool_4QNode_Bool_4QVal_Bool,Go) > [(lizzieLet0_4QNode_Bool_4QNode_Bool_4QVal_Bool_1,Go),
                                                                     (lizzieLet0_4QNode_Bool_4QNode_Bool_4QVal_Bool_2,Go)] */
  logic [1:0] lizzieLet0_4QNode_Bool_4QNode_Bool_4QVal_Bool_emitted;
  logic [1:0] lizzieLet0_4QNode_Bool_4QNode_Bool_4QVal_Bool_done;
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_4QVal_Bool_1_d = (lizzieLet0_4QNode_Bool_4QNode_Bool_4QVal_Bool_d[0] && (! lizzieLet0_4QNode_Bool_4QNode_Bool_4QVal_Bool_emitted[0]));
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_4QVal_Bool_2_d = (lizzieLet0_4QNode_Bool_4QNode_Bool_4QVal_Bool_d[0] && (! lizzieLet0_4QNode_Bool_4QNode_Bool_4QVal_Bool_emitted[1]));
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_4QVal_Bool_done = (lizzieLet0_4QNode_Bool_4QNode_Bool_4QVal_Bool_emitted | ({lizzieLet0_4QNode_Bool_4QNode_Bool_4QVal_Bool_2_d[0],
                                                                                                                         lizzieLet0_4QNode_Bool_4QNode_Bool_4QVal_Bool_1_d[0]} & {lizzieLet0_4QNode_Bool_4QNode_Bool_4QVal_Bool_2_r,
                                                                                                                                                                                  lizzieLet0_4QNode_Bool_4QNode_Bool_4QVal_Bool_1_r}));
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_4QVal_Bool_r = (& lizzieLet0_4QNode_Bool_4QNode_Bool_4QVal_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNode_Bool_4QNode_Bool_4QVal_Bool_emitted <= 2'd0;
    else
      lizzieLet0_4QNode_Bool_4QNode_Bool_4QVal_Bool_emitted <= (lizzieLet0_4QNode_Bool_4QNode_Bool_4QVal_Bool_r ? 2'd0 :
                                                                lizzieLet0_4QNode_Bool_4QNode_Bool_4QVal_Bool_done);
  
  /* dcon (Ty QTree_Bool,
      Dcon QError_Bool) : [(lizzieLet0_4QNode_Bool_4QNode_Bool_4QVal_Bool_1,Go)] > (lizzieLet0_4QNode_Bool_4QNode_Bool_4QVal_Bool_1QError_Bool,QTree_Bool) */
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_4QVal_Bool_1QError_Bool_d = QError_Bool_dc((& {lizzieLet0_4QNode_Bool_4QNode_Bool_4QVal_Bool_1_d[0]}), lizzieLet0_4QNode_Bool_4QNode_Bool_4QVal_Bool_1_d);
  assign {lizzieLet0_4QNode_Bool_4QNode_Bool_4QVal_Bool_1_r} = {1 {(lizzieLet0_4QNode_Bool_4QNode_Bool_4QVal_Bool_1QError_Bool_r && lizzieLet0_4QNode_Bool_4QNode_Bool_4QVal_Bool_1QError_Bool_d[0])}};
  
  /* buf (Ty QTree_Bool) : (lizzieLet0_4QNode_Bool_4QNode_Bool_4QVal_Bool_1QError_Bool,QTree_Bool) > (lizzieLet40_1_argbuf,QTree_Bool) */
  QTree_Bool_t lizzieLet0_4QNode_Bool_4QNode_Bool_4QVal_Bool_1QError_Bool_bufchan_d;
  logic lizzieLet0_4QNode_Bool_4QNode_Bool_4QVal_Bool_1QError_Bool_bufchan_r;
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_4QVal_Bool_1QError_Bool_r = ((! lizzieLet0_4QNode_Bool_4QNode_Bool_4QVal_Bool_1QError_Bool_bufchan_d[0]) || lizzieLet0_4QNode_Bool_4QNode_Bool_4QVal_Bool_1QError_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNode_Bool_4QNode_Bool_4QVal_Bool_1QError_Bool_bufchan_d <= {66'd0,
                                                                               1'd0};
    else
      if (lizzieLet0_4QNode_Bool_4QNode_Bool_4QVal_Bool_1QError_Bool_r)
        lizzieLet0_4QNode_Bool_4QNode_Bool_4QVal_Bool_1QError_Bool_bufchan_d <= lizzieLet0_4QNode_Bool_4QNode_Bool_4QVal_Bool_1QError_Bool_d;
  QTree_Bool_t lizzieLet0_4QNode_Bool_4QNode_Bool_4QVal_Bool_1QError_Bool_bufchan_buf;
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_4QVal_Bool_1QError_Bool_bufchan_r = (! lizzieLet0_4QNode_Bool_4QNode_Bool_4QVal_Bool_1QError_Bool_bufchan_buf[0]);
  assign lizzieLet40_1_argbuf_d = (lizzieLet0_4QNode_Bool_4QNode_Bool_4QVal_Bool_1QError_Bool_bufchan_buf[0] ? lizzieLet0_4QNode_Bool_4QNode_Bool_4QVal_Bool_1QError_Bool_bufchan_buf :
                                   lizzieLet0_4QNode_Bool_4QNode_Bool_4QVal_Bool_1QError_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNode_Bool_4QNode_Bool_4QVal_Bool_1QError_Bool_bufchan_buf <= {66'd0,
                                                                                 1'd0};
    else
      if ((lizzieLet40_1_argbuf_r && lizzieLet0_4QNode_Bool_4QNode_Bool_4QVal_Bool_1QError_Bool_bufchan_buf[0]))
        lizzieLet0_4QNode_Bool_4QNode_Bool_4QVal_Bool_1QError_Bool_bufchan_buf <= {66'd0,
                                                                                   1'd0};
      else if (((! lizzieLet40_1_argbuf_r) && (! lizzieLet0_4QNode_Bool_4QNode_Bool_4QVal_Bool_1QError_Bool_bufchan_buf[0])))
        lizzieLet0_4QNode_Bool_4QNode_Bool_4QVal_Bool_1QError_Bool_bufchan_buf <= lizzieLet0_4QNode_Bool_4QNode_Bool_4QVal_Bool_1QError_Bool_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet0_4QNode_Bool_4QNode_Bool_4QVal_Bool_2,Go) > (lizzieLet0_4QNode_Bool_4QNode_Bool_4QVal_Bool_2_argbuf,Go) */
  Go_t lizzieLet0_4QNode_Bool_4QNode_Bool_4QVal_Bool_2_bufchan_d;
  logic lizzieLet0_4QNode_Bool_4QNode_Bool_4QVal_Bool_2_bufchan_r;
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_4QVal_Bool_2_r = ((! lizzieLet0_4QNode_Bool_4QNode_Bool_4QVal_Bool_2_bufchan_d[0]) || lizzieLet0_4QNode_Bool_4QNode_Bool_4QVal_Bool_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNode_Bool_4QNode_Bool_4QVal_Bool_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet0_4QNode_Bool_4QNode_Bool_4QVal_Bool_2_r)
        lizzieLet0_4QNode_Bool_4QNode_Bool_4QVal_Bool_2_bufchan_d <= lizzieLet0_4QNode_Bool_4QNode_Bool_4QVal_Bool_2_d;
  Go_t lizzieLet0_4QNode_Bool_4QNode_Bool_4QVal_Bool_2_bufchan_buf;
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_4QVal_Bool_2_bufchan_r = (! lizzieLet0_4QNode_Bool_4QNode_Bool_4QVal_Bool_2_bufchan_buf[0]);
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_4QVal_Bool_2_argbuf_d = (lizzieLet0_4QNode_Bool_4QNode_Bool_4QVal_Bool_2_bufchan_buf[0] ? lizzieLet0_4QNode_Bool_4QNode_Bool_4QVal_Bool_2_bufchan_buf :
                                                                     lizzieLet0_4QNode_Bool_4QNode_Bool_4QVal_Bool_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNode_Bool_4QNode_Bool_4QVal_Bool_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet0_4QNode_Bool_4QNode_Bool_4QVal_Bool_2_argbuf_r && lizzieLet0_4QNode_Bool_4QNode_Bool_4QVal_Bool_2_bufchan_buf[0]))
        lizzieLet0_4QNode_Bool_4QNode_Bool_4QVal_Bool_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet0_4QNode_Bool_4QNode_Bool_4QVal_Bool_2_argbuf_r) && (! lizzieLet0_4QNode_Bool_4QNode_Bool_4QVal_Bool_2_bufchan_buf[0])))
        lizzieLet0_4QNode_Bool_4QNode_Bool_4QVal_Bool_2_bufchan_buf <= lizzieLet0_4QNode_Bool_4QNode_Bool_4QVal_Bool_2_bufchan_d;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_CTf) : (lizzieLet0_4QNode_Bool_4QNode_Bool_5,QTree_Bool) (lizzieLet0_4QNode_Bool_6QNode_Bool,Pointer_CTf) > [(lizzieLet0_4QNode_Bool_4QNode_Bool_5QNone_Bool,Pointer_CTf),
                                                                                                                               (lizzieLet0_4QNode_Bool_4QNode_Bool_5QVal_Bool,Pointer_CTf),
                                                                                                                               (lizzieLet0_4QNode_Bool_4QNode_Bool_5QNode_Bool,Pointer_CTf),
                                                                                                                               (lizzieLet0_4QNode_Bool_4QNode_Bool_5QError_Bool,Pointer_CTf)] */
  logic [3:0] lizzieLet0_4QNode_Bool_6QNode_Bool_onehotd;
  always_comb
    if ((lizzieLet0_4QNode_Bool_4QNode_Bool_5_d[0] && lizzieLet0_4QNode_Bool_6QNode_Bool_d[0]))
      unique case (lizzieLet0_4QNode_Bool_4QNode_Bool_5_d[2:1])
        2'd0: lizzieLet0_4QNode_Bool_6QNode_Bool_onehotd = 4'd1;
        2'd1: lizzieLet0_4QNode_Bool_6QNode_Bool_onehotd = 4'd2;
        2'd2: lizzieLet0_4QNode_Bool_6QNode_Bool_onehotd = 4'd4;
        2'd3: lizzieLet0_4QNode_Bool_6QNode_Bool_onehotd = 4'd8;
        default: lizzieLet0_4QNode_Bool_6QNode_Bool_onehotd = 4'd0;
      endcase
    else lizzieLet0_4QNode_Bool_6QNode_Bool_onehotd = 4'd0;
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_5QNone_Bool_d = {lizzieLet0_4QNode_Bool_6QNode_Bool_d[16:1],
                                                             lizzieLet0_4QNode_Bool_6QNode_Bool_onehotd[0]};
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_5QVal_Bool_d = {lizzieLet0_4QNode_Bool_6QNode_Bool_d[16:1],
                                                            lizzieLet0_4QNode_Bool_6QNode_Bool_onehotd[1]};
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_5QNode_Bool_d = {lizzieLet0_4QNode_Bool_6QNode_Bool_d[16:1],
                                                             lizzieLet0_4QNode_Bool_6QNode_Bool_onehotd[2]};
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_5QError_Bool_d = {lizzieLet0_4QNode_Bool_6QNode_Bool_d[16:1],
                                                              lizzieLet0_4QNode_Bool_6QNode_Bool_onehotd[3]};
  assign lizzieLet0_4QNode_Bool_6QNode_Bool_r = (| (lizzieLet0_4QNode_Bool_6QNode_Bool_onehotd & {lizzieLet0_4QNode_Bool_4QNode_Bool_5QError_Bool_r,
                                                                                                  lizzieLet0_4QNode_Bool_4QNode_Bool_5QNode_Bool_r,
                                                                                                  lizzieLet0_4QNode_Bool_4QNode_Bool_5QVal_Bool_r,
                                                                                                  lizzieLet0_4QNode_Bool_4QNode_Bool_5QNone_Bool_r}));
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_5_r = lizzieLet0_4QNode_Bool_6QNode_Bool_r;
  
  /* buf (Ty Pointer_CTf) : (lizzieLet0_4QNode_Bool_4QNode_Bool_5QError_Bool,Pointer_CTf) > (lizzieLet0_4QNode_Bool_4QNode_Bool_5QError_Bool_1_argbuf,Pointer_CTf) */
  Pointer_CTf_t lizzieLet0_4QNode_Bool_4QNode_Bool_5QError_Bool_bufchan_d;
  logic lizzieLet0_4QNode_Bool_4QNode_Bool_5QError_Bool_bufchan_r;
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_5QError_Bool_r = ((! lizzieLet0_4QNode_Bool_4QNode_Bool_5QError_Bool_bufchan_d[0]) || lizzieLet0_4QNode_Bool_4QNode_Bool_5QError_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNode_Bool_4QNode_Bool_5QError_Bool_bufchan_d <= {16'd0,
                                                                    1'd0};
    else
      if (lizzieLet0_4QNode_Bool_4QNode_Bool_5QError_Bool_r)
        lizzieLet0_4QNode_Bool_4QNode_Bool_5QError_Bool_bufchan_d <= lizzieLet0_4QNode_Bool_4QNode_Bool_5QError_Bool_d;
  Pointer_CTf_t lizzieLet0_4QNode_Bool_4QNode_Bool_5QError_Bool_bufchan_buf;
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_5QError_Bool_bufchan_r = (! lizzieLet0_4QNode_Bool_4QNode_Bool_5QError_Bool_bufchan_buf[0]);
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_5QError_Bool_1_argbuf_d = (lizzieLet0_4QNode_Bool_4QNode_Bool_5QError_Bool_bufchan_buf[0] ? lizzieLet0_4QNode_Bool_4QNode_Bool_5QError_Bool_bufchan_buf :
                                                                       lizzieLet0_4QNode_Bool_4QNode_Bool_5QError_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNode_Bool_4QNode_Bool_5QError_Bool_bufchan_buf <= {16'd0,
                                                                      1'd0};
    else
      if ((lizzieLet0_4QNode_Bool_4QNode_Bool_5QError_Bool_1_argbuf_r && lizzieLet0_4QNode_Bool_4QNode_Bool_5QError_Bool_bufchan_buf[0]))
        lizzieLet0_4QNode_Bool_4QNode_Bool_5QError_Bool_bufchan_buf <= {16'd0,
                                                                        1'd0};
      else if (((! lizzieLet0_4QNode_Bool_4QNode_Bool_5QError_Bool_1_argbuf_r) && (! lizzieLet0_4QNode_Bool_4QNode_Bool_5QError_Bool_bufchan_buf[0])))
        lizzieLet0_4QNode_Bool_4QNode_Bool_5QError_Bool_bufchan_buf <= lizzieLet0_4QNode_Bool_4QNode_Bool_5QError_Bool_bufchan_d;
  
  /* dcon (Ty CTf,
      Dcon Lcall_f3) : [(lizzieLet0_4QNode_Bool_4QNode_Bool_5QNode_Bool,Pointer_CTf),
                        (lizzieLet0_4QNode_Bool_4QNode_Bool_6QNode_Bool,Pointer_QTree_Bool),
                        (lizzieLet0_4QNode_Bool_4QNode_Bool_9QNode_Bool,Pointer_QTree_Bool),
                        (t1'a8W_destruct,Pointer_QTree_Bool),
                        (lizzieLet0_4QNode_Bool_4QNode_Bool_7QNode_Bool,Pointer_QTree_Bool),
                        (lizzieLet0_4QNode_Bool_4QNode_Bool_10QNode_Bool,Pointer_QTree_Bool),
                        (t2'a8X_destruct,Pointer_QTree_Bool),
                        (lizzieLet0_4QNode_Bool_4QNode_Bool_8QNode_Bool,Pointer_QTree_Bool),
                        (lizzieLet0_4QNode_Bool_4QNode_Bool_11QNode_Bool,Pointer_QTree_Bool),
                        (t3'a8Y_destruct,Pointer_QTree_Bool)] > (lizzieLet0_4QNode_Bool_4QNode_Bool_5QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_6QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_9QNode_Bool_1t1'a8W_1lizzieLet0_4QNode_Bool_4QNode_Bool_7QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_10QNode_Bool_1t2'a8X_1lizzieLet0_4QNode_Bool_4QNode_Bool_8QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_11QNode_Bool_1t3'a8Y_1Lcall_f3,CTf) */
  assign \lizzieLet0_4QNode_Bool_4QNode_Bool_5QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_6QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_9QNode_Bool_1t1'a8W_1lizzieLet0_4QNode_Bool_4QNode_Bool_7QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_10QNode_Bool_1t2'a8X_1lizzieLet0_4QNode_Bool_4QNode_Bool_8QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_11QNode_Bool_1t3'a8Y_1Lcall_f3_d  = Lcall_f3_dc((& {lizzieLet0_4QNode_Bool_4QNode_Bool_5QNode_Bool_d[0],
                                                                                                                                                                                                                                                                                                                                                                                                                  lizzieLet0_4QNode_Bool_4QNode_Bool_6QNode_Bool_d[0],
                                                                                                                                                                                                                                                                                                                                                                                                                  lizzieLet0_4QNode_Bool_4QNode_Bool_9QNode_Bool_d[0],
                                                                                                                                                                                                                                                                                                                                                                                                                  \t1'a8W_destruct_d [0],
                                                                                                                                                                                                                                                                                                                                                                                                                  lizzieLet0_4QNode_Bool_4QNode_Bool_7QNode_Bool_d[0],
                                                                                                                                                                                                                                                                                                                                                                                                                  lizzieLet0_4QNode_Bool_4QNode_Bool_10QNode_Bool_d[0],
                                                                                                                                                                                                                                                                                                                                                                                                                  \t2'a8X_destruct_d [0],
                                                                                                                                                                                                                                                                                                                                                                                                                  lizzieLet0_4QNode_Bool_4QNode_Bool_8QNode_Bool_d[0],
                                                                                                                                                                                                                                                                                                                                                                                                                  lizzieLet0_4QNode_Bool_4QNode_Bool_11QNode_Bool_d[0],
                                                                                                                                                                                                                                                                                                                                                                                                                  \t3'a8Y_destruct_d [0]}), lizzieLet0_4QNode_Bool_4QNode_Bool_5QNode_Bool_d, lizzieLet0_4QNode_Bool_4QNode_Bool_6QNode_Bool_d, lizzieLet0_4QNode_Bool_4QNode_Bool_9QNode_Bool_d, \t1'a8W_destruct_d , lizzieLet0_4QNode_Bool_4QNode_Bool_7QNode_Bool_d, lizzieLet0_4QNode_Bool_4QNode_Bool_10QNode_Bool_d, \t2'a8X_destruct_d , lizzieLet0_4QNode_Bool_4QNode_Bool_8QNode_Bool_d, lizzieLet0_4QNode_Bool_4QNode_Bool_11QNode_Bool_d, \t3'a8Y_destruct_d );
  assign {lizzieLet0_4QNode_Bool_4QNode_Bool_5QNode_Bool_r,
          lizzieLet0_4QNode_Bool_4QNode_Bool_6QNode_Bool_r,
          lizzieLet0_4QNode_Bool_4QNode_Bool_9QNode_Bool_r,
          \t1'a8W_destruct_r ,
          lizzieLet0_4QNode_Bool_4QNode_Bool_7QNode_Bool_r,
          lizzieLet0_4QNode_Bool_4QNode_Bool_10QNode_Bool_r,
          \t2'a8X_destruct_r ,
          lizzieLet0_4QNode_Bool_4QNode_Bool_8QNode_Bool_r,
          lizzieLet0_4QNode_Bool_4QNode_Bool_11QNode_Bool_r,
          \t3'a8Y_destruct_r } = {10 {(\lizzieLet0_4QNode_Bool_4QNode_Bool_5QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_6QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_9QNode_Bool_1t1'a8W_1lizzieLet0_4QNode_Bool_4QNode_Bool_7QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_10QNode_Bool_1t2'a8X_1lizzieLet0_4QNode_Bool_4QNode_Bool_8QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_11QNode_Bool_1t3'a8Y_1Lcall_f3_r  && \lizzieLet0_4QNode_Bool_4QNode_Bool_5QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_6QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_9QNode_Bool_1t1'a8W_1lizzieLet0_4QNode_Bool_4QNode_Bool_7QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_10QNode_Bool_1t2'a8X_1lizzieLet0_4QNode_Bool_4QNode_Bool_8QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_11QNode_Bool_1t3'a8Y_1Lcall_f3_d [0])}};
  
  /* buf (Ty CTf) : (lizzieLet0_4QNode_Bool_4QNode_Bool_5QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_6QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_9QNode_Bool_1t1'a8W_1lizzieLet0_4QNode_Bool_4QNode_Bool_7QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_10QNode_Bool_1t2'a8X_1lizzieLet0_4QNode_Bool_4QNode_Bool_8QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_11QNode_Bool_1t3'a8Y_1Lcall_f3,CTf) > (lizzieLet41_1_argbuf,CTf) */
  CTf_t \lizzieLet0_4QNode_Bool_4QNode_Bool_5QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_6QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_9QNode_Bool_1t1'a8W_1lizzieLet0_4QNode_Bool_4QNode_Bool_7QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_10QNode_Bool_1t2'a8X_1lizzieLet0_4QNode_Bool_4QNode_Bool_8QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_11QNode_Bool_1t3'a8Y_1Lcall_f3_bufchan_d ;
  logic \lizzieLet0_4QNode_Bool_4QNode_Bool_5QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_6QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_9QNode_Bool_1t1'a8W_1lizzieLet0_4QNode_Bool_4QNode_Bool_7QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_10QNode_Bool_1t2'a8X_1lizzieLet0_4QNode_Bool_4QNode_Bool_8QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_11QNode_Bool_1t3'a8Y_1Lcall_f3_bufchan_r ;
  assign \lizzieLet0_4QNode_Bool_4QNode_Bool_5QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_6QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_9QNode_Bool_1t1'a8W_1lizzieLet0_4QNode_Bool_4QNode_Bool_7QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_10QNode_Bool_1t2'a8X_1lizzieLet0_4QNode_Bool_4QNode_Bool_8QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_11QNode_Bool_1t3'a8Y_1Lcall_f3_r  = ((! \lizzieLet0_4QNode_Bool_4QNode_Bool_5QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_6QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_9QNode_Bool_1t1'a8W_1lizzieLet0_4QNode_Bool_4QNode_Bool_7QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_10QNode_Bool_1t2'a8X_1lizzieLet0_4QNode_Bool_4QNode_Bool_8QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_11QNode_Bool_1t3'a8Y_1Lcall_f3_bufchan_d [0]) || \lizzieLet0_4QNode_Bool_4QNode_Bool_5QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_6QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_9QNode_Bool_1t1'a8W_1lizzieLet0_4QNode_Bool_4QNode_Bool_7QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_10QNode_Bool_1t2'a8X_1lizzieLet0_4QNode_Bool_4QNode_Bool_8QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_11QNode_Bool_1t3'a8Y_1Lcall_f3_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet0_4QNode_Bool_4QNode_Bool_5QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_6QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_9QNode_Bool_1t1'a8W_1lizzieLet0_4QNode_Bool_4QNode_Bool_7QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_10QNode_Bool_1t2'a8X_1lizzieLet0_4QNode_Bool_4QNode_Bool_8QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_11QNode_Bool_1t3'a8Y_1Lcall_f3_bufchan_d  <= {163'd0,
                                                                                                                                                                                                                                                                                                                                                                                                         1'd0};
    else
      if (\lizzieLet0_4QNode_Bool_4QNode_Bool_5QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_6QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_9QNode_Bool_1t1'a8W_1lizzieLet0_4QNode_Bool_4QNode_Bool_7QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_10QNode_Bool_1t2'a8X_1lizzieLet0_4QNode_Bool_4QNode_Bool_8QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_11QNode_Bool_1t3'a8Y_1Lcall_f3_r )
        \lizzieLet0_4QNode_Bool_4QNode_Bool_5QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_6QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_9QNode_Bool_1t1'a8W_1lizzieLet0_4QNode_Bool_4QNode_Bool_7QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_10QNode_Bool_1t2'a8X_1lizzieLet0_4QNode_Bool_4QNode_Bool_8QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_11QNode_Bool_1t3'a8Y_1Lcall_f3_bufchan_d  <= \lizzieLet0_4QNode_Bool_4QNode_Bool_5QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_6QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_9QNode_Bool_1t1'a8W_1lizzieLet0_4QNode_Bool_4QNode_Bool_7QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_10QNode_Bool_1t2'a8X_1lizzieLet0_4QNode_Bool_4QNode_Bool_8QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_11QNode_Bool_1t3'a8Y_1Lcall_f3_d ;
  CTf_t \lizzieLet0_4QNode_Bool_4QNode_Bool_5QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_6QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_9QNode_Bool_1t1'a8W_1lizzieLet0_4QNode_Bool_4QNode_Bool_7QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_10QNode_Bool_1t2'a8X_1lizzieLet0_4QNode_Bool_4QNode_Bool_8QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_11QNode_Bool_1t3'a8Y_1Lcall_f3_bufchan_buf ;
  assign \lizzieLet0_4QNode_Bool_4QNode_Bool_5QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_6QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_9QNode_Bool_1t1'a8W_1lizzieLet0_4QNode_Bool_4QNode_Bool_7QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_10QNode_Bool_1t2'a8X_1lizzieLet0_4QNode_Bool_4QNode_Bool_8QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_11QNode_Bool_1t3'a8Y_1Lcall_f3_bufchan_r  = (! \lizzieLet0_4QNode_Bool_4QNode_Bool_5QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_6QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_9QNode_Bool_1t1'a8W_1lizzieLet0_4QNode_Bool_4QNode_Bool_7QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_10QNode_Bool_1t2'a8X_1lizzieLet0_4QNode_Bool_4QNode_Bool_8QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_11QNode_Bool_1t3'a8Y_1Lcall_f3_bufchan_buf [0]);
  assign lizzieLet41_1_argbuf_d = (\lizzieLet0_4QNode_Bool_4QNode_Bool_5QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_6QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_9QNode_Bool_1t1'a8W_1lizzieLet0_4QNode_Bool_4QNode_Bool_7QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_10QNode_Bool_1t2'a8X_1lizzieLet0_4QNode_Bool_4QNode_Bool_8QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_11QNode_Bool_1t3'a8Y_1Lcall_f3_bufchan_buf [0] ? \lizzieLet0_4QNode_Bool_4QNode_Bool_5QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_6QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_9QNode_Bool_1t1'a8W_1lizzieLet0_4QNode_Bool_4QNode_Bool_7QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_10QNode_Bool_1t2'a8X_1lizzieLet0_4QNode_Bool_4QNode_Bool_8QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_11QNode_Bool_1t3'a8Y_1Lcall_f3_bufchan_buf  :
                                   \lizzieLet0_4QNode_Bool_4QNode_Bool_5QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_6QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_9QNode_Bool_1t1'a8W_1lizzieLet0_4QNode_Bool_4QNode_Bool_7QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_10QNode_Bool_1t2'a8X_1lizzieLet0_4QNode_Bool_4QNode_Bool_8QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_11QNode_Bool_1t3'a8Y_1Lcall_f3_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet0_4QNode_Bool_4QNode_Bool_5QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_6QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_9QNode_Bool_1t1'a8W_1lizzieLet0_4QNode_Bool_4QNode_Bool_7QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_10QNode_Bool_1t2'a8X_1lizzieLet0_4QNode_Bool_4QNode_Bool_8QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_11QNode_Bool_1t3'a8Y_1Lcall_f3_bufchan_buf  <= {163'd0,
                                                                                                                                                                                                                                                                                                                                                                                                           1'd0};
    else
      if ((lizzieLet41_1_argbuf_r && \lizzieLet0_4QNode_Bool_4QNode_Bool_5QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_6QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_9QNode_Bool_1t1'a8W_1lizzieLet0_4QNode_Bool_4QNode_Bool_7QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_10QNode_Bool_1t2'a8X_1lizzieLet0_4QNode_Bool_4QNode_Bool_8QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_11QNode_Bool_1t3'a8Y_1Lcall_f3_bufchan_buf [0]))
        \lizzieLet0_4QNode_Bool_4QNode_Bool_5QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_6QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_9QNode_Bool_1t1'a8W_1lizzieLet0_4QNode_Bool_4QNode_Bool_7QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_10QNode_Bool_1t2'a8X_1lizzieLet0_4QNode_Bool_4QNode_Bool_8QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_11QNode_Bool_1t3'a8Y_1Lcall_f3_bufchan_buf  <= {163'd0,
                                                                                                                                                                                                                                                                                                                                                                                                             1'd0};
      else if (((! lizzieLet41_1_argbuf_r) && (! \lizzieLet0_4QNode_Bool_4QNode_Bool_5QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_6QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_9QNode_Bool_1t1'a8W_1lizzieLet0_4QNode_Bool_4QNode_Bool_7QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_10QNode_Bool_1t2'a8X_1lizzieLet0_4QNode_Bool_4QNode_Bool_8QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_11QNode_Bool_1t3'a8Y_1Lcall_f3_bufchan_buf [0])))
        \lizzieLet0_4QNode_Bool_4QNode_Bool_5QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_6QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_9QNode_Bool_1t1'a8W_1lizzieLet0_4QNode_Bool_4QNode_Bool_7QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_10QNode_Bool_1t2'a8X_1lizzieLet0_4QNode_Bool_4QNode_Bool_8QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_11QNode_Bool_1t3'a8Y_1Lcall_f3_bufchan_buf  <= \lizzieLet0_4QNode_Bool_4QNode_Bool_5QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_6QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_9QNode_Bool_1t1'a8W_1lizzieLet0_4QNode_Bool_4QNode_Bool_7QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_10QNode_Bool_1t2'a8X_1lizzieLet0_4QNode_Bool_4QNode_Bool_8QNode_Bool_1lizzieLet0_4QNode_Bool_4QNode_Bool_11QNode_Bool_1t3'a8Y_1Lcall_f3_bufchan_d ;
  
  /* buf (Ty Pointer_CTf) : (lizzieLet0_4QNode_Bool_4QNode_Bool_5QNone_Bool,Pointer_CTf) > (lizzieLet0_4QNode_Bool_4QNode_Bool_5QNone_Bool_1_argbuf,Pointer_CTf) */
  Pointer_CTf_t lizzieLet0_4QNode_Bool_4QNode_Bool_5QNone_Bool_bufchan_d;
  logic lizzieLet0_4QNode_Bool_4QNode_Bool_5QNone_Bool_bufchan_r;
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_5QNone_Bool_r = ((! lizzieLet0_4QNode_Bool_4QNode_Bool_5QNone_Bool_bufchan_d[0]) || lizzieLet0_4QNode_Bool_4QNode_Bool_5QNone_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNode_Bool_4QNode_Bool_5QNone_Bool_bufchan_d <= {16'd0,
                                                                   1'd0};
    else
      if (lizzieLet0_4QNode_Bool_4QNode_Bool_5QNone_Bool_r)
        lizzieLet0_4QNode_Bool_4QNode_Bool_5QNone_Bool_bufchan_d <= lizzieLet0_4QNode_Bool_4QNode_Bool_5QNone_Bool_d;
  Pointer_CTf_t lizzieLet0_4QNode_Bool_4QNode_Bool_5QNone_Bool_bufchan_buf;
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_5QNone_Bool_bufchan_r = (! lizzieLet0_4QNode_Bool_4QNode_Bool_5QNone_Bool_bufchan_buf[0]);
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_5QNone_Bool_1_argbuf_d = (lizzieLet0_4QNode_Bool_4QNode_Bool_5QNone_Bool_bufchan_buf[0] ? lizzieLet0_4QNode_Bool_4QNode_Bool_5QNone_Bool_bufchan_buf :
                                                                      lizzieLet0_4QNode_Bool_4QNode_Bool_5QNone_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNode_Bool_4QNode_Bool_5QNone_Bool_bufchan_buf <= {16'd0,
                                                                     1'd0};
    else
      if ((lizzieLet0_4QNode_Bool_4QNode_Bool_5QNone_Bool_1_argbuf_r && lizzieLet0_4QNode_Bool_4QNode_Bool_5QNone_Bool_bufchan_buf[0]))
        lizzieLet0_4QNode_Bool_4QNode_Bool_5QNone_Bool_bufchan_buf <= {16'd0,
                                                                       1'd0};
      else if (((! lizzieLet0_4QNode_Bool_4QNode_Bool_5QNone_Bool_1_argbuf_r) && (! lizzieLet0_4QNode_Bool_4QNode_Bool_5QNone_Bool_bufchan_buf[0])))
        lizzieLet0_4QNode_Bool_4QNode_Bool_5QNone_Bool_bufchan_buf <= lizzieLet0_4QNode_Bool_4QNode_Bool_5QNone_Bool_bufchan_d;
  
  /* buf (Ty Pointer_CTf) : (lizzieLet0_4QNode_Bool_4QNode_Bool_5QVal_Bool,Pointer_CTf) > (lizzieLet0_4QNode_Bool_4QNode_Bool_5QVal_Bool_1_argbuf,Pointer_CTf) */
  Pointer_CTf_t lizzieLet0_4QNode_Bool_4QNode_Bool_5QVal_Bool_bufchan_d;
  logic lizzieLet0_4QNode_Bool_4QNode_Bool_5QVal_Bool_bufchan_r;
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_5QVal_Bool_r = ((! lizzieLet0_4QNode_Bool_4QNode_Bool_5QVal_Bool_bufchan_d[0]) || lizzieLet0_4QNode_Bool_4QNode_Bool_5QVal_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNode_Bool_4QNode_Bool_5QVal_Bool_bufchan_d <= {16'd0,
                                                                  1'd0};
    else
      if (lizzieLet0_4QNode_Bool_4QNode_Bool_5QVal_Bool_r)
        lizzieLet0_4QNode_Bool_4QNode_Bool_5QVal_Bool_bufchan_d <= lizzieLet0_4QNode_Bool_4QNode_Bool_5QVal_Bool_d;
  Pointer_CTf_t lizzieLet0_4QNode_Bool_4QNode_Bool_5QVal_Bool_bufchan_buf;
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_5QVal_Bool_bufchan_r = (! lizzieLet0_4QNode_Bool_4QNode_Bool_5QVal_Bool_bufchan_buf[0]);
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_5QVal_Bool_1_argbuf_d = (lizzieLet0_4QNode_Bool_4QNode_Bool_5QVal_Bool_bufchan_buf[0] ? lizzieLet0_4QNode_Bool_4QNode_Bool_5QVal_Bool_bufchan_buf :
                                                                     lizzieLet0_4QNode_Bool_4QNode_Bool_5QVal_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNode_Bool_4QNode_Bool_5QVal_Bool_bufchan_buf <= {16'd0,
                                                                    1'd0};
    else
      if ((lizzieLet0_4QNode_Bool_4QNode_Bool_5QVal_Bool_1_argbuf_r && lizzieLet0_4QNode_Bool_4QNode_Bool_5QVal_Bool_bufchan_buf[0]))
        lizzieLet0_4QNode_Bool_4QNode_Bool_5QVal_Bool_bufchan_buf <= {16'd0,
                                                                      1'd0};
      else if (((! lizzieLet0_4QNode_Bool_4QNode_Bool_5QVal_Bool_1_argbuf_r) && (! lizzieLet0_4QNode_Bool_4QNode_Bool_5QVal_Bool_bufchan_buf[0])))
        lizzieLet0_4QNode_Bool_4QNode_Bool_5QVal_Bool_bufchan_buf <= lizzieLet0_4QNode_Bool_4QNode_Bool_5QVal_Bool_bufchan_d;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_QTree_Bool) : (lizzieLet0_4QNode_Bool_4QNode_Bool_6,QTree_Bool) (lizzieLet0_4QNode_Bool_7QNode_Bool,Pointer_QTree_Bool) > [(lizzieLet0_4QNode_Bool_4QNode_Bool_6QNone_Bool,Pointer_QTree_Bool),
                                                                                                                                             (_147,Pointer_QTree_Bool),
                                                                                                                                             (lizzieLet0_4QNode_Bool_4QNode_Bool_6QNode_Bool,Pointer_QTree_Bool),
                                                                                                                                             (_146,Pointer_QTree_Bool)] */
  logic [3:0] lizzieLet0_4QNode_Bool_7QNode_Bool_onehotd;
  always_comb
    if ((lizzieLet0_4QNode_Bool_4QNode_Bool_6_d[0] && lizzieLet0_4QNode_Bool_7QNode_Bool_d[0]))
      unique case (lizzieLet0_4QNode_Bool_4QNode_Bool_6_d[2:1])
        2'd0: lizzieLet0_4QNode_Bool_7QNode_Bool_onehotd = 4'd1;
        2'd1: lizzieLet0_4QNode_Bool_7QNode_Bool_onehotd = 4'd2;
        2'd2: lizzieLet0_4QNode_Bool_7QNode_Bool_onehotd = 4'd4;
        2'd3: lizzieLet0_4QNode_Bool_7QNode_Bool_onehotd = 4'd8;
        default: lizzieLet0_4QNode_Bool_7QNode_Bool_onehotd = 4'd0;
      endcase
    else lizzieLet0_4QNode_Bool_7QNode_Bool_onehotd = 4'd0;
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_6QNone_Bool_d = {lizzieLet0_4QNode_Bool_7QNode_Bool_d[16:1],
                                                             lizzieLet0_4QNode_Bool_7QNode_Bool_onehotd[0]};
  assign _147_d = {lizzieLet0_4QNode_Bool_7QNode_Bool_d[16:1],
                   lizzieLet0_4QNode_Bool_7QNode_Bool_onehotd[1]};
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_6QNode_Bool_d = {lizzieLet0_4QNode_Bool_7QNode_Bool_d[16:1],
                                                             lizzieLet0_4QNode_Bool_7QNode_Bool_onehotd[2]};
  assign _146_d = {lizzieLet0_4QNode_Bool_7QNode_Bool_d[16:1],
                   lizzieLet0_4QNode_Bool_7QNode_Bool_onehotd[3]};
  assign lizzieLet0_4QNode_Bool_7QNode_Bool_r = (| (lizzieLet0_4QNode_Bool_7QNode_Bool_onehotd & {_146_r,
                                                                                                  lizzieLet0_4QNode_Bool_4QNode_Bool_6QNode_Bool_r,
                                                                                                  _147_r,
                                                                                                  lizzieLet0_4QNode_Bool_4QNode_Bool_6QNone_Bool_r}));
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_6_r = lizzieLet0_4QNode_Bool_7QNode_Bool_r;
  
  /* buf (Ty Pointer_QTree_Bool) : (lizzieLet0_4QNode_Bool_4QNode_Bool_6QNone_Bool,Pointer_QTree_Bool) > (lizzieLet0_4QNode_Bool_4QNode_Bool_6QNone_Bool_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t lizzieLet0_4QNode_Bool_4QNode_Bool_6QNone_Bool_bufchan_d;
  logic lizzieLet0_4QNode_Bool_4QNode_Bool_6QNone_Bool_bufchan_r;
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_6QNone_Bool_r = ((! lizzieLet0_4QNode_Bool_4QNode_Bool_6QNone_Bool_bufchan_d[0]) || lizzieLet0_4QNode_Bool_4QNode_Bool_6QNone_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNode_Bool_4QNode_Bool_6QNone_Bool_bufchan_d <= {16'd0,
                                                                   1'd0};
    else
      if (lizzieLet0_4QNode_Bool_4QNode_Bool_6QNone_Bool_r)
        lizzieLet0_4QNode_Bool_4QNode_Bool_6QNone_Bool_bufchan_d <= lizzieLet0_4QNode_Bool_4QNode_Bool_6QNone_Bool_d;
  Pointer_QTree_Bool_t lizzieLet0_4QNode_Bool_4QNode_Bool_6QNone_Bool_bufchan_buf;
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_6QNone_Bool_bufchan_r = (! lizzieLet0_4QNode_Bool_4QNode_Bool_6QNone_Bool_bufchan_buf[0]);
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_6QNone_Bool_1_argbuf_d = (lizzieLet0_4QNode_Bool_4QNode_Bool_6QNone_Bool_bufchan_buf[0] ? lizzieLet0_4QNode_Bool_4QNode_Bool_6QNone_Bool_bufchan_buf :
                                                                      lizzieLet0_4QNode_Bool_4QNode_Bool_6QNone_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNode_Bool_4QNode_Bool_6QNone_Bool_bufchan_buf <= {16'd0,
                                                                     1'd0};
    else
      if ((lizzieLet0_4QNode_Bool_4QNode_Bool_6QNone_Bool_1_argbuf_r && lizzieLet0_4QNode_Bool_4QNode_Bool_6QNone_Bool_bufchan_buf[0]))
        lizzieLet0_4QNode_Bool_4QNode_Bool_6QNone_Bool_bufchan_buf <= {16'd0,
                                                                       1'd0};
      else if (((! lizzieLet0_4QNode_Bool_4QNode_Bool_6QNone_Bool_1_argbuf_r) && (! lizzieLet0_4QNode_Bool_4QNode_Bool_6QNone_Bool_bufchan_buf[0])))
        lizzieLet0_4QNode_Bool_4QNode_Bool_6QNone_Bool_bufchan_buf <= lizzieLet0_4QNode_Bool_4QNode_Bool_6QNone_Bool_bufchan_d;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_QTree_Bool) : (lizzieLet0_4QNode_Bool_4QNode_Bool_7,QTree_Bool) (lizzieLet0_4QNode_Bool_8QNode_Bool,Pointer_QTree_Bool) > [(lizzieLet0_4QNode_Bool_4QNode_Bool_7QNone_Bool,Pointer_QTree_Bool),
                                                                                                                                             (_145,Pointer_QTree_Bool),
                                                                                                                                             (lizzieLet0_4QNode_Bool_4QNode_Bool_7QNode_Bool,Pointer_QTree_Bool),
                                                                                                                                             (_144,Pointer_QTree_Bool)] */
  logic [3:0] lizzieLet0_4QNode_Bool_8QNode_Bool_onehotd;
  always_comb
    if ((lizzieLet0_4QNode_Bool_4QNode_Bool_7_d[0] && lizzieLet0_4QNode_Bool_8QNode_Bool_d[0]))
      unique case (lizzieLet0_4QNode_Bool_4QNode_Bool_7_d[2:1])
        2'd0: lizzieLet0_4QNode_Bool_8QNode_Bool_onehotd = 4'd1;
        2'd1: lizzieLet0_4QNode_Bool_8QNode_Bool_onehotd = 4'd2;
        2'd2: lizzieLet0_4QNode_Bool_8QNode_Bool_onehotd = 4'd4;
        2'd3: lizzieLet0_4QNode_Bool_8QNode_Bool_onehotd = 4'd8;
        default: lizzieLet0_4QNode_Bool_8QNode_Bool_onehotd = 4'd0;
      endcase
    else lizzieLet0_4QNode_Bool_8QNode_Bool_onehotd = 4'd0;
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_7QNone_Bool_d = {lizzieLet0_4QNode_Bool_8QNode_Bool_d[16:1],
                                                             lizzieLet0_4QNode_Bool_8QNode_Bool_onehotd[0]};
  assign _145_d = {lizzieLet0_4QNode_Bool_8QNode_Bool_d[16:1],
                   lizzieLet0_4QNode_Bool_8QNode_Bool_onehotd[1]};
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_7QNode_Bool_d = {lizzieLet0_4QNode_Bool_8QNode_Bool_d[16:1],
                                                             lizzieLet0_4QNode_Bool_8QNode_Bool_onehotd[2]};
  assign _144_d = {lizzieLet0_4QNode_Bool_8QNode_Bool_d[16:1],
                   lizzieLet0_4QNode_Bool_8QNode_Bool_onehotd[3]};
  assign lizzieLet0_4QNode_Bool_8QNode_Bool_r = (| (lizzieLet0_4QNode_Bool_8QNode_Bool_onehotd & {_144_r,
                                                                                                  lizzieLet0_4QNode_Bool_4QNode_Bool_7QNode_Bool_r,
                                                                                                  _145_r,
                                                                                                  lizzieLet0_4QNode_Bool_4QNode_Bool_7QNone_Bool_r}));
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_7_r = lizzieLet0_4QNode_Bool_8QNode_Bool_r;
  
  /* buf (Ty Pointer_QTree_Bool) : (lizzieLet0_4QNode_Bool_4QNode_Bool_7QNone_Bool,Pointer_QTree_Bool) > (lizzieLet0_4QNode_Bool_4QNode_Bool_7QNone_Bool_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t lizzieLet0_4QNode_Bool_4QNode_Bool_7QNone_Bool_bufchan_d;
  logic lizzieLet0_4QNode_Bool_4QNode_Bool_7QNone_Bool_bufchan_r;
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_7QNone_Bool_r = ((! lizzieLet0_4QNode_Bool_4QNode_Bool_7QNone_Bool_bufchan_d[0]) || lizzieLet0_4QNode_Bool_4QNode_Bool_7QNone_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNode_Bool_4QNode_Bool_7QNone_Bool_bufchan_d <= {16'd0,
                                                                   1'd0};
    else
      if (lizzieLet0_4QNode_Bool_4QNode_Bool_7QNone_Bool_r)
        lizzieLet0_4QNode_Bool_4QNode_Bool_7QNone_Bool_bufchan_d <= lizzieLet0_4QNode_Bool_4QNode_Bool_7QNone_Bool_d;
  Pointer_QTree_Bool_t lizzieLet0_4QNode_Bool_4QNode_Bool_7QNone_Bool_bufchan_buf;
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_7QNone_Bool_bufchan_r = (! lizzieLet0_4QNode_Bool_4QNode_Bool_7QNone_Bool_bufchan_buf[0]);
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_7QNone_Bool_1_argbuf_d = (lizzieLet0_4QNode_Bool_4QNode_Bool_7QNone_Bool_bufchan_buf[0] ? lizzieLet0_4QNode_Bool_4QNode_Bool_7QNone_Bool_bufchan_buf :
                                                                      lizzieLet0_4QNode_Bool_4QNode_Bool_7QNone_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNode_Bool_4QNode_Bool_7QNone_Bool_bufchan_buf <= {16'd0,
                                                                     1'd0};
    else
      if ((lizzieLet0_4QNode_Bool_4QNode_Bool_7QNone_Bool_1_argbuf_r && lizzieLet0_4QNode_Bool_4QNode_Bool_7QNone_Bool_bufchan_buf[0]))
        lizzieLet0_4QNode_Bool_4QNode_Bool_7QNone_Bool_bufchan_buf <= {16'd0,
                                                                       1'd0};
      else if (((! lizzieLet0_4QNode_Bool_4QNode_Bool_7QNone_Bool_1_argbuf_r) && (! lizzieLet0_4QNode_Bool_4QNode_Bool_7QNone_Bool_bufchan_buf[0])))
        lizzieLet0_4QNode_Bool_4QNode_Bool_7QNone_Bool_bufchan_buf <= lizzieLet0_4QNode_Bool_4QNode_Bool_7QNone_Bool_bufchan_d;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_QTree_Bool) : (lizzieLet0_4QNode_Bool_4QNode_Bool_8,QTree_Bool) (lizzieLet0_4QNode_Bool_9QNode_Bool,Pointer_QTree_Bool) > [(lizzieLet0_4QNode_Bool_4QNode_Bool_8QNone_Bool,Pointer_QTree_Bool),
                                                                                                                                             (_143,Pointer_QTree_Bool),
                                                                                                                                             (lizzieLet0_4QNode_Bool_4QNode_Bool_8QNode_Bool,Pointer_QTree_Bool),
                                                                                                                                             (_142,Pointer_QTree_Bool)] */
  logic [3:0] lizzieLet0_4QNode_Bool_9QNode_Bool_onehotd;
  always_comb
    if ((lizzieLet0_4QNode_Bool_4QNode_Bool_8_d[0] && lizzieLet0_4QNode_Bool_9QNode_Bool_d[0]))
      unique case (lizzieLet0_4QNode_Bool_4QNode_Bool_8_d[2:1])
        2'd0: lizzieLet0_4QNode_Bool_9QNode_Bool_onehotd = 4'd1;
        2'd1: lizzieLet0_4QNode_Bool_9QNode_Bool_onehotd = 4'd2;
        2'd2: lizzieLet0_4QNode_Bool_9QNode_Bool_onehotd = 4'd4;
        2'd3: lizzieLet0_4QNode_Bool_9QNode_Bool_onehotd = 4'd8;
        default: lizzieLet0_4QNode_Bool_9QNode_Bool_onehotd = 4'd0;
      endcase
    else lizzieLet0_4QNode_Bool_9QNode_Bool_onehotd = 4'd0;
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_8QNone_Bool_d = {lizzieLet0_4QNode_Bool_9QNode_Bool_d[16:1],
                                                             lizzieLet0_4QNode_Bool_9QNode_Bool_onehotd[0]};
  assign _143_d = {lizzieLet0_4QNode_Bool_9QNode_Bool_d[16:1],
                   lizzieLet0_4QNode_Bool_9QNode_Bool_onehotd[1]};
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_8QNode_Bool_d = {lizzieLet0_4QNode_Bool_9QNode_Bool_d[16:1],
                                                             lizzieLet0_4QNode_Bool_9QNode_Bool_onehotd[2]};
  assign _142_d = {lizzieLet0_4QNode_Bool_9QNode_Bool_d[16:1],
                   lizzieLet0_4QNode_Bool_9QNode_Bool_onehotd[3]};
  assign lizzieLet0_4QNode_Bool_9QNode_Bool_r = (| (lizzieLet0_4QNode_Bool_9QNode_Bool_onehotd & {_142_r,
                                                                                                  lizzieLet0_4QNode_Bool_4QNode_Bool_8QNode_Bool_r,
                                                                                                  _143_r,
                                                                                                  lizzieLet0_4QNode_Bool_4QNode_Bool_8QNone_Bool_r}));
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_8_r = lizzieLet0_4QNode_Bool_9QNode_Bool_r;
  
  /* buf (Ty Pointer_QTree_Bool) : (lizzieLet0_4QNode_Bool_4QNode_Bool_8QNone_Bool,Pointer_QTree_Bool) > (lizzieLet0_4QNode_Bool_4QNode_Bool_8QNone_Bool_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t lizzieLet0_4QNode_Bool_4QNode_Bool_8QNone_Bool_bufchan_d;
  logic lizzieLet0_4QNode_Bool_4QNode_Bool_8QNone_Bool_bufchan_r;
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_8QNone_Bool_r = ((! lizzieLet0_4QNode_Bool_4QNode_Bool_8QNone_Bool_bufchan_d[0]) || lizzieLet0_4QNode_Bool_4QNode_Bool_8QNone_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNode_Bool_4QNode_Bool_8QNone_Bool_bufchan_d <= {16'd0,
                                                                   1'd0};
    else
      if (lizzieLet0_4QNode_Bool_4QNode_Bool_8QNone_Bool_r)
        lizzieLet0_4QNode_Bool_4QNode_Bool_8QNone_Bool_bufchan_d <= lizzieLet0_4QNode_Bool_4QNode_Bool_8QNone_Bool_d;
  Pointer_QTree_Bool_t lizzieLet0_4QNode_Bool_4QNode_Bool_8QNone_Bool_bufchan_buf;
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_8QNone_Bool_bufchan_r = (! lizzieLet0_4QNode_Bool_4QNode_Bool_8QNone_Bool_bufchan_buf[0]);
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_8QNone_Bool_1_argbuf_d = (lizzieLet0_4QNode_Bool_4QNode_Bool_8QNone_Bool_bufchan_buf[0] ? lizzieLet0_4QNode_Bool_4QNode_Bool_8QNone_Bool_bufchan_buf :
                                                                      lizzieLet0_4QNode_Bool_4QNode_Bool_8QNone_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNode_Bool_4QNode_Bool_8QNone_Bool_bufchan_buf <= {16'd0,
                                                                     1'd0};
    else
      if ((lizzieLet0_4QNode_Bool_4QNode_Bool_8QNone_Bool_1_argbuf_r && lizzieLet0_4QNode_Bool_4QNode_Bool_8QNone_Bool_bufchan_buf[0]))
        lizzieLet0_4QNode_Bool_4QNode_Bool_8QNone_Bool_bufchan_buf <= {16'd0,
                                                                       1'd0};
      else if (((! lizzieLet0_4QNode_Bool_4QNode_Bool_8QNone_Bool_1_argbuf_r) && (! lizzieLet0_4QNode_Bool_4QNode_Bool_8QNone_Bool_bufchan_buf[0])))
        lizzieLet0_4QNode_Bool_4QNode_Bool_8QNone_Bool_bufchan_buf <= lizzieLet0_4QNode_Bool_4QNode_Bool_8QNone_Bool_bufchan_d;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_QTree_Bool) : (lizzieLet0_4QNode_Bool_4QNode_Bool_9,QTree_Bool) (t1a8R_destruct,Pointer_QTree_Bool) > [(lizzieLet0_4QNode_Bool_4QNode_Bool_9QNone_Bool,Pointer_QTree_Bool),
                                                                                                                         (_141,Pointer_QTree_Bool),
                                                                                                                         (lizzieLet0_4QNode_Bool_4QNode_Bool_9QNode_Bool,Pointer_QTree_Bool),
                                                                                                                         (_140,Pointer_QTree_Bool)] */
  logic [3:0] t1a8R_destruct_onehotd;
  always_comb
    if ((lizzieLet0_4QNode_Bool_4QNode_Bool_9_d[0] && t1a8R_destruct_d[0]))
      unique case (lizzieLet0_4QNode_Bool_4QNode_Bool_9_d[2:1])
        2'd0: t1a8R_destruct_onehotd = 4'd1;
        2'd1: t1a8R_destruct_onehotd = 4'd2;
        2'd2: t1a8R_destruct_onehotd = 4'd4;
        2'd3: t1a8R_destruct_onehotd = 4'd8;
        default: t1a8R_destruct_onehotd = 4'd0;
      endcase
    else t1a8R_destruct_onehotd = 4'd0;
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_9QNone_Bool_d = {t1a8R_destruct_d[16:1],
                                                             t1a8R_destruct_onehotd[0]};
  assign _141_d = {t1a8R_destruct_d[16:1],
                   t1a8R_destruct_onehotd[1]};
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_9QNode_Bool_d = {t1a8R_destruct_d[16:1],
                                                             t1a8R_destruct_onehotd[2]};
  assign _140_d = {t1a8R_destruct_d[16:1],
                   t1a8R_destruct_onehotd[3]};
  assign t1a8R_destruct_r = (| (t1a8R_destruct_onehotd & {_140_r,
                                                          lizzieLet0_4QNode_Bool_4QNode_Bool_9QNode_Bool_r,
                                                          _141_r,
                                                          lizzieLet0_4QNode_Bool_4QNode_Bool_9QNone_Bool_r}));
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_9_r = t1a8R_destruct_r;
  
  /* buf (Ty Pointer_QTree_Bool) : (lizzieLet0_4QNode_Bool_4QNode_Bool_9QNone_Bool,Pointer_QTree_Bool) > (lizzieLet0_4QNode_Bool_4QNode_Bool_9QNone_Bool_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t lizzieLet0_4QNode_Bool_4QNode_Bool_9QNone_Bool_bufchan_d;
  logic lizzieLet0_4QNode_Bool_4QNode_Bool_9QNone_Bool_bufchan_r;
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_9QNone_Bool_r = ((! lizzieLet0_4QNode_Bool_4QNode_Bool_9QNone_Bool_bufchan_d[0]) || lizzieLet0_4QNode_Bool_4QNode_Bool_9QNone_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNode_Bool_4QNode_Bool_9QNone_Bool_bufchan_d <= {16'd0,
                                                                   1'd0};
    else
      if (lizzieLet0_4QNode_Bool_4QNode_Bool_9QNone_Bool_r)
        lizzieLet0_4QNode_Bool_4QNode_Bool_9QNone_Bool_bufchan_d <= lizzieLet0_4QNode_Bool_4QNode_Bool_9QNone_Bool_d;
  Pointer_QTree_Bool_t lizzieLet0_4QNode_Bool_4QNode_Bool_9QNone_Bool_bufchan_buf;
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_9QNone_Bool_bufchan_r = (! lizzieLet0_4QNode_Bool_4QNode_Bool_9QNone_Bool_bufchan_buf[0]);
  assign lizzieLet0_4QNode_Bool_4QNode_Bool_9QNone_Bool_1_argbuf_d = (lizzieLet0_4QNode_Bool_4QNode_Bool_9QNone_Bool_bufchan_buf[0] ? lizzieLet0_4QNode_Bool_4QNode_Bool_9QNone_Bool_bufchan_buf :
                                                                      lizzieLet0_4QNode_Bool_4QNode_Bool_9QNone_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNode_Bool_4QNode_Bool_9QNone_Bool_bufchan_buf <= {16'd0,
                                                                     1'd0};
    else
      if ((lizzieLet0_4QNode_Bool_4QNode_Bool_9QNone_Bool_1_argbuf_r && lizzieLet0_4QNode_Bool_4QNode_Bool_9QNone_Bool_bufchan_buf[0]))
        lizzieLet0_4QNode_Bool_4QNode_Bool_9QNone_Bool_bufchan_buf <= {16'd0,
                                                                       1'd0};
      else if (((! lizzieLet0_4QNode_Bool_4QNode_Bool_9QNone_Bool_1_argbuf_r) && (! lizzieLet0_4QNode_Bool_4QNode_Bool_9QNone_Bool_bufchan_buf[0])))
        lizzieLet0_4QNode_Bool_4QNode_Bool_9QNone_Bool_bufchan_buf <= lizzieLet0_4QNode_Bool_4QNode_Bool_9QNone_Bool_bufchan_d;
  
  /* fork (Ty QTree_Bool) : (lizzieLet0_4QNode_Bool_4QNone_Bool,QTree_Bool) > [(lizzieLet0_4QNode_Bool_4QNone_Bool_1,QTree_Bool),
                                                                          (lizzieLet0_4QNode_Bool_4QNone_Bool_2,QTree_Bool),
                                                                          (lizzieLet0_4QNode_Bool_4QNone_Bool_3,QTree_Bool),
                                                                          (lizzieLet0_4QNode_Bool_4QNone_Bool_4,QTree_Bool),
                                                                          (lizzieLet0_4QNode_Bool_4QNone_Bool_5,QTree_Bool),
                                                                          (lizzieLet0_4QNode_Bool_4QNone_Bool_6,QTree_Bool),
                                                                          (lizzieLet0_4QNode_Bool_4QNone_Bool_7,QTree_Bool),
                                                                          (lizzieLet0_4QNode_Bool_4QNone_Bool_8,QTree_Bool),
                                                                          (lizzieLet0_4QNode_Bool_4QNone_Bool_9,QTree_Bool)] */
  logic [8:0] lizzieLet0_4QNode_Bool_4QNone_Bool_emitted;
  logic [8:0] lizzieLet0_4QNode_Bool_4QNone_Bool_done;
  assign lizzieLet0_4QNode_Bool_4QNone_Bool_1_d = {lizzieLet0_4QNode_Bool_4QNone_Bool_d[66:1],
                                                   (lizzieLet0_4QNode_Bool_4QNone_Bool_d[0] && (! lizzieLet0_4QNode_Bool_4QNone_Bool_emitted[0]))};
  assign lizzieLet0_4QNode_Bool_4QNone_Bool_2_d = {lizzieLet0_4QNode_Bool_4QNone_Bool_d[66:1],
                                                   (lizzieLet0_4QNode_Bool_4QNone_Bool_d[0] && (! lizzieLet0_4QNode_Bool_4QNone_Bool_emitted[1]))};
  assign lizzieLet0_4QNode_Bool_4QNone_Bool_3_d = {lizzieLet0_4QNode_Bool_4QNone_Bool_d[66:1],
                                                   (lizzieLet0_4QNode_Bool_4QNone_Bool_d[0] && (! lizzieLet0_4QNode_Bool_4QNone_Bool_emitted[2]))};
  assign lizzieLet0_4QNode_Bool_4QNone_Bool_4_d = {lizzieLet0_4QNode_Bool_4QNone_Bool_d[66:1],
                                                   (lizzieLet0_4QNode_Bool_4QNone_Bool_d[0] && (! lizzieLet0_4QNode_Bool_4QNone_Bool_emitted[3]))};
  assign lizzieLet0_4QNode_Bool_4QNone_Bool_5_d = {lizzieLet0_4QNode_Bool_4QNone_Bool_d[66:1],
                                                   (lizzieLet0_4QNode_Bool_4QNone_Bool_d[0] && (! lizzieLet0_4QNode_Bool_4QNone_Bool_emitted[4]))};
  assign lizzieLet0_4QNode_Bool_4QNone_Bool_6_d = {lizzieLet0_4QNode_Bool_4QNone_Bool_d[66:1],
                                                   (lizzieLet0_4QNode_Bool_4QNone_Bool_d[0] && (! lizzieLet0_4QNode_Bool_4QNone_Bool_emitted[5]))};
  assign lizzieLet0_4QNode_Bool_4QNone_Bool_7_d = {lizzieLet0_4QNode_Bool_4QNone_Bool_d[66:1],
                                                   (lizzieLet0_4QNode_Bool_4QNone_Bool_d[0] && (! lizzieLet0_4QNode_Bool_4QNone_Bool_emitted[6]))};
  assign lizzieLet0_4QNode_Bool_4QNone_Bool_8_d = {lizzieLet0_4QNode_Bool_4QNone_Bool_d[66:1],
                                                   (lizzieLet0_4QNode_Bool_4QNone_Bool_d[0] && (! lizzieLet0_4QNode_Bool_4QNone_Bool_emitted[7]))};
  assign lizzieLet0_4QNode_Bool_4QNone_Bool_9_d = {lizzieLet0_4QNode_Bool_4QNone_Bool_d[66:1],
                                                   (lizzieLet0_4QNode_Bool_4QNone_Bool_d[0] && (! lizzieLet0_4QNode_Bool_4QNone_Bool_emitted[8]))};
  assign lizzieLet0_4QNode_Bool_4QNone_Bool_done = (lizzieLet0_4QNode_Bool_4QNone_Bool_emitted | ({lizzieLet0_4QNode_Bool_4QNone_Bool_9_d[0],
                                                                                                   lizzieLet0_4QNode_Bool_4QNone_Bool_8_d[0],
                                                                                                   lizzieLet0_4QNode_Bool_4QNone_Bool_7_d[0],
                                                                                                   lizzieLet0_4QNode_Bool_4QNone_Bool_6_d[0],
                                                                                                   lizzieLet0_4QNode_Bool_4QNone_Bool_5_d[0],
                                                                                                   lizzieLet0_4QNode_Bool_4QNone_Bool_4_d[0],
                                                                                                   lizzieLet0_4QNode_Bool_4QNone_Bool_3_d[0],
                                                                                                   lizzieLet0_4QNode_Bool_4QNone_Bool_2_d[0],
                                                                                                   lizzieLet0_4QNode_Bool_4QNone_Bool_1_d[0]} & {lizzieLet0_4QNode_Bool_4QNone_Bool_9_r,
                                                                                                                                                 lizzieLet0_4QNode_Bool_4QNone_Bool_8_r,
                                                                                                                                                 lizzieLet0_4QNode_Bool_4QNone_Bool_7_r,
                                                                                                                                                 lizzieLet0_4QNode_Bool_4QNone_Bool_6_r,
                                                                                                                                                 lizzieLet0_4QNode_Bool_4QNone_Bool_5_r,
                                                                                                                                                 lizzieLet0_4QNode_Bool_4QNone_Bool_4_r,
                                                                                                                                                 lizzieLet0_4QNode_Bool_4QNone_Bool_3_r,
                                                                                                                                                 lizzieLet0_4QNode_Bool_4QNone_Bool_2_r,
                                                                                                                                                 lizzieLet0_4QNode_Bool_4QNone_Bool_1_r}));
  assign lizzieLet0_4QNode_Bool_4QNone_Bool_r = (& lizzieLet0_4QNode_Bool_4QNone_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNode_Bool_4QNone_Bool_emitted <= 9'd0;
    else
      lizzieLet0_4QNode_Bool_4QNone_Bool_emitted <= (lizzieLet0_4QNode_Bool_4QNone_Bool_r ? 9'd0 :
                                                     lizzieLet0_4QNode_Bool_4QNone_Bool_done);
  
  /* destruct (Ty QTree_Bool,
          Dcon QNode_Bool) : (lizzieLet0_4QNode_Bool_4QNone_Bool_1QNode_Bool,QTree_Bool) > [(t1a8M_destruct,Pointer_QTree_Bool),
                                                                                            (t2a8N_destruct,Pointer_QTree_Bool),
                                                                                            (t3a8O_destruct,Pointer_QTree_Bool),
                                                                                            (t4a8P_destruct,Pointer_QTree_Bool)] */
  logic [3:0] lizzieLet0_4QNode_Bool_4QNone_Bool_1QNode_Bool_emitted;
  logic [3:0] lizzieLet0_4QNode_Bool_4QNone_Bool_1QNode_Bool_done;
  assign t1a8M_destruct_d = {lizzieLet0_4QNode_Bool_4QNone_Bool_1QNode_Bool_d[18:3],
                             (lizzieLet0_4QNode_Bool_4QNone_Bool_1QNode_Bool_d[0] && (! lizzieLet0_4QNode_Bool_4QNone_Bool_1QNode_Bool_emitted[0]))};
  assign t2a8N_destruct_d = {lizzieLet0_4QNode_Bool_4QNone_Bool_1QNode_Bool_d[34:19],
                             (lizzieLet0_4QNode_Bool_4QNone_Bool_1QNode_Bool_d[0] && (! lizzieLet0_4QNode_Bool_4QNone_Bool_1QNode_Bool_emitted[1]))};
  assign t3a8O_destruct_d = {lizzieLet0_4QNode_Bool_4QNone_Bool_1QNode_Bool_d[50:35],
                             (lizzieLet0_4QNode_Bool_4QNone_Bool_1QNode_Bool_d[0] && (! lizzieLet0_4QNode_Bool_4QNone_Bool_1QNode_Bool_emitted[2]))};
  assign t4a8P_destruct_d = {lizzieLet0_4QNode_Bool_4QNone_Bool_1QNode_Bool_d[66:51],
                             (lizzieLet0_4QNode_Bool_4QNone_Bool_1QNode_Bool_d[0] && (! lizzieLet0_4QNode_Bool_4QNone_Bool_1QNode_Bool_emitted[3]))};
  assign lizzieLet0_4QNode_Bool_4QNone_Bool_1QNode_Bool_done = (lizzieLet0_4QNode_Bool_4QNone_Bool_1QNode_Bool_emitted | ({t4a8P_destruct_d[0],
                                                                                                                           t3a8O_destruct_d[0],
                                                                                                                           t2a8N_destruct_d[0],
                                                                                                                           t1a8M_destruct_d[0]} & {t4a8P_destruct_r,
                                                                                                                                                   t3a8O_destruct_r,
                                                                                                                                                   t2a8N_destruct_r,
                                                                                                                                                   t1a8M_destruct_r}));
  assign lizzieLet0_4QNode_Bool_4QNone_Bool_1QNode_Bool_r = (& lizzieLet0_4QNode_Bool_4QNone_Bool_1QNode_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNode_Bool_4QNone_Bool_1QNode_Bool_emitted <= 4'd0;
    else
      lizzieLet0_4QNode_Bool_4QNone_Bool_1QNode_Bool_emitted <= (lizzieLet0_4QNode_Bool_4QNone_Bool_1QNode_Bool_r ? 4'd0 :
                                                                 lizzieLet0_4QNode_Bool_4QNone_Bool_1QNode_Bool_done);
  
  /* demux (Ty QTree_Bool,
       Ty QTree_Bool) : (lizzieLet0_4QNode_Bool_4QNone_Bool_2,QTree_Bool) (lizzieLet0_4QNode_Bool_4QNone_Bool_1,QTree_Bool) > [(_139,QTree_Bool),
                                                                                                                               (_138,QTree_Bool),
                                                                                                                               (lizzieLet0_4QNode_Bool_4QNone_Bool_1QNode_Bool,QTree_Bool),
                                                                                                                               (_137,QTree_Bool)] */
  logic [3:0] lizzieLet0_4QNode_Bool_4QNone_Bool_1_onehotd;
  always_comb
    if ((lizzieLet0_4QNode_Bool_4QNone_Bool_2_d[0] && lizzieLet0_4QNode_Bool_4QNone_Bool_1_d[0]))
      unique case (lizzieLet0_4QNode_Bool_4QNone_Bool_2_d[2:1])
        2'd0: lizzieLet0_4QNode_Bool_4QNone_Bool_1_onehotd = 4'd1;
        2'd1: lizzieLet0_4QNode_Bool_4QNone_Bool_1_onehotd = 4'd2;
        2'd2: lizzieLet0_4QNode_Bool_4QNone_Bool_1_onehotd = 4'd4;
        2'd3: lizzieLet0_4QNode_Bool_4QNone_Bool_1_onehotd = 4'd8;
        default: lizzieLet0_4QNode_Bool_4QNone_Bool_1_onehotd = 4'd0;
      endcase
    else lizzieLet0_4QNode_Bool_4QNone_Bool_1_onehotd = 4'd0;
  assign _139_d = {lizzieLet0_4QNode_Bool_4QNone_Bool_1_d[66:1],
                   lizzieLet0_4QNode_Bool_4QNone_Bool_1_onehotd[0]};
  assign _138_d = {lizzieLet0_4QNode_Bool_4QNone_Bool_1_d[66:1],
                   lizzieLet0_4QNode_Bool_4QNone_Bool_1_onehotd[1]};
  assign lizzieLet0_4QNode_Bool_4QNone_Bool_1QNode_Bool_d = {lizzieLet0_4QNode_Bool_4QNone_Bool_1_d[66:1],
                                                             lizzieLet0_4QNode_Bool_4QNone_Bool_1_onehotd[2]};
  assign _137_d = {lizzieLet0_4QNode_Bool_4QNone_Bool_1_d[66:1],
                   lizzieLet0_4QNode_Bool_4QNone_Bool_1_onehotd[3]};
  assign lizzieLet0_4QNode_Bool_4QNone_Bool_1_r = (| (lizzieLet0_4QNode_Bool_4QNone_Bool_1_onehotd & {_137_r,
                                                                                                      lizzieLet0_4QNode_Bool_4QNone_Bool_1QNode_Bool_r,
                                                                                                      _138_r,
                                                                                                      _139_r}));
  assign lizzieLet0_4QNode_Bool_4QNone_Bool_2_r = lizzieLet0_4QNode_Bool_4QNone_Bool_1_r;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_QTree_Bool) : (lizzieLet0_4QNode_Bool_4QNone_Bool_3,QTree_Bool) (lizzieLet0_4QNode_Bool_10QNone_Bool,Pointer_QTree_Bool) > [(_136,Pointer_QTree_Bool),
                                                                                                                                              (_135,Pointer_QTree_Bool),
                                                                                                                                              (lizzieLet0_4QNode_Bool_4QNone_Bool_3QNode_Bool,Pointer_QTree_Bool),
                                                                                                                                              (_134,Pointer_QTree_Bool)] */
  logic [3:0] lizzieLet0_4QNode_Bool_10QNone_Bool_onehotd;
  always_comb
    if ((lizzieLet0_4QNode_Bool_4QNone_Bool_3_d[0] && lizzieLet0_4QNode_Bool_10QNone_Bool_d[0]))
      unique case (lizzieLet0_4QNode_Bool_4QNone_Bool_3_d[2:1])
        2'd0: lizzieLet0_4QNode_Bool_10QNone_Bool_onehotd = 4'd1;
        2'd1: lizzieLet0_4QNode_Bool_10QNone_Bool_onehotd = 4'd2;
        2'd2: lizzieLet0_4QNode_Bool_10QNone_Bool_onehotd = 4'd4;
        2'd3: lizzieLet0_4QNode_Bool_10QNone_Bool_onehotd = 4'd8;
        default: lizzieLet0_4QNode_Bool_10QNone_Bool_onehotd = 4'd0;
      endcase
    else lizzieLet0_4QNode_Bool_10QNone_Bool_onehotd = 4'd0;
  assign _136_d = {lizzieLet0_4QNode_Bool_10QNone_Bool_d[16:1],
                   lizzieLet0_4QNode_Bool_10QNone_Bool_onehotd[0]};
  assign _135_d = {lizzieLet0_4QNode_Bool_10QNone_Bool_d[16:1],
                   lizzieLet0_4QNode_Bool_10QNone_Bool_onehotd[1]};
  assign lizzieLet0_4QNode_Bool_4QNone_Bool_3QNode_Bool_d = {lizzieLet0_4QNode_Bool_10QNone_Bool_d[16:1],
                                                             lizzieLet0_4QNode_Bool_10QNone_Bool_onehotd[2]};
  assign _134_d = {lizzieLet0_4QNode_Bool_10QNone_Bool_d[16:1],
                   lizzieLet0_4QNode_Bool_10QNone_Bool_onehotd[3]};
  assign lizzieLet0_4QNode_Bool_10QNone_Bool_r = (| (lizzieLet0_4QNode_Bool_10QNone_Bool_onehotd & {_134_r,
                                                                                                    lizzieLet0_4QNode_Bool_4QNone_Bool_3QNode_Bool_r,
                                                                                                    _135_r,
                                                                                                    _136_r}));
  assign lizzieLet0_4QNode_Bool_4QNone_Bool_3_r = lizzieLet0_4QNode_Bool_10QNone_Bool_r;
  
  /* buf (Ty Pointer_QTree_Bool) : (lizzieLet0_4QNode_Bool_4QNone_Bool_3QNode_Bool,Pointer_QTree_Bool) > (lizzieLet0_4QNode_Bool_4QNone_Bool_3QNode_Bool_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t lizzieLet0_4QNode_Bool_4QNone_Bool_3QNode_Bool_bufchan_d;
  logic lizzieLet0_4QNode_Bool_4QNone_Bool_3QNode_Bool_bufchan_r;
  assign lizzieLet0_4QNode_Bool_4QNone_Bool_3QNode_Bool_r = ((! lizzieLet0_4QNode_Bool_4QNone_Bool_3QNode_Bool_bufchan_d[0]) || lizzieLet0_4QNode_Bool_4QNone_Bool_3QNode_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNode_Bool_4QNone_Bool_3QNode_Bool_bufchan_d <= {16'd0,
                                                                   1'd0};
    else
      if (lizzieLet0_4QNode_Bool_4QNone_Bool_3QNode_Bool_r)
        lizzieLet0_4QNode_Bool_4QNone_Bool_3QNode_Bool_bufchan_d <= lizzieLet0_4QNode_Bool_4QNone_Bool_3QNode_Bool_d;
  Pointer_QTree_Bool_t lizzieLet0_4QNode_Bool_4QNone_Bool_3QNode_Bool_bufchan_buf;
  assign lizzieLet0_4QNode_Bool_4QNone_Bool_3QNode_Bool_bufchan_r = (! lizzieLet0_4QNode_Bool_4QNone_Bool_3QNode_Bool_bufchan_buf[0]);
  assign lizzieLet0_4QNode_Bool_4QNone_Bool_3QNode_Bool_1_argbuf_d = (lizzieLet0_4QNode_Bool_4QNone_Bool_3QNode_Bool_bufchan_buf[0] ? lizzieLet0_4QNode_Bool_4QNone_Bool_3QNode_Bool_bufchan_buf :
                                                                      lizzieLet0_4QNode_Bool_4QNone_Bool_3QNode_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNode_Bool_4QNone_Bool_3QNode_Bool_bufchan_buf <= {16'd0,
                                                                     1'd0};
    else
      if ((lizzieLet0_4QNode_Bool_4QNone_Bool_3QNode_Bool_1_argbuf_r && lizzieLet0_4QNode_Bool_4QNone_Bool_3QNode_Bool_bufchan_buf[0]))
        lizzieLet0_4QNode_Bool_4QNone_Bool_3QNode_Bool_bufchan_buf <= {16'd0,
                                                                       1'd0};
      else if (((! lizzieLet0_4QNode_Bool_4QNone_Bool_3QNode_Bool_1_argbuf_r) && (! lizzieLet0_4QNode_Bool_4QNone_Bool_3QNode_Bool_bufchan_buf[0])))
        lizzieLet0_4QNode_Bool_4QNone_Bool_3QNode_Bool_bufchan_buf <= lizzieLet0_4QNode_Bool_4QNone_Bool_3QNode_Bool_bufchan_d;
  
  /* demux (Ty QTree_Bool,
       Ty Go) : (lizzieLet0_4QNode_Bool_4QNone_Bool_4,QTree_Bool) (lizzieLet0_4QNode_Bool_3QNone_Bool,Go) > [(lizzieLet0_4QNode_Bool_4QNone_Bool_4QNone_Bool,Go),
                                                                                                             (lizzieLet0_4QNode_Bool_4QNone_Bool_4QVal_Bool,Go),
                                                                                                             (lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool,Go),
                                                                                                             (lizzieLet0_4QNode_Bool_4QNone_Bool_4QError_Bool,Go)] */
  logic [3:0] lizzieLet0_4QNode_Bool_3QNone_Bool_onehotd;
  always_comb
    if ((lizzieLet0_4QNode_Bool_4QNone_Bool_4_d[0] && lizzieLet0_4QNode_Bool_3QNone_Bool_d[0]))
      unique case (lizzieLet0_4QNode_Bool_4QNone_Bool_4_d[2:1])
        2'd0: lizzieLet0_4QNode_Bool_3QNone_Bool_onehotd = 4'd1;
        2'd1: lizzieLet0_4QNode_Bool_3QNone_Bool_onehotd = 4'd2;
        2'd2: lizzieLet0_4QNode_Bool_3QNone_Bool_onehotd = 4'd4;
        2'd3: lizzieLet0_4QNode_Bool_3QNone_Bool_onehotd = 4'd8;
        default: lizzieLet0_4QNode_Bool_3QNone_Bool_onehotd = 4'd0;
      endcase
    else lizzieLet0_4QNode_Bool_3QNone_Bool_onehotd = 4'd0;
  assign lizzieLet0_4QNode_Bool_4QNone_Bool_4QNone_Bool_d = lizzieLet0_4QNode_Bool_3QNone_Bool_onehotd[0];
  assign lizzieLet0_4QNode_Bool_4QNone_Bool_4QVal_Bool_d = lizzieLet0_4QNode_Bool_3QNone_Bool_onehotd[1];
  assign lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_d = lizzieLet0_4QNode_Bool_3QNone_Bool_onehotd[2];
  assign lizzieLet0_4QNode_Bool_4QNone_Bool_4QError_Bool_d = lizzieLet0_4QNode_Bool_3QNone_Bool_onehotd[3];
  assign lizzieLet0_4QNode_Bool_3QNone_Bool_r = (| (lizzieLet0_4QNode_Bool_3QNone_Bool_onehotd & {lizzieLet0_4QNode_Bool_4QNone_Bool_4QError_Bool_r,
                                                                                                  lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_r,
                                                                                                  lizzieLet0_4QNode_Bool_4QNone_Bool_4QVal_Bool_r,
                                                                                                  lizzieLet0_4QNode_Bool_4QNone_Bool_4QNone_Bool_r}));
  assign lizzieLet0_4QNode_Bool_4QNone_Bool_4_r = lizzieLet0_4QNode_Bool_3QNone_Bool_r;
  
  /* fork (Ty Go) : (lizzieLet0_4QNode_Bool_4QNone_Bool_4QError_Bool,Go) > [(lizzieLet0_4QNode_Bool_4QNone_Bool_4QError_Bool_1,Go),
                                                                       (lizzieLet0_4QNode_Bool_4QNone_Bool_4QError_Bool_2,Go)] */
  logic [1:0] lizzieLet0_4QNode_Bool_4QNone_Bool_4QError_Bool_emitted;
  logic [1:0] lizzieLet0_4QNode_Bool_4QNone_Bool_4QError_Bool_done;
  assign lizzieLet0_4QNode_Bool_4QNone_Bool_4QError_Bool_1_d = (lizzieLet0_4QNode_Bool_4QNone_Bool_4QError_Bool_d[0] && (! lizzieLet0_4QNode_Bool_4QNone_Bool_4QError_Bool_emitted[0]));
  assign lizzieLet0_4QNode_Bool_4QNone_Bool_4QError_Bool_2_d = (lizzieLet0_4QNode_Bool_4QNone_Bool_4QError_Bool_d[0] && (! lizzieLet0_4QNode_Bool_4QNone_Bool_4QError_Bool_emitted[1]));
  assign lizzieLet0_4QNode_Bool_4QNone_Bool_4QError_Bool_done = (lizzieLet0_4QNode_Bool_4QNone_Bool_4QError_Bool_emitted | ({lizzieLet0_4QNode_Bool_4QNone_Bool_4QError_Bool_2_d[0],
                                                                                                                             lizzieLet0_4QNode_Bool_4QNone_Bool_4QError_Bool_1_d[0]} & {lizzieLet0_4QNode_Bool_4QNone_Bool_4QError_Bool_2_r,
                                                                                                                                                                                        lizzieLet0_4QNode_Bool_4QNone_Bool_4QError_Bool_1_r}));
  assign lizzieLet0_4QNode_Bool_4QNone_Bool_4QError_Bool_r = (& lizzieLet0_4QNode_Bool_4QNone_Bool_4QError_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNode_Bool_4QNone_Bool_4QError_Bool_emitted <= 2'd0;
    else
      lizzieLet0_4QNode_Bool_4QNone_Bool_4QError_Bool_emitted <= (lizzieLet0_4QNode_Bool_4QNone_Bool_4QError_Bool_r ? 2'd0 :
                                                                  lizzieLet0_4QNode_Bool_4QNone_Bool_4QError_Bool_done);
  
  /* dcon (Ty QTree_Bool,
      Dcon QError_Bool) : [(lizzieLet0_4QNode_Bool_4QNone_Bool_4QError_Bool_1,Go)] > (lizzieLet0_4QNode_Bool_4QNone_Bool_4QError_Bool_1QError_Bool,QTree_Bool) */
  assign lizzieLet0_4QNode_Bool_4QNone_Bool_4QError_Bool_1QError_Bool_d = QError_Bool_dc((& {lizzieLet0_4QNode_Bool_4QNone_Bool_4QError_Bool_1_d[0]}), lizzieLet0_4QNode_Bool_4QNone_Bool_4QError_Bool_1_d);
  assign {lizzieLet0_4QNode_Bool_4QNone_Bool_4QError_Bool_1_r} = {1 {(lizzieLet0_4QNode_Bool_4QNone_Bool_4QError_Bool_1QError_Bool_r && lizzieLet0_4QNode_Bool_4QNone_Bool_4QError_Bool_1QError_Bool_d[0])}};
  
  /* buf (Ty QTree_Bool) : (lizzieLet0_4QNode_Bool_4QNone_Bool_4QError_Bool_1QError_Bool,QTree_Bool) > (lizzieLet36_1_argbuf,QTree_Bool) */
  QTree_Bool_t lizzieLet0_4QNode_Bool_4QNone_Bool_4QError_Bool_1QError_Bool_bufchan_d;
  logic lizzieLet0_4QNode_Bool_4QNone_Bool_4QError_Bool_1QError_Bool_bufchan_r;
  assign lizzieLet0_4QNode_Bool_4QNone_Bool_4QError_Bool_1QError_Bool_r = ((! lizzieLet0_4QNode_Bool_4QNone_Bool_4QError_Bool_1QError_Bool_bufchan_d[0]) || lizzieLet0_4QNode_Bool_4QNone_Bool_4QError_Bool_1QError_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNode_Bool_4QNone_Bool_4QError_Bool_1QError_Bool_bufchan_d <= {66'd0,
                                                                                 1'd0};
    else
      if (lizzieLet0_4QNode_Bool_4QNone_Bool_4QError_Bool_1QError_Bool_r)
        lizzieLet0_4QNode_Bool_4QNone_Bool_4QError_Bool_1QError_Bool_bufchan_d <= lizzieLet0_4QNode_Bool_4QNone_Bool_4QError_Bool_1QError_Bool_d;
  QTree_Bool_t lizzieLet0_4QNode_Bool_4QNone_Bool_4QError_Bool_1QError_Bool_bufchan_buf;
  assign lizzieLet0_4QNode_Bool_4QNone_Bool_4QError_Bool_1QError_Bool_bufchan_r = (! lizzieLet0_4QNode_Bool_4QNone_Bool_4QError_Bool_1QError_Bool_bufchan_buf[0]);
  assign lizzieLet36_1_argbuf_d = (lizzieLet0_4QNode_Bool_4QNone_Bool_4QError_Bool_1QError_Bool_bufchan_buf[0] ? lizzieLet0_4QNode_Bool_4QNone_Bool_4QError_Bool_1QError_Bool_bufchan_buf :
                                   lizzieLet0_4QNode_Bool_4QNone_Bool_4QError_Bool_1QError_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNode_Bool_4QNone_Bool_4QError_Bool_1QError_Bool_bufchan_buf <= {66'd0,
                                                                                   1'd0};
    else
      if ((lizzieLet36_1_argbuf_r && lizzieLet0_4QNode_Bool_4QNone_Bool_4QError_Bool_1QError_Bool_bufchan_buf[0]))
        lizzieLet0_4QNode_Bool_4QNone_Bool_4QError_Bool_1QError_Bool_bufchan_buf <= {66'd0,
                                                                                     1'd0};
      else if (((! lizzieLet36_1_argbuf_r) && (! lizzieLet0_4QNode_Bool_4QNone_Bool_4QError_Bool_1QError_Bool_bufchan_buf[0])))
        lizzieLet0_4QNode_Bool_4QNone_Bool_4QError_Bool_1QError_Bool_bufchan_buf <= lizzieLet0_4QNode_Bool_4QNone_Bool_4QError_Bool_1QError_Bool_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet0_4QNode_Bool_4QNone_Bool_4QError_Bool_2,Go) > (lizzieLet0_4QNode_Bool_4QNone_Bool_4QError_Bool_2_argbuf,Go) */
  Go_t lizzieLet0_4QNode_Bool_4QNone_Bool_4QError_Bool_2_bufchan_d;
  logic lizzieLet0_4QNode_Bool_4QNone_Bool_4QError_Bool_2_bufchan_r;
  assign lizzieLet0_4QNode_Bool_4QNone_Bool_4QError_Bool_2_r = ((! lizzieLet0_4QNode_Bool_4QNone_Bool_4QError_Bool_2_bufchan_d[0]) || lizzieLet0_4QNode_Bool_4QNone_Bool_4QError_Bool_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNode_Bool_4QNone_Bool_4QError_Bool_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet0_4QNode_Bool_4QNone_Bool_4QError_Bool_2_r)
        lizzieLet0_4QNode_Bool_4QNone_Bool_4QError_Bool_2_bufchan_d <= lizzieLet0_4QNode_Bool_4QNone_Bool_4QError_Bool_2_d;
  Go_t lizzieLet0_4QNode_Bool_4QNone_Bool_4QError_Bool_2_bufchan_buf;
  assign lizzieLet0_4QNode_Bool_4QNone_Bool_4QError_Bool_2_bufchan_r = (! lizzieLet0_4QNode_Bool_4QNone_Bool_4QError_Bool_2_bufchan_buf[0]);
  assign lizzieLet0_4QNode_Bool_4QNone_Bool_4QError_Bool_2_argbuf_d = (lizzieLet0_4QNode_Bool_4QNone_Bool_4QError_Bool_2_bufchan_buf[0] ? lizzieLet0_4QNode_Bool_4QNone_Bool_4QError_Bool_2_bufchan_buf :
                                                                       lizzieLet0_4QNode_Bool_4QNone_Bool_4QError_Bool_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNode_Bool_4QNone_Bool_4QError_Bool_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet0_4QNode_Bool_4QNone_Bool_4QError_Bool_2_argbuf_r && lizzieLet0_4QNode_Bool_4QNone_Bool_4QError_Bool_2_bufchan_buf[0]))
        lizzieLet0_4QNode_Bool_4QNone_Bool_4QError_Bool_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet0_4QNode_Bool_4QNone_Bool_4QError_Bool_2_argbuf_r) && (! lizzieLet0_4QNode_Bool_4QNone_Bool_4QError_Bool_2_bufchan_buf[0])))
        lizzieLet0_4QNode_Bool_4QNone_Bool_4QError_Bool_2_bufchan_buf <= lizzieLet0_4QNode_Bool_4QNone_Bool_4QError_Bool_2_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool,Go) > [(lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_1,Go),
                                                                      (lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_2,Go),
                                                                      (lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_3,Go),
                                                                      (lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_4,Go),
                                                                      (lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_5,Go)] */
  logic [4:0] lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_emitted;
  logic [4:0] lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_done;
  assign lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_1_d = (lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_d[0] && (! lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_emitted[0]));
  assign lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_2_d = (lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_d[0] && (! lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_emitted[1]));
  assign lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_3_d = (lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_d[0] && (! lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_emitted[2]));
  assign lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_4_d = (lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_d[0] && (! lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_emitted[3]));
  assign lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_5_d = (lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_d[0] && (! lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_emitted[4]));
  assign lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_done = (lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_emitted | ({lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_5_d[0],
                                                                                                                           lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_4_d[0],
                                                                                                                           lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_3_d[0],
                                                                                                                           lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_2_d[0],
                                                                                                                           lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_1_d[0]} & {lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_5_r,
                                                                                                                                                                                     lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_4_r,
                                                                                                                                                                                     lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_3_r,
                                                                                                                                                                                     lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_2_r,
                                                                                                                                                                                     lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_1_r}));
  assign lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_r = (& lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_emitted <= 5'd0;
    else
      lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_emitted <= (lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_r ? 5'd0 :
                                                                 lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_done);
  
  /* buf (Ty Go) : (lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_1,Go) > (lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_1_argbuf,Go) */
  Go_t lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_1_bufchan_d;
  logic lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_1_bufchan_r;
  assign lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_1_r = ((! lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_1_bufchan_d[0]) || lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_1_bufchan_d <= 1'd0;
    else
      if (lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_1_r)
        lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_1_bufchan_d <= lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_1_d;
  Go_t lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_1_bufchan_buf;
  assign lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_1_bufchan_r = (! lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_1_bufchan_buf[0]);
  assign lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_1_argbuf_d = (lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_1_bufchan_buf[0] ? lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_1_bufchan_buf :
                                                                      lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_1_argbuf_r && lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_1_bufchan_buf[0]))
        lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_1_argbuf_r) && (! lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_1_bufchan_buf[0])))
        lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_1_bufchan_buf <= lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_1_bufchan_d;
  
  /* dcon (Ty TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool,
      Dcon TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool) : [(lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_1_argbuf,Go),
                                                               (lizzieLet0_4QNode_Bool_4QNone_Bool_3QNode_Bool_1_argbuf,Pointer_QTree_Bool),
                                                               (t4a8P_1_argbuf,Pointer_QTree_Bool)] > (f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool5,TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool) */
  assign \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool5_d  = TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_dc((& {lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_1_argbuf_d[0],
                                                                                                                                    lizzieLet0_4QNode_Bool_4QNone_Bool_3QNode_Bool_1_argbuf_d[0],
                                                                                                                                    t4a8P_1_argbuf_d[0]}), lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_1_argbuf_d, lizzieLet0_4QNode_Bool_4QNone_Bool_3QNode_Bool_1_argbuf_d, t4a8P_1_argbuf_d);
  assign {lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_1_argbuf_r,
          lizzieLet0_4QNode_Bool_4QNone_Bool_3QNode_Bool_1_argbuf_r,
          t4a8P_1_argbuf_r} = {3 {(\f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool5_r  && \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool5_d [0])}};
  
  /* buf (Ty Go) : (lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_2,Go) > (lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_2_argbuf,Go) */
  Go_t lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_2_bufchan_d;
  logic lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_2_bufchan_r;
  assign lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_2_r = ((! lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_2_bufchan_d[0]) || lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_2_r)
        lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_2_bufchan_d <= lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_2_d;
  Go_t lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_2_bufchan_buf;
  assign lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_2_bufchan_r = (! lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_2_bufchan_buf[0]);
  assign lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_2_argbuf_d = (lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_2_bufchan_buf[0] ? lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_2_bufchan_buf :
                                                                      lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_2_argbuf_r && lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_2_bufchan_buf[0]))
        lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_2_argbuf_r) && (! lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_2_bufchan_buf[0])))
        lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_2_bufchan_buf <= lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_2_bufchan_d;
  
  /* dcon (Ty TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool,
      Dcon TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool) : [(lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_2_argbuf,Go),
                                                               (lizzieLet0_4QNode_Bool_4QNone_Bool_9QNode_Bool_1_argbuf,Pointer_QTree_Bool),
                                                               (t3a8O_1_argbuf,Pointer_QTree_Bool)] > (f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool6,TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool) */
  assign \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool6_d  = TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_dc((& {lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_2_argbuf_d[0],
                                                                                                                                    lizzieLet0_4QNode_Bool_4QNone_Bool_9QNode_Bool_1_argbuf_d[0],
                                                                                                                                    t3a8O_1_argbuf_d[0]}), lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_2_argbuf_d, lizzieLet0_4QNode_Bool_4QNone_Bool_9QNode_Bool_1_argbuf_d, t3a8O_1_argbuf_d);
  assign {lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_2_argbuf_r,
          lizzieLet0_4QNode_Bool_4QNone_Bool_9QNode_Bool_1_argbuf_r,
          t3a8O_1_argbuf_r} = {3 {(\f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool6_r  && \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool6_d [0])}};
  
  /* buf (Ty Go) : (lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_3,Go) > (lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_3_argbuf,Go) */
  Go_t lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_3_bufchan_d;
  logic lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_3_bufchan_r;
  assign lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_3_r = ((! lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_3_bufchan_d[0]) || lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_3_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_3_bufchan_d <= 1'd0;
    else
      if (lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_3_r)
        lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_3_bufchan_d <= lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_3_d;
  Go_t lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_3_bufchan_buf;
  assign lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_3_bufchan_r = (! lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_3_bufchan_buf[0]);
  assign lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_3_argbuf_d = (lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_3_bufchan_buf[0] ? lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_3_bufchan_buf :
                                                                      lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_3_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_3_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_3_argbuf_r && lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_3_bufchan_buf[0]))
        lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_3_bufchan_buf <= 1'd0;
      else if (((! lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_3_argbuf_r) && (! lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_3_bufchan_buf[0])))
        lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_3_bufchan_buf <= lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_3_bufchan_d;
  
  /* dcon (Ty TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool,
      Dcon TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool) : [(lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_3_argbuf,Go),
                                                               (lizzieLet0_4QNode_Bool_4QNone_Bool_8QNode_Bool_1_argbuf,Pointer_QTree_Bool),
                                                               (t2a8N_1_argbuf,Pointer_QTree_Bool)] > (f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool7,TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool) */
  assign \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool7_d  = TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_dc((& {lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_3_argbuf_d[0],
                                                                                                                                    lizzieLet0_4QNode_Bool_4QNone_Bool_8QNode_Bool_1_argbuf_d[0],
                                                                                                                                    t2a8N_1_argbuf_d[0]}), lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_3_argbuf_d, lizzieLet0_4QNode_Bool_4QNone_Bool_8QNode_Bool_1_argbuf_d, t2a8N_1_argbuf_d);
  assign {lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_3_argbuf_r,
          lizzieLet0_4QNode_Bool_4QNone_Bool_8QNode_Bool_1_argbuf_r,
          t2a8N_1_argbuf_r} = {3 {(\f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool7_r  && \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool7_d [0])}};
  
  /* buf (Ty Go) : (lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_4,Go) > (lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_4_argbuf,Go) */
  Go_t lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_4_bufchan_d;
  logic lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_4_bufchan_r;
  assign lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_4_r = ((! lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_4_bufchan_d[0]) || lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_4_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_4_bufchan_d <= 1'd0;
    else
      if (lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_4_r)
        lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_4_bufchan_d <= lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_4_d;
  Go_t lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_4_bufchan_buf;
  assign lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_4_bufchan_r = (! lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_4_bufchan_buf[0]);
  assign lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_4_argbuf_d = (lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_4_bufchan_buf[0] ? lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_4_bufchan_buf :
                                                                      lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_4_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_4_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_4_argbuf_r && lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_4_bufchan_buf[0]))
        lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_4_bufchan_buf <= 1'd0;
      else if (((! lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_4_argbuf_r) && (! lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_4_bufchan_buf[0])))
        lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_4_bufchan_buf <= lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_4_bufchan_d;
  
  /* dcon (Ty TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool,
      Dcon TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool) : [(lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_4_argbuf,Go),
                                                               (lizzieLet0_4QNode_Bool_4QNone_Bool_7QNode_Bool_1_argbuf,Pointer_QTree_Bool),
                                                               (t1a8M_1_argbuf,Pointer_QTree_Bool)] > (f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool8,TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool) */
  assign \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool8_d  = TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_dc((& {lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_4_argbuf_d[0],
                                                                                                                                    lizzieLet0_4QNode_Bool_4QNone_Bool_7QNode_Bool_1_argbuf_d[0],
                                                                                                                                    t1a8M_1_argbuf_d[0]}), lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_4_argbuf_d, lizzieLet0_4QNode_Bool_4QNone_Bool_7QNode_Bool_1_argbuf_d, t1a8M_1_argbuf_d);
  assign {lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_4_argbuf_r,
          lizzieLet0_4QNode_Bool_4QNone_Bool_7QNode_Bool_1_argbuf_r,
          t1a8M_1_argbuf_r} = {3 {(\f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool8_r  && \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool8_d [0])}};
  
  /* buf (Ty Go) : (lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_5,Go) > (lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_5_argbuf,Go) */
  Go_t lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_5_bufchan_d;
  logic lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_5_bufchan_r;
  assign lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_5_r = ((! lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_5_bufchan_d[0]) || lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_5_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_5_bufchan_d <= 1'd0;
    else
      if (lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_5_r)
        lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_5_bufchan_d <= lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_5_d;
  Go_t lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_5_bufchan_buf;
  assign lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_5_bufchan_r = (! lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_5_bufchan_buf[0]);
  assign lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_5_argbuf_d = (lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_5_bufchan_buf[0] ? lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_5_bufchan_buf :
                                                                      lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_5_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_5_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_5_argbuf_r && lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_5_bufchan_buf[0]))
        lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_5_bufchan_buf <= 1'd0;
      else if (((! lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_5_argbuf_r) && (! lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_5_bufchan_buf[0])))
        lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_5_bufchan_buf <= lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_5_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet0_4QNode_Bool_4QNone_Bool_4QNone_Bool,Go) > (lizzieLet0_4QNode_Bool_4QNone_Bool_4QNone_Bool_1_argbuf,Go) */
  Go_t lizzieLet0_4QNode_Bool_4QNone_Bool_4QNone_Bool_bufchan_d;
  logic lizzieLet0_4QNode_Bool_4QNone_Bool_4QNone_Bool_bufchan_r;
  assign lizzieLet0_4QNode_Bool_4QNone_Bool_4QNone_Bool_r = ((! lizzieLet0_4QNode_Bool_4QNone_Bool_4QNone_Bool_bufchan_d[0]) || lizzieLet0_4QNode_Bool_4QNone_Bool_4QNone_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNode_Bool_4QNone_Bool_4QNone_Bool_bufchan_d <= 1'd0;
    else
      if (lizzieLet0_4QNode_Bool_4QNone_Bool_4QNone_Bool_r)
        lizzieLet0_4QNode_Bool_4QNone_Bool_4QNone_Bool_bufchan_d <= lizzieLet0_4QNode_Bool_4QNone_Bool_4QNone_Bool_d;
  Go_t lizzieLet0_4QNode_Bool_4QNone_Bool_4QNone_Bool_bufchan_buf;
  assign lizzieLet0_4QNode_Bool_4QNone_Bool_4QNone_Bool_bufchan_r = (! lizzieLet0_4QNode_Bool_4QNone_Bool_4QNone_Bool_bufchan_buf[0]);
  assign lizzieLet0_4QNode_Bool_4QNone_Bool_4QNone_Bool_1_argbuf_d = (lizzieLet0_4QNode_Bool_4QNone_Bool_4QNone_Bool_bufchan_buf[0] ? lizzieLet0_4QNode_Bool_4QNone_Bool_4QNone_Bool_bufchan_buf :
                                                                      lizzieLet0_4QNode_Bool_4QNone_Bool_4QNone_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNode_Bool_4QNone_Bool_4QNone_Bool_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet0_4QNode_Bool_4QNone_Bool_4QNone_Bool_1_argbuf_r && lizzieLet0_4QNode_Bool_4QNone_Bool_4QNone_Bool_bufchan_buf[0]))
        lizzieLet0_4QNode_Bool_4QNone_Bool_4QNone_Bool_bufchan_buf <= 1'd0;
      else if (((! lizzieLet0_4QNode_Bool_4QNone_Bool_4QNone_Bool_1_argbuf_r) && (! lizzieLet0_4QNode_Bool_4QNone_Bool_4QNone_Bool_bufchan_buf[0])))
        lizzieLet0_4QNode_Bool_4QNone_Bool_4QNone_Bool_bufchan_buf <= lizzieLet0_4QNode_Bool_4QNone_Bool_4QNone_Bool_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet0_4QNode_Bool_4QNone_Bool_4QVal_Bool,Go) > [(lizzieLet0_4QNode_Bool_4QNone_Bool_4QVal_Bool_1,Go),
                                                                     (lizzieLet0_4QNode_Bool_4QNone_Bool_4QVal_Bool_2,Go)] */
  logic [1:0] lizzieLet0_4QNode_Bool_4QNone_Bool_4QVal_Bool_emitted;
  logic [1:0] lizzieLet0_4QNode_Bool_4QNone_Bool_4QVal_Bool_done;
  assign lizzieLet0_4QNode_Bool_4QNone_Bool_4QVal_Bool_1_d = (lizzieLet0_4QNode_Bool_4QNone_Bool_4QVal_Bool_d[0] && (! lizzieLet0_4QNode_Bool_4QNone_Bool_4QVal_Bool_emitted[0]));
  assign lizzieLet0_4QNode_Bool_4QNone_Bool_4QVal_Bool_2_d = (lizzieLet0_4QNode_Bool_4QNone_Bool_4QVal_Bool_d[0] && (! lizzieLet0_4QNode_Bool_4QNone_Bool_4QVal_Bool_emitted[1]));
  assign lizzieLet0_4QNode_Bool_4QNone_Bool_4QVal_Bool_done = (lizzieLet0_4QNode_Bool_4QNone_Bool_4QVal_Bool_emitted | ({lizzieLet0_4QNode_Bool_4QNone_Bool_4QVal_Bool_2_d[0],
                                                                                                                         lizzieLet0_4QNode_Bool_4QNone_Bool_4QVal_Bool_1_d[0]} & {lizzieLet0_4QNode_Bool_4QNone_Bool_4QVal_Bool_2_r,
                                                                                                                                                                                  lizzieLet0_4QNode_Bool_4QNone_Bool_4QVal_Bool_1_r}));
  assign lizzieLet0_4QNode_Bool_4QNone_Bool_4QVal_Bool_r = (& lizzieLet0_4QNode_Bool_4QNone_Bool_4QVal_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNode_Bool_4QNone_Bool_4QVal_Bool_emitted <= 2'd0;
    else
      lizzieLet0_4QNode_Bool_4QNone_Bool_4QVal_Bool_emitted <= (lizzieLet0_4QNode_Bool_4QNone_Bool_4QVal_Bool_r ? 2'd0 :
                                                                lizzieLet0_4QNode_Bool_4QNone_Bool_4QVal_Bool_done);
  
  /* dcon (Ty QTree_Bool,
      Dcon QError_Bool) : [(lizzieLet0_4QNode_Bool_4QNone_Bool_4QVal_Bool_1,Go)] > (lizzieLet0_4QNode_Bool_4QNone_Bool_4QVal_Bool_1QError_Bool,QTree_Bool) */
  assign lizzieLet0_4QNode_Bool_4QNone_Bool_4QVal_Bool_1QError_Bool_d = QError_Bool_dc((& {lizzieLet0_4QNode_Bool_4QNone_Bool_4QVal_Bool_1_d[0]}), lizzieLet0_4QNode_Bool_4QNone_Bool_4QVal_Bool_1_d);
  assign {lizzieLet0_4QNode_Bool_4QNone_Bool_4QVal_Bool_1_r} = {1 {(lizzieLet0_4QNode_Bool_4QNone_Bool_4QVal_Bool_1QError_Bool_r && lizzieLet0_4QNode_Bool_4QNone_Bool_4QVal_Bool_1QError_Bool_d[0])}};
  
  /* buf (Ty QTree_Bool) : (lizzieLet0_4QNode_Bool_4QNone_Bool_4QVal_Bool_1QError_Bool,QTree_Bool) > (lizzieLet34_1_argbuf,QTree_Bool) */
  QTree_Bool_t lizzieLet0_4QNode_Bool_4QNone_Bool_4QVal_Bool_1QError_Bool_bufchan_d;
  logic lizzieLet0_4QNode_Bool_4QNone_Bool_4QVal_Bool_1QError_Bool_bufchan_r;
  assign lizzieLet0_4QNode_Bool_4QNone_Bool_4QVal_Bool_1QError_Bool_r = ((! lizzieLet0_4QNode_Bool_4QNone_Bool_4QVal_Bool_1QError_Bool_bufchan_d[0]) || lizzieLet0_4QNode_Bool_4QNone_Bool_4QVal_Bool_1QError_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNode_Bool_4QNone_Bool_4QVal_Bool_1QError_Bool_bufchan_d <= {66'd0,
                                                                               1'd0};
    else
      if (lizzieLet0_4QNode_Bool_4QNone_Bool_4QVal_Bool_1QError_Bool_r)
        lizzieLet0_4QNode_Bool_4QNone_Bool_4QVal_Bool_1QError_Bool_bufchan_d <= lizzieLet0_4QNode_Bool_4QNone_Bool_4QVal_Bool_1QError_Bool_d;
  QTree_Bool_t lizzieLet0_4QNode_Bool_4QNone_Bool_4QVal_Bool_1QError_Bool_bufchan_buf;
  assign lizzieLet0_4QNode_Bool_4QNone_Bool_4QVal_Bool_1QError_Bool_bufchan_r = (! lizzieLet0_4QNode_Bool_4QNone_Bool_4QVal_Bool_1QError_Bool_bufchan_buf[0]);
  assign lizzieLet34_1_argbuf_d = (lizzieLet0_4QNode_Bool_4QNone_Bool_4QVal_Bool_1QError_Bool_bufchan_buf[0] ? lizzieLet0_4QNode_Bool_4QNone_Bool_4QVal_Bool_1QError_Bool_bufchan_buf :
                                   lizzieLet0_4QNode_Bool_4QNone_Bool_4QVal_Bool_1QError_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNode_Bool_4QNone_Bool_4QVal_Bool_1QError_Bool_bufchan_buf <= {66'd0,
                                                                                 1'd0};
    else
      if ((lizzieLet34_1_argbuf_r && lizzieLet0_4QNode_Bool_4QNone_Bool_4QVal_Bool_1QError_Bool_bufchan_buf[0]))
        lizzieLet0_4QNode_Bool_4QNone_Bool_4QVal_Bool_1QError_Bool_bufchan_buf <= {66'd0,
                                                                                   1'd0};
      else if (((! lizzieLet34_1_argbuf_r) && (! lizzieLet0_4QNode_Bool_4QNone_Bool_4QVal_Bool_1QError_Bool_bufchan_buf[0])))
        lizzieLet0_4QNode_Bool_4QNone_Bool_4QVal_Bool_1QError_Bool_bufchan_buf <= lizzieLet0_4QNode_Bool_4QNone_Bool_4QVal_Bool_1QError_Bool_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet0_4QNode_Bool_4QNone_Bool_4QVal_Bool_2,Go) > (lizzieLet0_4QNode_Bool_4QNone_Bool_4QVal_Bool_2_argbuf,Go) */
  Go_t lizzieLet0_4QNode_Bool_4QNone_Bool_4QVal_Bool_2_bufchan_d;
  logic lizzieLet0_4QNode_Bool_4QNone_Bool_4QVal_Bool_2_bufchan_r;
  assign lizzieLet0_4QNode_Bool_4QNone_Bool_4QVal_Bool_2_r = ((! lizzieLet0_4QNode_Bool_4QNone_Bool_4QVal_Bool_2_bufchan_d[0]) || lizzieLet0_4QNode_Bool_4QNone_Bool_4QVal_Bool_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNode_Bool_4QNone_Bool_4QVal_Bool_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet0_4QNode_Bool_4QNone_Bool_4QVal_Bool_2_r)
        lizzieLet0_4QNode_Bool_4QNone_Bool_4QVal_Bool_2_bufchan_d <= lizzieLet0_4QNode_Bool_4QNone_Bool_4QVal_Bool_2_d;
  Go_t lizzieLet0_4QNode_Bool_4QNone_Bool_4QVal_Bool_2_bufchan_buf;
  assign lizzieLet0_4QNode_Bool_4QNone_Bool_4QVal_Bool_2_bufchan_r = (! lizzieLet0_4QNode_Bool_4QNone_Bool_4QVal_Bool_2_bufchan_buf[0]);
  assign lizzieLet0_4QNode_Bool_4QNone_Bool_4QVal_Bool_2_argbuf_d = (lizzieLet0_4QNode_Bool_4QNone_Bool_4QVal_Bool_2_bufchan_buf[0] ? lizzieLet0_4QNode_Bool_4QNone_Bool_4QVal_Bool_2_bufchan_buf :
                                                                     lizzieLet0_4QNode_Bool_4QNone_Bool_4QVal_Bool_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNode_Bool_4QNone_Bool_4QVal_Bool_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet0_4QNode_Bool_4QNone_Bool_4QVal_Bool_2_argbuf_r && lizzieLet0_4QNode_Bool_4QNone_Bool_4QVal_Bool_2_bufchan_buf[0]))
        lizzieLet0_4QNode_Bool_4QNone_Bool_4QVal_Bool_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet0_4QNode_Bool_4QNone_Bool_4QVal_Bool_2_argbuf_r) && (! lizzieLet0_4QNode_Bool_4QNone_Bool_4QVal_Bool_2_bufchan_buf[0])))
        lizzieLet0_4QNode_Bool_4QNone_Bool_4QVal_Bool_2_bufchan_buf <= lizzieLet0_4QNode_Bool_4QNone_Bool_4QVal_Bool_2_bufchan_d;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_QTree_Bool) : (lizzieLet0_4QNode_Bool_4QNone_Bool_5,QTree_Bool) (lizzieLet0_4QNode_Bool_5QNone_Bool,Pointer_QTree_Bool) > [(lizzieLet0_4QNode_Bool_4QNone_Bool_5QNone_Bool,Pointer_QTree_Bool),
                                                                                                                                             (_133,Pointer_QTree_Bool),
                                                                                                                                             (_132,Pointer_QTree_Bool),
                                                                                                                                             (_131,Pointer_QTree_Bool)] */
  logic [3:0] lizzieLet0_4QNode_Bool_5QNone_Bool_onehotd;
  always_comb
    if ((lizzieLet0_4QNode_Bool_4QNone_Bool_5_d[0] && lizzieLet0_4QNode_Bool_5QNone_Bool_d[0]))
      unique case (lizzieLet0_4QNode_Bool_4QNone_Bool_5_d[2:1])
        2'd0: lizzieLet0_4QNode_Bool_5QNone_Bool_onehotd = 4'd1;
        2'd1: lizzieLet0_4QNode_Bool_5QNone_Bool_onehotd = 4'd2;
        2'd2: lizzieLet0_4QNode_Bool_5QNone_Bool_onehotd = 4'd4;
        2'd3: lizzieLet0_4QNode_Bool_5QNone_Bool_onehotd = 4'd8;
        default: lizzieLet0_4QNode_Bool_5QNone_Bool_onehotd = 4'd0;
      endcase
    else lizzieLet0_4QNode_Bool_5QNone_Bool_onehotd = 4'd0;
  assign lizzieLet0_4QNode_Bool_4QNone_Bool_5QNone_Bool_d = {lizzieLet0_4QNode_Bool_5QNone_Bool_d[16:1],
                                                             lizzieLet0_4QNode_Bool_5QNone_Bool_onehotd[0]};
  assign _133_d = {lizzieLet0_4QNode_Bool_5QNone_Bool_d[16:1],
                   lizzieLet0_4QNode_Bool_5QNone_Bool_onehotd[1]};
  assign _132_d = {lizzieLet0_4QNode_Bool_5QNone_Bool_d[16:1],
                   lizzieLet0_4QNode_Bool_5QNone_Bool_onehotd[2]};
  assign _131_d = {lizzieLet0_4QNode_Bool_5QNone_Bool_d[16:1],
                   lizzieLet0_4QNode_Bool_5QNone_Bool_onehotd[3]};
  assign lizzieLet0_4QNode_Bool_5QNone_Bool_r = (| (lizzieLet0_4QNode_Bool_5QNone_Bool_onehotd & {_131_r,
                                                                                                  _132_r,
                                                                                                  _133_r,
                                                                                                  lizzieLet0_4QNode_Bool_4QNone_Bool_5QNone_Bool_r}));
  assign lizzieLet0_4QNode_Bool_4QNone_Bool_5_r = lizzieLet0_4QNode_Bool_5QNone_Bool_r;
  
  /* buf (Ty Pointer_QTree_Bool) : (lizzieLet0_4QNode_Bool_4QNone_Bool_5QNone_Bool,Pointer_QTree_Bool) > (lizzieLet0_4QNode_Bool_4QNone_Bool_5QNone_Bool_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t lizzieLet0_4QNode_Bool_4QNone_Bool_5QNone_Bool_bufchan_d;
  logic lizzieLet0_4QNode_Bool_4QNone_Bool_5QNone_Bool_bufchan_r;
  assign lizzieLet0_4QNode_Bool_4QNone_Bool_5QNone_Bool_r = ((! lizzieLet0_4QNode_Bool_4QNone_Bool_5QNone_Bool_bufchan_d[0]) || lizzieLet0_4QNode_Bool_4QNone_Bool_5QNone_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNode_Bool_4QNone_Bool_5QNone_Bool_bufchan_d <= {16'd0,
                                                                   1'd0};
    else
      if (lizzieLet0_4QNode_Bool_4QNone_Bool_5QNone_Bool_r)
        lizzieLet0_4QNode_Bool_4QNone_Bool_5QNone_Bool_bufchan_d <= lizzieLet0_4QNode_Bool_4QNone_Bool_5QNone_Bool_d;
  Pointer_QTree_Bool_t lizzieLet0_4QNode_Bool_4QNone_Bool_5QNone_Bool_bufchan_buf;
  assign lizzieLet0_4QNode_Bool_4QNone_Bool_5QNone_Bool_bufchan_r = (! lizzieLet0_4QNode_Bool_4QNone_Bool_5QNone_Bool_bufchan_buf[0]);
  assign lizzieLet0_4QNode_Bool_4QNone_Bool_5QNone_Bool_1_argbuf_d = (lizzieLet0_4QNode_Bool_4QNone_Bool_5QNone_Bool_bufchan_buf[0] ? lizzieLet0_4QNode_Bool_4QNone_Bool_5QNone_Bool_bufchan_buf :
                                                                      lizzieLet0_4QNode_Bool_4QNone_Bool_5QNone_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNode_Bool_4QNone_Bool_5QNone_Bool_bufchan_buf <= {16'd0,
                                                                     1'd0};
    else
      if ((lizzieLet0_4QNode_Bool_4QNone_Bool_5QNone_Bool_1_argbuf_r && lizzieLet0_4QNode_Bool_4QNone_Bool_5QNone_Bool_bufchan_buf[0]))
        lizzieLet0_4QNode_Bool_4QNone_Bool_5QNone_Bool_bufchan_buf <= {16'd0,
                                                                       1'd0};
      else if (((! lizzieLet0_4QNode_Bool_4QNone_Bool_5QNone_Bool_1_argbuf_r) && (! lizzieLet0_4QNode_Bool_4QNone_Bool_5QNone_Bool_bufchan_buf[0])))
        lizzieLet0_4QNode_Bool_4QNone_Bool_5QNone_Bool_bufchan_buf <= lizzieLet0_4QNode_Bool_4QNone_Bool_5QNone_Bool_bufchan_d;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_CTf) : (lizzieLet0_4QNode_Bool_4QNone_Bool_6,QTree_Bool) (lizzieLet0_4QNode_Bool_6QNone_Bool,Pointer_CTf) > [(lizzieLet0_4QNode_Bool_4QNone_Bool_6QNone_Bool,Pointer_CTf),
                                                                                                                               (lizzieLet0_4QNode_Bool_4QNone_Bool_6QVal_Bool,Pointer_CTf),
                                                                                                                               (lizzieLet0_4QNode_Bool_4QNone_Bool_6QNode_Bool,Pointer_CTf),
                                                                                                                               (lizzieLet0_4QNode_Bool_4QNone_Bool_6QError_Bool,Pointer_CTf)] */
  logic [3:0] lizzieLet0_4QNode_Bool_6QNone_Bool_onehotd;
  always_comb
    if ((lizzieLet0_4QNode_Bool_4QNone_Bool_6_d[0] && lizzieLet0_4QNode_Bool_6QNone_Bool_d[0]))
      unique case (lizzieLet0_4QNode_Bool_4QNone_Bool_6_d[2:1])
        2'd0: lizzieLet0_4QNode_Bool_6QNone_Bool_onehotd = 4'd1;
        2'd1: lizzieLet0_4QNode_Bool_6QNone_Bool_onehotd = 4'd2;
        2'd2: lizzieLet0_4QNode_Bool_6QNone_Bool_onehotd = 4'd4;
        2'd3: lizzieLet0_4QNode_Bool_6QNone_Bool_onehotd = 4'd8;
        default: lizzieLet0_4QNode_Bool_6QNone_Bool_onehotd = 4'd0;
      endcase
    else lizzieLet0_4QNode_Bool_6QNone_Bool_onehotd = 4'd0;
  assign lizzieLet0_4QNode_Bool_4QNone_Bool_6QNone_Bool_d = {lizzieLet0_4QNode_Bool_6QNone_Bool_d[16:1],
                                                             lizzieLet0_4QNode_Bool_6QNone_Bool_onehotd[0]};
  assign lizzieLet0_4QNode_Bool_4QNone_Bool_6QVal_Bool_d = {lizzieLet0_4QNode_Bool_6QNone_Bool_d[16:1],
                                                            lizzieLet0_4QNode_Bool_6QNone_Bool_onehotd[1]};
  assign lizzieLet0_4QNode_Bool_4QNone_Bool_6QNode_Bool_d = {lizzieLet0_4QNode_Bool_6QNone_Bool_d[16:1],
                                                             lizzieLet0_4QNode_Bool_6QNone_Bool_onehotd[2]};
  assign lizzieLet0_4QNode_Bool_4QNone_Bool_6QError_Bool_d = {lizzieLet0_4QNode_Bool_6QNone_Bool_d[16:1],
                                                              lizzieLet0_4QNode_Bool_6QNone_Bool_onehotd[3]};
  assign lizzieLet0_4QNode_Bool_6QNone_Bool_r = (| (lizzieLet0_4QNode_Bool_6QNone_Bool_onehotd & {lizzieLet0_4QNode_Bool_4QNone_Bool_6QError_Bool_r,
                                                                                                  lizzieLet0_4QNode_Bool_4QNone_Bool_6QNode_Bool_r,
                                                                                                  lizzieLet0_4QNode_Bool_4QNone_Bool_6QVal_Bool_r,
                                                                                                  lizzieLet0_4QNode_Bool_4QNone_Bool_6QNone_Bool_r}));
  assign lizzieLet0_4QNode_Bool_4QNone_Bool_6_r = lizzieLet0_4QNode_Bool_6QNone_Bool_r;
  
  /* buf (Ty Pointer_CTf) : (lizzieLet0_4QNode_Bool_4QNone_Bool_6QError_Bool,Pointer_CTf) > (lizzieLet0_4QNode_Bool_4QNone_Bool_6QError_Bool_1_argbuf,Pointer_CTf) */
  Pointer_CTf_t lizzieLet0_4QNode_Bool_4QNone_Bool_6QError_Bool_bufchan_d;
  logic lizzieLet0_4QNode_Bool_4QNone_Bool_6QError_Bool_bufchan_r;
  assign lizzieLet0_4QNode_Bool_4QNone_Bool_6QError_Bool_r = ((! lizzieLet0_4QNode_Bool_4QNone_Bool_6QError_Bool_bufchan_d[0]) || lizzieLet0_4QNode_Bool_4QNone_Bool_6QError_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNode_Bool_4QNone_Bool_6QError_Bool_bufchan_d <= {16'd0,
                                                                    1'd0};
    else
      if (lizzieLet0_4QNode_Bool_4QNone_Bool_6QError_Bool_r)
        lizzieLet0_4QNode_Bool_4QNone_Bool_6QError_Bool_bufchan_d <= lizzieLet0_4QNode_Bool_4QNone_Bool_6QError_Bool_d;
  Pointer_CTf_t lizzieLet0_4QNode_Bool_4QNone_Bool_6QError_Bool_bufchan_buf;
  assign lizzieLet0_4QNode_Bool_4QNone_Bool_6QError_Bool_bufchan_r = (! lizzieLet0_4QNode_Bool_4QNone_Bool_6QError_Bool_bufchan_buf[0]);
  assign lizzieLet0_4QNode_Bool_4QNone_Bool_6QError_Bool_1_argbuf_d = (lizzieLet0_4QNode_Bool_4QNone_Bool_6QError_Bool_bufchan_buf[0] ? lizzieLet0_4QNode_Bool_4QNone_Bool_6QError_Bool_bufchan_buf :
                                                                       lizzieLet0_4QNode_Bool_4QNone_Bool_6QError_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNode_Bool_4QNone_Bool_6QError_Bool_bufchan_buf <= {16'd0,
                                                                      1'd0};
    else
      if ((lizzieLet0_4QNode_Bool_4QNone_Bool_6QError_Bool_1_argbuf_r && lizzieLet0_4QNode_Bool_4QNone_Bool_6QError_Bool_bufchan_buf[0]))
        lizzieLet0_4QNode_Bool_4QNone_Bool_6QError_Bool_bufchan_buf <= {16'd0,
                                                                        1'd0};
      else if (((! lizzieLet0_4QNode_Bool_4QNone_Bool_6QError_Bool_1_argbuf_r) && (! lizzieLet0_4QNode_Bool_4QNone_Bool_6QError_Bool_bufchan_buf[0])))
        lizzieLet0_4QNode_Bool_4QNone_Bool_6QError_Bool_bufchan_buf <= lizzieLet0_4QNode_Bool_4QNone_Bool_6QError_Bool_bufchan_d;
  
  /* buf (Ty Pointer_CTf) : (lizzieLet0_4QNode_Bool_4QNone_Bool_6QNode_Bool,Pointer_CTf) > (lizzieLet0_4QNode_Bool_4QNone_Bool_6QNode_Bool_1_argbuf,Pointer_CTf) */
  Pointer_CTf_t lizzieLet0_4QNode_Bool_4QNone_Bool_6QNode_Bool_bufchan_d;
  logic lizzieLet0_4QNode_Bool_4QNone_Bool_6QNode_Bool_bufchan_r;
  assign lizzieLet0_4QNode_Bool_4QNone_Bool_6QNode_Bool_r = ((! lizzieLet0_4QNode_Bool_4QNone_Bool_6QNode_Bool_bufchan_d[0]) || lizzieLet0_4QNode_Bool_4QNone_Bool_6QNode_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNode_Bool_4QNone_Bool_6QNode_Bool_bufchan_d <= {16'd0,
                                                                   1'd0};
    else
      if (lizzieLet0_4QNode_Bool_4QNone_Bool_6QNode_Bool_r)
        lizzieLet0_4QNode_Bool_4QNone_Bool_6QNode_Bool_bufchan_d <= lizzieLet0_4QNode_Bool_4QNone_Bool_6QNode_Bool_d;
  Pointer_CTf_t lizzieLet0_4QNode_Bool_4QNone_Bool_6QNode_Bool_bufchan_buf;
  assign lizzieLet0_4QNode_Bool_4QNone_Bool_6QNode_Bool_bufchan_r = (! lizzieLet0_4QNode_Bool_4QNone_Bool_6QNode_Bool_bufchan_buf[0]);
  assign lizzieLet0_4QNode_Bool_4QNone_Bool_6QNode_Bool_1_argbuf_d = (lizzieLet0_4QNode_Bool_4QNone_Bool_6QNode_Bool_bufchan_buf[0] ? lizzieLet0_4QNode_Bool_4QNone_Bool_6QNode_Bool_bufchan_buf :
                                                                      lizzieLet0_4QNode_Bool_4QNone_Bool_6QNode_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNode_Bool_4QNone_Bool_6QNode_Bool_bufchan_buf <= {16'd0,
                                                                     1'd0};
    else
      if ((lizzieLet0_4QNode_Bool_4QNone_Bool_6QNode_Bool_1_argbuf_r && lizzieLet0_4QNode_Bool_4QNone_Bool_6QNode_Bool_bufchan_buf[0]))
        lizzieLet0_4QNode_Bool_4QNone_Bool_6QNode_Bool_bufchan_buf <= {16'd0,
                                                                       1'd0};
      else if (((! lizzieLet0_4QNode_Bool_4QNone_Bool_6QNode_Bool_1_argbuf_r) && (! lizzieLet0_4QNode_Bool_4QNone_Bool_6QNode_Bool_bufchan_buf[0])))
        lizzieLet0_4QNode_Bool_4QNone_Bool_6QNode_Bool_bufchan_buf <= lizzieLet0_4QNode_Bool_4QNone_Bool_6QNode_Bool_bufchan_d;
  
  /* buf (Ty Pointer_CTf) : (lizzieLet0_4QNode_Bool_4QNone_Bool_6QNone_Bool,Pointer_CTf) > (lizzieLet0_4QNode_Bool_4QNone_Bool_6QNone_Bool_1_argbuf,Pointer_CTf) */
  Pointer_CTf_t lizzieLet0_4QNode_Bool_4QNone_Bool_6QNone_Bool_bufchan_d;
  logic lizzieLet0_4QNode_Bool_4QNone_Bool_6QNone_Bool_bufchan_r;
  assign lizzieLet0_4QNode_Bool_4QNone_Bool_6QNone_Bool_r = ((! lizzieLet0_4QNode_Bool_4QNone_Bool_6QNone_Bool_bufchan_d[0]) || lizzieLet0_4QNode_Bool_4QNone_Bool_6QNone_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNode_Bool_4QNone_Bool_6QNone_Bool_bufchan_d <= {16'd0,
                                                                   1'd0};
    else
      if (lizzieLet0_4QNode_Bool_4QNone_Bool_6QNone_Bool_r)
        lizzieLet0_4QNode_Bool_4QNone_Bool_6QNone_Bool_bufchan_d <= lizzieLet0_4QNode_Bool_4QNone_Bool_6QNone_Bool_d;
  Pointer_CTf_t lizzieLet0_4QNode_Bool_4QNone_Bool_6QNone_Bool_bufchan_buf;
  assign lizzieLet0_4QNode_Bool_4QNone_Bool_6QNone_Bool_bufchan_r = (! lizzieLet0_4QNode_Bool_4QNone_Bool_6QNone_Bool_bufchan_buf[0]);
  assign lizzieLet0_4QNode_Bool_4QNone_Bool_6QNone_Bool_1_argbuf_d = (lizzieLet0_4QNode_Bool_4QNone_Bool_6QNone_Bool_bufchan_buf[0] ? lizzieLet0_4QNode_Bool_4QNone_Bool_6QNone_Bool_bufchan_buf :
                                                                      lizzieLet0_4QNode_Bool_4QNone_Bool_6QNone_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNode_Bool_4QNone_Bool_6QNone_Bool_bufchan_buf <= {16'd0,
                                                                     1'd0};
    else
      if ((lizzieLet0_4QNode_Bool_4QNone_Bool_6QNone_Bool_1_argbuf_r && lizzieLet0_4QNode_Bool_4QNone_Bool_6QNone_Bool_bufchan_buf[0]))
        lizzieLet0_4QNode_Bool_4QNone_Bool_6QNone_Bool_bufchan_buf <= {16'd0,
                                                                       1'd0};
      else if (((! lizzieLet0_4QNode_Bool_4QNone_Bool_6QNone_Bool_1_argbuf_r) && (! lizzieLet0_4QNode_Bool_4QNone_Bool_6QNone_Bool_bufchan_buf[0])))
        lizzieLet0_4QNode_Bool_4QNone_Bool_6QNone_Bool_bufchan_buf <= lizzieLet0_4QNode_Bool_4QNone_Bool_6QNone_Bool_bufchan_d;
  
  /* buf (Ty Pointer_CTf) : (lizzieLet0_4QNode_Bool_4QNone_Bool_6QVal_Bool,Pointer_CTf) > (lizzieLet0_4QNode_Bool_4QNone_Bool_6QVal_Bool_1_argbuf,Pointer_CTf) */
  Pointer_CTf_t lizzieLet0_4QNode_Bool_4QNone_Bool_6QVal_Bool_bufchan_d;
  logic lizzieLet0_4QNode_Bool_4QNone_Bool_6QVal_Bool_bufchan_r;
  assign lizzieLet0_4QNode_Bool_4QNone_Bool_6QVal_Bool_r = ((! lizzieLet0_4QNode_Bool_4QNone_Bool_6QVal_Bool_bufchan_d[0]) || lizzieLet0_4QNode_Bool_4QNone_Bool_6QVal_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNode_Bool_4QNone_Bool_6QVal_Bool_bufchan_d <= {16'd0,
                                                                  1'd0};
    else
      if (lizzieLet0_4QNode_Bool_4QNone_Bool_6QVal_Bool_r)
        lizzieLet0_4QNode_Bool_4QNone_Bool_6QVal_Bool_bufchan_d <= lizzieLet0_4QNode_Bool_4QNone_Bool_6QVal_Bool_d;
  Pointer_CTf_t lizzieLet0_4QNode_Bool_4QNone_Bool_6QVal_Bool_bufchan_buf;
  assign lizzieLet0_4QNode_Bool_4QNone_Bool_6QVal_Bool_bufchan_r = (! lizzieLet0_4QNode_Bool_4QNone_Bool_6QVal_Bool_bufchan_buf[0]);
  assign lizzieLet0_4QNode_Bool_4QNone_Bool_6QVal_Bool_1_argbuf_d = (lizzieLet0_4QNode_Bool_4QNone_Bool_6QVal_Bool_bufchan_buf[0] ? lizzieLet0_4QNode_Bool_4QNone_Bool_6QVal_Bool_bufchan_buf :
                                                                     lizzieLet0_4QNode_Bool_4QNone_Bool_6QVal_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNode_Bool_4QNone_Bool_6QVal_Bool_bufchan_buf <= {16'd0,
                                                                    1'd0};
    else
      if ((lizzieLet0_4QNode_Bool_4QNone_Bool_6QVal_Bool_1_argbuf_r && lizzieLet0_4QNode_Bool_4QNone_Bool_6QVal_Bool_bufchan_buf[0]))
        lizzieLet0_4QNode_Bool_4QNone_Bool_6QVal_Bool_bufchan_buf <= {16'd0,
                                                                      1'd0};
      else if (((! lizzieLet0_4QNode_Bool_4QNone_Bool_6QVal_Bool_1_argbuf_r) && (! lizzieLet0_4QNode_Bool_4QNone_Bool_6QVal_Bool_bufchan_buf[0])))
        lizzieLet0_4QNode_Bool_4QNone_Bool_6QVal_Bool_bufchan_buf <= lizzieLet0_4QNode_Bool_4QNone_Bool_6QVal_Bool_bufchan_d;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_QTree_Bool) : (lizzieLet0_4QNode_Bool_4QNone_Bool_7,QTree_Bool) (lizzieLet0_4QNode_Bool_7QNone_Bool,Pointer_QTree_Bool) > [(_130,Pointer_QTree_Bool),
                                                                                                                                             (_129,Pointer_QTree_Bool),
                                                                                                                                             (lizzieLet0_4QNode_Bool_4QNone_Bool_7QNode_Bool,Pointer_QTree_Bool),
                                                                                                                                             (_128,Pointer_QTree_Bool)] */
  logic [3:0] lizzieLet0_4QNode_Bool_7QNone_Bool_onehotd;
  always_comb
    if ((lizzieLet0_4QNode_Bool_4QNone_Bool_7_d[0] && lizzieLet0_4QNode_Bool_7QNone_Bool_d[0]))
      unique case (lizzieLet0_4QNode_Bool_4QNone_Bool_7_d[2:1])
        2'd0: lizzieLet0_4QNode_Bool_7QNone_Bool_onehotd = 4'd1;
        2'd1: lizzieLet0_4QNode_Bool_7QNone_Bool_onehotd = 4'd2;
        2'd2: lizzieLet0_4QNode_Bool_7QNone_Bool_onehotd = 4'd4;
        2'd3: lizzieLet0_4QNode_Bool_7QNone_Bool_onehotd = 4'd8;
        default: lizzieLet0_4QNode_Bool_7QNone_Bool_onehotd = 4'd0;
      endcase
    else lizzieLet0_4QNode_Bool_7QNone_Bool_onehotd = 4'd0;
  assign _130_d = {lizzieLet0_4QNode_Bool_7QNone_Bool_d[16:1],
                   lizzieLet0_4QNode_Bool_7QNone_Bool_onehotd[0]};
  assign _129_d = {lizzieLet0_4QNode_Bool_7QNone_Bool_d[16:1],
                   lizzieLet0_4QNode_Bool_7QNone_Bool_onehotd[1]};
  assign lizzieLet0_4QNode_Bool_4QNone_Bool_7QNode_Bool_d = {lizzieLet0_4QNode_Bool_7QNone_Bool_d[16:1],
                                                             lizzieLet0_4QNode_Bool_7QNone_Bool_onehotd[2]};
  assign _128_d = {lizzieLet0_4QNode_Bool_7QNone_Bool_d[16:1],
                   lizzieLet0_4QNode_Bool_7QNone_Bool_onehotd[3]};
  assign lizzieLet0_4QNode_Bool_7QNone_Bool_r = (| (lizzieLet0_4QNode_Bool_7QNone_Bool_onehotd & {_128_r,
                                                                                                  lizzieLet0_4QNode_Bool_4QNone_Bool_7QNode_Bool_r,
                                                                                                  _129_r,
                                                                                                  _130_r}));
  assign lizzieLet0_4QNode_Bool_4QNone_Bool_7_r = lizzieLet0_4QNode_Bool_7QNone_Bool_r;
  
  /* buf (Ty Pointer_QTree_Bool) : (lizzieLet0_4QNode_Bool_4QNone_Bool_7QNode_Bool,Pointer_QTree_Bool) > (lizzieLet0_4QNode_Bool_4QNone_Bool_7QNode_Bool_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t lizzieLet0_4QNode_Bool_4QNone_Bool_7QNode_Bool_bufchan_d;
  logic lizzieLet0_4QNode_Bool_4QNone_Bool_7QNode_Bool_bufchan_r;
  assign lizzieLet0_4QNode_Bool_4QNone_Bool_7QNode_Bool_r = ((! lizzieLet0_4QNode_Bool_4QNone_Bool_7QNode_Bool_bufchan_d[0]) || lizzieLet0_4QNode_Bool_4QNone_Bool_7QNode_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNode_Bool_4QNone_Bool_7QNode_Bool_bufchan_d <= {16'd0,
                                                                   1'd0};
    else
      if (lizzieLet0_4QNode_Bool_4QNone_Bool_7QNode_Bool_r)
        lizzieLet0_4QNode_Bool_4QNone_Bool_7QNode_Bool_bufchan_d <= lizzieLet0_4QNode_Bool_4QNone_Bool_7QNode_Bool_d;
  Pointer_QTree_Bool_t lizzieLet0_4QNode_Bool_4QNone_Bool_7QNode_Bool_bufchan_buf;
  assign lizzieLet0_4QNode_Bool_4QNone_Bool_7QNode_Bool_bufchan_r = (! lizzieLet0_4QNode_Bool_4QNone_Bool_7QNode_Bool_bufchan_buf[0]);
  assign lizzieLet0_4QNode_Bool_4QNone_Bool_7QNode_Bool_1_argbuf_d = (lizzieLet0_4QNode_Bool_4QNone_Bool_7QNode_Bool_bufchan_buf[0] ? lizzieLet0_4QNode_Bool_4QNone_Bool_7QNode_Bool_bufchan_buf :
                                                                      lizzieLet0_4QNode_Bool_4QNone_Bool_7QNode_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNode_Bool_4QNone_Bool_7QNode_Bool_bufchan_buf <= {16'd0,
                                                                     1'd0};
    else
      if ((lizzieLet0_4QNode_Bool_4QNone_Bool_7QNode_Bool_1_argbuf_r && lizzieLet0_4QNode_Bool_4QNone_Bool_7QNode_Bool_bufchan_buf[0]))
        lizzieLet0_4QNode_Bool_4QNone_Bool_7QNode_Bool_bufchan_buf <= {16'd0,
                                                                       1'd0};
      else if (((! lizzieLet0_4QNode_Bool_4QNone_Bool_7QNode_Bool_1_argbuf_r) && (! lizzieLet0_4QNode_Bool_4QNone_Bool_7QNode_Bool_bufchan_buf[0])))
        lizzieLet0_4QNode_Bool_4QNone_Bool_7QNode_Bool_bufchan_buf <= lizzieLet0_4QNode_Bool_4QNone_Bool_7QNode_Bool_bufchan_d;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_QTree_Bool) : (lizzieLet0_4QNode_Bool_4QNone_Bool_8,QTree_Bool) (lizzieLet0_4QNode_Bool_8QNone_Bool,Pointer_QTree_Bool) > [(_127,Pointer_QTree_Bool),
                                                                                                                                             (_126,Pointer_QTree_Bool),
                                                                                                                                             (lizzieLet0_4QNode_Bool_4QNone_Bool_8QNode_Bool,Pointer_QTree_Bool),
                                                                                                                                             (_125,Pointer_QTree_Bool)] */
  logic [3:0] lizzieLet0_4QNode_Bool_8QNone_Bool_onehotd;
  always_comb
    if ((lizzieLet0_4QNode_Bool_4QNone_Bool_8_d[0] && lizzieLet0_4QNode_Bool_8QNone_Bool_d[0]))
      unique case (lizzieLet0_4QNode_Bool_4QNone_Bool_8_d[2:1])
        2'd0: lizzieLet0_4QNode_Bool_8QNone_Bool_onehotd = 4'd1;
        2'd1: lizzieLet0_4QNode_Bool_8QNone_Bool_onehotd = 4'd2;
        2'd2: lizzieLet0_4QNode_Bool_8QNone_Bool_onehotd = 4'd4;
        2'd3: lizzieLet0_4QNode_Bool_8QNone_Bool_onehotd = 4'd8;
        default: lizzieLet0_4QNode_Bool_8QNone_Bool_onehotd = 4'd0;
      endcase
    else lizzieLet0_4QNode_Bool_8QNone_Bool_onehotd = 4'd0;
  assign _127_d = {lizzieLet0_4QNode_Bool_8QNone_Bool_d[16:1],
                   lizzieLet0_4QNode_Bool_8QNone_Bool_onehotd[0]};
  assign _126_d = {lizzieLet0_4QNode_Bool_8QNone_Bool_d[16:1],
                   lizzieLet0_4QNode_Bool_8QNone_Bool_onehotd[1]};
  assign lizzieLet0_4QNode_Bool_4QNone_Bool_8QNode_Bool_d = {lizzieLet0_4QNode_Bool_8QNone_Bool_d[16:1],
                                                             lizzieLet0_4QNode_Bool_8QNone_Bool_onehotd[2]};
  assign _125_d = {lizzieLet0_4QNode_Bool_8QNone_Bool_d[16:1],
                   lizzieLet0_4QNode_Bool_8QNone_Bool_onehotd[3]};
  assign lizzieLet0_4QNode_Bool_8QNone_Bool_r = (| (lizzieLet0_4QNode_Bool_8QNone_Bool_onehotd & {_125_r,
                                                                                                  lizzieLet0_4QNode_Bool_4QNone_Bool_8QNode_Bool_r,
                                                                                                  _126_r,
                                                                                                  _127_r}));
  assign lizzieLet0_4QNode_Bool_4QNone_Bool_8_r = lizzieLet0_4QNode_Bool_8QNone_Bool_r;
  
  /* buf (Ty Pointer_QTree_Bool) : (lizzieLet0_4QNode_Bool_4QNone_Bool_8QNode_Bool,Pointer_QTree_Bool) > (lizzieLet0_4QNode_Bool_4QNone_Bool_8QNode_Bool_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t lizzieLet0_4QNode_Bool_4QNone_Bool_8QNode_Bool_bufchan_d;
  logic lizzieLet0_4QNode_Bool_4QNone_Bool_8QNode_Bool_bufchan_r;
  assign lizzieLet0_4QNode_Bool_4QNone_Bool_8QNode_Bool_r = ((! lizzieLet0_4QNode_Bool_4QNone_Bool_8QNode_Bool_bufchan_d[0]) || lizzieLet0_4QNode_Bool_4QNone_Bool_8QNode_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNode_Bool_4QNone_Bool_8QNode_Bool_bufchan_d <= {16'd0,
                                                                   1'd0};
    else
      if (lizzieLet0_4QNode_Bool_4QNone_Bool_8QNode_Bool_r)
        lizzieLet0_4QNode_Bool_4QNone_Bool_8QNode_Bool_bufchan_d <= lizzieLet0_4QNode_Bool_4QNone_Bool_8QNode_Bool_d;
  Pointer_QTree_Bool_t lizzieLet0_4QNode_Bool_4QNone_Bool_8QNode_Bool_bufchan_buf;
  assign lizzieLet0_4QNode_Bool_4QNone_Bool_8QNode_Bool_bufchan_r = (! lizzieLet0_4QNode_Bool_4QNone_Bool_8QNode_Bool_bufchan_buf[0]);
  assign lizzieLet0_4QNode_Bool_4QNone_Bool_8QNode_Bool_1_argbuf_d = (lizzieLet0_4QNode_Bool_4QNone_Bool_8QNode_Bool_bufchan_buf[0] ? lizzieLet0_4QNode_Bool_4QNone_Bool_8QNode_Bool_bufchan_buf :
                                                                      lizzieLet0_4QNode_Bool_4QNone_Bool_8QNode_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNode_Bool_4QNone_Bool_8QNode_Bool_bufchan_buf <= {16'd0,
                                                                     1'd0};
    else
      if ((lizzieLet0_4QNode_Bool_4QNone_Bool_8QNode_Bool_1_argbuf_r && lizzieLet0_4QNode_Bool_4QNone_Bool_8QNode_Bool_bufchan_buf[0]))
        lizzieLet0_4QNode_Bool_4QNone_Bool_8QNode_Bool_bufchan_buf <= {16'd0,
                                                                       1'd0};
      else if (((! lizzieLet0_4QNode_Bool_4QNone_Bool_8QNode_Bool_1_argbuf_r) && (! lizzieLet0_4QNode_Bool_4QNone_Bool_8QNode_Bool_bufchan_buf[0])))
        lizzieLet0_4QNode_Bool_4QNone_Bool_8QNode_Bool_bufchan_buf <= lizzieLet0_4QNode_Bool_4QNone_Bool_8QNode_Bool_bufchan_d;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_QTree_Bool) : (lizzieLet0_4QNode_Bool_4QNone_Bool_9,QTree_Bool) (lizzieLet0_4QNode_Bool_9QNone_Bool,Pointer_QTree_Bool) > [(_124,Pointer_QTree_Bool),
                                                                                                                                             (_123,Pointer_QTree_Bool),
                                                                                                                                             (lizzieLet0_4QNode_Bool_4QNone_Bool_9QNode_Bool,Pointer_QTree_Bool),
                                                                                                                                             (_122,Pointer_QTree_Bool)] */
  logic [3:0] lizzieLet0_4QNode_Bool_9QNone_Bool_onehotd;
  always_comb
    if ((lizzieLet0_4QNode_Bool_4QNone_Bool_9_d[0] && lizzieLet0_4QNode_Bool_9QNone_Bool_d[0]))
      unique case (lizzieLet0_4QNode_Bool_4QNone_Bool_9_d[2:1])
        2'd0: lizzieLet0_4QNode_Bool_9QNone_Bool_onehotd = 4'd1;
        2'd1: lizzieLet0_4QNode_Bool_9QNone_Bool_onehotd = 4'd2;
        2'd2: lizzieLet0_4QNode_Bool_9QNone_Bool_onehotd = 4'd4;
        2'd3: lizzieLet0_4QNode_Bool_9QNone_Bool_onehotd = 4'd8;
        default: lizzieLet0_4QNode_Bool_9QNone_Bool_onehotd = 4'd0;
      endcase
    else lizzieLet0_4QNode_Bool_9QNone_Bool_onehotd = 4'd0;
  assign _124_d = {lizzieLet0_4QNode_Bool_9QNone_Bool_d[16:1],
                   lizzieLet0_4QNode_Bool_9QNone_Bool_onehotd[0]};
  assign _123_d = {lizzieLet0_4QNode_Bool_9QNone_Bool_d[16:1],
                   lizzieLet0_4QNode_Bool_9QNone_Bool_onehotd[1]};
  assign lizzieLet0_4QNode_Bool_4QNone_Bool_9QNode_Bool_d = {lizzieLet0_4QNode_Bool_9QNone_Bool_d[16:1],
                                                             lizzieLet0_4QNode_Bool_9QNone_Bool_onehotd[2]};
  assign _122_d = {lizzieLet0_4QNode_Bool_9QNone_Bool_d[16:1],
                   lizzieLet0_4QNode_Bool_9QNone_Bool_onehotd[3]};
  assign lizzieLet0_4QNode_Bool_9QNone_Bool_r = (| (lizzieLet0_4QNode_Bool_9QNone_Bool_onehotd & {_122_r,
                                                                                                  lizzieLet0_4QNode_Bool_4QNone_Bool_9QNode_Bool_r,
                                                                                                  _123_r,
                                                                                                  _124_r}));
  assign lizzieLet0_4QNode_Bool_4QNone_Bool_9_r = lizzieLet0_4QNode_Bool_9QNone_Bool_r;
  
  /* buf (Ty Pointer_QTree_Bool) : (lizzieLet0_4QNode_Bool_4QNone_Bool_9QNode_Bool,Pointer_QTree_Bool) > (lizzieLet0_4QNode_Bool_4QNone_Bool_9QNode_Bool_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t lizzieLet0_4QNode_Bool_4QNone_Bool_9QNode_Bool_bufchan_d;
  logic lizzieLet0_4QNode_Bool_4QNone_Bool_9QNode_Bool_bufchan_r;
  assign lizzieLet0_4QNode_Bool_4QNone_Bool_9QNode_Bool_r = ((! lizzieLet0_4QNode_Bool_4QNone_Bool_9QNode_Bool_bufchan_d[0]) || lizzieLet0_4QNode_Bool_4QNone_Bool_9QNode_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNode_Bool_4QNone_Bool_9QNode_Bool_bufchan_d <= {16'd0,
                                                                   1'd0};
    else
      if (lizzieLet0_4QNode_Bool_4QNone_Bool_9QNode_Bool_r)
        lizzieLet0_4QNode_Bool_4QNone_Bool_9QNode_Bool_bufchan_d <= lizzieLet0_4QNode_Bool_4QNone_Bool_9QNode_Bool_d;
  Pointer_QTree_Bool_t lizzieLet0_4QNode_Bool_4QNone_Bool_9QNode_Bool_bufchan_buf;
  assign lizzieLet0_4QNode_Bool_4QNone_Bool_9QNode_Bool_bufchan_r = (! lizzieLet0_4QNode_Bool_4QNone_Bool_9QNode_Bool_bufchan_buf[0]);
  assign lizzieLet0_4QNode_Bool_4QNone_Bool_9QNode_Bool_1_argbuf_d = (lizzieLet0_4QNode_Bool_4QNone_Bool_9QNode_Bool_bufchan_buf[0] ? lizzieLet0_4QNode_Bool_4QNone_Bool_9QNode_Bool_bufchan_buf :
                                                                      lizzieLet0_4QNode_Bool_4QNone_Bool_9QNode_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNode_Bool_4QNone_Bool_9QNode_Bool_bufchan_buf <= {16'd0,
                                                                     1'd0};
    else
      if ((lizzieLet0_4QNode_Bool_4QNone_Bool_9QNode_Bool_1_argbuf_r && lizzieLet0_4QNode_Bool_4QNone_Bool_9QNode_Bool_bufchan_buf[0]))
        lizzieLet0_4QNode_Bool_4QNone_Bool_9QNode_Bool_bufchan_buf <= {16'd0,
                                                                       1'd0};
      else if (((! lizzieLet0_4QNode_Bool_4QNone_Bool_9QNode_Bool_1_argbuf_r) && (! lizzieLet0_4QNode_Bool_4QNone_Bool_9QNode_Bool_bufchan_buf[0])))
        lizzieLet0_4QNode_Bool_4QNone_Bool_9QNode_Bool_bufchan_buf <= lizzieLet0_4QNode_Bool_4QNone_Bool_9QNode_Bool_bufchan_d;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_QTree_Bool) : (lizzieLet0_4QNode_Bool_5,QTree_Bool) (lizzieLet0_6QNode_Bool,Pointer_QTree_Bool) > [(lizzieLet0_4QNode_Bool_5QNone_Bool,Pointer_QTree_Bool),
                                                                                                                     (_121,Pointer_QTree_Bool),
                                                                                                                     (_120,Pointer_QTree_Bool),
                                                                                                                     (_119,Pointer_QTree_Bool)] */
  logic [3:0] lizzieLet0_6QNode_Bool_onehotd;
  always_comb
    if ((lizzieLet0_4QNode_Bool_5_d[0] && lizzieLet0_6QNode_Bool_d[0]))
      unique case (lizzieLet0_4QNode_Bool_5_d[2:1])
        2'd0: lizzieLet0_6QNode_Bool_onehotd = 4'd1;
        2'd1: lizzieLet0_6QNode_Bool_onehotd = 4'd2;
        2'd2: lizzieLet0_6QNode_Bool_onehotd = 4'd4;
        2'd3: lizzieLet0_6QNode_Bool_onehotd = 4'd8;
        default: lizzieLet0_6QNode_Bool_onehotd = 4'd0;
      endcase
    else lizzieLet0_6QNode_Bool_onehotd = 4'd0;
  assign lizzieLet0_4QNode_Bool_5QNone_Bool_d = {lizzieLet0_6QNode_Bool_d[16:1],
                                                 lizzieLet0_6QNode_Bool_onehotd[0]};
  assign _121_d = {lizzieLet0_6QNode_Bool_d[16:1],
                   lizzieLet0_6QNode_Bool_onehotd[1]};
  assign _120_d = {lizzieLet0_6QNode_Bool_d[16:1],
                   lizzieLet0_6QNode_Bool_onehotd[2]};
  assign _119_d = {lizzieLet0_6QNode_Bool_d[16:1],
                   lizzieLet0_6QNode_Bool_onehotd[3]};
  assign lizzieLet0_6QNode_Bool_r = (| (lizzieLet0_6QNode_Bool_onehotd & {_119_r,
                                                                          _120_r,
                                                                          _121_r,
                                                                          lizzieLet0_4QNode_Bool_5QNone_Bool_r}));
  assign lizzieLet0_4QNode_Bool_5_r = lizzieLet0_6QNode_Bool_r;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_CTf) : (lizzieLet0_4QNode_Bool_6,QTree_Bool) (lizzieLet0_9QNode_Bool,Pointer_CTf) > [(lizzieLet0_4QNode_Bool_6QNone_Bool,Pointer_CTf),
                                                                                                       (lizzieLet0_4QNode_Bool_6QVal_Bool,Pointer_CTf),
                                                                                                       (lizzieLet0_4QNode_Bool_6QNode_Bool,Pointer_CTf),
                                                                                                       (lizzieLet0_4QNode_Bool_6QError_Bool,Pointer_CTf)] */
  logic [3:0] lizzieLet0_9QNode_Bool_onehotd;
  always_comb
    if ((lizzieLet0_4QNode_Bool_6_d[0] && lizzieLet0_9QNode_Bool_d[0]))
      unique case (lizzieLet0_4QNode_Bool_6_d[2:1])
        2'd0: lizzieLet0_9QNode_Bool_onehotd = 4'd1;
        2'd1: lizzieLet0_9QNode_Bool_onehotd = 4'd2;
        2'd2: lizzieLet0_9QNode_Bool_onehotd = 4'd4;
        2'd3: lizzieLet0_9QNode_Bool_onehotd = 4'd8;
        default: lizzieLet0_9QNode_Bool_onehotd = 4'd0;
      endcase
    else lizzieLet0_9QNode_Bool_onehotd = 4'd0;
  assign lizzieLet0_4QNode_Bool_6QNone_Bool_d = {lizzieLet0_9QNode_Bool_d[16:1],
                                                 lizzieLet0_9QNode_Bool_onehotd[0]};
  assign lizzieLet0_4QNode_Bool_6QVal_Bool_d = {lizzieLet0_9QNode_Bool_d[16:1],
                                                lizzieLet0_9QNode_Bool_onehotd[1]};
  assign lizzieLet0_4QNode_Bool_6QNode_Bool_d = {lizzieLet0_9QNode_Bool_d[16:1],
                                                 lizzieLet0_9QNode_Bool_onehotd[2]};
  assign lizzieLet0_4QNode_Bool_6QError_Bool_d = {lizzieLet0_9QNode_Bool_d[16:1],
                                                  lizzieLet0_9QNode_Bool_onehotd[3]};
  assign lizzieLet0_9QNode_Bool_r = (| (lizzieLet0_9QNode_Bool_onehotd & {lizzieLet0_4QNode_Bool_6QError_Bool_r,
                                                                          lizzieLet0_4QNode_Bool_6QNode_Bool_r,
                                                                          lizzieLet0_4QNode_Bool_6QVal_Bool_r,
                                                                          lizzieLet0_4QNode_Bool_6QNone_Bool_r}));
  assign lizzieLet0_4QNode_Bool_6_r = lizzieLet0_9QNode_Bool_r;
  
  /* buf (Ty Pointer_CTf) : (lizzieLet0_4QNode_Bool_6QError_Bool,Pointer_CTf) > (lizzieLet0_4QNode_Bool_6QError_Bool_1_argbuf,Pointer_CTf) */
  Pointer_CTf_t lizzieLet0_4QNode_Bool_6QError_Bool_bufchan_d;
  logic lizzieLet0_4QNode_Bool_6QError_Bool_bufchan_r;
  assign lizzieLet0_4QNode_Bool_6QError_Bool_r = ((! lizzieLet0_4QNode_Bool_6QError_Bool_bufchan_d[0]) || lizzieLet0_4QNode_Bool_6QError_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNode_Bool_6QError_Bool_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet0_4QNode_Bool_6QError_Bool_r)
        lizzieLet0_4QNode_Bool_6QError_Bool_bufchan_d <= lizzieLet0_4QNode_Bool_6QError_Bool_d;
  Pointer_CTf_t lizzieLet0_4QNode_Bool_6QError_Bool_bufchan_buf;
  assign lizzieLet0_4QNode_Bool_6QError_Bool_bufchan_r = (! lizzieLet0_4QNode_Bool_6QError_Bool_bufchan_buf[0]);
  assign lizzieLet0_4QNode_Bool_6QError_Bool_1_argbuf_d = (lizzieLet0_4QNode_Bool_6QError_Bool_bufchan_buf[0] ? lizzieLet0_4QNode_Bool_6QError_Bool_bufchan_buf :
                                                           lizzieLet0_4QNode_Bool_6QError_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNode_Bool_6QError_Bool_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet0_4QNode_Bool_6QError_Bool_1_argbuf_r && lizzieLet0_4QNode_Bool_6QError_Bool_bufchan_buf[0]))
        lizzieLet0_4QNode_Bool_6QError_Bool_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet0_4QNode_Bool_6QError_Bool_1_argbuf_r) && (! lizzieLet0_4QNode_Bool_6QError_Bool_bufchan_buf[0])))
        lizzieLet0_4QNode_Bool_6QError_Bool_bufchan_buf <= lizzieLet0_4QNode_Bool_6QError_Bool_bufchan_d;
  
  /* buf (Ty Pointer_CTf) : (lizzieLet0_4QNode_Bool_6QVal_Bool,Pointer_CTf) > (lizzieLet0_4QNode_Bool_6QVal_Bool_1_argbuf,Pointer_CTf) */
  Pointer_CTf_t lizzieLet0_4QNode_Bool_6QVal_Bool_bufchan_d;
  logic lizzieLet0_4QNode_Bool_6QVal_Bool_bufchan_r;
  assign lizzieLet0_4QNode_Bool_6QVal_Bool_r = ((! lizzieLet0_4QNode_Bool_6QVal_Bool_bufchan_d[0]) || lizzieLet0_4QNode_Bool_6QVal_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNode_Bool_6QVal_Bool_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet0_4QNode_Bool_6QVal_Bool_r)
        lizzieLet0_4QNode_Bool_6QVal_Bool_bufchan_d <= lizzieLet0_4QNode_Bool_6QVal_Bool_d;
  Pointer_CTf_t lizzieLet0_4QNode_Bool_6QVal_Bool_bufchan_buf;
  assign lizzieLet0_4QNode_Bool_6QVal_Bool_bufchan_r = (! lizzieLet0_4QNode_Bool_6QVal_Bool_bufchan_buf[0]);
  assign lizzieLet0_4QNode_Bool_6QVal_Bool_1_argbuf_d = (lizzieLet0_4QNode_Bool_6QVal_Bool_bufchan_buf[0] ? lizzieLet0_4QNode_Bool_6QVal_Bool_bufchan_buf :
                                                         lizzieLet0_4QNode_Bool_6QVal_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNode_Bool_6QVal_Bool_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet0_4QNode_Bool_6QVal_Bool_1_argbuf_r && lizzieLet0_4QNode_Bool_6QVal_Bool_bufchan_buf[0]))
        lizzieLet0_4QNode_Bool_6QVal_Bool_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet0_4QNode_Bool_6QVal_Bool_1_argbuf_r) && (! lizzieLet0_4QNode_Bool_6QVal_Bool_bufchan_buf[0])))
        lizzieLet0_4QNode_Bool_6QVal_Bool_bufchan_buf <= lizzieLet0_4QNode_Bool_6QVal_Bool_bufchan_d;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_QTree_Bool) : (lizzieLet0_4QNode_Bool_7,QTree_Bool) (q1a8H_destruct,Pointer_QTree_Bool) > [(lizzieLet0_4QNode_Bool_7QNone_Bool,Pointer_QTree_Bool),
                                                                                                             (_118,Pointer_QTree_Bool),
                                                                                                             (lizzieLet0_4QNode_Bool_7QNode_Bool,Pointer_QTree_Bool),
                                                                                                             (_117,Pointer_QTree_Bool)] */
  logic [3:0] q1a8H_destruct_onehotd;
  always_comb
    if ((lizzieLet0_4QNode_Bool_7_d[0] && q1a8H_destruct_d[0]))
      unique case (lizzieLet0_4QNode_Bool_7_d[2:1])
        2'd0: q1a8H_destruct_onehotd = 4'd1;
        2'd1: q1a8H_destruct_onehotd = 4'd2;
        2'd2: q1a8H_destruct_onehotd = 4'd4;
        2'd3: q1a8H_destruct_onehotd = 4'd8;
        default: q1a8H_destruct_onehotd = 4'd0;
      endcase
    else q1a8H_destruct_onehotd = 4'd0;
  assign lizzieLet0_4QNode_Bool_7QNone_Bool_d = {q1a8H_destruct_d[16:1],
                                                 q1a8H_destruct_onehotd[0]};
  assign _118_d = {q1a8H_destruct_d[16:1],
                   q1a8H_destruct_onehotd[1]};
  assign lizzieLet0_4QNode_Bool_7QNode_Bool_d = {q1a8H_destruct_d[16:1],
                                                 q1a8H_destruct_onehotd[2]};
  assign _117_d = {q1a8H_destruct_d[16:1],
                   q1a8H_destruct_onehotd[3]};
  assign q1a8H_destruct_r = (| (q1a8H_destruct_onehotd & {_117_r,
                                                          lizzieLet0_4QNode_Bool_7QNode_Bool_r,
                                                          _118_r,
                                                          lizzieLet0_4QNode_Bool_7QNone_Bool_r}));
  assign lizzieLet0_4QNode_Bool_7_r = q1a8H_destruct_r;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_QTree_Bool) : (lizzieLet0_4QNode_Bool_8,QTree_Bool) (q2a8I_destruct,Pointer_QTree_Bool) > [(lizzieLet0_4QNode_Bool_8QNone_Bool,Pointer_QTree_Bool),
                                                                                                             (_116,Pointer_QTree_Bool),
                                                                                                             (lizzieLet0_4QNode_Bool_8QNode_Bool,Pointer_QTree_Bool),
                                                                                                             (_115,Pointer_QTree_Bool)] */
  logic [3:0] q2a8I_destruct_onehotd;
  always_comb
    if ((lizzieLet0_4QNode_Bool_8_d[0] && q2a8I_destruct_d[0]))
      unique case (lizzieLet0_4QNode_Bool_8_d[2:1])
        2'd0: q2a8I_destruct_onehotd = 4'd1;
        2'd1: q2a8I_destruct_onehotd = 4'd2;
        2'd2: q2a8I_destruct_onehotd = 4'd4;
        2'd3: q2a8I_destruct_onehotd = 4'd8;
        default: q2a8I_destruct_onehotd = 4'd0;
      endcase
    else q2a8I_destruct_onehotd = 4'd0;
  assign lizzieLet0_4QNode_Bool_8QNone_Bool_d = {q2a8I_destruct_d[16:1],
                                                 q2a8I_destruct_onehotd[0]};
  assign _116_d = {q2a8I_destruct_d[16:1],
                   q2a8I_destruct_onehotd[1]};
  assign lizzieLet0_4QNode_Bool_8QNode_Bool_d = {q2a8I_destruct_d[16:1],
                                                 q2a8I_destruct_onehotd[2]};
  assign _115_d = {q2a8I_destruct_d[16:1],
                   q2a8I_destruct_onehotd[3]};
  assign q2a8I_destruct_r = (| (q2a8I_destruct_onehotd & {_115_r,
                                                          lizzieLet0_4QNode_Bool_8QNode_Bool_r,
                                                          _116_r,
                                                          lizzieLet0_4QNode_Bool_8QNone_Bool_r}));
  assign lizzieLet0_4QNode_Bool_8_r = q2a8I_destruct_r;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_QTree_Bool) : (lizzieLet0_4QNode_Bool_9,QTree_Bool) (q3a8J_destruct,Pointer_QTree_Bool) > [(lizzieLet0_4QNode_Bool_9QNone_Bool,Pointer_QTree_Bool),
                                                                                                             (_114,Pointer_QTree_Bool),
                                                                                                             (lizzieLet0_4QNode_Bool_9QNode_Bool,Pointer_QTree_Bool),
                                                                                                             (_113,Pointer_QTree_Bool)] */
  logic [3:0] q3a8J_destruct_onehotd;
  always_comb
    if ((lizzieLet0_4QNode_Bool_9_d[0] && q3a8J_destruct_d[0]))
      unique case (lizzieLet0_4QNode_Bool_9_d[2:1])
        2'd0: q3a8J_destruct_onehotd = 4'd1;
        2'd1: q3a8J_destruct_onehotd = 4'd2;
        2'd2: q3a8J_destruct_onehotd = 4'd4;
        2'd3: q3a8J_destruct_onehotd = 4'd8;
        default: q3a8J_destruct_onehotd = 4'd0;
      endcase
    else q3a8J_destruct_onehotd = 4'd0;
  assign lizzieLet0_4QNode_Bool_9QNone_Bool_d = {q3a8J_destruct_d[16:1],
                                                 q3a8J_destruct_onehotd[0]};
  assign _114_d = {q3a8J_destruct_d[16:1],
                   q3a8J_destruct_onehotd[1]};
  assign lizzieLet0_4QNode_Bool_9QNode_Bool_d = {q3a8J_destruct_d[16:1],
                                                 q3a8J_destruct_onehotd[2]};
  assign _113_d = {q3a8J_destruct_d[16:1],
                   q3a8J_destruct_onehotd[3]};
  assign q3a8J_destruct_r = (| (q3a8J_destruct_onehotd & {_113_r,
                                                          lizzieLet0_4QNode_Bool_9QNode_Bool_r,
                                                          _114_r,
                                                          lizzieLet0_4QNode_Bool_9QNone_Bool_r}));
  assign lizzieLet0_4QNode_Bool_9_r = q3a8J_destruct_r;
  
  /* fork (Ty QTree_Bool) : (lizzieLet0_4QNone_Bool,QTree_Bool) > [(lizzieLet0_4QNone_Bool_1,QTree_Bool),
                                                              (lizzieLet0_4QNone_Bool_2,QTree_Bool),
                                                              (lizzieLet0_4QNone_Bool_3,QTree_Bool),
                                                              (lizzieLet0_4QNone_Bool_4,QTree_Bool),
                                                              (lizzieLet0_4QNone_Bool_5,QTree_Bool),
                                                              (lizzieLet0_4QNone_Bool_6,QTree_Bool),
                                                              (lizzieLet0_4QNone_Bool_7,QTree_Bool)] */
  logic [6:0] lizzieLet0_4QNone_Bool_emitted;
  logic [6:0] lizzieLet0_4QNone_Bool_done;
  assign lizzieLet0_4QNone_Bool_1_d = {lizzieLet0_4QNone_Bool_d[66:1],
                                       (lizzieLet0_4QNone_Bool_d[0] && (! lizzieLet0_4QNone_Bool_emitted[0]))};
  assign lizzieLet0_4QNone_Bool_2_d = {lizzieLet0_4QNone_Bool_d[66:1],
                                       (lizzieLet0_4QNone_Bool_d[0] && (! lizzieLet0_4QNone_Bool_emitted[1]))};
  assign lizzieLet0_4QNone_Bool_3_d = {lizzieLet0_4QNone_Bool_d[66:1],
                                       (lizzieLet0_4QNone_Bool_d[0] && (! lizzieLet0_4QNone_Bool_emitted[2]))};
  assign lizzieLet0_4QNone_Bool_4_d = {lizzieLet0_4QNone_Bool_d[66:1],
                                       (lizzieLet0_4QNone_Bool_d[0] && (! lizzieLet0_4QNone_Bool_emitted[3]))};
  assign lizzieLet0_4QNone_Bool_5_d = {lizzieLet0_4QNone_Bool_d[66:1],
                                       (lizzieLet0_4QNone_Bool_d[0] && (! lizzieLet0_4QNone_Bool_emitted[4]))};
  assign lizzieLet0_4QNone_Bool_6_d = {lizzieLet0_4QNone_Bool_d[66:1],
                                       (lizzieLet0_4QNone_Bool_d[0] && (! lizzieLet0_4QNone_Bool_emitted[5]))};
  assign lizzieLet0_4QNone_Bool_7_d = {lizzieLet0_4QNone_Bool_d[66:1],
                                       (lizzieLet0_4QNone_Bool_d[0] && (! lizzieLet0_4QNone_Bool_emitted[6]))};
  assign lizzieLet0_4QNone_Bool_done = (lizzieLet0_4QNone_Bool_emitted | ({lizzieLet0_4QNone_Bool_7_d[0],
                                                                           lizzieLet0_4QNone_Bool_6_d[0],
                                                                           lizzieLet0_4QNone_Bool_5_d[0],
                                                                           lizzieLet0_4QNone_Bool_4_d[0],
                                                                           lizzieLet0_4QNone_Bool_3_d[0],
                                                                           lizzieLet0_4QNone_Bool_2_d[0],
                                                                           lizzieLet0_4QNone_Bool_1_d[0]} & {lizzieLet0_4QNone_Bool_7_r,
                                                                                                             lizzieLet0_4QNone_Bool_6_r,
                                                                                                             lizzieLet0_4QNone_Bool_5_r,
                                                                                                             lizzieLet0_4QNone_Bool_4_r,
                                                                                                             lizzieLet0_4QNone_Bool_3_r,
                                                                                                             lizzieLet0_4QNone_Bool_2_r,
                                                                                                             lizzieLet0_4QNone_Bool_1_r}));
  assign lizzieLet0_4QNone_Bool_r = (& lizzieLet0_4QNone_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet0_4QNone_Bool_emitted <= 7'd0;
    else
      lizzieLet0_4QNone_Bool_emitted <= (lizzieLet0_4QNone_Bool_r ? 7'd0 :
                                         lizzieLet0_4QNone_Bool_done);
  
  /* destruct (Ty QTree_Bool,
          Dcon QNode_Bool) : (lizzieLet0_4QNone_Bool_1QNode_Bool,QTree_Bool) > [(q1a8d_destruct,Pointer_QTree_Bool),
                                                                                (q2a8e_destruct,Pointer_QTree_Bool),
                                                                                (q3a8f_destruct,Pointer_QTree_Bool),
                                                                                (q4a8g_destruct,Pointer_QTree_Bool)] */
  logic [3:0] lizzieLet0_4QNone_Bool_1QNode_Bool_emitted;
  logic [3:0] lizzieLet0_4QNone_Bool_1QNode_Bool_done;
  assign q1a8d_destruct_d = {lizzieLet0_4QNone_Bool_1QNode_Bool_d[18:3],
                             (lizzieLet0_4QNone_Bool_1QNode_Bool_d[0] && (! lizzieLet0_4QNone_Bool_1QNode_Bool_emitted[0]))};
  assign q2a8e_destruct_d = {lizzieLet0_4QNone_Bool_1QNode_Bool_d[34:19],
                             (lizzieLet0_4QNone_Bool_1QNode_Bool_d[0] && (! lizzieLet0_4QNone_Bool_1QNode_Bool_emitted[1]))};
  assign q3a8f_destruct_d = {lizzieLet0_4QNone_Bool_1QNode_Bool_d[50:35],
                             (lizzieLet0_4QNone_Bool_1QNode_Bool_d[0] && (! lizzieLet0_4QNone_Bool_1QNode_Bool_emitted[2]))};
  assign q4a8g_destruct_d = {lizzieLet0_4QNone_Bool_1QNode_Bool_d[66:51],
                             (lizzieLet0_4QNone_Bool_1QNode_Bool_d[0] && (! lizzieLet0_4QNone_Bool_1QNode_Bool_emitted[3]))};
  assign lizzieLet0_4QNone_Bool_1QNode_Bool_done = (lizzieLet0_4QNone_Bool_1QNode_Bool_emitted | ({q4a8g_destruct_d[0],
                                                                                                   q3a8f_destruct_d[0],
                                                                                                   q2a8e_destruct_d[0],
                                                                                                   q1a8d_destruct_d[0]} & {q4a8g_destruct_r,
                                                                                                                           q3a8f_destruct_r,
                                                                                                                           q2a8e_destruct_r,
                                                                                                                           q1a8d_destruct_r}));
  assign lizzieLet0_4QNone_Bool_1QNode_Bool_r = (& lizzieLet0_4QNone_Bool_1QNode_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNone_Bool_1QNode_Bool_emitted <= 4'd0;
    else
      lizzieLet0_4QNone_Bool_1QNode_Bool_emitted <= (lizzieLet0_4QNone_Bool_1QNode_Bool_r ? 4'd0 :
                                                     lizzieLet0_4QNone_Bool_1QNode_Bool_done);
  
  /* destruct (Ty QTree_Bool,
          Dcon QVal_Bool) : (lizzieLet0_4QNone_Bool_1QVal_Bool,QTree_Bool) > [(v1a87_destruct,MyBool)] */
  assign v1a87_destruct_d = {lizzieLet0_4QNone_Bool_1QVal_Bool_d[3:3],
                             lizzieLet0_4QNone_Bool_1QVal_Bool_d[0]};
  assign lizzieLet0_4QNone_Bool_1QVal_Bool_r = v1a87_destruct_r;
  
  /* demux (Ty QTree_Bool,
       Ty QTree_Bool) : (lizzieLet0_4QNone_Bool_2,QTree_Bool) (lizzieLet0_4QNone_Bool_1,QTree_Bool) > [(_112,QTree_Bool),
                                                                                                       (lizzieLet0_4QNone_Bool_1QVal_Bool,QTree_Bool),
                                                                                                       (lizzieLet0_4QNone_Bool_1QNode_Bool,QTree_Bool),
                                                                                                       (_111,QTree_Bool)] */
  logic [3:0] lizzieLet0_4QNone_Bool_1_onehotd;
  always_comb
    if ((lizzieLet0_4QNone_Bool_2_d[0] && lizzieLet0_4QNone_Bool_1_d[0]))
      unique case (lizzieLet0_4QNone_Bool_2_d[2:1])
        2'd0: lizzieLet0_4QNone_Bool_1_onehotd = 4'd1;
        2'd1: lizzieLet0_4QNone_Bool_1_onehotd = 4'd2;
        2'd2: lizzieLet0_4QNone_Bool_1_onehotd = 4'd4;
        2'd3: lizzieLet0_4QNone_Bool_1_onehotd = 4'd8;
        default: lizzieLet0_4QNone_Bool_1_onehotd = 4'd0;
      endcase
    else lizzieLet0_4QNone_Bool_1_onehotd = 4'd0;
  assign _112_d = {lizzieLet0_4QNone_Bool_1_d[66:1],
                   lizzieLet0_4QNone_Bool_1_onehotd[0]};
  assign lizzieLet0_4QNone_Bool_1QVal_Bool_d = {lizzieLet0_4QNone_Bool_1_d[66:1],
                                                lizzieLet0_4QNone_Bool_1_onehotd[1]};
  assign lizzieLet0_4QNone_Bool_1QNode_Bool_d = {lizzieLet0_4QNone_Bool_1_d[66:1],
                                                 lizzieLet0_4QNone_Bool_1_onehotd[2]};
  assign _111_d = {lizzieLet0_4QNone_Bool_1_d[66:1],
                   lizzieLet0_4QNone_Bool_1_onehotd[3]};
  assign lizzieLet0_4QNone_Bool_1_r = (| (lizzieLet0_4QNone_Bool_1_onehotd & {_111_r,
                                                                              lizzieLet0_4QNone_Bool_1QNode_Bool_r,
                                                                              lizzieLet0_4QNone_Bool_1QVal_Bool_r,
                                                                              _112_r}));
  assign lizzieLet0_4QNone_Bool_2_r = lizzieLet0_4QNone_Bool_1_r;
  
  /* demux (Ty QTree_Bool,
       Ty Go) : (lizzieLet0_4QNone_Bool_3,QTree_Bool) (lizzieLet0_3QNone_Bool,Go) > [(lizzieLet0_4QNone_Bool_3QNone_Bool,Go),
                                                                                     (lizzieLet0_4QNone_Bool_3QVal_Bool,Go),
                                                                                     (lizzieLet0_4QNone_Bool_3QNode_Bool,Go),
                                                                                     (lizzieLet0_4QNone_Bool_3QError_Bool,Go)] */
  logic [3:0] lizzieLet0_3QNone_Bool_onehotd;
  always_comb
    if ((lizzieLet0_4QNone_Bool_3_d[0] && lizzieLet0_3QNone_Bool_d[0]))
      unique case (lizzieLet0_4QNone_Bool_3_d[2:1])
        2'd0: lizzieLet0_3QNone_Bool_onehotd = 4'd1;
        2'd1: lizzieLet0_3QNone_Bool_onehotd = 4'd2;
        2'd2: lizzieLet0_3QNone_Bool_onehotd = 4'd4;
        2'd3: lizzieLet0_3QNone_Bool_onehotd = 4'd8;
        default: lizzieLet0_3QNone_Bool_onehotd = 4'd0;
      endcase
    else lizzieLet0_3QNone_Bool_onehotd = 4'd0;
  assign lizzieLet0_4QNone_Bool_3QNone_Bool_d = lizzieLet0_3QNone_Bool_onehotd[0];
  assign lizzieLet0_4QNone_Bool_3QVal_Bool_d = lizzieLet0_3QNone_Bool_onehotd[1];
  assign lizzieLet0_4QNone_Bool_3QNode_Bool_d = lizzieLet0_3QNone_Bool_onehotd[2];
  assign lizzieLet0_4QNone_Bool_3QError_Bool_d = lizzieLet0_3QNone_Bool_onehotd[3];
  assign lizzieLet0_3QNone_Bool_r = (| (lizzieLet0_3QNone_Bool_onehotd & {lizzieLet0_4QNone_Bool_3QError_Bool_r,
                                                                          lizzieLet0_4QNone_Bool_3QNode_Bool_r,
                                                                          lizzieLet0_4QNone_Bool_3QVal_Bool_r,
                                                                          lizzieLet0_4QNone_Bool_3QNone_Bool_r}));
  assign lizzieLet0_4QNone_Bool_3_r = lizzieLet0_3QNone_Bool_r;
  
  /* fork (Ty Go) : (lizzieLet0_4QNone_Bool_3QError_Bool,Go) > [(lizzieLet0_4QNone_Bool_3QError_Bool_1,Go),
                                                           (lizzieLet0_4QNone_Bool_3QError_Bool_2,Go)] */
  logic [1:0] lizzieLet0_4QNone_Bool_3QError_Bool_emitted;
  logic [1:0] lizzieLet0_4QNone_Bool_3QError_Bool_done;
  assign lizzieLet0_4QNone_Bool_3QError_Bool_1_d = (lizzieLet0_4QNone_Bool_3QError_Bool_d[0] && (! lizzieLet0_4QNone_Bool_3QError_Bool_emitted[0]));
  assign lizzieLet0_4QNone_Bool_3QError_Bool_2_d = (lizzieLet0_4QNone_Bool_3QError_Bool_d[0] && (! lizzieLet0_4QNone_Bool_3QError_Bool_emitted[1]));
  assign lizzieLet0_4QNone_Bool_3QError_Bool_done = (lizzieLet0_4QNone_Bool_3QError_Bool_emitted | ({lizzieLet0_4QNone_Bool_3QError_Bool_2_d[0],
                                                                                                     lizzieLet0_4QNone_Bool_3QError_Bool_1_d[0]} & {lizzieLet0_4QNone_Bool_3QError_Bool_2_r,
                                                                                                                                                    lizzieLet0_4QNone_Bool_3QError_Bool_1_r}));
  assign lizzieLet0_4QNone_Bool_3QError_Bool_r = (& lizzieLet0_4QNone_Bool_3QError_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNone_Bool_3QError_Bool_emitted <= 2'd0;
    else
      lizzieLet0_4QNone_Bool_3QError_Bool_emitted <= (lizzieLet0_4QNone_Bool_3QError_Bool_r ? 2'd0 :
                                                      lizzieLet0_4QNone_Bool_3QError_Bool_done);
  
  /* dcon (Ty QTree_Bool,
      Dcon QError_Bool) : [(lizzieLet0_4QNone_Bool_3QError_Bool_1,Go)] > (lizzieLet0_4QNone_Bool_3QError_Bool_1QError_Bool,QTree_Bool) */
  assign lizzieLet0_4QNone_Bool_3QError_Bool_1QError_Bool_d = QError_Bool_dc((& {lizzieLet0_4QNone_Bool_3QError_Bool_1_d[0]}), lizzieLet0_4QNone_Bool_3QError_Bool_1_d);
  assign {lizzieLet0_4QNone_Bool_3QError_Bool_1_r} = {1 {(lizzieLet0_4QNone_Bool_3QError_Bool_1QError_Bool_r && lizzieLet0_4QNone_Bool_3QError_Bool_1QError_Bool_d[0])}};
  
  /* buf (Ty QTree_Bool) : (lizzieLet0_4QNone_Bool_3QError_Bool_1QError_Bool,QTree_Bool) > (lizzieLet12_1_1_argbuf,QTree_Bool) */
  QTree_Bool_t lizzieLet0_4QNone_Bool_3QError_Bool_1QError_Bool_bufchan_d;
  logic lizzieLet0_4QNone_Bool_3QError_Bool_1QError_Bool_bufchan_r;
  assign lizzieLet0_4QNone_Bool_3QError_Bool_1QError_Bool_r = ((! lizzieLet0_4QNone_Bool_3QError_Bool_1QError_Bool_bufchan_d[0]) || lizzieLet0_4QNone_Bool_3QError_Bool_1QError_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNone_Bool_3QError_Bool_1QError_Bool_bufchan_d <= {66'd0,
                                                                     1'd0};
    else
      if (lizzieLet0_4QNone_Bool_3QError_Bool_1QError_Bool_r)
        lizzieLet0_4QNone_Bool_3QError_Bool_1QError_Bool_bufchan_d <= lizzieLet0_4QNone_Bool_3QError_Bool_1QError_Bool_d;
  QTree_Bool_t lizzieLet0_4QNone_Bool_3QError_Bool_1QError_Bool_bufchan_buf;
  assign lizzieLet0_4QNone_Bool_3QError_Bool_1QError_Bool_bufchan_r = (! lizzieLet0_4QNone_Bool_3QError_Bool_1QError_Bool_bufchan_buf[0]);
  assign lizzieLet12_1_1_argbuf_d = (lizzieLet0_4QNone_Bool_3QError_Bool_1QError_Bool_bufchan_buf[0] ? lizzieLet0_4QNone_Bool_3QError_Bool_1QError_Bool_bufchan_buf :
                                     lizzieLet0_4QNone_Bool_3QError_Bool_1QError_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNone_Bool_3QError_Bool_1QError_Bool_bufchan_buf <= {66'd0,
                                                                       1'd0};
    else
      if ((lizzieLet12_1_1_argbuf_r && lizzieLet0_4QNone_Bool_3QError_Bool_1QError_Bool_bufchan_buf[0]))
        lizzieLet0_4QNone_Bool_3QError_Bool_1QError_Bool_bufchan_buf <= {66'd0,
                                                                         1'd0};
      else if (((! lizzieLet12_1_1_argbuf_r) && (! lizzieLet0_4QNone_Bool_3QError_Bool_1QError_Bool_bufchan_buf[0])))
        lizzieLet0_4QNone_Bool_3QError_Bool_1QError_Bool_bufchan_buf <= lizzieLet0_4QNone_Bool_3QError_Bool_1QError_Bool_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet0_4QNone_Bool_3QError_Bool_2,Go) > (lizzieLet0_4QNone_Bool_3QError_Bool_2_argbuf,Go) */
  Go_t lizzieLet0_4QNone_Bool_3QError_Bool_2_bufchan_d;
  logic lizzieLet0_4QNone_Bool_3QError_Bool_2_bufchan_r;
  assign lizzieLet0_4QNone_Bool_3QError_Bool_2_r = ((! lizzieLet0_4QNone_Bool_3QError_Bool_2_bufchan_d[0]) || lizzieLet0_4QNone_Bool_3QError_Bool_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNone_Bool_3QError_Bool_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet0_4QNone_Bool_3QError_Bool_2_r)
        lizzieLet0_4QNone_Bool_3QError_Bool_2_bufchan_d <= lizzieLet0_4QNone_Bool_3QError_Bool_2_d;
  Go_t lizzieLet0_4QNone_Bool_3QError_Bool_2_bufchan_buf;
  assign lizzieLet0_4QNone_Bool_3QError_Bool_2_bufchan_r = (! lizzieLet0_4QNone_Bool_3QError_Bool_2_bufchan_buf[0]);
  assign lizzieLet0_4QNone_Bool_3QError_Bool_2_argbuf_d = (lizzieLet0_4QNone_Bool_3QError_Bool_2_bufchan_buf[0] ? lizzieLet0_4QNone_Bool_3QError_Bool_2_bufchan_buf :
                                                           lizzieLet0_4QNone_Bool_3QError_Bool_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNone_Bool_3QError_Bool_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet0_4QNone_Bool_3QError_Bool_2_argbuf_r && lizzieLet0_4QNone_Bool_3QError_Bool_2_bufchan_buf[0]))
        lizzieLet0_4QNone_Bool_3QError_Bool_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet0_4QNone_Bool_3QError_Bool_2_argbuf_r) && (! lizzieLet0_4QNone_Bool_3QError_Bool_2_bufchan_buf[0])))
        lizzieLet0_4QNone_Bool_3QError_Bool_2_bufchan_buf <= lizzieLet0_4QNone_Bool_3QError_Bool_2_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet0_4QNone_Bool_3QNone_Bool,Go) > (lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf,Go) */
  Go_t lizzieLet0_4QNone_Bool_3QNone_Bool_bufchan_d;
  logic lizzieLet0_4QNone_Bool_3QNone_Bool_bufchan_r;
  assign lizzieLet0_4QNone_Bool_3QNone_Bool_r = ((! lizzieLet0_4QNone_Bool_3QNone_Bool_bufchan_d[0]) || lizzieLet0_4QNone_Bool_3QNone_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNone_Bool_3QNone_Bool_bufchan_d <= 1'd0;
    else
      if (lizzieLet0_4QNone_Bool_3QNone_Bool_r)
        lizzieLet0_4QNone_Bool_3QNone_Bool_bufchan_d <= lizzieLet0_4QNone_Bool_3QNone_Bool_d;
  Go_t lizzieLet0_4QNone_Bool_3QNone_Bool_bufchan_buf;
  assign lizzieLet0_4QNone_Bool_3QNone_Bool_bufchan_r = (! lizzieLet0_4QNone_Bool_3QNone_Bool_bufchan_buf[0]);
  assign lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_d = (lizzieLet0_4QNone_Bool_3QNone_Bool_bufchan_buf[0] ? lizzieLet0_4QNone_Bool_3QNone_Bool_bufchan_buf :
                                                          lizzieLet0_4QNone_Bool_3QNone_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNone_Bool_3QNone_Bool_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_r && lizzieLet0_4QNone_Bool_3QNone_Bool_bufchan_buf[0]))
        lizzieLet0_4QNone_Bool_3QNone_Bool_bufchan_buf <= 1'd0;
      else if (((! lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_r) && (! lizzieLet0_4QNone_Bool_3QNone_Bool_bufchan_buf[0])))
        lizzieLet0_4QNone_Bool_3QNone_Bool_bufchan_buf <= lizzieLet0_4QNone_Bool_3QNone_Bool_bufchan_d;
  
  /* mergectrl (Ty C40,
           Ty Go) : [(lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf,Go),
                     (lizzieLet60_3Lcall_f0_1_argbuf,Go),
                     (lizzieLet0_4QNone_Bool_4QVal_Bool_3QNone_Bool_1_argbuf,Go),
                     (lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_argbuf,Go),
                     (lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_argbuf,Go),
                     (lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyTrue_2_argbuf,Go),
                     (lizzieLet0_4QNone_Bool_4QVal_Bool_3QNode_Bool_2_argbuf,Go),
                     (lizzieLet0_4QNone_Bool_4QVal_Bool_3QError_Bool_2_argbuf,Go),
                     (lizzieLet0_4QNone_Bool_4QNode_Bool_3QNone_Bool_1_argbuf,Go),
                     (lizzieLet0_4QNone_Bool_4QNode_Bool_3QVal_Bool_2_argbuf,Go),
                     (lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_5_argbuf,Go),
                     (lizzieLet0_4QNone_Bool_4QNode_Bool_3QError_Bool_2_argbuf,Go),
                     (lizzieLet0_4QNone_Bool_3QError_Bool_2_argbuf,Go),
                     (lizzieLet0_4QVal_Bool_4QNone_Bool_3QNone_Bool_1_argbuf,Go),
                     (lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_argbuf,Go),
                     (lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_argbuf,Go),
                     (lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyTrue_2_argbuf,Go),
                     (lizzieLet0_4QVal_Bool_4QNone_Bool_3QNode_Bool_2_argbuf,Go),
                     (lizzieLet0_4QVal_Bool_4QNone_Bool_3QError_Bool_2_argbuf,Go),
                     (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_1MyFalse_1_argbuf,Go),
                     (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNone_Bool_2_argbuf,Go),
                     (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QVal_Bool_2_argbuf,Go),
                     (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNode_Bool_2_argbuf,Go),
                     (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QError_Bool_2_argbuf,Go),
                     (lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNone_Bool_2_argbuf,Go),
                     (lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QVal_Bool_2_argbuf,Go),
                     (lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNode_Bool_2_argbuf,Go),
                     (lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QError_Bool_2_argbuf,Go),
                     (lizzieLet0_4QVal_Bool_3QNode_Bool_2_argbuf,Go),
                     (lizzieLet0_4QVal_Bool_3QError_Bool_2_argbuf,Go),
                     (lizzieLet0_4QNode_Bool_4QNone_Bool_4QNone_Bool_1_argbuf,Go),
                     (lizzieLet0_4QNode_Bool_4QNone_Bool_4QVal_Bool_2_argbuf,Go),
                     (lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_5_argbuf,Go),
                     (lizzieLet0_4QNode_Bool_4QNone_Bool_4QError_Bool_2_argbuf,Go),
                     (lizzieLet0_4QNode_Bool_3QVal_Bool_2_argbuf,Go),
                     (lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_5_argbuf,Go),
                     (lizzieLet0_4QNode_Bool_4QNode_Bool_4QVal_Bool_2_argbuf,Go),
                     (lizzieLet0_4QNode_Bool_4QNode_Bool_4QError_Bool_2_argbuf,Go),
                     (lizzieLet0_4QNode_Bool_3QError_Bool_2_argbuf,Go),
                     (lizzieLet0_3QError_Bool_2_argbuf,Go)] > (go_7_goMux_choice,C40) (go_7_goMux_data,Go) */
  logic [39:0] lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_select_d;
  assign lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_select_d = ((| lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_select_q) ? lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_select_q :
                                                                 (lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_d[0] ? 40'd1 :
                                                                  (lizzieLet60_3Lcall_f0_1_argbuf_d[0] ? 40'd2 :
                                                                   (lizzieLet0_4QNone_Bool_4QVal_Bool_3QNone_Bool_1_argbuf_d[0] ? 40'd4 :
                                                                    (lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_argbuf_d[0] ? 40'd8 :
                                                                     (lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_argbuf_d[0] ? 40'd16 :
                                                                      (lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyTrue_2_argbuf_d[0] ? 40'd32 :
                                                                       (lizzieLet0_4QNone_Bool_4QVal_Bool_3QNode_Bool_2_argbuf_d[0] ? 40'd64 :
                                                                        (lizzieLet0_4QNone_Bool_4QVal_Bool_3QError_Bool_2_argbuf_d[0] ? 40'd128 :
                                                                         (lizzieLet0_4QNone_Bool_4QNode_Bool_3QNone_Bool_1_argbuf_d[0] ? 40'd256 :
                                                                          (lizzieLet0_4QNone_Bool_4QNode_Bool_3QVal_Bool_2_argbuf_d[0] ? 40'd512 :
                                                                           (lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_5_argbuf_d[0] ? 40'd1024 :
                                                                            (lizzieLet0_4QNone_Bool_4QNode_Bool_3QError_Bool_2_argbuf_d[0] ? 40'd2048 :
                                                                             (lizzieLet0_4QNone_Bool_3QError_Bool_2_argbuf_d[0] ? 40'd4096 :
                                                                              (lizzieLet0_4QVal_Bool_4QNone_Bool_3QNone_Bool_1_argbuf_d[0] ? 40'd8192 :
                                                                               (lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_argbuf_d[0] ? 40'd16384 :
                                                                                (lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_argbuf_d[0] ? 40'd32768 :
                                                                                 (lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyTrue_2_argbuf_d[0] ? 40'd65536 :
                                                                                  (lizzieLet0_4QVal_Bool_4QNone_Bool_3QNode_Bool_2_argbuf_d[0] ? 40'd131072 :
                                                                                   (lizzieLet0_4QVal_Bool_4QNone_Bool_3QError_Bool_2_argbuf_d[0] ? 40'd262144 :
                                                                                    (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_1MyFalse_1_argbuf_d[0] ? 40'd524288 :
                                                                                     (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNone_Bool_2_argbuf_d[0] ? 40'd1048576 :
                                                                                      (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QVal_Bool_2_argbuf_d[0] ? 40'd2097152 :
                                                                                       (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNode_Bool_2_argbuf_d[0] ? 40'd4194304 :
                                                                                        (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QError_Bool_2_argbuf_d[0] ? 40'd8388608 :
                                                                                         (lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNone_Bool_2_argbuf_d[0] ? 40'd16777216 :
                                                                                          (lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QVal_Bool_2_argbuf_d[0] ? 40'd33554432 :
                                                                                           (lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNode_Bool_2_argbuf_d[0] ? 40'd67108864 :
                                                                                            (lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QError_Bool_2_argbuf_d[0] ? 40'd134217728 :
                                                                                             (lizzieLet0_4QVal_Bool_3QNode_Bool_2_argbuf_d[0] ? 40'd268435456 :
                                                                                              (lizzieLet0_4QVal_Bool_3QError_Bool_2_argbuf_d[0] ? 40'd536870912 :
                                                                                               (lizzieLet0_4QNode_Bool_4QNone_Bool_4QNone_Bool_1_argbuf_d[0] ? 40'd1073741824 :
                                                                                                (lizzieLet0_4QNode_Bool_4QNone_Bool_4QVal_Bool_2_argbuf_d[0] ? 40'd2147483648 :
                                                                                                 (lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_5_argbuf_d[0] ? 40'd4294967296 :
                                                                                                  (lizzieLet0_4QNode_Bool_4QNone_Bool_4QError_Bool_2_argbuf_d[0] ? 40'd8589934592 :
                                                                                                   (lizzieLet0_4QNode_Bool_3QVal_Bool_2_argbuf_d[0] ? 40'd17179869184 :
                                                                                                    (lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_5_argbuf_d[0] ? 40'd34359738368 :
                                                                                                     (lizzieLet0_4QNode_Bool_4QNode_Bool_4QVal_Bool_2_argbuf_d[0] ? 40'd68719476736 :
                                                                                                      (lizzieLet0_4QNode_Bool_4QNode_Bool_4QError_Bool_2_argbuf_d[0] ? 40'd137438953472 :
                                                                                                       (lizzieLet0_4QNode_Bool_3QError_Bool_2_argbuf_d[0] ? 40'd274877906944 :
                                                                                                        (lizzieLet0_3QError_Bool_2_argbuf_d[0] ? 40'd549755813888 :
                                                                                                         40'd0)))))))))))))))))))))))))))))))))))))))));
  logic [39:0] lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_select_q <= 40'd0;
    else
      lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_select_q <= (lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_done ? 40'd0 :
                                                               lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_select_d);
  logic [1:0] lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_emit_q <= 2'd0;
    else
      lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_emit_q <= (lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_done ? 2'd0 :
                                                             lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_emit_d);
  logic [1:0] lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_emit_d;
  assign lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_emit_d = (lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_emit_q | ({go_7_goMux_choice_d[0],
                                                                                                                      go_7_goMux_data_d[0]} & {go_7_goMux_choice_r,
                                                                                                                                               go_7_goMux_data_r}));
  logic lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_done;
  assign lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_done = (& lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_emit_d);
  assign {lizzieLet0_3QError_Bool_2_argbuf_r,
          lizzieLet0_4QNode_Bool_3QError_Bool_2_argbuf_r,
          lizzieLet0_4QNode_Bool_4QNode_Bool_4QError_Bool_2_argbuf_r,
          lizzieLet0_4QNode_Bool_4QNode_Bool_4QVal_Bool_2_argbuf_r,
          lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_5_argbuf_r,
          lizzieLet0_4QNode_Bool_3QVal_Bool_2_argbuf_r,
          lizzieLet0_4QNode_Bool_4QNone_Bool_4QError_Bool_2_argbuf_r,
          lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_5_argbuf_r,
          lizzieLet0_4QNode_Bool_4QNone_Bool_4QVal_Bool_2_argbuf_r,
          lizzieLet0_4QNode_Bool_4QNone_Bool_4QNone_Bool_1_argbuf_r,
          lizzieLet0_4QVal_Bool_3QError_Bool_2_argbuf_r,
          lizzieLet0_4QVal_Bool_3QNode_Bool_2_argbuf_r,
          lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QError_Bool_2_argbuf_r,
          lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNode_Bool_2_argbuf_r,
          lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QVal_Bool_2_argbuf_r,
          lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNone_Bool_2_argbuf_r,
          lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QError_Bool_2_argbuf_r,
          lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNode_Bool_2_argbuf_r,
          lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QVal_Bool_2_argbuf_r,
          lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNone_Bool_2_argbuf_r,
          lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_1MyFalse_1_argbuf_r,
          lizzieLet0_4QVal_Bool_4QNone_Bool_3QError_Bool_2_argbuf_r,
          lizzieLet0_4QVal_Bool_4QNone_Bool_3QNode_Bool_2_argbuf_r,
          lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyTrue_2_argbuf_r,
          lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_argbuf_r,
          lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_argbuf_r,
          lizzieLet0_4QVal_Bool_4QNone_Bool_3QNone_Bool_1_argbuf_r,
          lizzieLet0_4QNone_Bool_3QError_Bool_2_argbuf_r,
          lizzieLet0_4QNone_Bool_4QNode_Bool_3QError_Bool_2_argbuf_r,
          lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_5_argbuf_r,
          lizzieLet0_4QNone_Bool_4QNode_Bool_3QVal_Bool_2_argbuf_r,
          lizzieLet0_4QNone_Bool_4QNode_Bool_3QNone_Bool_1_argbuf_r,
          lizzieLet0_4QNone_Bool_4QVal_Bool_3QError_Bool_2_argbuf_r,
          lizzieLet0_4QNone_Bool_4QVal_Bool_3QNode_Bool_2_argbuf_r,
          lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyTrue_2_argbuf_r,
          lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_argbuf_r,
          lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_argbuf_r,
          lizzieLet0_4QNone_Bool_4QVal_Bool_3QNone_Bool_1_argbuf_r,
          lizzieLet60_3Lcall_f0_1_argbuf_r,
          lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_r} = (lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_done ? lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_select_d :
                                                            40'd0);
  assign go_7_goMux_data_d = ((lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_select_d[0] && (! lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_emit_q[0])) ? lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_d :
                              ((lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_select_d[1] && (! lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_emit_q[0])) ? lizzieLet60_3Lcall_f0_1_argbuf_d :
                               ((lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_select_d[2] && (! lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_emit_q[0])) ? lizzieLet0_4QNone_Bool_4QVal_Bool_3QNone_Bool_1_argbuf_d :
                                ((lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_select_d[3] && (! lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_emit_q[0])) ? lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_argbuf_d :
                                 ((lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_select_d[4] && (! lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_emit_q[0])) ? lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_argbuf_d :
                                  ((lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_select_d[5] && (! lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_emit_q[0])) ? lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyTrue_2_argbuf_d :
                                   ((lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_select_d[6] && (! lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_emit_q[0])) ? lizzieLet0_4QNone_Bool_4QVal_Bool_3QNode_Bool_2_argbuf_d :
                                    ((lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_select_d[7] && (! lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_emit_q[0])) ? lizzieLet0_4QNone_Bool_4QVal_Bool_3QError_Bool_2_argbuf_d :
                                     ((lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_select_d[8] && (! lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_emit_q[0])) ? lizzieLet0_4QNone_Bool_4QNode_Bool_3QNone_Bool_1_argbuf_d :
                                      ((lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_select_d[9] && (! lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_emit_q[0])) ? lizzieLet0_4QNone_Bool_4QNode_Bool_3QVal_Bool_2_argbuf_d :
                                       ((lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_select_d[10] && (! lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_emit_q[0])) ? lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_5_argbuf_d :
                                        ((lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_select_d[11] && (! lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_emit_q[0])) ? lizzieLet0_4QNone_Bool_4QNode_Bool_3QError_Bool_2_argbuf_d :
                                         ((lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_select_d[12] && (! lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_emit_q[0])) ? lizzieLet0_4QNone_Bool_3QError_Bool_2_argbuf_d :
                                          ((lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_select_d[13] && (! lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_emit_q[0])) ? lizzieLet0_4QVal_Bool_4QNone_Bool_3QNone_Bool_1_argbuf_d :
                                           ((lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_select_d[14] && (! lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_emit_q[0])) ? lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_argbuf_d :
                                            ((lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_select_d[15] && (! lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_emit_q[0])) ? lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_argbuf_d :
                                             ((lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_select_d[16] && (! lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_emit_q[0])) ? lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyTrue_2_argbuf_d :
                                              ((lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_select_d[17] && (! lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_emit_q[0])) ? lizzieLet0_4QVal_Bool_4QNone_Bool_3QNode_Bool_2_argbuf_d :
                                               ((lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_select_d[18] && (! lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_emit_q[0])) ? lizzieLet0_4QVal_Bool_4QNone_Bool_3QError_Bool_2_argbuf_d :
                                                ((lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_select_d[19] && (! lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_emit_q[0])) ? lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_1MyFalse_1_argbuf_d :
                                                 ((lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_select_d[20] && (! lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_emit_q[0])) ? lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNone_Bool_2_argbuf_d :
                                                  ((lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_select_d[21] && (! lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_emit_q[0])) ? lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QVal_Bool_2_argbuf_d :
                                                   ((lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_select_d[22] && (! lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_emit_q[0])) ? lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNode_Bool_2_argbuf_d :
                                                    ((lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_select_d[23] && (! lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_emit_q[0])) ? lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QError_Bool_2_argbuf_d :
                                                     ((lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_select_d[24] && (! lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_emit_q[0])) ? lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNone_Bool_2_argbuf_d :
                                                      ((lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_select_d[25] && (! lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_emit_q[0])) ? lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QVal_Bool_2_argbuf_d :
                                                       ((lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_select_d[26] && (! lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_emit_q[0])) ? lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNode_Bool_2_argbuf_d :
                                                        ((lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_select_d[27] && (! lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_emit_q[0])) ? lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QError_Bool_2_argbuf_d :
                                                         ((lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_select_d[28] && (! lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_emit_q[0])) ? lizzieLet0_4QVal_Bool_3QNode_Bool_2_argbuf_d :
                                                          ((lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_select_d[29] && (! lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_emit_q[0])) ? lizzieLet0_4QVal_Bool_3QError_Bool_2_argbuf_d :
                                                           ((lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_select_d[30] && (! lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_emit_q[0])) ? lizzieLet0_4QNode_Bool_4QNone_Bool_4QNone_Bool_1_argbuf_d :
                                                            ((lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_select_d[31] && (! lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_emit_q[0])) ? lizzieLet0_4QNode_Bool_4QNone_Bool_4QVal_Bool_2_argbuf_d :
                                                             ((lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_select_d[32] && (! lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_emit_q[0])) ? lizzieLet0_4QNode_Bool_4QNone_Bool_4QNode_Bool_5_argbuf_d :
                                                              ((lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_select_d[33] && (! lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_emit_q[0])) ? lizzieLet0_4QNode_Bool_4QNone_Bool_4QError_Bool_2_argbuf_d :
                                                               ((lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_select_d[34] && (! lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_emit_q[0])) ? lizzieLet0_4QNode_Bool_3QVal_Bool_2_argbuf_d :
                                                                ((lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_select_d[35] && (! lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_emit_q[0])) ? lizzieLet0_4QNode_Bool_4QNode_Bool_4QNone_Bool_5_argbuf_d :
                                                                 ((lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_select_d[36] && (! lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_emit_q[0])) ? lizzieLet0_4QNode_Bool_4QNode_Bool_4QVal_Bool_2_argbuf_d :
                                                                  ((lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_select_d[37] && (! lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_emit_q[0])) ? lizzieLet0_4QNode_Bool_4QNode_Bool_4QError_Bool_2_argbuf_d :
                                                                   ((lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_select_d[38] && (! lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_emit_q[0])) ? lizzieLet0_4QNode_Bool_3QError_Bool_2_argbuf_d :
                                                                    ((lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_select_d[39] && (! lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_emit_q[0])) ? lizzieLet0_3QError_Bool_2_argbuf_d :
                                                                     1'd0))))))))))))))))))))))))))))))))))))))));
  assign go_7_goMux_choice_d = ((lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_select_d[0] && (! lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_emit_q[1])) ? C1_40_dc(1'd1) :
                                ((lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_select_d[1] && (! lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_emit_q[1])) ? C2_40_dc(1'd1) :
                                 ((lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_select_d[2] && (! lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_emit_q[1])) ? C3_40_dc(1'd1) :
                                  ((lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_select_d[3] && (! lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_emit_q[1])) ? C4_40_dc(1'd1) :
                                   ((lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_select_d[4] && (! lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_emit_q[1])) ? C5_40_dc(1'd1) :
                                    ((lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_select_d[5] && (! lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_emit_q[1])) ? C6_40_dc(1'd1) :
                                     ((lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_select_d[6] && (! lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_emit_q[1])) ? C7_40_dc(1'd1) :
                                      ((lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_select_d[7] && (! lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_emit_q[1])) ? C8_40_dc(1'd1) :
                                       ((lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_select_d[8] && (! lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_emit_q[1])) ? C9_40_dc(1'd1) :
                                        ((lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_select_d[9] && (! lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_emit_q[1])) ? C10_40_dc(1'd1) :
                                         ((lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_select_d[10] && (! lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_emit_q[1])) ? C11_40_dc(1'd1) :
                                          ((lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_select_d[11] && (! lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_emit_q[1])) ? C12_40_dc(1'd1) :
                                           ((lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_select_d[12] && (! lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_emit_q[1])) ? C13_40_dc(1'd1) :
                                            ((lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_select_d[13] && (! lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_emit_q[1])) ? C14_40_dc(1'd1) :
                                             ((lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_select_d[14] && (! lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_emit_q[1])) ? C15_40_dc(1'd1) :
                                              ((lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_select_d[15] && (! lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_emit_q[1])) ? C16_40_dc(1'd1) :
                                               ((lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_select_d[16] && (! lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_emit_q[1])) ? C17_40_dc(1'd1) :
                                                ((lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_select_d[17] && (! lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_emit_q[1])) ? C18_40_dc(1'd1) :
                                                 ((lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_select_d[18] && (! lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_emit_q[1])) ? C19_40_dc(1'd1) :
                                                  ((lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_select_d[19] && (! lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_emit_q[1])) ? C20_40_dc(1'd1) :
                                                   ((lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_select_d[20] && (! lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_emit_q[1])) ? C21_40_dc(1'd1) :
                                                    ((lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_select_d[21] && (! lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_emit_q[1])) ? C22_40_dc(1'd1) :
                                                     ((lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_select_d[22] && (! lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_emit_q[1])) ? C23_40_dc(1'd1) :
                                                      ((lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_select_d[23] && (! lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_emit_q[1])) ? C24_40_dc(1'd1) :
                                                       ((lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_select_d[24] && (! lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_emit_q[1])) ? C25_40_dc(1'd1) :
                                                        ((lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_select_d[25] && (! lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_emit_q[1])) ? C26_40_dc(1'd1) :
                                                         ((lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_select_d[26] && (! lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_emit_q[1])) ? C27_40_dc(1'd1) :
                                                          ((lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_select_d[27] && (! lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_emit_q[1])) ? C28_40_dc(1'd1) :
                                                           ((lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_select_d[28] && (! lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_emit_q[1])) ? C29_40_dc(1'd1) :
                                                            ((lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_select_d[29] && (! lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_emit_q[1])) ? C30_40_dc(1'd1) :
                                                             ((lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_select_d[30] && (! lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_emit_q[1])) ? C31_40_dc(1'd1) :
                                                              ((lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_select_d[31] && (! lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_emit_q[1])) ? C32_40_dc(1'd1) :
                                                               ((lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_select_d[32] && (! lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_emit_q[1])) ? C33_40_dc(1'd1) :
                                                                ((lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_select_d[33] && (! lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_emit_q[1])) ? C34_40_dc(1'd1) :
                                                                 ((lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_select_d[34] && (! lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_emit_q[1])) ? C35_40_dc(1'd1) :
                                                                  ((lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_select_d[35] && (! lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_emit_q[1])) ? C36_40_dc(1'd1) :
                                                                   ((lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_select_d[36] && (! lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_emit_q[1])) ? C37_40_dc(1'd1) :
                                                                    ((lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_select_d[37] && (! lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_emit_q[1])) ? C38_40_dc(1'd1) :
                                                                     ((lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_select_d[38] && (! lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_emit_q[1])) ? C39_40_dc(1'd1) :
                                                                      ((lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_select_d[39] && (! lizzieLet0_4QNone_Bool_3QNone_Bool_1_argbuf_emit_q[1])) ? C40_40_dc(1'd1) :
                                                                       {6'd0,
                                                                        1'd0}))))))))))))))))))))))))))))))))))))))));
  
  /* demux (Ty QTree_Bool,
       Ty QTree_Bool) : (lizzieLet0_4QNone_Bool_4,QTree_Bool) (lizzieLet0_5QNone_Bool,QTree_Bool) > [(_110,QTree_Bool),
                                                                                                     (lizzieLet0_4QNone_Bool_4QVal_Bool,QTree_Bool),
                                                                                                     (lizzieLet0_4QNone_Bool_4QNode_Bool,QTree_Bool),
                                                                                                     (_109,QTree_Bool)] */
  logic [3:0] lizzieLet0_5QNone_Bool_onehotd;
  always_comb
    if ((lizzieLet0_4QNone_Bool_4_d[0] && lizzieLet0_5QNone_Bool_d[0]))
      unique case (lizzieLet0_4QNone_Bool_4_d[2:1])
        2'd0: lizzieLet0_5QNone_Bool_onehotd = 4'd1;
        2'd1: lizzieLet0_5QNone_Bool_onehotd = 4'd2;
        2'd2: lizzieLet0_5QNone_Bool_onehotd = 4'd4;
        2'd3: lizzieLet0_5QNone_Bool_onehotd = 4'd8;
        default: lizzieLet0_5QNone_Bool_onehotd = 4'd0;
      endcase
    else lizzieLet0_5QNone_Bool_onehotd = 4'd0;
  assign _110_d = {lizzieLet0_5QNone_Bool_d[66:1],
                   lizzieLet0_5QNone_Bool_onehotd[0]};
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_d = {lizzieLet0_5QNone_Bool_d[66:1],
                                                lizzieLet0_5QNone_Bool_onehotd[1]};
  assign lizzieLet0_4QNone_Bool_4QNode_Bool_d = {lizzieLet0_5QNone_Bool_d[66:1],
                                                 lizzieLet0_5QNone_Bool_onehotd[2]};
  assign _109_d = {lizzieLet0_5QNone_Bool_d[66:1],
                   lizzieLet0_5QNone_Bool_onehotd[3]};
  assign lizzieLet0_5QNone_Bool_r = (| (lizzieLet0_5QNone_Bool_onehotd & {_109_r,
                                                                          lizzieLet0_4QNone_Bool_4QNode_Bool_r,
                                                                          lizzieLet0_4QNone_Bool_4QVal_Bool_r,
                                                                          _110_r}));
  assign lizzieLet0_4QNone_Bool_4_r = lizzieLet0_5QNone_Bool_r;
  
  /* fork (Ty QTree_Bool) : (lizzieLet0_4QNone_Bool_4QNode_Bool,QTree_Bool) > [(lizzieLet0_4QNone_Bool_4QNode_Bool_1,QTree_Bool),
                                                                          (lizzieLet0_4QNone_Bool_4QNode_Bool_2,QTree_Bool),
                                                                          (lizzieLet0_4QNone_Bool_4QNode_Bool_3,QTree_Bool),
                                                                          (lizzieLet0_4QNone_Bool_4QNode_Bool_4,QTree_Bool),
                                                                          (lizzieLet0_4QNone_Bool_4QNode_Bool_5,QTree_Bool),
                                                                          (lizzieLet0_4QNone_Bool_4QNode_Bool_6,QTree_Bool),
                                                                          (lizzieLet0_4QNone_Bool_4QNode_Bool_7,QTree_Bool),
                                                                          (lizzieLet0_4QNone_Bool_4QNode_Bool_8,QTree_Bool),
                                                                          (lizzieLet0_4QNone_Bool_4QNode_Bool_9,QTree_Bool)] */
  logic [8:0] lizzieLet0_4QNone_Bool_4QNode_Bool_emitted;
  logic [8:0] lizzieLet0_4QNone_Bool_4QNode_Bool_done;
  assign lizzieLet0_4QNone_Bool_4QNode_Bool_1_d = {lizzieLet0_4QNone_Bool_4QNode_Bool_d[66:1],
                                                   (lizzieLet0_4QNone_Bool_4QNode_Bool_d[0] && (! lizzieLet0_4QNone_Bool_4QNode_Bool_emitted[0]))};
  assign lizzieLet0_4QNone_Bool_4QNode_Bool_2_d = {lizzieLet0_4QNone_Bool_4QNode_Bool_d[66:1],
                                                   (lizzieLet0_4QNone_Bool_4QNode_Bool_d[0] && (! lizzieLet0_4QNone_Bool_4QNode_Bool_emitted[1]))};
  assign lizzieLet0_4QNone_Bool_4QNode_Bool_3_d = {lizzieLet0_4QNone_Bool_4QNode_Bool_d[66:1],
                                                   (lizzieLet0_4QNone_Bool_4QNode_Bool_d[0] && (! lizzieLet0_4QNone_Bool_4QNode_Bool_emitted[2]))};
  assign lizzieLet0_4QNone_Bool_4QNode_Bool_4_d = {lizzieLet0_4QNone_Bool_4QNode_Bool_d[66:1],
                                                   (lizzieLet0_4QNone_Bool_4QNode_Bool_d[0] && (! lizzieLet0_4QNone_Bool_4QNode_Bool_emitted[3]))};
  assign lizzieLet0_4QNone_Bool_4QNode_Bool_5_d = {lizzieLet0_4QNone_Bool_4QNode_Bool_d[66:1],
                                                   (lizzieLet0_4QNone_Bool_4QNode_Bool_d[0] && (! lizzieLet0_4QNone_Bool_4QNode_Bool_emitted[4]))};
  assign lizzieLet0_4QNone_Bool_4QNode_Bool_6_d = {lizzieLet0_4QNone_Bool_4QNode_Bool_d[66:1],
                                                   (lizzieLet0_4QNone_Bool_4QNode_Bool_d[0] && (! lizzieLet0_4QNone_Bool_4QNode_Bool_emitted[5]))};
  assign lizzieLet0_4QNone_Bool_4QNode_Bool_7_d = {lizzieLet0_4QNone_Bool_4QNode_Bool_d[66:1],
                                                   (lizzieLet0_4QNone_Bool_4QNode_Bool_d[0] && (! lizzieLet0_4QNone_Bool_4QNode_Bool_emitted[6]))};
  assign lizzieLet0_4QNone_Bool_4QNode_Bool_8_d = {lizzieLet0_4QNone_Bool_4QNode_Bool_d[66:1],
                                                   (lizzieLet0_4QNone_Bool_4QNode_Bool_d[0] && (! lizzieLet0_4QNone_Bool_4QNode_Bool_emitted[7]))};
  assign lizzieLet0_4QNone_Bool_4QNode_Bool_9_d = {lizzieLet0_4QNone_Bool_4QNode_Bool_d[66:1],
                                                   (lizzieLet0_4QNone_Bool_4QNode_Bool_d[0] && (! lizzieLet0_4QNone_Bool_4QNode_Bool_emitted[8]))};
  assign lizzieLet0_4QNone_Bool_4QNode_Bool_done = (lizzieLet0_4QNone_Bool_4QNode_Bool_emitted | ({lizzieLet0_4QNone_Bool_4QNode_Bool_9_d[0],
                                                                                                   lizzieLet0_4QNone_Bool_4QNode_Bool_8_d[0],
                                                                                                   lizzieLet0_4QNone_Bool_4QNode_Bool_7_d[0],
                                                                                                   lizzieLet0_4QNone_Bool_4QNode_Bool_6_d[0],
                                                                                                   lizzieLet0_4QNone_Bool_4QNode_Bool_5_d[0],
                                                                                                   lizzieLet0_4QNone_Bool_4QNode_Bool_4_d[0],
                                                                                                   lizzieLet0_4QNone_Bool_4QNode_Bool_3_d[0],
                                                                                                   lizzieLet0_4QNone_Bool_4QNode_Bool_2_d[0],
                                                                                                   lizzieLet0_4QNone_Bool_4QNode_Bool_1_d[0]} & {lizzieLet0_4QNone_Bool_4QNode_Bool_9_r,
                                                                                                                                                 lizzieLet0_4QNone_Bool_4QNode_Bool_8_r,
                                                                                                                                                 lizzieLet0_4QNone_Bool_4QNode_Bool_7_r,
                                                                                                                                                 lizzieLet0_4QNone_Bool_4QNode_Bool_6_r,
                                                                                                                                                 lizzieLet0_4QNone_Bool_4QNode_Bool_5_r,
                                                                                                                                                 lizzieLet0_4QNone_Bool_4QNode_Bool_4_r,
                                                                                                                                                 lizzieLet0_4QNone_Bool_4QNode_Bool_3_r,
                                                                                                                                                 lizzieLet0_4QNone_Bool_4QNode_Bool_2_r,
                                                                                                                                                 lizzieLet0_4QNone_Bool_4QNode_Bool_1_r}));
  assign lizzieLet0_4QNone_Bool_4QNode_Bool_r = (& lizzieLet0_4QNone_Bool_4QNode_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNone_Bool_4QNode_Bool_emitted <= 9'd0;
    else
      lizzieLet0_4QNone_Bool_4QNode_Bool_emitted <= (lizzieLet0_4QNone_Bool_4QNode_Bool_r ? 9'd0 :
                                                     lizzieLet0_4QNone_Bool_4QNode_Bool_done);
  
  /* destruct (Ty QTree_Bool,
          Dcon QNode_Bool) : (lizzieLet0_4QNone_Bool_4QNode_Bool_1QNode_Bool,QTree_Bool) > [(t1a8i_destruct,Pointer_QTree_Bool),
                                                                                            (t2a8j_destruct,Pointer_QTree_Bool),
                                                                                            (t3a8k_destruct,Pointer_QTree_Bool),
                                                                                            (t4a8l_destruct,Pointer_QTree_Bool)] */
  logic [3:0] lizzieLet0_4QNone_Bool_4QNode_Bool_1QNode_Bool_emitted;
  logic [3:0] lizzieLet0_4QNone_Bool_4QNode_Bool_1QNode_Bool_done;
  assign t1a8i_destruct_d = {lizzieLet0_4QNone_Bool_4QNode_Bool_1QNode_Bool_d[18:3],
                             (lizzieLet0_4QNone_Bool_4QNode_Bool_1QNode_Bool_d[0] && (! lizzieLet0_4QNone_Bool_4QNode_Bool_1QNode_Bool_emitted[0]))};
  assign t2a8j_destruct_d = {lizzieLet0_4QNone_Bool_4QNode_Bool_1QNode_Bool_d[34:19],
                             (lizzieLet0_4QNone_Bool_4QNode_Bool_1QNode_Bool_d[0] && (! lizzieLet0_4QNone_Bool_4QNode_Bool_1QNode_Bool_emitted[1]))};
  assign t3a8k_destruct_d = {lizzieLet0_4QNone_Bool_4QNode_Bool_1QNode_Bool_d[50:35],
                             (lizzieLet0_4QNone_Bool_4QNode_Bool_1QNode_Bool_d[0] && (! lizzieLet0_4QNone_Bool_4QNode_Bool_1QNode_Bool_emitted[2]))};
  assign t4a8l_destruct_d = {lizzieLet0_4QNone_Bool_4QNode_Bool_1QNode_Bool_d[66:51],
                             (lizzieLet0_4QNone_Bool_4QNode_Bool_1QNode_Bool_d[0] && (! lizzieLet0_4QNone_Bool_4QNode_Bool_1QNode_Bool_emitted[3]))};
  assign lizzieLet0_4QNone_Bool_4QNode_Bool_1QNode_Bool_done = (lizzieLet0_4QNone_Bool_4QNode_Bool_1QNode_Bool_emitted | ({t4a8l_destruct_d[0],
                                                                                                                           t3a8k_destruct_d[0],
                                                                                                                           t2a8j_destruct_d[0],
                                                                                                                           t1a8i_destruct_d[0]} & {t4a8l_destruct_r,
                                                                                                                                                   t3a8k_destruct_r,
                                                                                                                                                   t2a8j_destruct_r,
                                                                                                                                                   t1a8i_destruct_r}));
  assign lizzieLet0_4QNone_Bool_4QNode_Bool_1QNode_Bool_r = (& lizzieLet0_4QNone_Bool_4QNode_Bool_1QNode_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNone_Bool_4QNode_Bool_1QNode_Bool_emitted <= 4'd0;
    else
      lizzieLet0_4QNone_Bool_4QNode_Bool_1QNode_Bool_emitted <= (lizzieLet0_4QNone_Bool_4QNode_Bool_1QNode_Bool_r ? 4'd0 :
                                                                 lizzieLet0_4QNone_Bool_4QNode_Bool_1QNode_Bool_done);
  
  /* demux (Ty QTree_Bool,
       Ty QTree_Bool) : (lizzieLet0_4QNone_Bool_4QNode_Bool_2,QTree_Bool) (lizzieLet0_4QNone_Bool_4QNode_Bool_1,QTree_Bool) > [(_108,QTree_Bool),
                                                                                                                               (_107,QTree_Bool),
                                                                                                                               (lizzieLet0_4QNone_Bool_4QNode_Bool_1QNode_Bool,QTree_Bool),
                                                                                                                               (_106,QTree_Bool)] */
  logic [3:0] lizzieLet0_4QNone_Bool_4QNode_Bool_1_onehotd;
  always_comb
    if ((lizzieLet0_4QNone_Bool_4QNode_Bool_2_d[0] && lizzieLet0_4QNone_Bool_4QNode_Bool_1_d[0]))
      unique case (lizzieLet0_4QNone_Bool_4QNode_Bool_2_d[2:1])
        2'd0: lizzieLet0_4QNone_Bool_4QNode_Bool_1_onehotd = 4'd1;
        2'd1: lizzieLet0_4QNone_Bool_4QNode_Bool_1_onehotd = 4'd2;
        2'd2: lizzieLet0_4QNone_Bool_4QNode_Bool_1_onehotd = 4'd4;
        2'd3: lizzieLet0_4QNone_Bool_4QNode_Bool_1_onehotd = 4'd8;
        default: lizzieLet0_4QNone_Bool_4QNode_Bool_1_onehotd = 4'd0;
      endcase
    else lizzieLet0_4QNone_Bool_4QNode_Bool_1_onehotd = 4'd0;
  assign _108_d = {lizzieLet0_4QNone_Bool_4QNode_Bool_1_d[66:1],
                   lizzieLet0_4QNone_Bool_4QNode_Bool_1_onehotd[0]};
  assign _107_d = {lizzieLet0_4QNone_Bool_4QNode_Bool_1_d[66:1],
                   lizzieLet0_4QNone_Bool_4QNode_Bool_1_onehotd[1]};
  assign lizzieLet0_4QNone_Bool_4QNode_Bool_1QNode_Bool_d = {lizzieLet0_4QNone_Bool_4QNode_Bool_1_d[66:1],
                                                             lizzieLet0_4QNone_Bool_4QNode_Bool_1_onehotd[2]};
  assign _106_d = {lizzieLet0_4QNone_Bool_4QNode_Bool_1_d[66:1],
                   lizzieLet0_4QNone_Bool_4QNode_Bool_1_onehotd[3]};
  assign lizzieLet0_4QNone_Bool_4QNode_Bool_1_r = (| (lizzieLet0_4QNone_Bool_4QNode_Bool_1_onehotd & {_106_r,
                                                                                                      lizzieLet0_4QNone_Bool_4QNode_Bool_1QNode_Bool_r,
                                                                                                      _107_r,
                                                                                                      _108_r}));
  assign lizzieLet0_4QNone_Bool_4QNode_Bool_2_r = lizzieLet0_4QNone_Bool_4QNode_Bool_1_r;
  
  /* demux (Ty QTree_Bool,
       Ty Go) : (lizzieLet0_4QNone_Bool_4QNode_Bool_3,QTree_Bool) (lizzieLet0_4QNone_Bool_3QNode_Bool,Go) > [(lizzieLet0_4QNone_Bool_4QNode_Bool_3QNone_Bool,Go),
                                                                                                             (lizzieLet0_4QNone_Bool_4QNode_Bool_3QVal_Bool,Go),
                                                                                                             (lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool,Go),
                                                                                                             (lizzieLet0_4QNone_Bool_4QNode_Bool_3QError_Bool,Go)] */
  logic [3:0] lizzieLet0_4QNone_Bool_3QNode_Bool_onehotd;
  always_comb
    if ((lizzieLet0_4QNone_Bool_4QNode_Bool_3_d[0] && lizzieLet0_4QNone_Bool_3QNode_Bool_d[0]))
      unique case (lizzieLet0_4QNone_Bool_4QNode_Bool_3_d[2:1])
        2'd0: lizzieLet0_4QNone_Bool_3QNode_Bool_onehotd = 4'd1;
        2'd1: lizzieLet0_4QNone_Bool_3QNode_Bool_onehotd = 4'd2;
        2'd2: lizzieLet0_4QNone_Bool_3QNode_Bool_onehotd = 4'd4;
        2'd3: lizzieLet0_4QNone_Bool_3QNode_Bool_onehotd = 4'd8;
        default: lizzieLet0_4QNone_Bool_3QNode_Bool_onehotd = 4'd0;
      endcase
    else lizzieLet0_4QNone_Bool_3QNode_Bool_onehotd = 4'd0;
  assign lizzieLet0_4QNone_Bool_4QNode_Bool_3QNone_Bool_d = lizzieLet0_4QNone_Bool_3QNode_Bool_onehotd[0];
  assign lizzieLet0_4QNone_Bool_4QNode_Bool_3QVal_Bool_d = lizzieLet0_4QNone_Bool_3QNode_Bool_onehotd[1];
  assign lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_d = lizzieLet0_4QNone_Bool_3QNode_Bool_onehotd[2];
  assign lizzieLet0_4QNone_Bool_4QNode_Bool_3QError_Bool_d = lizzieLet0_4QNone_Bool_3QNode_Bool_onehotd[3];
  assign lizzieLet0_4QNone_Bool_3QNode_Bool_r = (| (lizzieLet0_4QNone_Bool_3QNode_Bool_onehotd & {lizzieLet0_4QNone_Bool_4QNode_Bool_3QError_Bool_r,
                                                                                                  lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_r,
                                                                                                  lizzieLet0_4QNone_Bool_4QNode_Bool_3QVal_Bool_r,
                                                                                                  lizzieLet0_4QNone_Bool_4QNode_Bool_3QNone_Bool_r}));
  assign lizzieLet0_4QNone_Bool_4QNode_Bool_3_r = lizzieLet0_4QNone_Bool_3QNode_Bool_r;
  
  /* fork (Ty Go) : (lizzieLet0_4QNone_Bool_4QNode_Bool_3QError_Bool,Go) > [(lizzieLet0_4QNone_Bool_4QNode_Bool_3QError_Bool_1,Go),
                                                                       (lizzieLet0_4QNone_Bool_4QNode_Bool_3QError_Bool_2,Go)] */
  logic [1:0] lizzieLet0_4QNone_Bool_4QNode_Bool_3QError_Bool_emitted;
  logic [1:0] lizzieLet0_4QNone_Bool_4QNode_Bool_3QError_Bool_done;
  assign lizzieLet0_4QNone_Bool_4QNode_Bool_3QError_Bool_1_d = (lizzieLet0_4QNone_Bool_4QNode_Bool_3QError_Bool_d[0] && (! lizzieLet0_4QNone_Bool_4QNode_Bool_3QError_Bool_emitted[0]));
  assign lizzieLet0_4QNone_Bool_4QNode_Bool_3QError_Bool_2_d = (lizzieLet0_4QNone_Bool_4QNode_Bool_3QError_Bool_d[0] && (! lizzieLet0_4QNone_Bool_4QNode_Bool_3QError_Bool_emitted[1]));
  assign lizzieLet0_4QNone_Bool_4QNode_Bool_3QError_Bool_done = (lizzieLet0_4QNone_Bool_4QNode_Bool_3QError_Bool_emitted | ({lizzieLet0_4QNone_Bool_4QNode_Bool_3QError_Bool_2_d[0],
                                                                                                                             lizzieLet0_4QNone_Bool_4QNode_Bool_3QError_Bool_1_d[0]} & {lizzieLet0_4QNone_Bool_4QNode_Bool_3QError_Bool_2_r,
                                                                                                                                                                                        lizzieLet0_4QNone_Bool_4QNode_Bool_3QError_Bool_1_r}));
  assign lizzieLet0_4QNone_Bool_4QNode_Bool_3QError_Bool_r = (& lizzieLet0_4QNone_Bool_4QNode_Bool_3QError_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNone_Bool_4QNode_Bool_3QError_Bool_emitted <= 2'd0;
    else
      lizzieLet0_4QNone_Bool_4QNode_Bool_3QError_Bool_emitted <= (lizzieLet0_4QNone_Bool_4QNode_Bool_3QError_Bool_r ? 2'd0 :
                                                                  lizzieLet0_4QNone_Bool_4QNode_Bool_3QError_Bool_done);
  
  /* dcon (Ty QTree_Bool,
      Dcon QError_Bool) : [(lizzieLet0_4QNone_Bool_4QNode_Bool_3QError_Bool_1,Go)] > (lizzieLet0_4QNone_Bool_4QNode_Bool_3QError_Bool_1QError_Bool,QTree_Bool) */
  assign lizzieLet0_4QNone_Bool_4QNode_Bool_3QError_Bool_1QError_Bool_d = QError_Bool_dc((& {lizzieLet0_4QNone_Bool_4QNode_Bool_3QError_Bool_1_d[0]}), lizzieLet0_4QNone_Bool_4QNode_Bool_3QError_Bool_1_d);
  assign {lizzieLet0_4QNone_Bool_4QNode_Bool_3QError_Bool_1_r} = {1 {(lizzieLet0_4QNone_Bool_4QNode_Bool_3QError_Bool_1QError_Bool_r && lizzieLet0_4QNone_Bool_4QNode_Bool_3QError_Bool_1QError_Bool_d[0])}};
  
  /* buf (Ty QTree_Bool) : (lizzieLet0_4QNone_Bool_4QNode_Bool_3QError_Bool_1QError_Bool,QTree_Bool) > (lizzieLet11_1_1_argbuf,QTree_Bool) */
  QTree_Bool_t lizzieLet0_4QNone_Bool_4QNode_Bool_3QError_Bool_1QError_Bool_bufchan_d;
  logic lizzieLet0_4QNone_Bool_4QNode_Bool_3QError_Bool_1QError_Bool_bufchan_r;
  assign lizzieLet0_4QNone_Bool_4QNode_Bool_3QError_Bool_1QError_Bool_r = ((! lizzieLet0_4QNone_Bool_4QNode_Bool_3QError_Bool_1QError_Bool_bufchan_d[0]) || lizzieLet0_4QNone_Bool_4QNode_Bool_3QError_Bool_1QError_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNone_Bool_4QNode_Bool_3QError_Bool_1QError_Bool_bufchan_d <= {66'd0,
                                                                                 1'd0};
    else
      if (lizzieLet0_4QNone_Bool_4QNode_Bool_3QError_Bool_1QError_Bool_r)
        lizzieLet0_4QNone_Bool_4QNode_Bool_3QError_Bool_1QError_Bool_bufchan_d <= lizzieLet0_4QNone_Bool_4QNode_Bool_3QError_Bool_1QError_Bool_d;
  QTree_Bool_t lizzieLet0_4QNone_Bool_4QNode_Bool_3QError_Bool_1QError_Bool_bufchan_buf;
  assign lizzieLet0_4QNone_Bool_4QNode_Bool_3QError_Bool_1QError_Bool_bufchan_r = (! lizzieLet0_4QNone_Bool_4QNode_Bool_3QError_Bool_1QError_Bool_bufchan_buf[0]);
  assign lizzieLet11_1_1_argbuf_d = (lizzieLet0_4QNone_Bool_4QNode_Bool_3QError_Bool_1QError_Bool_bufchan_buf[0] ? lizzieLet0_4QNone_Bool_4QNode_Bool_3QError_Bool_1QError_Bool_bufchan_buf :
                                     lizzieLet0_4QNone_Bool_4QNode_Bool_3QError_Bool_1QError_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNone_Bool_4QNode_Bool_3QError_Bool_1QError_Bool_bufchan_buf <= {66'd0,
                                                                                   1'd0};
    else
      if ((lizzieLet11_1_1_argbuf_r && lizzieLet0_4QNone_Bool_4QNode_Bool_3QError_Bool_1QError_Bool_bufchan_buf[0]))
        lizzieLet0_4QNone_Bool_4QNode_Bool_3QError_Bool_1QError_Bool_bufchan_buf <= {66'd0,
                                                                                     1'd0};
      else if (((! lizzieLet11_1_1_argbuf_r) && (! lizzieLet0_4QNone_Bool_4QNode_Bool_3QError_Bool_1QError_Bool_bufchan_buf[0])))
        lizzieLet0_4QNone_Bool_4QNode_Bool_3QError_Bool_1QError_Bool_bufchan_buf <= lizzieLet0_4QNone_Bool_4QNode_Bool_3QError_Bool_1QError_Bool_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet0_4QNone_Bool_4QNode_Bool_3QError_Bool_2,Go) > (lizzieLet0_4QNone_Bool_4QNode_Bool_3QError_Bool_2_argbuf,Go) */
  Go_t lizzieLet0_4QNone_Bool_4QNode_Bool_3QError_Bool_2_bufchan_d;
  logic lizzieLet0_4QNone_Bool_4QNode_Bool_3QError_Bool_2_bufchan_r;
  assign lizzieLet0_4QNone_Bool_4QNode_Bool_3QError_Bool_2_r = ((! lizzieLet0_4QNone_Bool_4QNode_Bool_3QError_Bool_2_bufchan_d[0]) || lizzieLet0_4QNone_Bool_4QNode_Bool_3QError_Bool_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNone_Bool_4QNode_Bool_3QError_Bool_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet0_4QNone_Bool_4QNode_Bool_3QError_Bool_2_r)
        lizzieLet0_4QNone_Bool_4QNode_Bool_3QError_Bool_2_bufchan_d <= lizzieLet0_4QNone_Bool_4QNode_Bool_3QError_Bool_2_d;
  Go_t lizzieLet0_4QNone_Bool_4QNode_Bool_3QError_Bool_2_bufchan_buf;
  assign lizzieLet0_4QNone_Bool_4QNode_Bool_3QError_Bool_2_bufchan_r = (! lizzieLet0_4QNone_Bool_4QNode_Bool_3QError_Bool_2_bufchan_buf[0]);
  assign lizzieLet0_4QNone_Bool_4QNode_Bool_3QError_Bool_2_argbuf_d = (lizzieLet0_4QNone_Bool_4QNode_Bool_3QError_Bool_2_bufchan_buf[0] ? lizzieLet0_4QNone_Bool_4QNode_Bool_3QError_Bool_2_bufchan_buf :
                                                                       lizzieLet0_4QNone_Bool_4QNode_Bool_3QError_Bool_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNone_Bool_4QNode_Bool_3QError_Bool_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet0_4QNone_Bool_4QNode_Bool_3QError_Bool_2_argbuf_r && lizzieLet0_4QNone_Bool_4QNode_Bool_3QError_Bool_2_bufchan_buf[0]))
        lizzieLet0_4QNone_Bool_4QNode_Bool_3QError_Bool_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet0_4QNone_Bool_4QNode_Bool_3QError_Bool_2_argbuf_r) && (! lizzieLet0_4QNone_Bool_4QNode_Bool_3QError_Bool_2_bufchan_buf[0])))
        lizzieLet0_4QNone_Bool_4QNode_Bool_3QError_Bool_2_bufchan_buf <= lizzieLet0_4QNone_Bool_4QNode_Bool_3QError_Bool_2_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool,Go) > [(lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_1,Go),
                                                                      (lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_2,Go),
                                                                      (lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_3,Go),
                                                                      (lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_4,Go),
                                                                      (lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_5,Go)] */
  logic [4:0] lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_emitted;
  logic [4:0] lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_done;
  assign lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_1_d = (lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_d[0] && (! lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_emitted[0]));
  assign lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_2_d = (lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_d[0] && (! lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_emitted[1]));
  assign lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_3_d = (lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_d[0] && (! lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_emitted[2]));
  assign lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_4_d = (lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_d[0] && (! lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_emitted[3]));
  assign lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_5_d = (lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_d[0] && (! lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_emitted[4]));
  assign lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_done = (lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_emitted | ({lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_5_d[0],
                                                                                                                           lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_4_d[0],
                                                                                                                           lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_3_d[0],
                                                                                                                           lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_2_d[0],
                                                                                                                           lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_1_d[0]} & {lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_5_r,
                                                                                                                                                                                     lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_4_r,
                                                                                                                                                                                     lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_3_r,
                                                                                                                                                                                     lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_2_r,
                                                                                                                                                                                     lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_1_r}));
  assign lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_r = (& lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_emitted <= 5'd0;
    else
      lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_emitted <= (lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_r ? 5'd0 :
                                                                 lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_done);
  
  /* buf (Ty Go) : (lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_1,Go) > (lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_1_argbuf,Go) */
  Go_t lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_1_bufchan_d;
  logic lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_1_bufchan_r;
  assign lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_1_r = ((! lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_1_bufchan_d[0]) || lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_1_bufchan_d <= 1'd0;
    else
      if (lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_1_r)
        lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_1_bufchan_d <= lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_1_d;
  Go_t lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_1_bufchan_buf;
  assign lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_1_bufchan_r = (! lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_1_bufchan_buf[0]);
  assign lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_1_argbuf_d = (lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_1_bufchan_buf[0] ? lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_1_bufchan_buf :
                                                                      lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_1_argbuf_r && lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_1_bufchan_buf[0]))
        lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_1_argbuf_r) && (! lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_1_bufchan_buf[0])))
        lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_1_bufchan_buf <= lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_1_bufchan_d;
  
  /* dcon (Ty TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool,
      Dcon TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool) : [(lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_1_argbuf,Go),
                                                               (lizzieLet0_4QNone_Bool_4QNode_Bool_9QNode_Bool_1_argbuf,Pointer_QTree_Bool),
                                                               (t4a8l_1_argbuf,Pointer_QTree_Bool)] > (f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_1,TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool) */
  assign \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_1_d  = TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_dc((& {lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_1_argbuf_d[0],
                                                                                                                                     lizzieLet0_4QNone_Bool_4QNode_Bool_9QNode_Bool_1_argbuf_d[0],
                                                                                                                                     t4a8l_1_argbuf_d[0]}), lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_1_argbuf_d, lizzieLet0_4QNone_Bool_4QNode_Bool_9QNode_Bool_1_argbuf_d, t4a8l_1_argbuf_d);
  assign {lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_1_argbuf_r,
          lizzieLet0_4QNone_Bool_4QNode_Bool_9QNode_Bool_1_argbuf_r,
          t4a8l_1_argbuf_r} = {3 {(\f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_1_r  && \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_1_d [0])}};
  
  /* buf (Ty Go) : (lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_2,Go) > (lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_2_argbuf,Go) */
  Go_t lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_2_bufchan_d;
  logic lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_2_bufchan_r;
  assign lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_2_r = ((! lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_2_bufchan_d[0]) || lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_2_r)
        lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_2_bufchan_d <= lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_2_d;
  Go_t lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_2_bufchan_buf;
  assign lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_2_bufchan_r = (! lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_2_bufchan_buf[0]);
  assign lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_2_argbuf_d = (lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_2_bufchan_buf[0] ? lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_2_bufchan_buf :
                                                                      lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_2_argbuf_r && lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_2_bufchan_buf[0]))
        lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_2_argbuf_r) && (! lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_2_bufchan_buf[0])))
        lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_2_bufchan_buf <= lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_2_bufchan_d;
  
  /* dcon (Ty TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool,
      Dcon TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool) : [(lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_2_argbuf,Go),
                                                               (lizzieLet0_4QNone_Bool_4QNode_Bool_8QNode_Bool_1_argbuf,Pointer_QTree_Bool),
                                                               (t3a8k_1_argbuf,Pointer_QTree_Bool)] > (f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool2,TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool) */
  assign \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool2_d  = TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_dc((& {lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_2_argbuf_d[0],
                                                                                                                                    lizzieLet0_4QNone_Bool_4QNode_Bool_8QNode_Bool_1_argbuf_d[0],
                                                                                                                                    t3a8k_1_argbuf_d[0]}), lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_2_argbuf_d, lizzieLet0_4QNone_Bool_4QNode_Bool_8QNode_Bool_1_argbuf_d, t3a8k_1_argbuf_d);
  assign {lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_2_argbuf_r,
          lizzieLet0_4QNone_Bool_4QNode_Bool_8QNode_Bool_1_argbuf_r,
          t3a8k_1_argbuf_r} = {3 {(\f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool2_r  && \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool2_d [0])}};
  
  /* buf (Ty Go) : (lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_3,Go) > (lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_3_argbuf,Go) */
  Go_t lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_3_bufchan_d;
  logic lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_3_bufchan_r;
  assign lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_3_r = ((! lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_3_bufchan_d[0]) || lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_3_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_3_bufchan_d <= 1'd0;
    else
      if (lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_3_r)
        lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_3_bufchan_d <= lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_3_d;
  Go_t lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_3_bufchan_buf;
  assign lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_3_bufchan_r = (! lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_3_bufchan_buf[0]);
  assign lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_3_argbuf_d = (lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_3_bufchan_buf[0] ? lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_3_bufchan_buf :
                                                                      lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_3_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_3_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_3_argbuf_r && lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_3_bufchan_buf[0]))
        lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_3_bufchan_buf <= 1'd0;
      else if (((! lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_3_argbuf_r) && (! lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_3_bufchan_buf[0])))
        lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_3_bufchan_buf <= lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_3_bufchan_d;
  
  /* dcon (Ty TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool,
      Dcon TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool) : [(lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_3_argbuf,Go),
                                                               (lizzieLet0_4QNone_Bool_4QNode_Bool_7QNode_Bool_1_argbuf,Pointer_QTree_Bool),
                                                               (t2a8j_1_argbuf,Pointer_QTree_Bool)] > (f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool3,TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool) */
  assign \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool3_d  = TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_dc((& {lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_3_argbuf_d[0],
                                                                                                                                    lizzieLet0_4QNone_Bool_4QNode_Bool_7QNode_Bool_1_argbuf_d[0],
                                                                                                                                    t2a8j_1_argbuf_d[0]}), lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_3_argbuf_d, lizzieLet0_4QNone_Bool_4QNode_Bool_7QNode_Bool_1_argbuf_d, t2a8j_1_argbuf_d);
  assign {lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_3_argbuf_r,
          lizzieLet0_4QNone_Bool_4QNode_Bool_7QNode_Bool_1_argbuf_r,
          t2a8j_1_argbuf_r} = {3 {(\f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool3_r  && \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool3_d [0])}};
  
  /* buf (Ty Go) : (lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_4,Go) > (lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_4_argbuf,Go) */
  Go_t lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_4_bufchan_d;
  logic lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_4_bufchan_r;
  assign lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_4_r = ((! lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_4_bufchan_d[0]) || lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_4_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_4_bufchan_d <= 1'd0;
    else
      if (lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_4_r)
        lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_4_bufchan_d <= lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_4_d;
  Go_t lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_4_bufchan_buf;
  assign lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_4_bufchan_r = (! lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_4_bufchan_buf[0]);
  assign lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_4_argbuf_d = (lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_4_bufchan_buf[0] ? lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_4_bufchan_buf :
                                                                      lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_4_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_4_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_4_argbuf_r && lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_4_bufchan_buf[0]))
        lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_4_bufchan_buf <= 1'd0;
      else if (((! lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_4_argbuf_r) && (! lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_4_bufchan_buf[0])))
        lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_4_bufchan_buf <= lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_4_bufchan_d;
  
  /* dcon (Ty TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool,
      Dcon TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool) : [(lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_4_argbuf,Go),
                                                               (lizzieLet0_4QNone_Bool_4QNode_Bool_6QNode_Bool_1_argbuf,Pointer_QTree_Bool),
                                                               (t1a8i_1_argbuf,Pointer_QTree_Bool)] > (f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool4,TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool) */
  assign \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool4_d  = TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_dc((& {lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_4_argbuf_d[0],
                                                                                                                                    lizzieLet0_4QNone_Bool_4QNode_Bool_6QNode_Bool_1_argbuf_d[0],
                                                                                                                                    t1a8i_1_argbuf_d[0]}), lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_4_argbuf_d, lizzieLet0_4QNone_Bool_4QNode_Bool_6QNode_Bool_1_argbuf_d, t1a8i_1_argbuf_d);
  assign {lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_4_argbuf_r,
          lizzieLet0_4QNone_Bool_4QNode_Bool_6QNode_Bool_1_argbuf_r,
          t1a8i_1_argbuf_r} = {3 {(\f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool4_r  && \f''''''''''''TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool4_d [0])}};
  
  /* buf (Ty Go) : (lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_5,Go) > (lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_5_argbuf,Go) */
  Go_t lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_5_bufchan_d;
  logic lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_5_bufchan_r;
  assign lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_5_r = ((! lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_5_bufchan_d[0]) || lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_5_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_5_bufchan_d <= 1'd0;
    else
      if (lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_5_r)
        lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_5_bufchan_d <= lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_5_d;
  Go_t lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_5_bufchan_buf;
  assign lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_5_bufchan_r = (! lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_5_bufchan_buf[0]);
  assign lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_5_argbuf_d = (lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_5_bufchan_buf[0] ? lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_5_bufchan_buf :
                                                                      lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_5_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_5_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_5_argbuf_r && lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_5_bufchan_buf[0]))
        lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_5_bufchan_buf <= 1'd0;
      else if (((! lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_5_argbuf_r) && (! lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_5_bufchan_buf[0])))
        lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_5_bufchan_buf <= lizzieLet0_4QNone_Bool_4QNode_Bool_3QNode_Bool_5_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet0_4QNone_Bool_4QNode_Bool_3QNone_Bool,Go) > (lizzieLet0_4QNone_Bool_4QNode_Bool_3QNone_Bool_1_argbuf,Go) */
  Go_t lizzieLet0_4QNone_Bool_4QNode_Bool_3QNone_Bool_bufchan_d;
  logic lizzieLet0_4QNone_Bool_4QNode_Bool_3QNone_Bool_bufchan_r;
  assign lizzieLet0_4QNone_Bool_4QNode_Bool_3QNone_Bool_r = ((! lizzieLet0_4QNone_Bool_4QNode_Bool_3QNone_Bool_bufchan_d[0]) || lizzieLet0_4QNone_Bool_4QNode_Bool_3QNone_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNone_Bool_4QNode_Bool_3QNone_Bool_bufchan_d <= 1'd0;
    else
      if (lizzieLet0_4QNone_Bool_4QNode_Bool_3QNone_Bool_r)
        lizzieLet0_4QNone_Bool_4QNode_Bool_3QNone_Bool_bufchan_d <= lizzieLet0_4QNone_Bool_4QNode_Bool_3QNone_Bool_d;
  Go_t lizzieLet0_4QNone_Bool_4QNode_Bool_3QNone_Bool_bufchan_buf;
  assign lizzieLet0_4QNone_Bool_4QNode_Bool_3QNone_Bool_bufchan_r = (! lizzieLet0_4QNone_Bool_4QNode_Bool_3QNone_Bool_bufchan_buf[0]);
  assign lizzieLet0_4QNone_Bool_4QNode_Bool_3QNone_Bool_1_argbuf_d = (lizzieLet0_4QNone_Bool_4QNode_Bool_3QNone_Bool_bufchan_buf[0] ? lizzieLet0_4QNone_Bool_4QNode_Bool_3QNone_Bool_bufchan_buf :
                                                                      lizzieLet0_4QNone_Bool_4QNode_Bool_3QNone_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNone_Bool_4QNode_Bool_3QNone_Bool_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet0_4QNone_Bool_4QNode_Bool_3QNone_Bool_1_argbuf_r && lizzieLet0_4QNone_Bool_4QNode_Bool_3QNone_Bool_bufchan_buf[0]))
        lizzieLet0_4QNone_Bool_4QNode_Bool_3QNone_Bool_bufchan_buf <= 1'd0;
      else if (((! lizzieLet0_4QNone_Bool_4QNode_Bool_3QNone_Bool_1_argbuf_r) && (! lizzieLet0_4QNone_Bool_4QNode_Bool_3QNone_Bool_bufchan_buf[0])))
        lizzieLet0_4QNone_Bool_4QNode_Bool_3QNone_Bool_bufchan_buf <= lizzieLet0_4QNone_Bool_4QNode_Bool_3QNone_Bool_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet0_4QNone_Bool_4QNode_Bool_3QVal_Bool,Go) > [(lizzieLet0_4QNone_Bool_4QNode_Bool_3QVal_Bool_1,Go),
                                                                     (lizzieLet0_4QNone_Bool_4QNode_Bool_3QVal_Bool_2,Go)] */
  logic [1:0] lizzieLet0_4QNone_Bool_4QNode_Bool_3QVal_Bool_emitted;
  logic [1:0] lizzieLet0_4QNone_Bool_4QNode_Bool_3QVal_Bool_done;
  assign lizzieLet0_4QNone_Bool_4QNode_Bool_3QVal_Bool_1_d = (lizzieLet0_4QNone_Bool_4QNode_Bool_3QVal_Bool_d[0] && (! lizzieLet0_4QNone_Bool_4QNode_Bool_3QVal_Bool_emitted[0]));
  assign lizzieLet0_4QNone_Bool_4QNode_Bool_3QVal_Bool_2_d = (lizzieLet0_4QNone_Bool_4QNode_Bool_3QVal_Bool_d[0] && (! lizzieLet0_4QNone_Bool_4QNode_Bool_3QVal_Bool_emitted[1]));
  assign lizzieLet0_4QNone_Bool_4QNode_Bool_3QVal_Bool_done = (lizzieLet0_4QNone_Bool_4QNode_Bool_3QVal_Bool_emitted | ({lizzieLet0_4QNone_Bool_4QNode_Bool_3QVal_Bool_2_d[0],
                                                                                                                         lizzieLet0_4QNone_Bool_4QNode_Bool_3QVal_Bool_1_d[0]} & {lizzieLet0_4QNone_Bool_4QNode_Bool_3QVal_Bool_2_r,
                                                                                                                                                                                  lizzieLet0_4QNone_Bool_4QNode_Bool_3QVal_Bool_1_r}));
  assign lizzieLet0_4QNone_Bool_4QNode_Bool_3QVal_Bool_r = (& lizzieLet0_4QNone_Bool_4QNode_Bool_3QVal_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNone_Bool_4QNode_Bool_3QVal_Bool_emitted <= 2'd0;
    else
      lizzieLet0_4QNone_Bool_4QNode_Bool_3QVal_Bool_emitted <= (lizzieLet0_4QNone_Bool_4QNode_Bool_3QVal_Bool_r ? 2'd0 :
                                                                lizzieLet0_4QNone_Bool_4QNode_Bool_3QVal_Bool_done);
  
  /* dcon (Ty QTree_Bool,
      Dcon QError_Bool) : [(lizzieLet0_4QNone_Bool_4QNode_Bool_3QVal_Bool_1,Go)] > (lizzieLet0_4QNone_Bool_4QNode_Bool_3QVal_Bool_1QError_Bool,QTree_Bool) */
  assign lizzieLet0_4QNone_Bool_4QNode_Bool_3QVal_Bool_1QError_Bool_d = QError_Bool_dc((& {lizzieLet0_4QNone_Bool_4QNode_Bool_3QVal_Bool_1_d[0]}), lizzieLet0_4QNone_Bool_4QNode_Bool_3QVal_Bool_1_d);
  assign {lizzieLet0_4QNone_Bool_4QNode_Bool_3QVal_Bool_1_r} = {1 {(lizzieLet0_4QNone_Bool_4QNode_Bool_3QVal_Bool_1QError_Bool_r && lizzieLet0_4QNone_Bool_4QNode_Bool_3QVal_Bool_1QError_Bool_d[0])}};
  
  /* buf (Ty QTree_Bool) : (lizzieLet0_4QNone_Bool_4QNode_Bool_3QVal_Bool_1QError_Bool,QTree_Bool) > (lizzieLet9_1_1_argbuf,QTree_Bool) */
  QTree_Bool_t lizzieLet0_4QNone_Bool_4QNode_Bool_3QVal_Bool_1QError_Bool_bufchan_d;
  logic lizzieLet0_4QNone_Bool_4QNode_Bool_3QVal_Bool_1QError_Bool_bufchan_r;
  assign lizzieLet0_4QNone_Bool_4QNode_Bool_3QVal_Bool_1QError_Bool_r = ((! lizzieLet0_4QNone_Bool_4QNode_Bool_3QVal_Bool_1QError_Bool_bufchan_d[0]) || lizzieLet0_4QNone_Bool_4QNode_Bool_3QVal_Bool_1QError_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNone_Bool_4QNode_Bool_3QVal_Bool_1QError_Bool_bufchan_d <= {66'd0,
                                                                               1'd0};
    else
      if (lizzieLet0_4QNone_Bool_4QNode_Bool_3QVal_Bool_1QError_Bool_r)
        lizzieLet0_4QNone_Bool_4QNode_Bool_3QVal_Bool_1QError_Bool_bufchan_d <= lizzieLet0_4QNone_Bool_4QNode_Bool_3QVal_Bool_1QError_Bool_d;
  QTree_Bool_t lizzieLet0_4QNone_Bool_4QNode_Bool_3QVal_Bool_1QError_Bool_bufchan_buf;
  assign lizzieLet0_4QNone_Bool_4QNode_Bool_3QVal_Bool_1QError_Bool_bufchan_r = (! lizzieLet0_4QNone_Bool_4QNode_Bool_3QVal_Bool_1QError_Bool_bufchan_buf[0]);
  assign lizzieLet9_1_1_argbuf_d = (lizzieLet0_4QNone_Bool_4QNode_Bool_3QVal_Bool_1QError_Bool_bufchan_buf[0] ? lizzieLet0_4QNone_Bool_4QNode_Bool_3QVal_Bool_1QError_Bool_bufchan_buf :
                                    lizzieLet0_4QNone_Bool_4QNode_Bool_3QVal_Bool_1QError_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNone_Bool_4QNode_Bool_3QVal_Bool_1QError_Bool_bufchan_buf <= {66'd0,
                                                                                 1'd0};
    else
      if ((lizzieLet9_1_1_argbuf_r && lizzieLet0_4QNone_Bool_4QNode_Bool_3QVal_Bool_1QError_Bool_bufchan_buf[0]))
        lizzieLet0_4QNone_Bool_4QNode_Bool_3QVal_Bool_1QError_Bool_bufchan_buf <= {66'd0,
                                                                                   1'd0};
      else if (((! lizzieLet9_1_1_argbuf_r) && (! lizzieLet0_4QNone_Bool_4QNode_Bool_3QVal_Bool_1QError_Bool_bufchan_buf[0])))
        lizzieLet0_4QNone_Bool_4QNode_Bool_3QVal_Bool_1QError_Bool_bufchan_buf <= lizzieLet0_4QNone_Bool_4QNode_Bool_3QVal_Bool_1QError_Bool_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet0_4QNone_Bool_4QNode_Bool_3QVal_Bool_2,Go) > (lizzieLet0_4QNone_Bool_4QNode_Bool_3QVal_Bool_2_argbuf,Go) */
  Go_t lizzieLet0_4QNone_Bool_4QNode_Bool_3QVal_Bool_2_bufchan_d;
  logic lizzieLet0_4QNone_Bool_4QNode_Bool_3QVal_Bool_2_bufchan_r;
  assign lizzieLet0_4QNone_Bool_4QNode_Bool_3QVal_Bool_2_r = ((! lizzieLet0_4QNone_Bool_4QNode_Bool_3QVal_Bool_2_bufchan_d[0]) || lizzieLet0_4QNone_Bool_4QNode_Bool_3QVal_Bool_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNone_Bool_4QNode_Bool_3QVal_Bool_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet0_4QNone_Bool_4QNode_Bool_3QVal_Bool_2_r)
        lizzieLet0_4QNone_Bool_4QNode_Bool_3QVal_Bool_2_bufchan_d <= lizzieLet0_4QNone_Bool_4QNode_Bool_3QVal_Bool_2_d;
  Go_t lizzieLet0_4QNone_Bool_4QNode_Bool_3QVal_Bool_2_bufchan_buf;
  assign lizzieLet0_4QNone_Bool_4QNode_Bool_3QVal_Bool_2_bufchan_r = (! lizzieLet0_4QNone_Bool_4QNode_Bool_3QVal_Bool_2_bufchan_buf[0]);
  assign lizzieLet0_4QNone_Bool_4QNode_Bool_3QVal_Bool_2_argbuf_d = (lizzieLet0_4QNone_Bool_4QNode_Bool_3QVal_Bool_2_bufchan_buf[0] ? lizzieLet0_4QNone_Bool_4QNode_Bool_3QVal_Bool_2_bufchan_buf :
                                                                     lizzieLet0_4QNone_Bool_4QNode_Bool_3QVal_Bool_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNone_Bool_4QNode_Bool_3QVal_Bool_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet0_4QNone_Bool_4QNode_Bool_3QVal_Bool_2_argbuf_r && lizzieLet0_4QNone_Bool_4QNode_Bool_3QVal_Bool_2_bufchan_buf[0]))
        lizzieLet0_4QNone_Bool_4QNode_Bool_3QVal_Bool_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet0_4QNone_Bool_4QNode_Bool_3QVal_Bool_2_argbuf_r) && (! lizzieLet0_4QNone_Bool_4QNode_Bool_3QVal_Bool_2_bufchan_buf[0])))
        lizzieLet0_4QNone_Bool_4QNode_Bool_3QVal_Bool_2_bufchan_buf <= lizzieLet0_4QNone_Bool_4QNode_Bool_3QVal_Bool_2_bufchan_d;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_QTree_Bool) : (lizzieLet0_4QNone_Bool_4QNode_Bool_4,QTree_Bool) (lizzieLet0_4QNone_Bool_5QNode_Bool,Pointer_QTree_Bool) > [(lizzieLet0_4QNone_Bool_4QNode_Bool_4QNone_Bool,Pointer_QTree_Bool),
                                                                                                                                             (_105,Pointer_QTree_Bool),
                                                                                                                                             (_104,Pointer_QTree_Bool),
                                                                                                                                             (_103,Pointer_QTree_Bool)] */
  logic [3:0] lizzieLet0_4QNone_Bool_5QNode_Bool_onehotd;
  always_comb
    if ((lizzieLet0_4QNone_Bool_4QNode_Bool_4_d[0] && lizzieLet0_4QNone_Bool_5QNode_Bool_d[0]))
      unique case (lizzieLet0_4QNone_Bool_4QNode_Bool_4_d[2:1])
        2'd0: lizzieLet0_4QNone_Bool_5QNode_Bool_onehotd = 4'd1;
        2'd1: lizzieLet0_4QNone_Bool_5QNode_Bool_onehotd = 4'd2;
        2'd2: lizzieLet0_4QNone_Bool_5QNode_Bool_onehotd = 4'd4;
        2'd3: lizzieLet0_4QNone_Bool_5QNode_Bool_onehotd = 4'd8;
        default: lizzieLet0_4QNone_Bool_5QNode_Bool_onehotd = 4'd0;
      endcase
    else lizzieLet0_4QNone_Bool_5QNode_Bool_onehotd = 4'd0;
  assign lizzieLet0_4QNone_Bool_4QNode_Bool_4QNone_Bool_d = {lizzieLet0_4QNone_Bool_5QNode_Bool_d[16:1],
                                                             lizzieLet0_4QNone_Bool_5QNode_Bool_onehotd[0]};
  assign _105_d = {lizzieLet0_4QNone_Bool_5QNode_Bool_d[16:1],
                   lizzieLet0_4QNone_Bool_5QNode_Bool_onehotd[1]};
  assign _104_d = {lizzieLet0_4QNone_Bool_5QNode_Bool_d[16:1],
                   lizzieLet0_4QNone_Bool_5QNode_Bool_onehotd[2]};
  assign _103_d = {lizzieLet0_4QNone_Bool_5QNode_Bool_d[16:1],
                   lizzieLet0_4QNone_Bool_5QNode_Bool_onehotd[3]};
  assign lizzieLet0_4QNone_Bool_5QNode_Bool_r = (| (lizzieLet0_4QNone_Bool_5QNode_Bool_onehotd & {_103_r,
                                                                                                  _104_r,
                                                                                                  _105_r,
                                                                                                  lizzieLet0_4QNone_Bool_4QNode_Bool_4QNone_Bool_r}));
  assign lizzieLet0_4QNone_Bool_4QNode_Bool_4_r = lizzieLet0_4QNone_Bool_5QNode_Bool_r;
  
  /* buf (Ty Pointer_QTree_Bool) : (lizzieLet0_4QNone_Bool_4QNode_Bool_4QNone_Bool,Pointer_QTree_Bool) > (lizzieLet0_4QNone_Bool_4QNode_Bool_4QNone_Bool_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t lizzieLet0_4QNone_Bool_4QNode_Bool_4QNone_Bool_bufchan_d;
  logic lizzieLet0_4QNone_Bool_4QNode_Bool_4QNone_Bool_bufchan_r;
  assign lizzieLet0_4QNone_Bool_4QNode_Bool_4QNone_Bool_r = ((! lizzieLet0_4QNone_Bool_4QNode_Bool_4QNone_Bool_bufchan_d[0]) || lizzieLet0_4QNone_Bool_4QNode_Bool_4QNone_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNone_Bool_4QNode_Bool_4QNone_Bool_bufchan_d <= {16'd0,
                                                                   1'd0};
    else
      if (lizzieLet0_4QNone_Bool_4QNode_Bool_4QNone_Bool_r)
        lizzieLet0_4QNone_Bool_4QNode_Bool_4QNone_Bool_bufchan_d <= lizzieLet0_4QNone_Bool_4QNode_Bool_4QNone_Bool_d;
  Pointer_QTree_Bool_t lizzieLet0_4QNone_Bool_4QNode_Bool_4QNone_Bool_bufchan_buf;
  assign lizzieLet0_4QNone_Bool_4QNode_Bool_4QNone_Bool_bufchan_r = (! lizzieLet0_4QNone_Bool_4QNode_Bool_4QNone_Bool_bufchan_buf[0]);
  assign lizzieLet0_4QNone_Bool_4QNode_Bool_4QNone_Bool_1_argbuf_d = (lizzieLet0_4QNone_Bool_4QNode_Bool_4QNone_Bool_bufchan_buf[0] ? lizzieLet0_4QNone_Bool_4QNode_Bool_4QNone_Bool_bufchan_buf :
                                                                      lizzieLet0_4QNone_Bool_4QNode_Bool_4QNone_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNone_Bool_4QNode_Bool_4QNone_Bool_bufchan_buf <= {16'd0,
                                                                     1'd0};
    else
      if ((lizzieLet0_4QNone_Bool_4QNode_Bool_4QNone_Bool_1_argbuf_r && lizzieLet0_4QNone_Bool_4QNode_Bool_4QNone_Bool_bufchan_buf[0]))
        lizzieLet0_4QNone_Bool_4QNode_Bool_4QNone_Bool_bufchan_buf <= {16'd0,
                                                                       1'd0};
      else if (((! lizzieLet0_4QNone_Bool_4QNode_Bool_4QNone_Bool_1_argbuf_r) && (! lizzieLet0_4QNone_Bool_4QNode_Bool_4QNone_Bool_bufchan_buf[0])))
        lizzieLet0_4QNone_Bool_4QNode_Bool_4QNone_Bool_bufchan_buf <= lizzieLet0_4QNone_Bool_4QNode_Bool_4QNone_Bool_bufchan_d;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_CTf) : (lizzieLet0_4QNone_Bool_4QNode_Bool_5,QTree_Bool) (lizzieLet0_4QNone_Bool_7QNode_Bool,Pointer_CTf) > [(lizzieLet0_4QNone_Bool_4QNode_Bool_5QNone_Bool,Pointer_CTf),
                                                                                                                               (lizzieLet0_4QNone_Bool_4QNode_Bool_5QVal_Bool,Pointer_CTf),
                                                                                                                               (lizzieLet0_4QNone_Bool_4QNode_Bool_5QNode_Bool,Pointer_CTf),
                                                                                                                               (lizzieLet0_4QNone_Bool_4QNode_Bool_5QError_Bool,Pointer_CTf)] */
  logic [3:0] lizzieLet0_4QNone_Bool_7QNode_Bool_onehotd;
  always_comb
    if ((lizzieLet0_4QNone_Bool_4QNode_Bool_5_d[0] && lizzieLet0_4QNone_Bool_7QNode_Bool_d[0]))
      unique case (lizzieLet0_4QNone_Bool_4QNode_Bool_5_d[2:1])
        2'd0: lizzieLet0_4QNone_Bool_7QNode_Bool_onehotd = 4'd1;
        2'd1: lizzieLet0_4QNone_Bool_7QNode_Bool_onehotd = 4'd2;
        2'd2: lizzieLet0_4QNone_Bool_7QNode_Bool_onehotd = 4'd4;
        2'd3: lizzieLet0_4QNone_Bool_7QNode_Bool_onehotd = 4'd8;
        default: lizzieLet0_4QNone_Bool_7QNode_Bool_onehotd = 4'd0;
      endcase
    else lizzieLet0_4QNone_Bool_7QNode_Bool_onehotd = 4'd0;
  assign lizzieLet0_4QNone_Bool_4QNode_Bool_5QNone_Bool_d = {lizzieLet0_4QNone_Bool_7QNode_Bool_d[16:1],
                                                             lizzieLet0_4QNone_Bool_7QNode_Bool_onehotd[0]};
  assign lizzieLet0_4QNone_Bool_4QNode_Bool_5QVal_Bool_d = {lizzieLet0_4QNone_Bool_7QNode_Bool_d[16:1],
                                                            lizzieLet0_4QNone_Bool_7QNode_Bool_onehotd[1]};
  assign lizzieLet0_4QNone_Bool_4QNode_Bool_5QNode_Bool_d = {lizzieLet0_4QNone_Bool_7QNode_Bool_d[16:1],
                                                             lizzieLet0_4QNone_Bool_7QNode_Bool_onehotd[2]};
  assign lizzieLet0_4QNone_Bool_4QNode_Bool_5QError_Bool_d = {lizzieLet0_4QNone_Bool_7QNode_Bool_d[16:1],
                                                              lizzieLet0_4QNone_Bool_7QNode_Bool_onehotd[3]};
  assign lizzieLet0_4QNone_Bool_7QNode_Bool_r = (| (lizzieLet0_4QNone_Bool_7QNode_Bool_onehotd & {lizzieLet0_4QNone_Bool_4QNode_Bool_5QError_Bool_r,
                                                                                                  lizzieLet0_4QNone_Bool_4QNode_Bool_5QNode_Bool_r,
                                                                                                  lizzieLet0_4QNone_Bool_4QNode_Bool_5QVal_Bool_r,
                                                                                                  lizzieLet0_4QNone_Bool_4QNode_Bool_5QNone_Bool_r}));
  assign lizzieLet0_4QNone_Bool_4QNode_Bool_5_r = lizzieLet0_4QNone_Bool_7QNode_Bool_r;
  
  /* buf (Ty Pointer_CTf) : (lizzieLet0_4QNone_Bool_4QNode_Bool_5QError_Bool,Pointer_CTf) > (lizzieLet0_4QNone_Bool_4QNode_Bool_5QError_Bool_1_argbuf,Pointer_CTf) */
  Pointer_CTf_t lizzieLet0_4QNone_Bool_4QNode_Bool_5QError_Bool_bufchan_d;
  logic lizzieLet0_4QNone_Bool_4QNode_Bool_5QError_Bool_bufchan_r;
  assign lizzieLet0_4QNone_Bool_4QNode_Bool_5QError_Bool_r = ((! lizzieLet0_4QNone_Bool_4QNode_Bool_5QError_Bool_bufchan_d[0]) || lizzieLet0_4QNone_Bool_4QNode_Bool_5QError_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNone_Bool_4QNode_Bool_5QError_Bool_bufchan_d <= {16'd0,
                                                                    1'd0};
    else
      if (lizzieLet0_4QNone_Bool_4QNode_Bool_5QError_Bool_r)
        lizzieLet0_4QNone_Bool_4QNode_Bool_5QError_Bool_bufchan_d <= lizzieLet0_4QNone_Bool_4QNode_Bool_5QError_Bool_d;
  Pointer_CTf_t lizzieLet0_4QNone_Bool_4QNode_Bool_5QError_Bool_bufchan_buf;
  assign lizzieLet0_4QNone_Bool_4QNode_Bool_5QError_Bool_bufchan_r = (! lizzieLet0_4QNone_Bool_4QNode_Bool_5QError_Bool_bufchan_buf[0]);
  assign lizzieLet0_4QNone_Bool_4QNode_Bool_5QError_Bool_1_argbuf_d = (lizzieLet0_4QNone_Bool_4QNode_Bool_5QError_Bool_bufchan_buf[0] ? lizzieLet0_4QNone_Bool_4QNode_Bool_5QError_Bool_bufchan_buf :
                                                                       lizzieLet0_4QNone_Bool_4QNode_Bool_5QError_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNone_Bool_4QNode_Bool_5QError_Bool_bufchan_buf <= {16'd0,
                                                                      1'd0};
    else
      if ((lizzieLet0_4QNone_Bool_4QNode_Bool_5QError_Bool_1_argbuf_r && lizzieLet0_4QNone_Bool_4QNode_Bool_5QError_Bool_bufchan_buf[0]))
        lizzieLet0_4QNone_Bool_4QNode_Bool_5QError_Bool_bufchan_buf <= {16'd0,
                                                                        1'd0};
      else if (((! lizzieLet0_4QNone_Bool_4QNode_Bool_5QError_Bool_1_argbuf_r) && (! lizzieLet0_4QNone_Bool_4QNode_Bool_5QError_Bool_bufchan_buf[0])))
        lizzieLet0_4QNone_Bool_4QNode_Bool_5QError_Bool_bufchan_buf <= lizzieLet0_4QNone_Bool_4QNode_Bool_5QError_Bool_bufchan_d;
  
  /* buf (Ty Pointer_CTf) : (lizzieLet0_4QNone_Bool_4QNode_Bool_5QNode_Bool,Pointer_CTf) > (lizzieLet0_4QNone_Bool_4QNode_Bool_5QNode_Bool_1_argbuf,Pointer_CTf) */
  Pointer_CTf_t lizzieLet0_4QNone_Bool_4QNode_Bool_5QNode_Bool_bufchan_d;
  logic lizzieLet0_4QNone_Bool_4QNode_Bool_5QNode_Bool_bufchan_r;
  assign lizzieLet0_4QNone_Bool_4QNode_Bool_5QNode_Bool_r = ((! lizzieLet0_4QNone_Bool_4QNode_Bool_5QNode_Bool_bufchan_d[0]) || lizzieLet0_4QNone_Bool_4QNode_Bool_5QNode_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNone_Bool_4QNode_Bool_5QNode_Bool_bufchan_d <= {16'd0,
                                                                   1'd0};
    else
      if (lizzieLet0_4QNone_Bool_4QNode_Bool_5QNode_Bool_r)
        lizzieLet0_4QNone_Bool_4QNode_Bool_5QNode_Bool_bufchan_d <= lizzieLet0_4QNone_Bool_4QNode_Bool_5QNode_Bool_d;
  Pointer_CTf_t lizzieLet0_4QNone_Bool_4QNode_Bool_5QNode_Bool_bufchan_buf;
  assign lizzieLet0_4QNone_Bool_4QNode_Bool_5QNode_Bool_bufchan_r = (! lizzieLet0_4QNone_Bool_4QNode_Bool_5QNode_Bool_bufchan_buf[0]);
  assign lizzieLet0_4QNone_Bool_4QNode_Bool_5QNode_Bool_1_argbuf_d = (lizzieLet0_4QNone_Bool_4QNode_Bool_5QNode_Bool_bufchan_buf[0] ? lizzieLet0_4QNone_Bool_4QNode_Bool_5QNode_Bool_bufchan_buf :
                                                                      lizzieLet0_4QNone_Bool_4QNode_Bool_5QNode_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNone_Bool_4QNode_Bool_5QNode_Bool_bufchan_buf <= {16'd0,
                                                                     1'd0};
    else
      if ((lizzieLet0_4QNone_Bool_4QNode_Bool_5QNode_Bool_1_argbuf_r && lizzieLet0_4QNone_Bool_4QNode_Bool_5QNode_Bool_bufchan_buf[0]))
        lizzieLet0_4QNone_Bool_4QNode_Bool_5QNode_Bool_bufchan_buf <= {16'd0,
                                                                       1'd0};
      else if (((! lizzieLet0_4QNone_Bool_4QNode_Bool_5QNode_Bool_1_argbuf_r) && (! lizzieLet0_4QNone_Bool_4QNode_Bool_5QNode_Bool_bufchan_buf[0])))
        lizzieLet0_4QNone_Bool_4QNode_Bool_5QNode_Bool_bufchan_buf <= lizzieLet0_4QNone_Bool_4QNode_Bool_5QNode_Bool_bufchan_d;
  
  /* buf (Ty Pointer_CTf) : (lizzieLet0_4QNone_Bool_4QNode_Bool_5QNone_Bool,Pointer_CTf) > (lizzieLet0_4QNone_Bool_4QNode_Bool_5QNone_Bool_1_argbuf,Pointer_CTf) */
  Pointer_CTf_t lizzieLet0_4QNone_Bool_4QNode_Bool_5QNone_Bool_bufchan_d;
  logic lizzieLet0_4QNone_Bool_4QNode_Bool_5QNone_Bool_bufchan_r;
  assign lizzieLet0_4QNone_Bool_4QNode_Bool_5QNone_Bool_r = ((! lizzieLet0_4QNone_Bool_4QNode_Bool_5QNone_Bool_bufchan_d[0]) || lizzieLet0_4QNone_Bool_4QNode_Bool_5QNone_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNone_Bool_4QNode_Bool_5QNone_Bool_bufchan_d <= {16'd0,
                                                                   1'd0};
    else
      if (lizzieLet0_4QNone_Bool_4QNode_Bool_5QNone_Bool_r)
        lizzieLet0_4QNone_Bool_4QNode_Bool_5QNone_Bool_bufchan_d <= lizzieLet0_4QNone_Bool_4QNode_Bool_5QNone_Bool_d;
  Pointer_CTf_t lizzieLet0_4QNone_Bool_4QNode_Bool_5QNone_Bool_bufchan_buf;
  assign lizzieLet0_4QNone_Bool_4QNode_Bool_5QNone_Bool_bufchan_r = (! lizzieLet0_4QNone_Bool_4QNode_Bool_5QNone_Bool_bufchan_buf[0]);
  assign lizzieLet0_4QNone_Bool_4QNode_Bool_5QNone_Bool_1_argbuf_d = (lizzieLet0_4QNone_Bool_4QNode_Bool_5QNone_Bool_bufchan_buf[0] ? lizzieLet0_4QNone_Bool_4QNode_Bool_5QNone_Bool_bufchan_buf :
                                                                      lizzieLet0_4QNone_Bool_4QNode_Bool_5QNone_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNone_Bool_4QNode_Bool_5QNone_Bool_bufchan_buf <= {16'd0,
                                                                     1'd0};
    else
      if ((lizzieLet0_4QNone_Bool_4QNode_Bool_5QNone_Bool_1_argbuf_r && lizzieLet0_4QNone_Bool_4QNode_Bool_5QNone_Bool_bufchan_buf[0]))
        lizzieLet0_4QNone_Bool_4QNode_Bool_5QNone_Bool_bufchan_buf <= {16'd0,
                                                                       1'd0};
      else if (((! lizzieLet0_4QNone_Bool_4QNode_Bool_5QNone_Bool_1_argbuf_r) && (! lizzieLet0_4QNone_Bool_4QNode_Bool_5QNone_Bool_bufchan_buf[0])))
        lizzieLet0_4QNone_Bool_4QNode_Bool_5QNone_Bool_bufchan_buf <= lizzieLet0_4QNone_Bool_4QNode_Bool_5QNone_Bool_bufchan_d;
  
  /* buf (Ty Pointer_CTf) : (lizzieLet0_4QNone_Bool_4QNode_Bool_5QVal_Bool,Pointer_CTf) > (lizzieLet0_4QNone_Bool_4QNode_Bool_5QVal_Bool_1_argbuf,Pointer_CTf) */
  Pointer_CTf_t lizzieLet0_4QNone_Bool_4QNode_Bool_5QVal_Bool_bufchan_d;
  logic lizzieLet0_4QNone_Bool_4QNode_Bool_5QVal_Bool_bufchan_r;
  assign lizzieLet0_4QNone_Bool_4QNode_Bool_5QVal_Bool_r = ((! lizzieLet0_4QNone_Bool_4QNode_Bool_5QVal_Bool_bufchan_d[0]) || lizzieLet0_4QNone_Bool_4QNode_Bool_5QVal_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNone_Bool_4QNode_Bool_5QVal_Bool_bufchan_d <= {16'd0,
                                                                  1'd0};
    else
      if (lizzieLet0_4QNone_Bool_4QNode_Bool_5QVal_Bool_r)
        lizzieLet0_4QNone_Bool_4QNode_Bool_5QVal_Bool_bufchan_d <= lizzieLet0_4QNone_Bool_4QNode_Bool_5QVal_Bool_d;
  Pointer_CTf_t lizzieLet0_4QNone_Bool_4QNode_Bool_5QVal_Bool_bufchan_buf;
  assign lizzieLet0_4QNone_Bool_4QNode_Bool_5QVal_Bool_bufchan_r = (! lizzieLet0_4QNone_Bool_4QNode_Bool_5QVal_Bool_bufchan_buf[0]);
  assign lizzieLet0_4QNone_Bool_4QNode_Bool_5QVal_Bool_1_argbuf_d = (lizzieLet0_4QNone_Bool_4QNode_Bool_5QVal_Bool_bufchan_buf[0] ? lizzieLet0_4QNone_Bool_4QNode_Bool_5QVal_Bool_bufchan_buf :
                                                                     lizzieLet0_4QNone_Bool_4QNode_Bool_5QVal_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNone_Bool_4QNode_Bool_5QVal_Bool_bufchan_buf <= {16'd0,
                                                                    1'd0};
    else
      if ((lizzieLet0_4QNone_Bool_4QNode_Bool_5QVal_Bool_1_argbuf_r && lizzieLet0_4QNone_Bool_4QNode_Bool_5QVal_Bool_bufchan_buf[0]))
        lizzieLet0_4QNone_Bool_4QNode_Bool_5QVal_Bool_bufchan_buf <= {16'd0,
                                                                      1'd0};
      else if (((! lizzieLet0_4QNone_Bool_4QNode_Bool_5QVal_Bool_1_argbuf_r) && (! lizzieLet0_4QNone_Bool_4QNode_Bool_5QVal_Bool_bufchan_buf[0])))
        lizzieLet0_4QNone_Bool_4QNode_Bool_5QVal_Bool_bufchan_buf <= lizzieLet0_4QNone_Bool_4QNode_Bool_5QVal_Bool_bufchan_d;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_QTree_Bool) : (lizzieLet0_4QNone_Bool_4QNode_Bool_6,QTree_Bool) (q1a8d_destruct,Pointer_QTree_Bool) > [(_102,Pointer_QTree_Bool),
                                                                                                                         (_101,Pointer_QTree_Bool),
                                                                                                                         (lizzieLet0_4QNone_Bool_4QNode_Bool_6QNode_Bool,Pointer_QTree_Bool),
                                                                                                                         (_100,Pointer_QTree_Bool)] */
  logic [3:0] q1a8d_destruct_onehotd;
  always_comb
    if ((lizzieLet0_4QNone_Bool_4QNode_Bool_6_d[0] && q1a8d_destruct_d[0]))
      unique case (lizzieLet0_4QNone_Bool_4QNode_Bool_6_d[2:1])
        2'd0: q1a8d_destruct_onehotd = 4'd1;
        2'd1: q1a8d_destruct_onehotd = 4'd2;
        2'd2: q1a8d_destruct_onehotd = 4'd4;
        2'd3: q1a8d_destruct_onehotd = 4'd8;
        default: q1a8d_destruct_onehotd = 4'd0;
      endcase
    else q1a8d_destruct_onehotd = 4'd0;
  assign _102_d = {q1a8d_destruct_d[16:1],
                   q1a8d_destruct_onehotd[0]};
  assign _101_d = {q1a8d_destruct_d[16:1],
                   q1a8d_destruct_onehotd[1]};
  assign lizzieLet0_4QNone_Bool_4QNode_Bool_6QNode_Bool_d = {q1a8d_destruct_d[16:1],
                                                             q1a8d_destruct_onehotd[2]};
  assign _100_d = {q1a8d_destruct_d[16:1],
                   q1a8d_destruct_onehotd[3]};
  assign q1a8d_destruct_r = (| (q1a8d_destruct_onehotd & {_100_r,
                                                          lizzieLet0_4QNone_Bool_4QNode_Bool_6QNode_Bool_r,
                                                          _101_r,
                                                          _102_r}));
  assign lizzieLet0_4QNone_Bool_4QNode_Bool_6_r = q1a8d_destruct_r;
  
  /* buf (Ty Pointer_QTree_Bool) : (lizzieLet0_4QNone_Bool_4QNode_Bool_6QNode_Bool,Pointer_QTree_Bool) > (lizzieLet0_4QNone_Bool_4QNode_Bool_6QNode_Bool_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t lizzieLet0_4QNone_Bool_4QNode_Bool_6QNode_Bool_bufchan_d;
  logic lizzieLet0_4QNone_Bool_4QNode_Bool_6QNode_Bool_bufchan_r;
  assign lizzieLet0_4QNone_Bool_4QNode_Bool_6QNode_Bool_r = ((! lizzieLet0_4QNone_Bool_4QNode_Bool_6QNode_Bool_bufchan_d[0]) || lizzieLet0_4QNone_Bool_4QNode_Bool_6QNode_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNone_Bool_4QNode_Bool_6QNode_Bool_bufchan_d <= {16'd0,
                                                                   1'd0};
    else
      if (lizzieLet0_4QNone_Bool_4QNode_Bool_6QNode_Bool_r)
        lizzieLet0_4QNone_Bool_4QNode_Bool_6QNode_Bool_bufchan_d <= lizzieLet0_4QNone_Bool_4QNode_Bool_6QNode_Bool_d;
  Pointer_QTree_Bool_t lizzieLet0_4QNone_Bool_4QNode_Bool_6QNode_Bool_bufchan_buf;
  assign lizzieLet0_4QNone_Bool_4QNode_Bool_6QNode_Bool_bufchan_r = (! lizzieLet0_4QNone_Bool_4QNode_Bool_6QNode_Bool_bufchan_buf[0]);
  assign lizzieLet0_4QNone_Bool_4QNode_Bool_6QNode_Bool_1_argbuf_d = (lizzieLet0_4QNone_Bool_4QNode_Bool_6QNode_Bool_bufchan_buf[0] ? lizzieLet0_4QNone_Bool_4QNode_Bool_6QNode_Bool_bufchan_buf :
                                                                      lizzieLet0_4QNone_Bool_4QNode_Bool_6QNode_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNone_Bool_4QNode_Bool_6QNode_Bool_bufchan_buf <= {16'd0,
                                                                     1'd0};
    else
      if ((lizzieLet0_4QNone_Bool_4QNode_Bool_6QNode_Bool_1_argbuf_r && lizzieLet0_4QNone_Bool_4QNode_Bool_6QNode_Bool_bufchan_buf[0]))
        lizzieLet0_4QNone_Bool_4QNode_Bool_6QNode_Bool_bufchan_buf <= {16'd0,
                                                                       1'd0};
      else if (((! lizzieLet0_4QNone_Bool_4QNode_Bool_6QNode_Bool_1_argbuf_r) && (! lizzieLet0_4QNone_Bool_4QNode_Bool_6QNode_Bool_bufchan_buf[0])))
        lizzieLet0_4QNone_Bool_4QNode_Bool_6QNode_Bool_bufchan_buf <= lizzieLet0_4QNone_Bool_4QNode_Bool_6QNode_Bool_bufchan_d;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_QTree_Bool) : (lizzieLet0_4QNone_Bool_4QNode_Bool_7,QTree_Bool) (q2a8e_destruct,Pointer_QTree_Bool) > [(_99,Pointer_QTree_Bool),
                                                                                                                         (_98,Pointer_QTree_Bool),
                                                                                                                         (lizzieLet0_4QNone_Bool_4QNode_Bool_7QNode_Bool,Pointer_QTree_Bool),
                                                                                                                         (_97,Pointer_QTree_Bool)] */
  logic [3:0] q2a8e_destruct_onehotd;
  always_comb
    if ((lizzieLet0_4QNone_Bool_4QNode_Bool_7_d[0] && q2a8e_destruct_d[0]))
      unique case (lizzieLet0_4QNone_Bool_4QNode_Bool_7_d[2:1])
        2'd0: q2a8e_destruct_onehotd = 4'd1;
        2'd1: q2a8e_destruct_onehotd = 4'd2;
        2'd2: q2a8e_destruct_onehotd = 4'd4;
        2'd3: q2a8e_destruct_onehotd = 4'd8;
        default: q2a8e_destruct_onehotd = 4'd0;
      endcase
    else q2a8e_destruct_onehotd = 4'd0;
  assign _99_d = {q2a8e_destruct_d[16:1], q2a8e_destruct_onehotd[0]};
  assign _98_d = {q2a8e_destruct_d[16:1], q2a8e_destruct_onehotd[1]};
  assign lizzieLet0_4QNone_Bool_4QNode_Bool_7QNode_Bool_d = {q2a8e_destruct_d[16:1],
                                                             q2a8e_destruct_onehotd[2]};
  assign _97_d = {q2a8e_destruct_d[16:1], q2a8e_destruct_onehotd[3]};
  assign q2a8e_destruct_r = (| (q2a8e_destruct_onehotd & {_97_r,
                                                          lizzieLet0_4QNone_Bool_4QNode_Bool_7QNode_Bool_r,
                                                          _98_r,
                                                          _99_r}));
  assign lizzieLet0_4QNone_Bool_4QNode_Bool_7_r = q2a8e_destruct_r;
  
  /* buf (Ty Pointer_QTree_Bool) : (lizzieLet0_4QNone_Bool_4QNode_Bool_7QNode_Bool,Pointer_QTree_Bool) > (lizzieLet0_4QNone_Bool_4QNode_Bool_7QNode_Bool_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t lizzieLet0_4QNone_Bool_4QNode_Bool_7QNode_Bool_bufchan_d;
  logic lizzieLet0_4QNone_Bool_4QNode_Bool_7QNode_Bool_bufchan_r;
  assign lizzieLet0_4QNone_Bool_4QNode_Bool_7QNode_Bool_r = ((! lizzieLet0_4QNone_Bool_4QNode_Bool_7QNode_Bool_bufchan_d[0]) || lizzieLet0_4QNone_Bool_4QNode_Bool_7QNode_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNone_Bool_4QNode_Bool_7QNode_Bool_bufchan_d <= {16'd0,
                                                                   1'd0};
    else
      if (lizzieLet0_4QNone_Bool_4QNode_Bool_7QNode_Bool_r)
        lizzieLet0_4QNone_Bool_4QNode_Bool_7QNode_Bool_bufchan_d <= lizzieLet0_4QNone_Bool_4QNode_Bool_7QNode_Bool_d;
  Pointer_QTree_Bool_t lizzieLet0_4QNone_Bool_4QNode_Bool_7QNode_Bool_bufchan_buf;
  assign lizzieLet0_4QNone_Bool_4QNode_Bool_7QNode_Bool_bufchan_r = (! lizzieLet0_4QNone_Bool_4QNode_Bool_7QNode_Bool_bufchan_buf[0]);
  assign lizzieLet0_4QNone_Bool_4QNode_Bool_7QNode_Bool_1_argbuf_d = (lizzieLet0_4QNone_Bool_4QNode_Bool_7QNode_Bool_bufchan_buf[0] ? lizzieLet0_4QNone_Bool_4QNode_Bool_7QNode_Bool_bufchan_buf :
                                                                      lizzieLet0_4QNone_Bool_4QNode_Bool_7QNode_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNone_Bool_4QNode_Bool_7QNode_Bool_bufchan_buf <= {16'd0,
                                                                     1'd0};
    else
      if ((lizzieLet0_4QNone_Bool_4QNode_Bool_7QNode_Bool_1_argbuf_r && lizzieLet0_4QNone_Bool_4QNode_Bool_7QNode_Bool_bufchan_buf[0]))
        lizzieLet0_4QNone_Bool_4QNode_Bool_7QNode_Bool_bufchan_buf <= {16'd0,
                                                                       1'd0};
      else if (((! lizzieLet0_4QNone_Bool_4QNode_Bool_7QNode_Bool_1_argbuf_r) && (! lizzieLet0_4QNone_Bool_4QNode_Bool_7QNode_Bool_bufchan_buf[0])))
        lizzieLet0_4QNone_Bool_4QNode_Bool_7QNode_Bool_bufchan_buf <= lizzieLet0_4QNone_Bool_4QNode_Bool_7QNode_Bool_bufchan_d;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_QTree_Bool) : (lizzieLet0_4QNone_Bool_4QNode_Bool_8,QTree_Bool) (q3a8f_destruct,Pointer_QTree_Bool) > [(_96,Pointer_QTree_Bool),
                                                                                                                         (_95,Pointer_QTree_Bool),
                                                                                                                         (lizzieLet0_4QNone_Bool_4QNode_Bool_8QNode_Bool,Pointer_QTree_Bool),
                                                                                                                         (_94,Pointer_QTree_Bool)] */
  logic [3:0] q3a8f_destruct_onehotd;
  always_comb
    if ((lizzieLet0_4QNone_Bool_4QNode_Bool_8_d[0] && q3a8f_destruct_d[0]))
      unique case (lizzieLet0_4QNone_Bool_4QNode_Bool_8_d[2:1])
        2'd0: q3a8f_destruct_onehotd = 4'd1;
        2'd1: q3a8f_destruct_onehotd = 4'd2;
        2'd2: q3a8f_destruct_onehotd = 4'd4;
        2'd3: q3a8f_destruct_onehotd = 4'd8;
        default: q3a8f_destruct_onehotd = 4'd0;
      endcase
    else q3a8f_destruct_onehotd = 4'd0;
  assign _96_d = {q3a8f_destruct_d[16:1], q3a8f_destruct_onehotd[0]};
  assign _95_d = {q3a8f_destruct_d[16:1], q3a8f_destruct_onehotd[1]};
  assign lizzieLet0_4QNone_Bool_4QNode_Bool_8QNode_Bool_d = {q3a8f_destruct_d[16:1],
                                                             q3a8f_destruct_onehotd[2]};
  assign _94_d = {q3a8f_destruct_d[16:1], q3a8f_destruct_onehotd[3]};
  assign q3a8f_destruct_r = (| (q3a8f_destruct_onehotd & {_94_r,
                                                          lizzieLet0_4QNone_Bool_4QNode_Bool_8QNode_Bool_r,
                                                          _95_r,
                                                          _96_r}));
  assign lizzieLet0_4QNone_Bool_4QNode_Bool_8_r = q3a8f_destruct_r;
  
  /* buf (Ty Pointer_QTree_Bool) : (lizzieLet0_4QNone_Bool_4QNode_Bool_8QNode_Bool,Pointer_QTree_Bool) > (lizzieLet0_4QNone_Bool_4QNode_Bool_8QNode_Bool_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t lizzieLet0_4QNone_Bool_4QNode_Bool_8QNode_Bool_bufchan_d;
  logic lizzieLet0_4QNone_Bool_4QNode_Bool_8QNode_Bool_bufchan_r;
  assign lizzieLet0_4QNone_Bool_4QNode_Bool_8QNode_Bool_r = ((! lizzieLet0_4QNone_Bool_4QNode_Bool_8QNode_Bool_bufchan_d[0]) || lizzieLet0_4QNone_Bool_4QNode_Bool_8QNode_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNone_Bool_4QNode_Bool_8QNode_Bool_bufchan_d <= {16'd0,
                                                                   1'd0};
    else
      if (lizzieLet0_4QNone_Bool_4QNode_Bool_8QNode_Bool_r)
        lizzieLet0_4QNone_Bool_4QNode_Bool_8QNode_Bool_bufchan_d <= lizzieLet0_4QNone_Bool_4QNode_Bool_8QNode_Bool_d;
  Pointer_QTree_Bool_t lizzieLet0_4QNone_Bool_4QNode_Bool_8QNode_Bool_bufchan_buf;
  assign lizzieLet0_4QNone_Bool_4QNode_Bool_8QNode_Bool_bufchan_r = (! lizzieLet0_4QNone_Bool_4QNode_Bool_8QNode_Bool_bufchan_buf[0]);
  assign lizzieLet0_4QNone_Bool_4QNode_Bool_8QNode_Bool_1_argbuf_d = (lizzieLet0_4QNone_Bool_4QNode_Bool_8QNode_Bool_bufchan_buf[0] ? lizzieLet0_4QNone_Bool_4QNode_Bool_8QNode_Bool_bufchan_buf :
                                                                      lizzieLet0_4QNone_Bool_4QNode_Bool_8QNode_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNone_Bool_4QNode_Bool_8QNode_Bool_bufchan_buf <= {16'd0,
                                                                     1'd0};
    else
      if ((lizzieLet0_4QNone_Bool_4QNode_Bool_8QNode_Bool_1_argbuf_r && lizzieLet0_4QNone_Bool_4QNode_Bool_8QNode_Bool_bufchan_buf[0]))
        lizzieLet0_4QNone_Bool_4QNode_Bool_8QNode_Bool_bufchan_buf <= {16'd0,
                                                                       1'd0};
      else if (((! lizzieLet0_4QNone_Bool_4QNode_Bool_8QNode_Bool_1_argbuf_r) && (! lizzieLet0_4QNone_Bool_4QNode_Bool_8QNode_Bool_bufchan_buf[0])))
        lizzieLet0_4QNone_Bool_4QNode_Bool_8QNode_Bool_bufchan_buf <= lizzieLet0_4QNone_Bool_4QNode_Bool_8QNode_Bool_bufchan_d;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_QTree_Bool) : (lizzieLet0_4QNone_Bool_4QNode_Bool_9,QTree_Bool) (q4a8g_destruct,Pointer_QTree_Bool) > [(_93,Pointer_QTree_Bool),
                                                                                                                         (_92,Pointer_QTree_Bool),
                                                                                                                         (lizzieLet0_4QNone_Bool_4QNode_Bool_9QNode_Bool,Pointer_QTree_Bool),
                                                                                                                         (_91,Pointer_QTree_Bool)] */
  logic [3:0] q4a8g_destruct_onehotd;
  always_comb
    if ((lizzieLet0_4QNone_Bool_4QNode_Bool_9_d[0] && q4a8g_destruct_d[0]))
      unique case (lizzieLet0_4QNone_Bool_4QNode_Bool_9_d[2:1])
        2'd0: q4a8g_destruct_onehotd = 4'd1;
        2'd1: q4a8g_destruct_onehotd = 4'd2;
        2'd2: q4a8g_destruct_onehotd = 4'd4;
        2'd3: q4a8g_destruct_onehotd = 4'd8;
        default: q4a8g_destruct_onehotd = 4'd0;
      endcase
    else q4a8g_destruct_onehotd = 4'd0;
  assign _93_d = {q4a8g_destruct_d[16:1], q4a8g_destruct_onehotd[0]};
  assign _92_d = {q4a8g_destruct_d[16:1], q4a8g_destruct_onehotd[1]};
  assign lizzieLet0_4QNone_Bool_4QNode_Bool_9QNode_Bool_d = {q4a8g_destruct_d[16:1],
                                                             q4a8g_destruct_onehotd[2]};
  assign _91_d = {q4a8g_destruct_d[16:1], q4a8g_destruct_onehotd[3]};
  assign q4a8g_destruct_r = (| (q4a8g_destruct_onehotd & {_91_r,
                                                          lizzieLet0_4QNone_Bool_4QNode_Bool_9QNode_Bool_r,
                                                          _92_r,
                                                          _93_r}));
  assign lizzieLet0_4QNone_Bool_4QNode_Bool_9_r = q4a8g_destruct_r;
  
  /* buf (Ty Pointer_QTree_Bool) : (lizzieLet0_4QNone_Bool_4QNode_Bool_9QNode_Bool,Pointer_QTree_Bool) > (lizzieLet0_4QNone_Bool_4QNode_Bool_9QNode_Bool_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t lizzieLet0_4QNone_Bool_4QNode_Bool_9QNode_Bool_bufchan_d;
  logic lizzieLet0_4QNone_Bool_4QNode_Bool_9QNode_Bool_bufchan_r;
  assign lizzieLet0_4QNone_Bool_4QNode_Bool_9QNode_Bool_r = ((! lizzieLet0_4QNone_Bool_4QNode_Bool_9QNode_Bool_bufchan_d[0]) || lizzieLet0_4QNone_Bool_4QNode_Bool_9QNode_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNone_Bool_4QNode_Bool_9QNode_Bool_bufchan_d <= {16'd0,
                                                                   1'd0};
    else
      if (lizzieLet0_4QNone_Bool_4QNode_Bool_9QNode_Bool_r)
        lizzieLet0_4QNone_Bool_4QNode_Bool_9QNode_Bool_bufchan_d <= lizzieLet0_4QNone_Bool_4QNode_Bool_9QNode_Bool_d;
  Pointer_QTree_Bool_t lizzieLet0_4QNone_Bool_4QNode_Bool_9QNode_Bool_bufchan_buf;
  assign lizzieLet0_4QNone_Bool_4QNode_Bool_9QNode_Bool_bufchan_r = (! lizzieLet0_4QNone_Bool_4QNode_Bool_9QNode_Bool_bufchan_buf[0]);
  assign lizzieLet0_4QNone_Bool_4QNode_Bool_9QNode_Bool_1_argbuf_d = (lizzieLet0_4QNone_Bool_4QNode_Bool_9QNode_Bool_bufchan_buf[0] ? lizzieLet0_4QNone_Bool_4QNode_Bool_9QNode_Bool_bufchan_buf :
                                                                      lizzieLet0_4QNone_Bool_4QNode_Bool_9QNode_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNone_Bool_4QNode_Bool_9QNode_Bool_bufchan_buf <= {16'd0,
                                                                     1'd0};
    else
      if ((lizzieLet0_4QNone_Bool_4QNode_Bool_9QNode_Bool_1_argbuf_r && lizzieLet0_4QNone_Bool_4QNode_Bool_9QNode_Bool_bufchan_buf[0]))
        lizzieLet0_4QNone_Bool_4QNode_Bool_9QNode_Bool_bufchan_buf <= {16'd0,
                                                                       1'd0};
      else if (((! lizzieLet0_4QNone_Bool_4QNode_Bool_9QNode_Bool_1_argbuf_r) && (! lizzieLet0_4QNone_Bool_4QNode_Bool_9QNode_Bool_bufchan_buf[0])))
        lizzieLet0_4QNone_Bool_4QNode_Bool_9QNode_Bool_bufchan_buf <= lizzieLet0_4QNone_Bool_4QNode_Bool_9QNode_Bool_bufchan_d;
  
  /* fork (Ty QTree_Bool) : (lizzieLet0_4QNone_Bool_4QVal_Bool,QTree_Bool) > [(lizzieLet0_4QNone_Bool_4QVal_Bool_1,QTree_Bool),
                                                                         (lizzieLet0_4QNone_Bool_4QVal_Bool_2,QTree_Bool),
                                                                         (lizzieLet0_4QNone_Bool_4QVal_Bool_3,QTree_Bool),
                                                                         (lizzieLet0_4QNone_Bool_4QVal_Bool_4,QTree_Bool),
                                                                         (lizzieLet0_4QNone_Bool_4QVal_Bool_5,QTree_Bool),
                                                                         (lizzieLet0_4QNone_Bool_4QVal_Bool_6,QTree_Bool)] */
  logic [5:0] lizzieLet0_4QNone_Bool_4QVal_Bool_emitted;
  logic [5:0] lizzieLet0_4QNone_Bool_4QVal_Bool_done;
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_1_d = {lizzieLet0_4QNone_Bool_4QVal_Bool_d[66:1],
                                                  (lizzieLet0_4QNone_Bool_4QVal_Bool_d[0] && (! lizzieLet0_4QNone_Bool_4QVal_Bool_emitted[0]))};
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_2_d = {lizzieLet0_4QNone_Bool_4QVal_Bool_d[66:1],
                                                  (lizzieLet0_4QNone_Bool_4QVal_Bool_d[0] && (! lizzieLet0_4QNone_Bool_4QVal_Bool_emitted[1]))};
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_3_d = {lizzieLet0_4QNone_Bool_4QVal_Bool_d[66:1],
                                                  (lizzieLet0_4QNone_Bool_4QVal_Bool_d[0] && (! lizzieLet0_4QNone_Bool_4QVal_Bool_emitted[2]))};
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_4_d = {lizzieLet0_4QNone_Bool_4QVal_Bool_d[66:1],
                                                  (lizzieLet0_4QNone_Bool_4QVal_Bool_d[0] && (! lizzieLet0_4QNone_Bool_4QVal_Bool_emitted[3]))};
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_5_d = {lizzieLet0_4QNone_Bool_4QVal_Bool_d[66:1],
                                                  (lizzieLet0_4QNone_Bool_4QVal_Bool_d[0] && (! lizzieLet0_4QNone_Bool_4QVal_Bool_emitted[4]))};
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_6_d = {lizzieLet0_4QNone_Bool_4QVal_Bool_d[66:1],
                                                  (lizzieLet0_4QNone_Bool_4QVal_Bool_d[0] && (! lizzieLet0_4QNone_Bool_4QVal_Bool_emitted[5]))};
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_done = (lizzieLet0_4QNone_Bool_4QVal_Bool_emitted | ({lizzieLet0_4QNone_Bool_4QVal_Bool_6_d[0],
                                                                                                 lizzieLet0_4QNone_Bool_4QVal_Bool_5_d[0],
                                                                                                 lizzieLet0_4QNone_Bool_4QVal_Bool_4_d[0],
                                                                                                 lizzieLet0_4QNone_Bool_4QVal_Bool_3_d[0],
                                                                                                 lizzieLet0_4QNone_Bool_4QVal_Bool_2_d[0],
                                                                                                 lizzieLet0_4QNone_Bool_4QVal_Bool_1_d[0]} & {lizzieLet0_4QNone_Bool_4QVal_Bool_6_r,
                                                                                                                                              lizzieLet0_4QNone_Bool_4QVal_Bool_5_r,
                                                                                                                                              lizzieLet0_4QNone_Bool_4QVal_Bool_4_r,
                                                                                                                                              lizzieLet0_4QNone_Bool_4QVal_Bool_3_r,
                                                                                                                                              lizzieLet0_4QNone_Bool_4QVal_Bool_2_r,
                                                                                                                                              lizzieLet0_4QNone_Bool_4QVal_Bool_1_r}));
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_r = (& lizzieLet0_4QNone_Bool_4QVal_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNone_Bool_4QVal_Bool_emitted <= 6'd0;
    else
      lizzieLet0_4QNone_Bool_4QVal_Bool_emitted <= (lizzieLet0_4QNone_Bool_4QVal_Bool_r ? 6'd0 :
                                                    lizzieLet0_4QNone_Bool_4QVal_Bool_done);
  
  /* destruct (Ty QTree_Bool,
          Dcon QVal_Bool) : (lizzieLet0_4QNone_Bool_4QVal_Bool_1QVal_Bool,QTree_Bool) > [(va88_destruct,MyBool)] */
  assign va88_destruct_d = {lizzieLet0_4QNone_Bool_4QVal_Bool_1QVal_Bool_d[3:3],
                            lizzieLet0_4QNone_Bool_4QVal_Bool_1QVal_Bool_d[0]};
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_1QVal_Bool_r = va88_destruct_r;
  
  /* demux (Ty QTree_Bool,
       Ty QTree_Bool) : (lizzieLet0_4QNone_Bool_4QVal_Bool_2,QTree_Bool) (lizzieLet0_4QNone_Bool_4QVal_Bool_1,QTree_Bool) > [(_90,QTree_Bool),
                                                                                                                             (lizzieLet0_4QNone_Bool_4QVal_Bool_1QVal_Bool,QTree_Bool),
                                                                                                                             (_89,QTree_Bool),
                                                                                                                             (_88,QTree_Bool)] */
  logic [3:0] lizzieLet0_4QNone_Bool_4QVal_Bool_1_onehotd;
  always_comb
    if ((lizzieLet0_4QNone_Bool_4QVal_Bool_2_d[0] && lizzieLet0_4QNone_Bool_4QVal_Bool_1_d[0]))
      unique case (lizzieLet0_4QNone_Bool_4QVal_Bool_2_d[2:1])
        2'd0: lizzieLet0_4QNone_Bool_4QVal_Bool_1_onehotd = 4'd1;
        2'd1: lizzieLet0_4QNone_Bool_4QVal_Bool_1_onehotd = 4'd2;
        2'd2: lizzieLet0_4QNone_Bool_4QVal_Bool_1_onehotd = 4'd4;
        2'd3: lizzieLet0_4QNone_Bool_4QVal_Bool_1_onehotd = 4'd8;
        default: lizzieLet0_4QNone_Bool_4QVal_Bool_1_onehotd = 4'd0;
      endcase
    else lizzieLet0_4QNone_Bool_4QVal_Bool_1_onehotd = 4'd0;
  assign _90_d = {lizzieLet0_4QNone_Bool_4QVal_Bool_1_d[66:1],
                  lizzieLet0_4QNone_Bool_4QVal_Bool_1_onehotd[0]};
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_1QVal_Bool_d = {lizzieLet0_4QNone_Bool_4QVal_Bool_1_d[66:1],
                                                           lizzieLet0_4QNone_Bool_4QVal_Bool_1_onehotd[1]};
  assign _89_d = {lizzieLet0_4QNone_Bool_4QVal_Bool_1_d[66:1],
                  lizzieLet0_4QNone_Bool_4QVal_Bool_1_onehotd[2]};
  assign _88_d = {lizzieLet0_4QNone_Bool_4QVal_Bool_1_d[66:1],
                  lizzieLet0_4QNone_Bool_4QVal_Bool_1_onehotd[3]};
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_1_r = (| (lizzieLet0_4QNone_Bool_4QVal_Bool_1_onehotd & {_88_r,
                                                                                                    _89_r,
                                                                                                    lizzieLet0_4QNone_Bool_4QVal_Bool_1QVal_Bool_r,
                                                                                                    _90_r}));
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_2_r = lizzieLet0_4QNone_Bool_4QVal_Bool_1_r;
  
  /* demux (Ty QTree_Bool,
       Ty Go) : (lizzieLet0_4QNone_Bool_4QVal_Bool_3,QTree_Bool) (lizzieLet0_4QNone_Bool_3QVal_Bool,Go) > [(lizzieLet0_4QNone_Bool_4QVal_Bool_3QNone_Bool,Go),
                                                                                                           (lizzieLet0_4QNone_Bool_4QVal_Bool_3QVal_Bool,Go),
                                                                                                           (lizzieLet0_4QNone_Bool_4QVal_Bool_3QNode_Bool,Go),
                                                                                                           (lizzieLet0_4QNone_Bool_4QVal_Bool_3QError_Bool,Go)] */
  logic [3:0] lizzieLet0_4QNone_Bool_3QVal_Bool_onehotd;
  always_comb
    if ((lizzieLet0_4QNone_Bool_4QVal_Bool_3_d[0] && lizzieLet0_4QNone_Bool_3QVal_Bool_d[0]))
      unique case (lizzieLet0_4QNone_Bool_4QVal_Bool_3_d[2:1])
        2'd0: lizzieLet0_4QNone_Bool_3QVal_Bool_onehotd = 4'd1;
        2'd1: lizzieLet0_4QNone_Bool_3QVal_Bool_onehotd = 4'd2;
        2'd2: lizzieLet0_4QNone_Bool_3QVal_Bool_onehotd = 4'd4;
        2'd3: lizzieLet0_4QNone_Bool_3QVal_Bool_onehotd = 4'd8;
        default: lizzieLet0_4QNone_Bool_3QVal_Bool_onehotd = 4'd0;
      endcase
    else lizzieLet0_4QNone_Bool_3QVal_Bool_onehotd = 4'd0;
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_3QNone_Bool_d = lizzieLet0_4QNone_Bool_3QVal_Bool_onehotd[0];
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_3QVal_Bool_d = lizzieLet0_4QNone_Bool_3QVal_Bool_onehotd[1];
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_3QNode_Bool_d = lizzieLet0_4QNone_Bool_3QVal_Bool_onehotd[2];
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_3QError_Bool_d = lizzieLet0_4QNone_Bool_3QVal_Bool_onehotd[3];
  assign lizzieLet0_4QNone_Bool_3QVal_Bool_r = (| (lizzieLet0_4QNone_Bool_3QVal_Bool_onehotd & {lizzieLet0_4QNone_Bool_4QVal_Bool_3QError_Bool_r,
                                                                                                lizzieLet0_4QNone_Bool_4QVal_Bool_3QNode_Bool_r,
                                                                                                lizzieLet0_4QNone_Bool_4QVal_Bool_3QVal_Bool_r,
                                                                                                lizzieLet0_4QNone_Bool_4QVal_Bool_3QNone_Bool_r}));
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_3_r = lizzieLet0_4QNone_Bool_3QVal_Bool_r;
  
  /* fork (Ty Go) : (lizzieLet0_4QNone_Bool_4QVal_Bool_3QError_Bool,Go) > [(lizzieLet0_4QNone_Bool_4QVal_Bool_3QError_Bool_1,Go),
                                                                      (lizzieLet0_4QNone_Bool_4QVal_Bool_3QError_Bool_2,Go)] */
  logic [1:0] lizzieLet0_4QNone_Bool_4QVal_Bool_3QError_Bool_emitted;
  logic [1:0] lizzieLet0_4QNone_Bool_4QVal_Bool_3QError_Bool_done;
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_3QError_Bool_1_d = (lizzieLet0_4QNone_Bool_4QVal_Bool_3QError_Bool_d[0] && (! lizzieLet0_4QNone_Bool_4QVal_Bool_3QError_Bool_emitted[0]));
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_3QError_Bool_2_d = (lizzieLet0_4QNone_Bool_4QVal_Bool_3QError_Bool_d[0] && (! lizzieLet0_4QNone_Bool_4QVal_Bool_3QError_Bool_emitted[1]));
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_3QError_Bool_done = (lizzieLet0_4QNone_Bool_4QVal_Bool_3QError_Bool_emitted | ({lizzieLet0_4QNone_Bool_4QVal_Bool_3QError_Bool_2_d[0],
                                                                                                                           lizzieLet0_4QNone_Bool_4QVal_Bool_3QError_Bool_1_d[0]} & {lizzieLet0_4QNone_Bool_4QVal_Bool_3QError_Bool_2_r,
                                                                                                                                                                                     lizzieLet0_4QNone_Bool_4QVal_Bool_3QError_Bool_1_r}));
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_3QError_Bool_r = (& lizzieLet0_4QNone_Bool_4QVal_Bool_3QError_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNone_Bool_4QVal_Bool_3QError_Bool_emitted <= 2'd0;
    else
      lizzieLet0_4QNone_Bool_4QVal_Bool_3QError_Bool_emitted <= (lizzieLet0_4QNone_Bool_4QVal_Bool_3QError_Bool_r ? 2'd0 :
                                                                 lizzieLet0_4QNone_Bool_4QVal_Bool_3QError_Bool_done);
  
  /* dcon (Ty QTree_Bool,
      Dcon QError_Bool) : [(lizzieLet0_4QNone_Bool_4QVal_Bool_3QError_Bool_1,Go)] > (lizzieLet0_4QNone_Bool_4QVal_Bool_3QError_Bool_1QError_Bool,QTree_Bool) */
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_3QError_Bool_1QError_Bool_d = QError_Bool_dc((& {lizzieLet0_4QNone_Bool_4QVal_Bool_3QError_Bool_1_d[0]}), lizzieLet0_4QNone_Bool_4QVal_Bool_3QError_Bool_1_d);
  assign {lizzieLet0_4QNone_Bool_4QVal_Bool_3QError_Bool_1_r} = {1 {(lizzieLet0_4QNone_Bool_4QVal_Bool_3QError_Bool_1QError_Bool_r && lizzieLet0_4QNone_Bool_4QVal_Bool_3QError_Bool_1QError_Bool_d[0])}};
  
  /* buf (Ty QTree_Bool) : (lizzieLet0_4QNone_Bool_4QVal_Bool_3QError_Bool_1QError_Bool,QTree_Bool) > (lizzieLet7_1_argbuf,QTree_Bool) */
  QTree_Bool_t lizzieLet0_4QNone_Bool_4QVal_Bool_3QError_Bool_1QError_Bool_bufchan_d;
  logic lizzieLet0_4QNone_Bool_4QVal_Bool_3QError_Bool_1QError_Bool_bufchan_r;
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_3QError_Bool_1QError_Bool_r = ((! lizzieLet0_4QNone_Bool_4QVal_Bool_3QError_Bool_1QError_Bool_bufchan_d[0]) || lizzieLet0_4QNone_Bool_4QVal_Bool_3QError_Bool_1QError_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNone_Bool_4QVal_Bool_3QError_Bool_1QError_Bool_bufchan_d <= {66'd0,
                                                                                1'd0};
    else
      if (lizzieLet0_4QNone_Bool_4QVal_Bool_3QError_Bool_1QError_Bool_r)
        lizzieLet0_4QNone_Bool_4QVal_Bool_3QError_Bool_1QError_Bool_bufchan_d <= lizzieLet0_4QNone_Bool_4QVal_Bool_3QError_Bool_1QError_Bool_d;
  QTree_Bool_t lizzieLet0_4QNone_Bool_4QVal_Bool_3QError_Bool_1QError_Bool_bufchan_buf;
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_3QError_Bool_1QError_Bool_bufchan_r = (! lizzieLet0_4QNone_Bool_4QVal_Bool_3QError_Bool_1QError_Bool_bufchan_buf[0]);
  assign lizzieLet7_1_argbuf_d = (lizzieLet0_4QNone_Bool_4QVal_Bool_3QError_Bool_1QError_Bool_bufchan_buf[0] ? lizzieLet0_4QNone_Bool_4QVal_Bool_3QError_Bool_1QError_Bool_bufchan_buf :
                                  lizzieLet0_4QNone_Bool_4QVal_Bool_3QError_Bool_1QError_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNone_Bool_4QVal_Bool_3QError_Bool_1QError_Bool_bufchan_buf <= {66'd0,
                                                                                  1'd0};
    else
      if ((lizzieLet7_1_argbuf_r && lizzieLet0_4QNone_Bool_4QVal_Bool_3QError_Bool_1QError_Bool_bufchan_buf[0]))
        lizzieLet0_4QNone_Bool_4QVal_Bool_3QError_Bool_1QError_Bool_bufchan_buf <= {66'd0,
                                                                                    1'd0};
      else if (((! lizzieLet7_1_argbuf_r) && (! lizzieLet0_4QNone_Bool_4QVal_Bool_3QError_Bool_1QError_Bool_bufchan_buf[0])))
        lizzieLet0_4QNone_Bool_4QVal_Bool_3QError_Bool_1QError_Bool_bufchan_buf <= lizzieLet0_4QNone_Bool_4QVal_Bool_3QError_Bool_1QError_Bool_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet0_4QNone_Bool_4QVal_Bool_3QError_Bool_2,Go) > (lizzieLet0_4QNone_Bool_4QVal_Bool_3QError_Bool_2_argbuf,Go) */
  Go_t lizzieLet0_4QNone_Bool_4QVal_Bool_3QError_Bool_2_bufchan_d;
  logic lizzieLet0_4QNone_Bool_4QVal_Bool_3QError_Bool_2_bufchan_r;
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_3QError_Bool_2_r = ((! lizzieLet0_4QNone_Bool_4QVal_Bool_3QError_Bool_2_bufchan_d[0]) || lizzieLet0_4QNone_Bool_4QVal_Bool_3QError_Bool_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNone_Bool_4QVal_Bool_3QError_Bool_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet0_4QNone_Bool_4QVal_Bool_3QError_Bool_2_r)
        lizzieLet0_4QNone_Bool_4QVal_Bool_3QError_Bool_2_bufchan_d <= lizzieLet0_4QNone_Bool_4QVal_Bool_3QError_Bool_2_d;
  Go_t lizzieLet0_4QNone_Bool_4QVal_Bool_3QError_Bool_2_bufchan_buf;
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_3QError_Bool_2_bufchan_r = (! lizzieLet0_4QNone_Bool_4QVal_Bool_3QError_Bool_2_bufchan_buf[0]);
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_3QError_Bool_2_argbuf_d = (lizzieLet0_4QNone_Bool_4QVal_Bool_3QError_Bool_2_bufchan_buf[0] ? lizzieLet0_4QNone_Bool_4QVal_Bool_3QError_Bool_2_bufchan_buf :
                                                                      lizzieLet0_4QNone_Bool_4QVal_Bool_3QError_Bool_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNone_Bool_4QVal_Bool_3QError_Bool_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet0_4QNone_Bool_4QVal_Bool_3QError_Bool_2_argbuf_r && lizzieLet0_4QNone_Bool_4QVal_Bool_3QError_Bool_2_bufchan_buf[0]))
        lizzieLet0_4QNone_Bool_4QVal_Bool_3QError_Bool_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet0_4QNone_Bool_4QVal_Bool_3QError_Bool_2_argbuf_r) && (! lizzieLet0_4QNone_Bool_4QVal_Bool_3QError_Bool_2_bufchan_buf[0])))
        lizzieLet0_4QNone_Bool_4QVal_Bool_3QError_Bool_2_bufchan_buf <= lizzieLet0_4QNone_Bool_4QVal_Bool_3QError_Bool_2_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet0_4QNone_Bool_4QVal_Bool_3QNode_Bool,Go) > [(lizzieLet0_4QNone_Bool_4QVal_Bool_3QNode_Bool_1,Go),
                                                                     (lizzieLet0_4QNone_Bool_4QVal_Bool_3QNode_Bool_2,Go)] */
  logic [1:0] lizzieLet0_4QNone_Bool_4QVal_Bool_3QNode_Bool_emitted;
  logic [1:0] lizzieLet0_4QNone_Bool_4QVal_Bool_3QNode_Bool_done;
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_3QNode_Bool_1_d = (lizzieLet0_4QNone_Bool_4QVal_Bool_3QNode_Bool_d[0] && (! lizzieLet0_4QNone_Bool_4QVal_Bool_3QNode_Bool_emitted[0]));
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_3QNode_Bool_2_d = (lizzieLet0_4QNone_Bool_4QVal_Bool_3QNode_Bool_d[0] && (! lizzieLet0_4QNone_Bool_4QVal_Bool_3QNode_Bool_emitted[1]));
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_3QNode_Bool_done = (lizzieLet0_4QNone_Bool_4QVal_Bool_3QNode_Bool_emitted | ({lizzieLet0_4QNone_Bool_4QVal_Bool_3QNode_Bool_2_d[0],
                                                                                                                         lizzieLet0_4QNone_Bool_4QVal_Bool_3QNode_Bool_1_d[0]} & {lizzieLet0_4QNone_Bool_4QVal_Bool_3QNode_Bool_2_r,
                                                                                                                                                                                  lizzieLet0_4QNone_Bool_4QVal_Bool_3QNode_Bool_1_r}));
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_3QNode_Bool_r = (& lizzieLet0_4QNone_Bool_4QVal_Bool_3QNode_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNone_Bool_4QVal_Bool_3QNode_Bool_emitted <= 2'd0;
    else
      lizzieLet0_4QNone_Bool_4QVal_Bool_3QNode_Bool_emitted <= (lizzieLet0_4QNone_Bool_4QVal_Bool_3QNode_Bool_r ? 2'd0 :
                                                                lizzieLet0_4QNone_Bool_4QVal_Bool_3QNode_Bool_done);
  
  /* dcon (Ty QTree_Bool,
      Dcon QError_Bool) : [(lizzieLet0_4QNone_Bool_4QVal_Bool_3QNode_Bool_1,Go)] > (lizzieLet0_4QNone_Bool_4QVal_Bool_3QNode_Bool_1QError_Bool,QTree_Bool) */
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_3QNode_Bool_1QError_Bool_d = QError_Bool_dc((& {lizzieLet0_4QNone_Bool_4QVal_Bool_3QNode_Bool_1_d[0]}), lizzieLet0_4QNone_Bool_4QVal_Bool_3QNode_Bool_1_d);
  assign {lizzieLet0_4QNone_Bool_4QVal_Bool_3QNode_Bool_1_r} = {1 {(lizzieLet0_4QNone_Bool_4QVal_Bool_3QNode_Bool_1QError_Bool_r && lizzieLet0_4QNone_Bool_4QVal_Bool_3QNode_Bool_1QError_Bool_d[0])}};
  
  /* buf (Ty QTree_Bool) : (lizzieLet0_4QNone_Bool_4QVal_Bool_3QNode_Bool_1QError_Bool,QTree_Bool) > (lizzieLet6_1_argbuf,QTree_Bool) */
  QTree_Bool_t lizzieLet0_4QNone_Bool_4QVal_Bool_3QNode_Bool_1QError_Bool_bufchan_d;
  logic lizzieLet0_4QNone_Bool_4QVal_Bool_3QNode_Bool_1QError_Bool_bufchan_r;
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_3QNode_Bool_1QError_Bool_r = ((! lizzieLet0_4QNone_Bool_4QVal_Bool_3QNode_Bool_1QError_Bool_bufchan_d[0]) || lizzieLet0_4QNone_Bool_4QVal_Bool_3QNode_Bool_1QError_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNone_Bool_4QVal_Bool_3QNode_Bool_1QError_Bool_bufchan_d <= {66'd0,
                                                                               1'd0};
    else
      if (lizzieLet0_4QNone_Bool_4QVal_Bool_3QNode_Bool_1QError_Bool_r)
        lizzieLet0_4QNone_Bool_4QVal_Bool_3QNode_Bool_1QError_Bool_bufchan_d <= lizzieLet0_4QNone_Bool_4QVal_Bool_3QNode_Bool_1QError_Bool_d;
  QTree_Bool_t lizzieLet0_4QNone_Bool_4QVal_Bool_3QNode_Bool_1QError_Bool_bufchan_buf;
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_3QNode_Bool_1QError_Bool_bufchan_r = (! lizzieLet0_4QNone_Bool_4QVal_Bool_3QNode_Bool_1QError_Bool_bufchan_buf[0]);
  assign lizzieLet6_1_argbuf_d = (lizzieLet0_4QNone_Bool_4QVal_Bool_3QNode_Bool_1QError_Bool_bufchan_buf[0] ? lizzieLet0_4QNone_Bool_4QVal_Bool_3QNode_Bool_1QError_Bool_bufchan_buf :
                                  lizzieLet0_4QNone_Bool_4QVal_Bool_3QNode_Bool_1QError_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNone_Bool_4QVal_Bool_3QNode_Bool_1QError_Bool_bufchan_buf <= {66'd0,
                                                                                 1'd0};
    else
      if ((lizzieLet6_1_argbuf_r && lizzieLet0_4QNone_Bool_4QVal_Bool_3QNode_Bool_1QError_Bool_bufchan_buf[0]))
        lizzieLet0_4QNone_Bool_4QVal_Bool_3QNode_Bool_1QError_Bool_bufchan_buf <= {66'd0,
                                                                                   1'd0};
      else if (((! lizzieLet6_1_argbuf_r) && (! lizzieLet0_4QNone_Bool_4QVal_Bool_3QNode_Bool_1QError_Bool_bufchan_buf[0])))
        lizzieLet0_4QNone_Bool_4QVal_Bool_3QNode_Bool_1QError_Bool_bufchan_buf <= lizzieLet0_4QNone_Bool_4QVal_Bool_3QNode_Bool_1QError_Bool_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet0_4QNone_Bool_4QVal_Bool_3QNode_Bool_2,Go) > (lizzieLet0_4QNone_Bool_4QVal_Bool_3QNode_Bool_2_argbuf,Go) */
  Go_t lizzieLet0_4QNone_Bool_4QVal_Bool_3QNode_Bool_2_bufchan_d;
  logic lizzieLet0_4QNone_Bool_4QVal_Bool_3QNode_Bool_2_bufchan_r;
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_3QNode_Bool_2_r = ((! lizzieLet0_4QNone_Bool_4QVal_Bool_3QNode_Bool_2_bufchan_d[0]) || lizzieLet0_4QNone_Bool_4QVal_Bool_3QNode_Bool_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNone_Bool_4QVal_Bool_3QNode_Bool_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet0_4QNone_Bool_4QVal_Bool_3QNode_Bool_2_r)
        lizzieLet0_4QNone_Bool_4QVal_Bool_3QNode_Bool_2_bufchan_d <= lizzieLet0_4QNone_Bool_4QVal_Bool_3QNode_Bool_2_d;
  Go_t lizzieLet0_4QNone_Bool_4QVal_Bool_3QNode_Bool_2_bufchan_buf;
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_3QNode_Bool_2_bufchan_r = (! lizzieLet0_4QNone_Bool_4QVal_Bool_3QNode_Bool_2_bufchan_buf[0]);
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_3QNode_Bool_2_argbuf_d = (lizzieLet0_4QNone_Bool_4QVal_Bool_3QNode_Bool_2_bufchan_buf[0] ? lizzieLet0_4QNone_Bool_4QVal_Bool_3QNode_Bool_2_bufchan_buf :
                                                                     lizzieLet0_4QNone_Bool_4QVal_Bool_3QNode_Bool_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNone_Bool_4QVal_Bool_3QNode_Bool_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet0_4QNone_Bool_4QVal_Bool_3QNode_Bool_2_argbuf_r && lizzieLet0_4QNone_Bool_4QVal_Bool_3QNode_Bool_2_bufchan_buf[0]))
        lizzieLet0_4QNone_Bool_4QVal_Bool_3QNode_Bool_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet0_4QNone_Bool_4QVal_Bool_3QNode_Bool_2_argbuf_r) && (! lizzieLet0_4QNone_Bool_4QVal_Bool_3QNode_Bool_2_bufchan_buf[0])))
        lizzieLet0_4QNone_Bool_4QVal_Bool_3QNode_Bool_2_bufchan_buf <= lizzieLet0_4QNone_Bool_4QVal_Bool_3QNode_Bool_2_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet0_4QNone_Bool_4QVal_Bool_3QNone_Bool,Go) > (lizzieLet0_4QNone_Bool_4QVal_Bool_3QNone_Bool_1_argbuf,Go) */
  Go_t lizzieLet0_4QNone_Bool_4QVal_Bool_3QNone_Bool_bufchan_d;
  logic lizzieLet0_4QNone_Bool_4QVal_Bool_3QNone_Bool_bufchan_r;
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_3QNone_Bool_r = ((! lizzieLet0_4QNone_Bool_4QVal_Bool_3QNone_Bool_bufchan_d[0]) || lizzieLet0_4QNone_Bool_4QVal_Bool_3QNone_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNone_Bool_4QVal_Bool_3QNone_Bool_bufchan_d <= 1'd0;
    else
      if (lizzieLet0_4QNone_Bool_4QVal_Bool_3QNone_Bool_r)
        lizzieLet0_4QNone_Bool_4QVal_Bool_3QNone_Bool_bufchan_d <= lizzieLet0_4QNone_Bool_4QVal_Bool_3QNone_Bool_d;
  Go_t lizzieLet0_4QNone_Bool_4QVal_Bool_3QNone_Bool_bufchan_buf;
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_3QNone_Bool_bufchan_r = (! lizzieLet0_4QNone_Bool_4QVal_Bool_3QNone_Bool_bufchan_buf[0]);
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_3QNone_Bool_1_argbuf_d = (lizzieLet0_4QNone_Bool_4QVal_Bool_3QNone_Bool_bufchan_buf[0] ? lizzieLet0_4QNone_Bool_4QVal_Bool_3QNone_Bool_bufchan_buf :
                                                                     lizzieLet0_4QNone_Bool_4QVal_Bool_3QNone_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNone_Bool_4QVal_Bool_3QNone_Bool_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet0_4QNone_Bool_4QVal_Bool_3QNone_Bool_1_argbuf_r && lizzieLet0_4QNone_Bool_4QVal_Bool_3QNone_Bool_bufchan_buf[0]))
        lizzieLet0_4QNone_Bool_4QVal_Bool_3QNone_Bool_bufchan_buf <= 1'd0;
      else if (((! lizzieLet0_4QNone_Bool_4QVal_Bool_3QNone_Bool_1_argbuf_r) && (! lizzieLet0_4QNone_Bool_4QVal_Bool_3QNone_Bool_bufchan_buf[0])))
        lizzieLet0_4QNone_Bool_4QVal_Bool_3QNone_Bool_bufchan_buf <= lizzieLet0_4QNone_Bool_4QVal_Bool_3QNone_Bool_bufchan_d;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_QTree_Bool) : (lizzieLet0_4QNone_Bool_4QVal_Bool_4,QTree_Bool) (lizzieLet0_4QNone_Bool_5QVal_Bool,Pointer_QTree_Bool) > [(lizzieLet0_4QNone_Bool_4QVal_Bool_4QNone_Bool,Pointer_QTree_Bool),
                                                                                                                                           (_87,Pointer_QTree_Bool),
                                                                                                                                           (_86,Pointer_QTree_Bool),
                                                                                                                                           (_85,Pointer_QTree_Bool)] */
  logic [3:0] lizzieLet0_4QNone_Bool_5QVal_Bool_onehotd;
  always_comb
    if ((lizzieLet0_4QNone_Bool_4QVal_Bool_4_d[0] && lizzieLet0_4QNone_Bool_5QVal_Bool_d[0]))
      unique case (lizzieLet0_4QNone_Bool_4QVal_Bool_4_d[2:1])
        2'd0: lizzieLet0_4QNone_Bool_5QVal_Bool_onehotd = 4'd1;
        2'd1: lizzieLet0_4QNone_Bool_5QVal_Bool_onehotd = 4'd2;
        2'd2: lizzieLet0_4QNone_Bool_5QVal_Bool_onehotd = 4'd4;
        2'd3: lizzieLet0_4QNone_Bool_5QVal_Bool_onehotd = 4'd8;
        default: lizzieLet0_4QNone_Bool_5QVal_Bool_onehotd = 4'd0;
      endcase
    else lizzieLet0_4QNone_Bool_5QVal_Bool_onehotd = 4'd0;
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_4QNone_Bool_d = {lizzieLet0_4QNone_Bool_5QVal_Bool_d[16:1],
                                                            lizzieLet0_4QNone_Bool_5QVal_Bool_onehotd[0]};
  assign _87_d = {lizzieLet0_4QNone_Bool_5QVal_Bool_d[16:1],
                  lizzieLet0_4QNone_Bool_5QVal_Bool_onehotd[1]};
  assign _86_d = {lizzieLet0_4QNone_Bool_5QVal_Bool_d[16:1],
                  lizzieLet0_4QNone_Bool_5QVal_Bool_onehotd[2]};
  assign _85_d = {lizzieLet0_4QNone_Bool_5QVal_Bool_d[16:1],
                  lizzieLet0_4QNone_Bool_5QVal_Bool_onehotd[3]};
  assign lizzieLet0_4QNone_Bool_5QVal_Bool_r = (| (lizzieLet0_4QNone_Bool_5QVal_Bool_onehotd & {_85_r,
                                                                                                _86_r,
                                                                                                _87_r,
                                                                                                lizzieLet0_4QNone_Bool_4QVal_Bool_4QNone_Bool_r}));
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_4_r = lizzieLet0_4QNone_Bool_5QVal_Bool_r;
  
  /* buf (Ty Pointer_QTree_Bool) : (lizzieLet0_4QNone_Bool_4QVal_Bool_4QNone_Bool,Pointer_QTree_Bool) > (lizzieLet0_4QNone_Bool_4QVal_Bool_4QNone_Bool_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t lizzieLet0_4QNone_Bool_4QVal_Bool_4QNone_Bool_bufchan_d;
  logic lizzieLet0_4QNone_Bool_4QVal_Bool_4QNone_Bool_bufchan_r;
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_4QNone_Bool_r = ((! lizzieLet0_4QNone_Bool_4QVal_Bool_4QNone_Bool_bufchan_d[0]) || lizzieLet0_4QNone_Bool_4QVal_Bool_4QNone_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNone_Bool_4QVal_Bool_4QNone_Bool_bufchan_d <= {16'd0,
                                                                  1'd0};
    else
      if (lizzieLet0_4QNone_Bool_4QVal_Bool_4QNone_Bool_r)
        lizzieLet0_4QNone_Bool_4QVal_Bool_4QNone_Bool_bufchan_d <= lizzieLet0_4QNone_Bool_4QVal_Bool_4QNone_Bool_d;
  Pointer_QTree_Bool_t lizzieLet0_4QNone_Bool_4QVal_Bool_4QNone_Bool_bufchan_buf;
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_4QNone_Bool_bufchan_r = (! lizzieLet0_4QNone_Bool_4QVal_Bool_4QNone_Bool_bufchan_buf[0]);
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_4QNone_Bool_1_argbuf_d = (lizzieLet0_4QNone_Bool_4QVal_Bool_4QNone_Bool_bufchan_buf[0] ? lizzieLet0_4QNone_Bool_4QVal_Bool_4QNone_Bool_bufchan_buf :
                                                                     lizzieLet0_4QNone_Bool_4QVal_Bool_4QNone_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNone_Bool_4QVal_Bool_4QNone_Bool_bufchan_buf <= {16'd0,
                                                                    1'd0};
    else
      if ((lizzieLet0_4QNone_Bool_4QVal_Bool_4QNone_Bool_1_argbuf_r && lizzieLet0_4QNone_Bool_4QVal_Bool_4QNone_Bool_bufchan_buf[0]))
        lizzieLet0_4QNone_Bool_4QVal_Bool_4QNone_Bool_bufchan_buf <= {16'd0,
                                                                      1'd0};
      else if (((! lizzieLet0_4QNone_Bool_4QVal_Bool_4QNone_Bool_1_argbuf_r) && (! lizzieLet0_4QNone_Bool_4QVal_Bool_4QNone_Bool_bufchan_buf[0])))
        lizzieLet0_4QNone_Bool_4QVal_Bool_4QNone_Bool_bufchan_buf <= lizzieLet0_4QNone_Bool_4QVal_Bool_4QNone_Bool_bufchan_d;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_CTf) : (lizzieLet0_4QNone_Bool_4QVal_Bool_5,QTree_Bool) (lizzieLet0_4QNone_Bool_7QVal_Bool,Pointer_CTf) > [(lizzieLet0_4QNone_Bool_4QVal_Bool_5QNone_Bool,Pointer_CTf),
                                                                                                                             (lizzieLet0_4QNone_Bool_4QVal_Bool_5QVal_Bool,Pointer_CTf),
                                                                                                                             (lizzieLet0_4QNone_Bool_4QVal_Bool_5QNode_Bool,Pointer_CTf),
                                                                                                                             (lizzieLet0_4QNone_Bool_4QVal_Bool_5QError_Bool,Pointer_CTf)] */
  logic [3:0] lizzieLet0_4QNone_Bool_7QVal_Bool_onehotd;
  always_comb
    if ((lizzieLet0_4QNone_Bool_4QVal_Bool_5_d[0] && lizzieLet0_4QNone_Bool_7QVal_Bool_d[0]))
      unique case (lizzieLet0_4QNone_Bool_4QVal_Bool_5_d[2:1])
        2'd0: lizzieLet0_4QNone_Bool_7QVal_Bool_onehotd = 4'd1;
        2'd1: lizzieLet0_4QNone_Bool_7QVal_Bool_onehotd = 4'd2;
        2'd2: lizzieLet0_4QNone_Bool_7QVal_Bool_onehotd = 4'd4;
        2'd3: lizzieLet0_4QNone_Bool_7QVal_Bool_onehotd = 4'd8;
        default: lizzieLet0_4QNone_Bool_7QVal_Bool_onehotd = 4'd0;
      endcase
    else lizzieLet0_4QNone_Bool_7QVal_Bool_onehotd = 4'd0;
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_5QNone_Bool_d = {lizzieLet0_4QNone_Bool_7QVal_Bool_d[16:1],
                                                            lizzieLet0_4QNone_Bool_7QVal_Bool_onehotd[0]};
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_5QVal_Bool_d = {lizzieLet0_4QNone_Bool_7QVal_Bool_d[16:1],
                                                           lizzieLet0_4QNone_Bool_7QVal_Bool_onehotd[1]};
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_5QNode_Bool_d = {lizzieLet0_4QNone_Bool_7QVal_Bool_d[16:1],
                                                            lizzieLet0_4QNone_Bool_7QVal_Bool_onehotd[2]};
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_5QError_Bool_d = {lizzieLet0_4QNone_Bool_7QVal_Bool_d[16:1],
                                                             lizzieLet0_4QNone_Bool_7QVal_Bool_onehotd[3]};
  assign lizzieLet0_4QNone_Bool_7QVal_Bool_r = (| (lizzieLet0_4QNone_Bool_7QVal_Bool_onehotd & {lizzieLet0_4QNone_Bool_4QVal_Bool_5QError_Bool_r,
                                                                                                lizzieLet0_4QNone_Bool_4QVal_Bool_5QNode_Bool_r,
                                                                                                lizzieLet0_4QNone_Bool_4QVal_Bool_5QVal_Bool_r,
                                                                                                lizzieLet0_4QNone_Bool_4QVal_Bool_5QNone_Bool_r}));
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_5_r = lizzieLet0_4QNone_Bool_7QVal_Bool_r;
  
  /* buf (Ty Pointer_CTf) : (lizzieLet0_4QNone_Bool_4QVal_Bool_5QError_Bool,Pointer_CTf) > (lizzieLet0_4QNone_Bool_4QVal_Bool_5QError_Bool_1_argbuf,Pointer_CTf) */
  Pointer_CTf_t lizzieLet0_4QNone_Bool_4QVal_Bool_5QError_Bool_bufchan_d;
  logic lizzieLet0_4QNone_Bool_4QVal_Bool_5QError_Bool_bufchan_r;
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_5QError_Bool_r = ((! lizzieLet0_4QNone_Bool_4QVal_Bool_5QError_Bool_bufchan_d[0]) || lizzieLet0_4QNone_Bool_4QVal_Bool_5QError_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNone_Bool_4QVal_Bool_5QError_Bool_bufchan_d <= {16'd0,
                                                                   1'd0};
    else
      if (lizzieLet0_4QNone_Bool_4QVal_Bool_5QError_Bool_r)
        lizzieLet0_4QNone_Bool_4QVal_Bool_5QError_Bool_bufchan_d <= lizzieLet0_4QNone_Bool_4QVal_Bool_5QError_Bool_d;
  Pointer_CTf_t lizzieLet0_4QNone_Bool_4QVal_Bool_5QError_Bool_bufchan_buf;
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_5QError_Bool_bufchan_r = (! lizzieLet0_4QNone_Bool_4QVal_Bool_5QError_Bool_bufchan_buf[0]);
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_5QError_Bool_1_argbuf_d = (lizzieLet0_4QNone_Bool_4QVal_Bool_5QError_Bool_bufchan_buf[0] ? lizzieLet0_4QNone_Bool_4QVal_Bool_5QError_Bool_bufchan_buf :
                                                                      lizzieLet0_4QNone_Bool_4QVal_Bool_5QError_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNone_Bool_4QVal_Bool_5QError_Bool_bufchan_buf <= {16'd0,
                                                                     1'd0};
    else
      if ((lizzieLet0_4QNone_Bool_4QVal_Bool_5QError_Bool_1_argbuf_r && lizzieLet0_4QNone_Bool_4QVal_Bool_5QError_Bool_bufchan_buf[0]))
        lizzieLet0_4QNone_Bool_4QVal_Bool_5QError_Bool_bufchan_buf <= {16'd0,
                                                                       1'd0};
      else if (((! lizzieLet0_4QNone_Bool_4QVal_Bool_5QError_Bool_1_argbuf_r) && (! lizzieLet0_4QNone_Bool_4QVal_Bool_5QError_Bool_bufchan_buf[0])))
        lizzieLet0_4QNone_Bool_4QVal_Bool_5QError_Bool_bufchan_buf <= lizzieLet0_4QNone_Bool_4QVal_Bool_5QError_Bool_bufchan_d;
  
  /* buf (Ty Pointer_CTf) : (lizzieLet0_4QNone_Bool_4QVal_Bool_5QNode_Bool,Pointer_CTf) > (lizzieLet0_4QNone_Bool_4QVal_Bool_5QNode_Bool_1_argbuf,Pointer_CTf) */
  Pointer_CTf_t lizzieLet0_4QNone_Bool_4QVal_Bool_5QNode_Bool_bufchan_d;
  logic lizzieLet0_4QNone_Bool_4QVal_Bool_5QNode_Bool_bufchan_r;
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_5QNode_Bool_r = ((! lizzieLet0_4QNone_Bool_4QVal_Bool_5QNode_Bool_bufchan_d[0]) || lizzieLet0_4QNone_Bool_4QVal_Bool_5QNode_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNone_Bool_4QVal_Bool_5QNode_Bool_bufchan_d <= {16'd0,
                                                                  1'd0};
    else
      if (lizzieLet0_4QNone_Bool_4QVal_Bool_5QNode_Bool_r)
        lizzieLet0_4QNone_Bool_4QVal_Bool_5QNode_Bool_bufchan_d <= lizzieLet0_4QNone_Bool_4QVal_Bool_5QNode_Bool_d;
  Pointer_CTf_t lizzieLet0_4QNone_Bool_4QVal_Bool_5QNode_Bool_bufchan_buf;
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_5QNode_Bool_bufchan_r = (! lizzieLet0_4QNone_Bool_4QVal_Bool_5QNode_Bool_bufchan_buf[0]);
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_5QNode_Bool_1_argbuf_d = (lizzieLet0_4QNone_Bool_4QVal_Bool_5QNode_Bool_bufchan_buf[0] ? lizzieLet0_4QNone_Bool_4QVal_Bool_5QNode_Bool_bufchan_buf :
                                                                     lizzieLet0_4QNone_Bool_4QVal_Bool_5QNode_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNone_Bool_4QVal_Bool_5QNode_Bool_bufchan_buf <= {16'd0,
                                                                    1'd0};
    else
      if ((lizzieLet0_4QNone_Bool_4QVal_Bool_5QNode_Bool_1_argbuf_r && lizzieLet0_4QNone_Bool_4QVal_Bool_5QNode_Bool_bufchan_buf[0]))
        lizzieLet0_4QNone_Bool_4QVal_Bool_5QNode_Bool_bufchan_buf <= {16'd0,
                                                                      1'd0};
      else if (((! lizzieLet0_4QNone_Bool_4QVal_Bool_5QNode_Bool_1_argbuf_r) && (! lizzieLet0_4QNone_Bool_4QVal_Bool_5QNode_Bool_bufchan_buf[0])))
        lizzieLet0_4QNone_Bool_4QVal_Bool_5QNode_Bool_bufchan_buf <= lizzieLet0_4QNone_Bool_4QVal_Bool_5QNode_Bool_bufchan_d;
  
  /* buf (Ty Pointer_CTf) : (lizzieLet0_4QNone_Bool_4QVal_Bool_5QNone_Bool,Pointer_CTf) > (lizzieLet0_4QNone_Bool_4QVal_Bool_5QNone_Bool_1_argbuf,Pointer_CTf) */
  Pointer_CTf_t lizzieLet0_4QNone_Bool_4QVal_Bool_5QNone_Bool_bufchan_d;
  logic lizzieLet0_4QNone_Bool_4QVal_Bool_5QNone_Bool_bufchan_r;
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_5QNone_Bool_r = ((! lizzieLet0_4QNone_Bool_4QVal_Bool_5QNone_Bool_bufchan_d[0]) || lizzieLet0_4QNone_Bool_4QVal_Bool_5QNone_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNone_Bool_4QVal_Bool_5QNone_Bool_bufchan_d <= {16'd0,
                                                                  1'd0};
    else
      if (lizzieLet0_4QNone_Bool_4QVal_Bool_5QNone_Bool_r)
        lizzieLet0_4QNone_Bool_4QVal_Bool_5QNone_Bool_bufchan_d <= lizzieLet0_4QNone_Bool_4QVal_Bool_5QNone_Bool_d;
  Pointer_CTf_t lizzieLet0_4QNone_Bool_4QVal_Bool_5QNone_Bool_bufchan_buf;
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_5QNone_Bool_bufchan_r = (! lizzieLet0_4QNone_Bool_4QVal_Bool_5QNone_Bool_bufchan_buf[0]);
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_5QNone_Bool_1_argbuf_d = (lizzieLet0_4QNone_Bool_4QVal_Bool_5QNone_Bool_bufchan_buf[0] ? lizzieLet0_4QNone_Bool_4QVal_Bool_5QNone_Bool_bufchan_buf :
                                                                     lizzieLet0_4QNone_Bool_4QVal_Bool_5QNone_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNone_Bool_4QVal_Bool_5QNone_Bool_bufchan_buf <= {16'd0,
                                                                    1'd0};
    else
      if ((lizzieLet0_4QNone_Bool_4QVal_Bool_5QNone_Bool_1_argbuf_r && lizzieLet0_4QNone_Bool_4QVal_Bool_5QNone_Bool_bufchan_buf[0]))
        lizzieLet0_4QNone_Bool_4QVal_Bool_5QNone_Bool_bufchan_buf <= {16'd0,
                                                                      1'd0};
      else if (((! lizzieLet0_4QNone_Bool_4QVal_Bool_5QNone_Bool_1_argbuf_r) && (! lizzieLet0_4QNone_Bool_4QVal_Bool_5QNone_Bool_bufchan_buf[0])))
        lizzieLet0_4QNone_Bool_4QVal_Bool_5QNone_Bool_bufchan_buf <= lizzieLet0_4QNone_Bool_4QVal_Bool_5QNone_Bool_bufchan_d;
  
  /* demux (Ty QTree_Bool,
       Ty MyBool) : (lizzieLet0_4QNone_Bool_4QVal_Bool_6,QTree_Bool) (v1a87_destruct,MyBool) > [(_84,MyBool),
                                                                                                (lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool,MyBool),
                                                                                                (_83,MyBool),
                                                                                                (_82,MyBool)] */
  logic [3:0] v1a87_destruct_onehotd;
  always_comb
    if ((lizzieLet0_4QNone_Bool_4QVal_Bool_6_d[0] && v1a87_destruct_d[0]))
      unique case (lizzieLet0_4QNone_Bool_4QVal_Bool_6_d[2:1])
        2'd0: v1a87_destruct_onehotd = 4'd1;
        2'd1: v1a87_destruct_onehotd = 4'd2;
        2'd2: v1a87_destruct_onehotd = 4'd4;
        2'd3: v1a87_destruct_onehotd = 4'd8;
        default: v1a87_destruct_onehotd = 4'd0;
      endcase
    else v1a87_destruct_onehotd = 4'd0;
  assign _84_d = {v1a87_destruct_d[1:1], v1a87_destruct_onehotd[0]};
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_d = {v1a87_destruct_d[1:1],
                                                           v1a87_destruct_onehotd[1]};
  assign _83_d = {v1a87_destruct_d[1:1], v1a87_destruct_onehotd[2]};
  assign _82_d = {v1a87_destruct_d[1:1], v1a87_destruct_onehotd[3]};
  assign v1a87_destruct_r = (| (v1a87_destruct_onehotd & {_82_r,
                                                          _83_r,
                                                          lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_r,
                                                          _84_r}));
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_6_r = v1a87_destruct_r;
  
  /* fork (Ty MyBool) : (lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool,MyBool) > [(lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1,MyBool),
                                                                            (lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_2,MyBool),
                                                                            (lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3,MyBool)] */
  logic [2:0] lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_emitted;
  logic [2:0] lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_done;
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1_d = {lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_d[1:1],
                                                             (lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_d[0] && (! lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_emitted[0]))};
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_2_d = {lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_d[1:1],
                                                             (lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_d[0] && (! lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_emitted[1]))};
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3_d = {lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_d[1:1],
                                                             (lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_d[0] && (! lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_emitted[2]))};
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_done = (lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_emitted | ({lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3_d[0],
                                                                                                                       lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_2_d[0],
                                                                                                                       lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1_d[0]} & {lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3_r,
                                                                                                                                                                               lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_2_r,
                                                                                                                                                                               lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1_r}));
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_r = (& lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_emitted <= 3'd0;
    else
      lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_emitted <= (lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_r ? 3'd0 :
                                                               lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_done);
  
  /* demux (Ty MyBool,
       Ty Go) : (lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1,MyBool) (lizzieLet0_4QNone_Bool_4QVal_Bool_3QVal_Bool,Go) > [(lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyFalse,Go),
                                                                                                                             (lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyTrue,Go)] */
  logic [1:0] lizzieLet0_4QNone_Bool_4QVal_Bool_3QVal_Bool_onehotd;
  always_comb
    if ((lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1_d[0] && lizzieLet0_4QNone_Bool_4QVal_Bool_3QVal_Bool_d[0]))
      unique case (lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1_d[1:1])
        1'd0: lizzieLet0_4QNone_Bool_4QVal_Bool_3QVal_Bool_onehotd = 2'd1;
        1'd1: lizzieLet0_4QNone_Bool_4QVal_Bool_3QVal_Bool_onehotd = 2'd2;
        default:
          lizzieLet0_4QNone_Bool_4QVal_Bool_3QVal_Bool_onehotd = 2'd0;
      endcase
    else lizzieLet0_4QNone_Bool_4QVal_Bool_3QVal_Bool_onehotd = 2'd0;
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyFalse_d = lizzieLet0_4QNone_Bool_4QVal_Bool_3QVal_Bool_onehotd[0];
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyTrue_d = lizzieLet0_4QNone_Bool_4QVal_Bool_3QVal_Bool_onehotd[1];
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_3QVal_Bool_r = (| (lizzieLet0_4QNone_Bool_4QVal_Bool_3QVal_Bool_onehotd & {lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyTrue_r,
                                                                                                                      lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyFalse_r}));
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1_r = lizzieLet0_4QNone_Bool_4QVal_Bool_3QVal_Bool_r;
  
  /* fork (Ty Go) : (lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyTrue,Go) > [(lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyTrue_1,Go),
                                                                            (lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyTrue_2,Go)] */
  logic [1:0] lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyTrue_emitted;
  logic [1:0] lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyTrue_done;
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyTrue_1_d = (lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyTrue_d[0] && (! lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyTrue_emitted[0]));
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyTrue_2_d = (lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyTrue_d[0] && (! lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyTrue_emitted[1]));
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyTrue_done = (lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyTrue_emitted | ({lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyTrue_2_d[0],
                                                                                                                                       lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyTrue_1_d[0]} & {lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyTrue_2_r,
                                                                                                                                                                                                       lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyTrue_1_r}));
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyTrue_r = (& lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyTrue_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyTrue_emitted <= 2'd0;
    else
      lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyTrue_emitted <= (lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyTrue_r ? 2'd0 :
                                                                       lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyTrue_done);
  
  /* buf (Ty Go) : (lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyTrue_1,Go) > (lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyTrue_1_argbuf,Go) */
  Go_t lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyTrue_1_bufchan_d;
  logic lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyTrue_1_bufchan_r;
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyTrue_1_r = ((! lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyTrue_1_bufchan_d[0]) || lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyTrue_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyTrue_1_bufchan_d <= 1'd0;
    else
      if (lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyTrue_1_r)
        lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyTrue_1_bufchan_d <= lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyTrue_1_d;
  Go_t lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyTrue_1_bufchan_buf;
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyTrue_1_bufchan_r = (! lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyTrue_1_bufchan_buf[0]);
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyTrue_1_argbuf_d = (lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyTrue_1_bufchan_buf[0] ? lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyTrue_1_bufchan_buf :
                                                                            lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyTrue_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyTrue_1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyTrue_1_argbuf_r && lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyTrue_1_bufchan_buf[0]))
        lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyTrue_1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyTrue_1_argbuf_r) && (! lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyTrue_1_bufchan_buf[0])))
        lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyTrue_1_bufchan_buf <= lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyTrue_1_bufchan_d;
  
  /* dcon (Ty TupGo,
      Dcon TupGo) : [(lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyTrue_1_argbuf,Go)] > (lvlrf2-0TupGo2,TupGo) */
  assign \lvlrf2-0TupGo2_d  = TupGo_dc((& {lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyTrue_1_argbuf_d[0]}), lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyTrue_1_argbuf_d);
  assign {lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyTrue_1_argbuf_r} = {1 {(\lvlrf2-0TupGo2_r  && \lvlrf2-0TupGo2_d [0])}};
  
  /* buf (Ty Go) : (lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyTrue_2,Go) > (lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyTrue_2_argbuf,Go) */
  Go_t lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyTrue_2_bufchan_d;
  logic lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyTrue_2_bufchan_r;
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyTrue_2_r = ((! lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyTrue_2_bufchan_d[0]) || lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyTrue_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyTrue_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyTrue_2_r)
        lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyTrue_2_bufchan_d <= lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyTrue_2_d;
  Go_t lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyTrue_2_bufchan_buf;
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyTrue_2_bufchan_r = (! lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyTrue_2_bufchan_buf[0]);
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyTrue_2_argbuf_d = (lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyTrue_2_bufchan_buf[0] ? lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyTrue_2_bufchan_buf :
                                                                            lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyTrue_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyTrue_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyTrue_2_argbuf_r && lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyTrue_2_bufchan_buf[0]))
        lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyTrue_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyTrue_2_argbuf_r) && (! lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyTrue_2_bufchan_buf[0])))
        lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyTrue_2_bufchan_buf <= lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyTrue_2_bufchan_d;
  
  /* demux (Ty MyBool,
       Ty Pointer_CTf) : (lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_2,MyBool) (lizzieLet0_4QNone_Bool_4QVal_Bool_5QVal_Bool,Pointer_CTf) > [(lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_2MyFalse,Pointer_CTf),
                                                                                                                                               (lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_2MyTrue,Pointer_CTf)] */
  logic [1:0] lizzieLet0_4QNone_Bool_4QVal_Bool_5QVal_Bool_onehotd;
  always_comb
    if ((lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_2_d[0] && lizzieLet0_4QNone_Bool_4QVal_Bool_5QVal_Bool_d[0]))
      unique case (lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_2_d[1:1])
        1'd0: lizzieLet0_4QNone_Bool_4QVal_Bool_5QVal_Bool_onehotd = 2'd1;
        1'd1: lizzieLet0_4QNone_Bool_4QVal_Bool_5QVal_Bool_onehotd = 2'd2;
        default:
          lizzieLet0_4QNone_Bool_4QVal_Bool_5QVal_Bool_onehotd = 2'd0;
      endcase
    else lizzieLet0_4QNone_Bool_4QVal_Bool_5QVal_Bool_onehotd = 2'd0;
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_2MyFalse_d = {lizzieLet0_4QNone_Bool_4QVal_Bool_5QVal_Bool_d[16:1],
                                                                    lizzieLet0_4QNone_Bool_4QVal_Bool_5QVal_Bool_onehotd[0]};
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_2MyTrue_d = {lizzieLet0_4QNone_Bool_4QVal_Bool_5QVal_Bool_d[16:1],
                                                                   lizzieLet0_4QNone_Bool_4QVal_Bool_5QVal_Bool_onehotd[1]};
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_5QVal_Bool_r = (| (lizzieLet0_4QNone_Bool_4QVal_Bool_5QVal_Bool_onehotd & {lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_2MyTrue_r,
                                                                                                                      lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_2MyFalse_r}));
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_2_r = lizzieLet0_4QNone_Bool_4QVal_Bool_5QVal_Bool_r;
  
  /* buf (Ty Pointer_CTf) : (lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_2MyTrue,Pointer_CTf) > (lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_2MyTrue_1_argbuf,Pointer_CTf) */
  Pointer_CTf_t lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_2MyTrue_bufchan_d;
  logic lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_2MyTrue_bufchan_r;
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_2MyTrue_r = ((! lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_2MyTrue_bufchan_d[0]) || lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_2MyTrue_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_2MyTrue_bufchan_d <= {16'd0,
                                                                         1'd0};
    else
      if (lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_2MyTrue_r)
        lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_2MyTrue_bufchan_d <= lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_2MyTrue_d;
  Pointer_CTf_t lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_2MyTrue_bufchan_buf;
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_2MyTrue_bufchan_r = (! lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_2MyTrue_bufchan_buf[0]);
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_2MyTrue_1_argbuf_d = (lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_2MyTrue_bufchan_buf[0] ? lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_2MyTrue_bufchan_buf :
                                                                            lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_2MyTrue_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_2MyTrue_bufchan_buf <= {16'd0,
                                                                           1'd0};
    else
      if ((lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_2MyTrue_1_argbuf_r && lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_2MyTrue_bufchan_buf[0]))
        lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_2MyTrue_bufchan_buf <= {16'd0,
                                                                             1'd0};
      else if (((! lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_2MyTrue_1_argbuf_r) && (! lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_2MyTrue_bufchan_buf[0])))
        lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_2MyTrue_bufchan_buf <= lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_2MyTrue_bufchan_d;
  
  /* demux (Ty MyBool,
       Ty MyBool) : (lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3,MyBool) (va88_destruct,MyBool) > [(lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse,MyBool),
                                                                                                      (_81,MyBool)] */
  logic [1:0] va88_destruct_onehotd;
  always_comb
    if ((lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3_d[0] && va88_destruct_d[0]))
      unique case (lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3_d[1:1])
        1'd0: va88_destruct_onehotd = 2'd1;
        1'd1: va88_destruct_onehotd = 2'd2;
        default: va88_destruct_onehotd = 2'd0;
      endcase
    else va88_destruct_onehotd = 2'd0;
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_d = {va88_destruct_d[1:1],
                                                                    va88_destruct_onehotd[0]};
  assign _81_d = {va88_destruct_d[1:1], va88_destruct_onehotd[1]};
  assign va88_destruct_r = (| (va88_destruct_onehotd & {_81_r,
                                                        lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_r}));
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3_r = va88_destruct_r;
  
  /* fork (Ty MyBool) : (lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse,MyBool) > [(lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1,MyBool),
                                                                                     (lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_2,MyBool)] */
  logic [1:0] lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_emitted;
  logic [1:0] lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_done;
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1_d = {lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_d[1:1],
                                                                      (lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_d[0] && (! lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_emitted[0]))};
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_2_d = {lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_d[1:1],
                                                                      (lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_d[0] && (! lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_emitted[1]))};
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_done = (lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_emitted | ({lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_2_d[0],
                                                                                                                                         lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1_d[0]} & {lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_2_r,
                                                                                                                                                                                                          lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1_r}));
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_r = (& lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_emitted <= 2'd0;
    else
      lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_emitted <= (lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_r ? 2'd0 :
                                                                        lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_done);
  
  /* demux (Ty MyBool,
       Ty Go) : (lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1,MyBool) (lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyFalse,Go) > [(lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse,Go),
                                                                                                                                               (lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue,Go)] */
  logic [1:0] lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyFalse_onehotd;
  always_comb
    if ((lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1_d[0] && lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyFalse_d[0]))
      unique case (lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1_d[1:1])
        1'd0:
          lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyFalse_onehotd = 2'd1;
        1'd1:
          lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyFalse_onehotd = 2'd2;
        default:
          lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyFalse_onehotd = 2'd0;
      endcase
    else
      lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyFalse_onehotd = 2'd0;
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_d = lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyFalse_onehotd[0];
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_d = lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyFalse_onehotd[1];
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyFalse_r = (| (lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyFalse_onehotd & {lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_r,
                                                                                                                                        lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_r}));
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1_r = lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_1MyFalse_r;
  
  /* fork (Ty Go) : (lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse,Go) > [(lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1,Go),
                                                                                      (lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2,Go)] */
  logic [1:0] lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_emitted;
  logic [1:0] lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_done;
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1_d = (lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_d[0] && (! lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_emitted[0]));
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_d = (lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_d[0] && (! lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_emitted[1]));
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_done = (lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_emitted | ({lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_d[0],
                                                                                                                                                           lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1_d[0]} & {lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_r,
                                                                                                                                                                                                                                     lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1_r}));
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_r = (& lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_emitted <= 2'd0;
    else
      lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_emitted <= (lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_r ? 2'd0 :
                                                                                 lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_done);
  
  /* dcon (Ty QTree_Bool,
      Dcon QNone_Bool) : [(lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1,Go)] > (lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool,QTree_Bool) */
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_d = QNone_Bool_dc((& {lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1_d[0]}), lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1_d);
  assign {lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1_r} = {1 {(lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_r && lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_d[0])}};
  
  /* buf (Ty QTree_Bool) : (lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool,QTree_Bool) > (lizzieLet3_1_argbuf,QTree_Bool) */
  QTree_Bool_t lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_bufchan_d;
  logic lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_bufchan_r;
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_r = ((! lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_bufchan_d[0]) || lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_bufchan_d <= {66'd0,
                                                                                               1'd0};
    else
      if (lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_r)
        lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_bufchan_d <= lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_d;
  QTree_Bool_t lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_bufchan_buf;
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_bufchan_r = (! lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_bufchan_buf[0]);
  assign lizzieLet3_1_argbuf_d = (lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_bufchan_buf[0] ? lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_bufchan_buf :
                                  lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_bufchan_buf <= {66'd0,
                                                                                                 1'd0};
    else
      if ((lizzieLet3_1_argbuf_r && lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_bufchan_buf[0]))
        lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_bufchan_buf <= {66'd0,
                                                                                                   1'd0};
      else if (((! lizzieLet3_1_argbuf_r) && (! lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_bufchan_buf[0])))
        lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_bufchan_buf <= lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2,Go) > (lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_argbuf,Go) */
  Go_t lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_bufchan_d;
  logic lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_bufchan_r;
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_r = ((! lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_bufchan_d[0]) || lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_r)
        lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_bufchan_d <= lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_d;
  Go_t lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_bufchan_buf;
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_bufchan_r = (! lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_bufchan_buf[0]);
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_argbuf_d = (lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_bufchan_buf[0] ? lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_bufchan_buf :
                                                                                      lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_argbuf_r && lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_bufchan_buf[0]))
        lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_argbuf_r) && (! lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_bufchan_buf[0])))
        lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_bufchan_buf <= lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue,Go) > [(lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1,Go),
                                                                                     (lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2,Go)] */
  logic [1:0] lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_emitted;
  logic [1:0] lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_done;
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_d = (lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_d[0] && (! lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_emitted[0]));
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_d = (lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_d[0] && (! lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_emitted[1]));
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_done = (lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_emitted | ({lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_d[0],
                                                                                                                                                         lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_d[0]} & {lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_r,
                                                                                                                                                                                                                                  lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_r}));
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_r = (& lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_emitted <= 2'd0;
    else
      lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_emitted <= (lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_r ? 2'd0 :
                                                                                lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_done);
  
  /* buf (Ty Go) : (lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1,Go) > (lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_argbuf,Go) */
  Go_t lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_bufchan_d;
  logic lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_bufchan_r;
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_r = ((! lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_bufchan_d[0]) || lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_bufchan_d <= 1'd0;
    else
      if (lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_r)
        lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_bufchan_d <= lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_d;
  Go_t lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_bufchan_buf;
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_bufchan_r = (! lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_bufchan_buf[0]);
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_argbuf_d = (lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_bufchan_buf[0] ? lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_bufchan_buf :
                                                                                     lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_argbuf_r && lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_bufchan_buf[0]))
        lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_argbuf_r) && (! lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_bufchan_buf[0])))
        lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_bufchan_buf <= lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_bufchan_d;
  
  /* dcon (Ty TupGo,
      Dcon TupGo) : [(lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_argbuf,Go)] > (lvlrf2-0TupGo_1,TupGo) */
  assign \lvlrf2-0TupGo_1_d  = TupGo_dc((& {lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_argbuf_d[0]}), lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_argbuf_d);
  assign {lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_argbuf_r} = {1 {(\lvlrf2-0TupGo_1_r  && \lvlrf2-0TupGo_1_d [0])}};
  
  /* buf (Ty Go) : (lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2,Go) > (lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_argbuf,Go) */
  Go_t lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_bufchan_d;
  logic lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_bufchan_r;
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_r = ((! lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_bufchan_d[0]) || lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_r)
        lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_bufchan_d <= lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_d;
  Go_t lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_bufchan_buf;
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_bufchan_r = (! lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_bufchan_buf[0]);
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_argbuf_d = (lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_bufchan_buf[0] ? lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_bufchan_buf :
                                                                                     lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_argbuf_r && lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_bufchan_buf[0]))
        lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_argbuf_r) && (! lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_bufchan_buf[0])))
        lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_bufchan_buf <= lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_bufchan_d;
  
  /* demux (Ty MyBool,
       Ty Pointer_CTf) : (lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_2,MyBool) (lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_2MyFalse,Pointer_CTf) > [(lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_2MyFalse,Pointer_CTf),
                                                                                                                                                                 (lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_2MyTrue,Pointer_CTf)] */
  logic [1:0] lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_2MyFalse_onehotd;
  always_comb
    if ((lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_2_d[0] && lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_2MyFalse_d[0]))
      unique case (lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_2_d[1:1])
        1'd0:
          lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_2MyFalse_onehotd = 2'd1;
        1'd1:
          lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_2MyFalse_onehotd = 2'd2;
        default:
          lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_2MyFalse_onehotd = 2'd0;
      endcase
    else
      lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_2MyFalse_onehotd = 2'd0;
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_2MyFalse_d = {lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_2MyFalse_d[16:1],
                                                                             lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_2MyFalse_onehotd[0]};
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_2MyTrue_d = {lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_2MyFalse_d[16:1],
                                                                            lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_2MyFalse_onehotd[1]};
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_2MyFalse_r = (| (lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_2MyFalse_onehotd & {lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_2MyTrue_r,
                                                                                                                                        lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_2MyFalse_r}));
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_2_r = lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_2MyFalse_r;
  
  /* buf (Ty Pointer_CTf) : (lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_2MyFalse,Pointer_CTf) > (lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_2MyFalse_1_argbuf,Pointer_CTf) */
  Pointer_CTf_t lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_2MyFalse_bufchan_d;
  logic lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_2MyFalse_bufchan_r;
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_2MyFalse_r = ((! lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_2MyFalse_bufchan_d[0]) || lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_2MyFalse_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_2MyFalse_bufchan_d <= {16'd0,
                                                                                   1'd0};
    else
      if (lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_2MyFalse_r)
        lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_2MyFalse_bufchan_d <= lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_2MyFalse_d;
  Pointer_CTf_t lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_2MyFalse_bufchan_buf;
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_2MyFalse_bufchan_r = (! lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_2MyFalse_bufchan_buf[0]);
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_2MyFalse_1_argbuf_d = (lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_2MyFalse_bufchan_buf[0] ? lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_2MyFalse_bufchan_buf :
                                                                                      lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_2MyFalse_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_2MyFalse_bufchan_buf <= {16'd0,
                                                                                     1'd0};
    else
      if ((lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_2MyFalse_1_argbuf_r && lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_2MyFalse_bufchan_buf[0]))
        lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_2MyFalse_bufchan_buf <= {16'd0,
                                                                                       1'd0};
      else if (((! lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_2MyFalse_1_argbuf_r) && (! lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_2MyFalse_bufchan_buf[0])))
        lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_2MyFalse_bufchan_buf <= lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_2MyFalse_bufchan_d;
  
  /* buf (Ty Pointer_CTf) : (lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_2MyTrue,Pointer_CTf) > (lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_2MyTrue_1_argbuf,Pointer_CTf) */
  Pointer_CTf_t lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_2MyTrue_bufchan_d;
  logic lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_2MyTrue_bufchan_r;
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_2MyTrue_r = ((! lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_2MyTrue_bufchan_d[0]) || lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_2MyTrue_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_2MyTrue_bufchan_d <= {16'd0,
                                                                                  1'd0};
    else
      if (lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_2MyTrue_r)
        lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_2MyTrue_bufchan_d <= lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_2MyTrue_d;
  Pointer_CTf_t lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_2MyTrue_bufchan_buf;
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_2MyTrue_bufchan_r = (! lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_2MyTrue_bufchan_buf[0]);
  assign lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_2MyTrue_1_argbuf_d = (lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_2MyTrue_bufchan_buf[0] ? lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_2MyTrue_bufchan_buf :
                                                                                     lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_2MyTrue_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_2MyTrue_bufchan_buf <= {16'd0,
                                                                                    1'd0};
    else
      if ((lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_2MyTrue_1_argbuf_r && lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_2MyTrue_bufchan_buf[0]))
        lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_2MyTrue_bufchan_buf <= {16'd0,
                                                                                      1'd0};
      else if (((! lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_2MyTrue_1_argbuf_r) && (! lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_2MyTrue_bufchan_buf[0])))
        lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_2MyTrue_bufchan_buf <= lizzieLet0_4QNone_Bool_4QVal_Bool_6QVal_Bool_3MyFalse_2MyTrue_bufchan_d;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_QTree_Bool) : (lizzieLet0_4QNone_Bool_5,QTree_Bool) (lizzieLet0_7QNone_Bool,Pointer_QTree_Bool) > [(_80,Pointer_QTree_Bool),
                                                                                                                     (lizzieLet0_4QNone_Bool_5QVal_Bool,Pointer_QTree_Bool),
                                                                                                                     (lizzieLet0_4QNone_Bool_5QNode_Bool,Pointer_QTree_Bool),
                                                                                                                     (_79,Pointer_QTree_Bool)] */
  logic [3:0] lizzieLet0_7QNone_Bool_onehotd;
  always_comb
    if ((lizzieLet0_4QNone_Bool_5_d[0] && lizzieLet0_7QNone_Bool_d[0]))
      unique case (lizzieLet0_4QNone_Bool_5_d[2:1])
        2'd0: lizzieLet0_7QNone_Bool_onehotd = 4'd1;
        2'd1: lizzieLet0_7QNone_Bool_onehotd = 4'd2;
        2'd2: lizzieLet0_7QNone_Bool_onehotd = 4'd4;
        2'd3: lizzieLet0_7QNone_Bool_onehotd = 4'd8;
        default: lizzieLet0_7QNone_Bool_onehotd = 4'd0;
      endcase
    else lizzieLet0_7QNone_Bool_onehotd = 4'd0;
  assign _80_d = {lizzieLet0_7QNone_Bool_d[16:1],
                  lizzieLet0_7QNone_Bool_onehotd[0]};
  assign lizzieLet0_4QNone_Bool_5QVal_Bool_d = {lizzieLet0_7QNone_Bool_d[16:1],
                                                lizzieLet0_7QNone_Bool_onehotd[1]};
  assign lizzieLet0_4QNone_Bool_5QNode_Bool_d = {lizzieLet0_7QNone_Bool_d[16:1],
                                                 lizzieLet0_7QNone_Bool_onehotd[2]};
  assign _79_d = {lizzieLet0_7QNone_Bool_d[16:1],
                  lizzieLet0_7QNone_Bool_onehotd[3]};
  assign lizzieLet0_7QNone_Bool_r = (| (lizzieLet0_7QNone_Bool_onehotd & {_79_r,
                                                                          lizzieLet0_4QNone_Bool_5QNode_Bool_r,
                                                                          lizzieLet0_4QNone_Bool_5QVal_Bool_r,
                                                                          _80_r}));
  assign lizzieLet0_4QNone_Bool_5_r = lizzieLet0_7QNone_Bool_r;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_QTree_Bool) : (lizzieLet0_4QNone_Bool_6,QTree_Bool) (lizzieLet0_8QNone_Bool,Pointer_QTree_Bool) > [(lizzieLet0_4QNone_Bool_6QNone_Bool,Pointer_QTree_Bool),
                                                                                                                     (_78,Pointer_QTree_Bool),
                                                                                                                     (_77,Pointer_QTree_Bool),
                                                                                                                     (_76,Pointer_QTree_Bool)] */
  logic [3:0] lizzieLet0_8QNone_Bool_onehotd;
  always_comb
    if ((lizzieLet0_4QNone_Bool_6_d[0] && lizzieLet0_8QNone_Bool_d[0]))
      unique case (lizzieLet0_4QNone_Bool_6_d[2:1])
        2'd0: lizzieLet0_8QNone_Bool_onehotd = 4'd1;
        2'd1: lizzieLet0_8QNone_Bool_onehotd = 4'd2;
        2'd2: lizzieLet0_8QNone_Bool_onehotd = 4'd4;
        2'd3: lizzieLet0_8QNone_Bool_onehotd = 4'd8;
        default: lizzieLet0_8QNone_Bool_onehotd = 4'd0;
      endcase
    else lizzieLet0_8QNone_Bool_onehotd = 4'd0;
  assign lizzieLet0_4QNone_Bool_6QNone_Bool_d = {lizzieLet0_8QNone_Bool_d[16:1],
                                                 lizzieLet0_8QNone_Bool_onehotd[0]};
  assign _78_d = {lizzieLet0_8QNone_Bool_d[16:1],
                  lizzieLet0_8QNone_Bool_onehotd[1]};
  assign _77_d = {lizzieLet0_8QNone_Bool_d[16:1],
                  lizzieLet0_8QNone_Bool_onehotd[2]};
  assign _76_d = {lizzieLet0_8QNone_Bool_d[16:1],
                  lizzieLet0_8QNone_Bool_onehotd[3]};
  assign lizzieLet0_8QNone_Bool_r = (| (lizzieLet0_8QNone_Bool_onehotd & {_76_r,
                                                                          _77_r,
                                                                          _78_r,
                                                                          lizzieLet0_4QNone_Bool_6QNone_Bool_r}));
  assign lizzieLet0_4QNone_Bool_6_r = lizzieLet0_8QNone_Bool_r;
  
  /* buf (Ty Pointer_QTree_Bool) : (lizzieLet0_4QNone_Bool_6QNone_Bool,Pointer_QTree_Bool) > (lizzieLet0_4QNone_Bool_6QNone_Bool_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t lizzieLet0_4QNone_Bool_6QNone_Bool_bufchan_d;
  logic lizzieLet0_4QNone_Bool_6QNone_Bool_bufchan_r;
  assign lizzieLet0_4QNone_Bool_6QNone_Bool_r = ((! lizzieLet0_4QNone_Bool_6QNone_Bool_bufchan_d[0]) || lizzieLet0_4QNone_Bool_6QNone_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNone_Bool_6QNone_Bool_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet0_4QNone_Bool_6QNone_Bool_r)
        lizzieLet0_4QNone_Bool_6QNone_Bool_bufchan_d <= lizzieLet0_4QNone_Bool_6QNone_Bool_d;
  Pointer_QTree_Bool_t lizzieLet0_4QNone_Bool_6QNone_Bool_bufchan_buf;
  assign lizzieLet0_4QNone_Bool_6QNone_Bool_bufchan_r = (! lizzieLet0_4QNone_Bool_6QNone_Bool_bufchan_buf[0]);
  assign lizzieLet0_4QNone_Bool_6QNone_Bool_1_argbuf_d = (lizzieLet0_4QNone_Bool_6QNone_Bool_bufchan_buf[0] ? lizzieLet0_4QNone_Bool_6QNone_Bool_bufchan_buf :
                                                          lizzieLet0_4QNone_Bool_6QNone_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNone_Bool_6QNone_Bool_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet0_4QNone_Bool_6QNone_Bool_1_argbuf_r && lizzieLet0_4QNone_Bool_6QNone_Bool_bufchan_buf[0]))
        lizzieLet0_4QNone_Bool_6QNone_Bool_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet0_4QNone_Bool_6QNone_Bool_1_argbuf_r) && (! lizzieLet0_4QNone_Bool_6QNone_Bool_bufchan_buf[0])))
        lizzieLet0_4QNone_Bool_6QNone_Bool_bufchan_buf <= lizzieLet0_4QNone_Bool_6QNone_Bool_bufchan_d;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_CTf) : (lizzieLet0_4QNone_Bool_7,QTree_Bool) (lizzieLet0_9QNone_Bool,Pointer_CTf) > [(lizzieLet0_4QNone_Bool_7QNone_Bool,Pointer_CTf),
                                                                                                       (lizzieLet0_4QNone_Bool_7QVal_Bool,Pointer_CTf),
                                                                                                       (lizzieLet0_4QNone_Bool_7QNode_Bool,Pointer_CTf),
                                                                                                       (lizzieLet0_4QNone_Bool_7QError_Bool,Pointer_CTf)] */
  logic [3:0] lizzieLet0_9QNone_Bool_onehotd;
  always_comb
    if ((lizzieLet0_4QNone_Bool_7_d[0] && lizzieLet0_9QNone_Bool_d[0]))
      unique case (lizzieLet0_4QNone_Bool_7_d[2:1])
        2'd0: lizzieLet0_9QNone_Bool_onehotd = 4'd1;
        2'd1: lizzieLet0_9QNone_Bool_onehotd = 4'd2;
        2'd2: lizzieLet0_9QNone_Bool_onehotd = 4'd4;
        2'd3: lizzieLet0_9QNone_Bool_onehotd = 4'd8;
        default: lizzieLet0_9QNone_Bool_onehotd = 4'd0;
      endcase
    else lizzieLet0_9QNone_Bool_onehotd = 4'd0;
  assign lizzieLet0_4QNone_Bool_7QNone_Bool_d = {lizzieLet0_9QNone_Bool_d[16:1],
                                                 lizzieLet0_9QNone_Bool_onehotd[0]};
  assign lizzieLet0_4QNone_Bool_7QVal_Bool_d = {lizzieLet0_9QNone_Bool_d[16:1],
                                                lizzieLet0_9QNone_Bool_onehotd[1]};
  assign lizzieLet0_4QNone_Bool_7QNode_Bool_d = {lizzieLet0_9QNone_Bool_d[16:1],
                                                 lizzieLet0_9QNone_Bool_onehotd[2]};
  assign lizzieLet0_4QNone_Bool_7QError_Bool_d = {lizzieLet0_9QNone_Bool_d[16:1],
                                                  lizzieLet0_9QNone_Bool_onehotd[3]};
  assign lizzieLet0_9QNone_Bool_r = (| (lizzieLet0_9QNone_Bool_onehotd & {lizzieLet0_4QNone_Bool_7QError_Bool_r,
                                                                          lizzieLet0_4QNone_Bool_7QNode_Bool_r,
                                                                          lizzieLet0_4QNone_Bool_7QVal_Bool_r,
                                                                          lizzieLet0_4QNone_Bool_7QNone_Bool_r}));
  assign lizzieLet0_4QNone_Bool_7_r = lizzieLet0_9QNone_Bool_r;
  
  /* buf (Ty Pointer_CTf) : (lizzieLet0_4QNone_Bool_7QError_Bool,Pointer_CTf) > (lizzieLet0_4QNone_Bool_7QError_Bool_1_argbuf,Pointer_CTf) */
  Pointer_CTf_t lizzieLet0_4QNone_Bool_7QError_Bool_bufchan_d;
  logic lizzieLet0_4QNone_Bool_7QError_Bool_bufchan_r;
  assign lizzieLet0_4QNone_Bool_7QError_Bool_r = ((! lizzieLet0_4QNone_Bool_7QError_Bool_bufchan_d[0]) || lizzieLet0_4QNone_Bool_7QError_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNone_Bool_7QError_Bool_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet0_4QNone_Bool_7QError_Bool_r)
        lizzieLet0_4QNone_Bool_7QError_Bool_bufchan_d <= lizzieLet0_4QNone_Bool_7QError_Bool_d;
  Pointer_CTf_t lizzieLet0_4QNone_Bool_7QError_Bool_bufchan_buf;
  assign lizzieLet0_4QNone_Bool_7QError_Bool_bufchan_r = (! lizzieLet0_4QNone_Bool_7QError_Bool_bufchan_buf[0]);
  assign lizzieLet0_4QNone_Bool_7QError_Bool_1_argbuf_d = (lizzieLet0_4QNone_Bool_7QError_Bool_bufchan_buf[0] ? lizzieLet0_4QNone_Bool_7QError_Bool_bufchan_buf :
                                                           lizzieLet0_4QNone_Bool_7QError_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNone_Bool_7QError_Bool_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet0_4QNone_Bool_7QError_Bool_1_argbuf_r && lizzieLet0_4QNone_Bool_7QError_Bool_bufchan_buf[0]))
        lizzieLet0_4QNone_Bool_7QError_Bool_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet0_4QNone_Bool_7QError_Bool_1_argbuf_r) && (! lizzieLet0_4QNone_Bool_7QError_Bool_bufchan_buf[0])))
        lizzieLet0_4QNone_Bool_7QError_Bool_bufchan_buf <= lizzieLet0_4QNone_Bool_7QError_Bool_bufchan_d;
  
  /* buf (Ty Pointer_CTf) : (lizzieLet0_4QNone_Bool_7QNone_Bool,Pointer_CTf) > (lizzieLet0_4QNone_Bool_7QNone_Bool_1_argbuf,Pointer_CTf) */
  Pointer_CTf_t lizzieLet0_4QNone_Bool_7QNone_Bool_bufchan_d;
  logic lizzieLet0_4QNone_Bool_7QNone_Bool_bufchan_r;
  assign lizzieLet0_4QNone_Bool_7QNone_Bool_r = ((! lizzieLet0_4QNone_Bool_7QNone_Bool_bufchan_d[0]) || lizzieLet0_4QNone_Bool_7QNone_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNone_Bool_7QNone_Bool_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet0_4QNone_Bool_7QNone_Bool_r)
        lizzieLet0_4QNone_Bool_7QNone_Bool_bufchan_d <= lizzieLet0_4QNone_Bool_7QNone_Bool_d;
  Pointer_CTf_t lizzieLet0_4QNone_Bool_7QNone_Bool_bufchan_buf;
  assign lizzieLet0_4QNone_Bool_7QNone_Bool_bufchan_r = (! lizzieLet0_4QNone_Bool_7QNone_Bool_bufchan_buf[0]);
  assign lizzieLet0_4QNone_Bool_7QNone_Bool_1_argbuf_d = (lizzieLet0_4QNone_Bool_7QNone_Bool_bufchan_buf[0] ? lizzieLet0_4QNone_Bool_7QNone_Bool_bufchan_buf :
                                                          lizzieLet0_4QNone_Bool_7QNone_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNone_Bool_7QNone_Bool_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet0_4QNone_Bool_7QNone_Bool_1_argbuf_r && lizzieLet0_4QNone_Bool_7QNone_Bool_bufchan_buf[0]))
        lizzieLet0_4QNone_Bool_7QNone_Bool_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet0_4QNone_Bool_7QNone_Bool_1_argbuf_r) && (! lizzieLet0_4QNone_Bool_7QNone_Bool_bufchan_buf[0])))
        lizzieLet0_4QNone_Bool_7QNone_Bool_bufchan_buf <= lizzieLet0_4QNone_Bool_7QNone_Bool_bufchan_d;
  
  /* fork (Ty QTree_Bool) : (lizzieLet0_4QVal_Bool,QTree_Bool) > [(lizzieLet0_4QVal_Bool_1,QTree_Bool),
                                                             (lizzieLet0_4QVal_Bool_2,QTree_Bool),
                                                             (lizzieLet0_4QVal_Bool_3,QTree_Bool),
                                                             (lizzieLet0_4QVal_Bool_4,QTree_Bool),
                                                             (lizzieLet0_4QVal_Bool_5,QTree_Bool),
                                                             (lizzieLet0_4QVal_Bool_6,QTree_Bool),
                                                             (lizzieLet0_4QVal_Bool_7,QTree_Bool),
                                                             (lizzieLet0_4QVal_Bool_8,QTree_Bool)] */
  logic [7:0] lizzieLet0_4QVal_Bool_emitted;
  logic [7:0] lizzieLet0_4QVal_Bool_done;
  assign lizzieLet0_4QVal_Bool_1_d = {lizzieLet0_4QVal_Bool_d[66:1],
                                      (lizzieLet0_4QVal_Bool_d[0] && (! lizzieLet0_4QVal_Bool_emitted[0]))};
  assign lizzieLet0_4QVal_Bool_2_d = {lizzieLet0_4QVal_Bool_d[66:1],
                                      (lizzieLet0_4QVal_Bool_d[0] && (! lizzieLet0_4QVal_Bool_emitted[1]))};
  assign lizzieLet0_4QVal_Bool_3_d = {lizzieLet0_4QVal_Bool_d[66:1],
                                      (lizzieLet0_4QVal_Bool_d[0] && (! lizzieLet0_4QVal_Bool_emitted[2]))};
  assign lizzieLet0_4QVal_Bool_4_d = {lizzieLet0_4QVal_Bool_d[66:1],
                                      (lizzieLet0_4QVal_Bool_d[0] && (! lizzieLet0_4QVal_Bool_emitted[3]))};
  assign lizzieLet0_4QVal_Bool_5_d = {lizzieLet0_4QVal_Bool_d[66:1],
                                      (lizzieLet0_4QVal_Bool_d[0] && (! lizzieLet0_4QVal_Bool_emitted[4]))};
  assign lizzieLet0_4QVal_Bool_6_d = {lizzieLet0_4QVal_Bool_d[66:1],
                                      (lizzieLet0_4QVal_Bool_d[0] && (! lizzieLet0_4QVal_Bool_emitted[5]))};
  assign lizzieLet0_4QVal_Bool_7_d = {lizzieLet0_4QVal_Bool_d[66:1],
                                      (lizzieLet0_4QVal_Bool_d[0] && (! lizzieLet0_4QVal_Bool_emitted[6]))};
  assign lizzieLet0_4QVal_Bool_8_d = {lizzieLet0_4QVal_Bool_d[66:1],
                                      (lizzieLet0_4QVal_Bool_d[0] && (! lizzieLet0_4QVal_Bool_emitted[7]))};
  assign lizzieLet0_4QVal_Bool_done = (lizzieLet0_4QVal_Bool_emitted | ({lizzieLet0_4QVal_Bool_8_d[0],
                                                                         lizzieLet0_4QVal_Bool_7_d[0],
                                                                         lizzieLet0_4QVal_Bool_6_d[0],
                                                                         lizzieLet0_4QVal_Bool_5_d[0],
                                                                         lizzieLet0_4QVal_Bool_4_d[0],
                                                                         lizzieLet0_4QVal_Bool_3_d[0],
                                                                         lizzieLet0_4QVal_Bool_2_d[0],
                                                                         lizzieLet0_4QVal_Bool_1_d[0]} & {lizzieLet0_4QVal_Bool_8_r,
                                                                                                          lizzieLet0_4QVal_Bool_7_r,
                                                                                                          lizzieLet0_4QVal_Bool_6_r,
                                                                                                          lizzieLet0_4QVal_Bool_5_r,
                                                                                                          lizzieLet0_4QVal_Bool_4_r,
                                                                                                          lizzieLet0_4QVal_Bool_3_r,
                                                                                                          lizzieLet0_4QVal_Bool_2_r,
                                                                                                          lizzieLet0_4QVal_Bool_1_r}));
  assign lizzieLet0_4QVal_Bool_r = (& lizzieLet0_4QVal_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet0_4QVal_Bool_emitted <= 8'd0;
    else
      lizzieLet0_4QVal_Bool_emitted <= (lizzieLet0_4QVal_Bool_r ? 8'd0 :
                                        lizzieLet0_4QVal_Bool_done);
  
  /* destruct (Ty QTree_Bool,
          Dcon QVal_Bool) : (lizzieLet0_4QVal_Bool_1QVal_Bool,QTree_Bool) > [(va8s_destruct,MyBool)] */
  assign va8s_destruct_d = {lizzieLet0_4QVal_Bool_1QVal_Bool_d[3:3],
                            lizzieLet0_4QVal_Bool_1QVal_Bool_d[0]};
  assign lizzieLet0_4QVal_Bool_1QVal_Bool_r = va8s_destruct_r;
  
  /* demux (Ty QTree_Bool,
       Ty QTree_Bool) : (lizzieLet0_4QVal_Bool_2,QTree_Bool) (lizzieLet0_4QVal_Bool_1,QTree_Bool) > [(_75,QTree_Bool),
                                                                                                     (lizzieLet0_4QVal_Bool_1QVal_Bool,QTree_Bool),
                                                                                                     (_74,QTree_Bool),
                                                                                                     (_73,QTree_Bool)] */
  logic [3:0] lizzieLet0_4QVal_Bool_1_onehotd;
  always_comb
    if ((lizzieLet0_4QVal_Bool_2_d[0] && lizzieLet0_4QVal_Bool_1_d[0]))
      unique case (lizzieLet0_4QVal_Bool_2_d[2:1])
        2'd0: lizzieLet0_4QVal_Bool_1_onehotd = 4'd1;
        2'd1: lizzieLet0_4QVal_Bool_1_onehotd = 4'd2;
        2'd2: lizzieLet0_4QVal_Bool_1_onehotd = 4'd4;
        2'd3: lizzieLet0_4QVal_Bool_1_onehotd = 4'd8;
        default: lizzieLet0_4QVal_Bool_1_onehotd = 4'd0;
      endcase
    else lizzieLet0_4QVal_Bool_1_onehotd = 4'd0;
  assign _75_d = {lizzieLet0_4QVal_Bool_1_d[66:1],
                  lizzieLet0_4QVal_Bool_1_onehotd[0]};
  assign lizzieLet0_4QVal_Bool_1QVal_Bool_d = {lizzieLet0_4QVal_Bool_1_d[66:1],
                                               lizzieLet0_4QVal_Bool_1_onehotd[1]};
  assign _74_d = {lizzieLet0_4QVal_Bool_1_d[66:1],
                  lizzieLet0_4QVal_Bool_1_onehotd[2]};
  assign _73_d = {lizzieLet0_4QVal_Bool_1_d[66:1],
                  lizzieLet0_4QVal_Bool_1_onehotd[3]};
  assign lizzieLet0_4QVal_Bool_1_r = (| (lizzieLet0_4QVal_Bool_1_onehotd & {_73_r,
                                                                            _74_r,
                                                                            lizzieLet0_4QVal_Bool_1QVal_Bool_r,
                                                                            _75_r}));
  assign lizzieLet0_4QVal_Bool_2_r = lizzieLet0_4QVal_Bool_1_r;
  
  /* demux (Ty QTree_Bool,
       Ty Go) : (lizzieLet0_4QVal_Bool_3,QTree_Bool) (lizzieLet0_3QVal_Bool,Go) > [(lizzieLet0_4QVal_Bool_3QNone_Bool,Go),
                                                                                   (lizzieLet0_4QVal_Bool_3QVal_Bool,Go),
                                                                                   (lizzieLet0_4QVal_Bool_3QNode_Bool,Go),
                                                                                   (lizzieLet0_4QVal_Bool_3QError_Bool,Go)] */
  logic [3:0] lizzieLet0_3QVal_Bool_onehotd;
  always_comb
    if ((lizzieLet0_4QVal_Bool_3_d[0] && lizzieLet0_3QVal_Bool_d[0]))
      unique case (lizzieLet0_4QVal_Bool_3_d[2:1])
        2'd0: lizzieLet0_3QVal_Bool_onehotd = 4'd1;
        2'd1: lizzieLet0_3QVal_Bool_onehotd = 4'd2;
        2'd2: lizzieLet0_3QVal_Bool_onehotd = 4'd4;
        2'd3: lizzieLet0_3QVal_Bool_onehotd = 4'd8;
        default: lizzieLet0_3QVal_Bool_onehotd = 4'd0;
      endcase
    else lizzieLet0_3QVal_Bool_onehotd = 4'd0;
  assign lizzieLet0_4QVal_Bool_3QNone_Bool_d = lizzieLet0_3QVal_Bool_onehotd[0];
  assign lizzieLet0_4QVal_Bool_3QVal_Bool_d = lizzieLet0_3QVal_Bool_onehotd[1];
  assign lizzieLet0_4QVal_Bool_3QNode_Bool_d = lizzieLet0_3QVal_Bool_onehotd[2];
  assign lizzieLet0_4QVal_Bool_3QError_Bool_d = lizzieLet0_3QVal_Bool_onehotd[3];
  assign lizzieLet0_3QVal_Bool_r = (| (lizzieLet0_3QVal_Bool_onehotd & {lizzieLet0_4QVal_Bool_3QError_Bool_r,
                                                                        lizzieLet0_4QVal_Bool_3QNode_Bool_r,
                                                                        lizzieLet0_4QVal_Bool_3QVal_Bool_r,
                                                                        lizzieLet0_4QVal_Bool_3QNone_Bool_r}));
  assign lizzieLet0_4QVal_Bool_3_r = lizzieLet0_3QVal_Bool_r;
  
  /* fork (Ty Go) : (lizzieLet0_4QVal_Bool_3QError_Bool,Go) > [(lizzieLet0_4QVal_Bool_3QError_Bool_1,Go),
                                                          (lizzieLet0_4QVal_Bool_3QError_Bool_2,Go)] */
  logic [1:0] lizzieLet0_4QVal_Bool_3QError_Bool_emitted;
  logic [1:0] lizzieLet0_4QVal_Bool_3QError_Bool_done;
  assign lizzieLet0_4QVal_Bool_3QError_Bool_1_d = (lizzieLet0_4QVal_Bool_3QError_Bool_d[0] && (! lizzieLet0_4QVal_Bool_3QError_Bool_emitted[0]));
  assign lizzieLet0_4QVal_Bool_3QError_Bool_2_d = (lizzieLet0_4QVal_Bool_3QError_Bool_d[0] && (! lizzieLet0_4QVal_Bool_3QError_Bool_emitted[1]));
  assign lizzieLet0_4QVal_Bool_3QError_Bool_done = (lizzieLet0_4QVal_Bool_3QError_Bool_emitted | ({lizzieLet0_4QVal_Bool_3QError_Bool_2_d[0],
                                                                                                   lizzieLet0_4QVal_Bool_3QError_Bool_1_d[0]} & {lizzieLet0_4QVal_Bool_3QError_Bool_2_r,
                                                                                                                                                 lizzieLet0_4QVal_Bool_3QError_Bool_1_r}));
  assign lizzieLet0_4QVal_Bool_3QError_Bool_r = (& lizzieLet0_4QVal_Bool_3QError_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_3QError_Bool_emitted <= 2'd0;
    else
      lizzieLet0_4QVal_Bool_3QError_Bool_emitted <= (lizzieLet0_4QVal_Bool_3QError_Bool_r ? 2'd0 :
                                                     lizzieLet0_4QVal_Bool_3QError_Bool_done);
  
  /* dcon (Ty QTree_Bool,
      Dcon QError_Bool) : [(lizzieLet0_4QVal_Bool_3QError_Bool_1,Go)] > (lizzieLet0_4QVal_Bool_3QError_Bool_1QError_Bool,QTree_Bool) */
  assign lizzieLet0_4QVal_Bool_3QError_Bool_1QError_Bool_d = QError_Bool_dc((& {lizzieLet0_4QVal_Bool_3QError_Bool_1_d[0]}), lizzieLet0_4QVal_Bool_3QError_Bool_1_d);
  assign {lizzieLet0_4QVal_Bool_3QError_Bool_1_r} = {1 {(lizzieLet0_4QVal_Bool_3QError_Bool_1QError_Bool_r && lizzieLet0_4QVal_Bool_3QError_Bool_1QError_Bool_d[0])}};
  
  /* buf (Ty QTree_Bool) : (lizzieLet0_4QVal_Bool_3QError_Bool_1QError_Bool,QTree_Bool) > (lizzieLet31_1_argbuf,QTree_Bool) */
  QTree_Bool_t lizzieLet0_4QVal_Bool_3QError_Bool_1QError_Bool_bufchan_d;
  logic lizzieLet0_4QVal_Bool_3QError_Bool_1QError_Bool_bufchan_r;
  assign lizzieLet0_4QVal_Bool_3QError_Bool_1QError_Bool_r = ((! lizzieLet0_4QVal_Bool_3QError_Bool_1QError_Bool_bufchan_d[0]) || lizzieLet0_4QVal_Bool_3QError_Bool_1QError_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_3QError_Bool_1QError_Bool_bufchan_d <= {66'd0,
                                                                    1'd0};
    else
      if (lizzieLet0_4QVal_Bool_3QError_Bool_1QError_Bool_r)
        lizzieLet0_4QVal_Bool_3QError_Bool_1QError_Bool_bufchan_d <= lizzieLet0_4QVal_Bool_3QError_Bool_1QError_Bool_d;
  QTree_Bool_t lizzieLet0_4QVal_Bool_3QError_Bool_1QError_Bool_bufchan_buf;
  assign lizzieLet0_4QVal_Bool_3QError_Bool_1QError_Bool_bufchan_r = (! lizzieLet0_4QVal_Bool_3QError_Bool_1QError_Bool_bufchan_buf[0]);
  assign lizzieLet31_1_argbuf_d = (lizzieLet0_4QVal_Bool_3QError_Bool_1QError_Bool_bufchan_buf[0] ? lizzieLet0_4QVal_Bool_3QError_Bool_1QError_Bool_bufchan_buf :
                                   lizzieLet0_4QVal_Bool_3QError_Bool_1QError_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_3QError_Bool_1QError_Bool_bufchan_buf <= {66'd0,
                                                                      1'd0};
    else
      if ((lizzieLet31_1_argbuf_r && lizzieLet0_4QVal_Bool_3QError_Bool_1QError_Bool_bufchan_buf[0]))
        lizzieLet0_4QVal_Bool_3QError_Bool_1QError_Bool_bufchan_buf <= {66'd0,
                                                                        1'd0};
      else if (((! lizzieLet31_1_argbuf_r) && (! lizzieLet0_4QVal_Bool_3QError_Bool_1QError_Bool_bufchan_buf[0])))
        lizzieLet0_4QVal_Bool_3QError_Bool_1QError_Bool_bufchan_buf <= lizzieLet0_4QVal_Bool_3QError_Bool_1QError_Bool_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet0_4QVal_Bool_3QError_Bool_2,Go) > (lizzieLet0_4QVal_Bool_3QError_Bool_2_argbuf,Go) */
  Go_t lizzieLet0_4QVal_Bool_3QError_Bool_2_bufchan_d;
  logic lizzieLet0_4QVal_Bool_3QError_Bool_2_bufchan_r;
  assign lizzieLet0_4QVal_Bool_3QError_Bool_2_r = ((! lizzieLet0_4QVal_Bool_3QError_Bool_2_bufchan_d[0]) || lizzieLet0_4QVal_Bool_3QError_Bool_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_3QError_Bool_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet0_4QVal_Bool_3QError_Bool_2_r)
        lizzieLet0_4QVal_Bool_3QError_Bool_2_bufchan_d <= lizzieLet0_4QVal_Bool_3QError_Bool_2_d;
  Go_t lizzieLet0_4QVal_Bool_3QError_Bool_2_bufchan_buf;
  assign lizzieLet0_4QVal_Bool_3QError_Bool_2_bufchan_r = (! lizzieLet0_4QVal_Bool_3QError_Bool_2_bufchan_buf[0]);
  assign lizzieLet0_4QVal_Bool_3QError_Bool_2_argbuf_d = (lizzieLet0_4QVal_Bool_3QError_Bool_2_bufchan_buf[0] ? lizzieLet0_4QVal_Bool_3QError_Bool_2_bufchan_buf :
                                                          lizzieLet0_4QVal_Bool_3QError_Bool_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_3QError_Bool_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet0_4QVal_Bool_3QError_Bool_2_argbuf_r && lizzieLet0_4QVal_Bool_3QError_Bool_2_bufchan_buf[0]))
        lizzieLet0_4QVal_Bool_3QError_Bool_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet0_4QVal_Bool_3QError_Bool_2_argbuf_r) && (! lizzieLet0_4QVal_Bool_3QError_Bool_2_bufchan_buf[0])))
        lizzieLet0_4QVal_Bool_3QError_Bool_2_bufchan_buf <= lizzieLet0_4QVal_Bool_3QError_Bool_2_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet0_4QVal_Bool_3QNode_Bool,Go) > [(lizzieLet0_4QVal_Bool_3QNode_Bool_1,Go),
                                                         (lizzieLet0_4QVal_Bool_3QNode_Bool_2,Go)] */
  logic [1:0] lizzieLet0_4QVal_Bool_3QNode_Bool_emitted;
  logic [1:0] lizzieLet0_4QVal_Bool_3QNode_Bool_done;
  assign lizzieLet0_4QVal_Bool_3QNode_Bool_1_d = (lizzieLet0_4QVal_Bool_3QNode_Bool_d[0] && (! lizzieLet0_4QVal_Bool_3QNode_Bool_emitted[0]));
  assign lizzieLet0_4QVal_Bool_3QNode_Bool_2_d = (lizzieLet0_4QVal_Bool_3QNode_Bool_d[0] && (! lizzieLet0_4QVal_Bool_3QNode_Bool_emitted[1]));
  assign lizzieLet0_4QVal_Bool_3QNode_Bool_done = (lizzieLet0_4QVal_Bool_3QNode_Bool_emitted | ({lizzieLet0_4QVal_Bool_3QNode_Bool_2_d[0],
                                                                                                 lizzieLet0_4QVal_Bool_3QNode_Bool_1_d[0]} & {lizzieLet0_4QVal_Bool_3QNode_Bool_2_r,
                                                                                                                                              lizzieLet0_4QVal_Bool_3QNode_Bool_1_r}));
  assign lizzieLet0_4QVal_Bool_3QNode_Bool_r = (& lizzieLet0_4QVal_Bool_3QNode_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_3QNode_Bool_emitted <= 2'd0;
    else
      lizzieLet0_4QVal_Bool_3QNode_Bool_emitted <= (lizzieLet0_4QVal_Bool_3QNode_Bool_r ? 2'd0 :
                                                    lizzieLet0_4QVal_Bool_3QNode_Bool_done);
  
  /* dcon (Ty QTree_Bool,
      Dcon QError_Bool) : [(lizzieLet0_4QVal_Bool_3QNode_Bool_1,Go)] > (lizzieLet0_4QVal_Bool_3QNode_Bool_1QError_Bool,QTree_Bool) */
  assign lizzieLet0_4QVal_Bool_3QNode_Bool_1QError_Bool_d = QError_Bool_dc((& {lizzieLet0_4QVal_Bool_3QNode_Bool_1_d[0]}), lizzieLet0_4QVal_Bool_3QNode_Bool_1_d);
  assign {lizzieLet0_4QVal_Bool_3QNode_Bool_1_r} = {1 {(lizzieLet0_4QVal_Bool_3QNode_Bool_1QError_Bool_r && lizzieLet0_4QVal_Bool_3QNode_Bool_1QError_Bool_d[0])}};
  
  /* buf (Ty QTree_Bool) : (lizzieLet0_4QVal_Bool_3QNode_Bool_1QError_Bool,QTree_Bool) > (lizzieLet30_1_argbuf,QTree_Bool) */
  QTree_Bool_t lizzieLet0_4QVal_Bool_3QNode_Bool_1QError_Bool_bufchan_d;
  logic lizzieLet0_4QVal_Bool_3QNode_Bool_1QError_Bool_bufchan_r;
  assign lizzieLet0_4QVal_Bool_3QNode_Bool_1QError_Bool_r = ((! lizzieLet0_4QVal_Bool_3QNode_Bool_1QError_Bool_bufchan_d[0]) || lizzieLet0_4QVal_Bool_3QNode_Bool_1QError_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_3QNode_Bool_1QError_Bool_bufchan_d <= {66'd0,
                                                                   1'd0};
    else
      if (lizzieLet0_4QVal_Bool_3QNode_Bool_1QError_Bool_r)
        lizzieLet0_4QVal_Bool_3QNode_Bool_1QError_Bool_bufchan_d <= lizzieLet0_4QVal_Bool_3QNode_Bool_1QError_Bool_d;
  QTree_Bool_t lizzieLet0_4QVal_Bool_3QNode_Bool_1QError_Bool_bufchan_buf;
  assign lizzieLet0_4QVal_Bool_3QNode_Bool_1QError_Bool_bufchan_r = (! lizzieLet0_4QVal_Bool_3QNode_Bool_1QError_Bool_bufchan_buf[0]);
  assign lizzieLet30_1_argbuf_d = (lizzieLet0_4QVal_Bool_3QNode_Bool_1QError_Bool_bufchan_buf[0] ? lizzieLet0_4QVal_Bool_3QNode_Bool_1QError_Bool_bufchan_buf :
                                   lizzieLet0_4QVal_Bool_3QNode_Bool_1QError_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_3QNode_Bool_1QError_Bool_bufchan_buf <= {66'd0,
                                                                     1'd0};
    else
      if ((lizzieLet30_1_argbuf_r && lizzieLet0_4QVal_Bool_3QNode_Bool_1QError_Bool_bufchan_buf[0]))
        lizzieLet0_4QVal_Bool_3QNode_Bool_1QError_Bool_bufchan_buf <= {66'd0,
                                                                       1'd0};
      else if (((! lizzieLet30_1_argbuf_r) && (! lizzieLet0_4QVal_Bool_3QNode_Bool_1QError_Bool_bufchan_buf[0])))
        lizzieLet0_4QVal_Bool_3QNode_Bool_1QError_Bool_bufchan_buf <= lizzieLet0_4QVal_Bool_3QNode_Bool_1QError_Bool_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet0_4QVal_Bool_3QNode_Bool_2,Go) > (lizzieLet0_4QVal_Bool_3QNode_Bool_2_argbuf,Go) */
  Go_t lizzieLet0_4QVal_Bool_3QNode_Bool_2_bufchan_d;
  logic lizzieLet0_4QVal_Bool_3QNode_Bool_2_bufchan_r;
  assign lizzieLet0_4QVal_Bool_3QNode_Bool_2_r = ((! lizzieLet0_4QVal_Bool_3QNode_Bool_2_bufchan_d[0]) || lizzieLet0_4QVal_Bool_3QNode_Bool_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_3QNode_Bool_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet0_4QVal_Bool_3QNode_Bool_2_r)
        lizzieLet0_4QVal_Bool_3QNode_Bool_2_bufchan_d <= lizzieLet0_4QVal_Bool_3QNode_Bool_2_d;
  Go_t lizzieLet0_4QVal_Bool_3QNode_Bool_2_bufchan_buf;
  assign lizzieLet0_4QVal_Bool_3QNode_Bool_2_bufchan_r = (! lizzieLet0_4QVal_Bool_3QNode_Bool_2_bufchan_buf[0]);
  assign lizzieLet0_4QVal_Bool_3QNode_Bool_2_argbuf_d = (lizzieLet0_4QVal_Bool_3QNode_Bool_2_bufchan_buf[0] ? lizzieLet0_4QVal_Bool_3QNode_Bool_2_bufchan_buf :
                                                         lizzieLet0_4QVal_Bool_3QNode_Bool_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_3QNode_Bool_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet0_4QVal_Bool_3QNode_Bool_2_argbuf_r && lizzieLet0_4QVal_Bool_3QNode_Bool_2_bufchan_buf[0]))
        lizzieLet0_4QVal_Bool_3QNode_Bool_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet0_4QVal_Bool_3QNode_Bool_2_argbuf_r) && (! lizzieLet0_4QVal_Bool_3QNode_Bool_2_bufchan_buf[0])))
        lizzieLet0_4QVal_Bool_3QNode_Bool_2_bufchan_buf <= lizzieLet0_4QVal_Bool_3QNode_Bool_2_bufchan_d;
  
  /* demux (Ty QTree_Bool,
       Ty QTree_Bool) : (lizzieLet0_4QVal_Bool_4,QTree_Bool) (lizzieLet0_5QVal_Bool,QTree_Bool) > [(lizzieLet0_4QVal_Bool_4QNone_Bool,QTree_Bool),
                                                                                                   (lizzieLet0_4QVal_Bool_4QVal_Bool,QTree_Bool),
                                                                                                   (_72,QTree_Bool),
                                                                                                   (_71,QTree_Bool)] */
  logic [3:0] lizzieLet0_5QVal_Bool_onehotd;
  always_comb
    if ((lizzieLet0_4QVal_Bool_4_d[0] && lizzieLet0_5QVal_Bool_d[0]))
      unique case (lizzieLet0_4QVal_Bool_4_d[2:1])
        2'd0: lizzieLet0_5QVal_Bool_onehotd = 4'd1;
        2'd1: lizzieLet0_5QVal_Bool_onehotd = 4'd2;
        2'd2: lizzieLet0_5QVal_Bool_onehotd = 4'd4;
        2'd3: lizzieLet0_5QVal_Bool_onehotd = 4'd8;
        default: lizzieLet0_5QVal_Bool_onehotd = 4'd0;
      endcase
    else lizzieLet0_5QVal_Bool_onehotd = 4'd0;
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_d = {lizzieLet0_5QVal_Bool_d[66:1],
                                                lizzieLet0_5QVal_Bool_onehotd[0]};
  assign lizzieLet0_4QVal_Bool_4QVal_Bool_d = {lizzieLet0_5QVal_Bool_d[66:1],
                                               lizzieLet0_5QVal_Bool_onehotd[1]};
  assign _72_d = {lizzieLet0_5QVal_Bool_d[66:1],
                  lizzieLet0_5QVal_Bool_onehotd[2]};
  assign _71_d = {lizzieLet0_5QVal_Bool_d[66:1],
                  lizzieLet0_5QVal_Bool_onehotd[3]};
  assign lizzieLet0_5QVal_Bool_r = (| (lizzieLet0_5QVal_Bool_onehotd & {_71_r,
                                                                        _72_r,
                                                                        lizzieLet0_4QVal_Bool_4QVal_Bool_r,
                                                                        lizzieLet0_4QVal_Bool_4QNone_Bool_r}));
  assign lizzieLet0_4QVal_Bool_4_r = lizzieLet0_5QVal_Bool_r;
  
  /* fork (Ty QTree_Bool) : (lizzieLet0_4QVal_Bool_4QNone_Bool,QTree_Bool) > [(lizzieLet0_4QVal_Bool_4QNone_Bool_1,QTree_Bool),
                                                                         (lizzieLet0_4QVal_Bool_4QNone_Bool_2,QTree_Bool),
                                                                         (lizzieLet0_4QVal_Bool_4QNone_Bool_3,QTree_Bool),
                                                                         (lizzieLet0_4QVal_Bool_4QNone_Bool_4,QTree_Bool),
                                                                         (lizzieLet0_4QVal_Bool_4QNone_Bool_5,QTree_Bool),
                                                                         (lizzieLet0_4QVal_Bool_4QNone_Bool_6,QTree_Bool)] */
  logic [5:0] lizzieLet0_4QVal_Bool_4QNone_Bool_emitted;
  logic [5:0] lizzieLet0_4QVal_Bool_4QNone_Bool_done;
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_1_d = {lizzieLet0_4QVal_Bool_4QNone_Bool_d[66:1],
                                                  (lizzieLet0_4QVal_Bool_4QNone_Bool_d[0] && (! lizzieLet0_4QVal_Bool_4QNone_Bool_emitted[0]))};
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_2_d = {lizzieLet0_4QVal_Bool_4QNone_Bool_d[66:1],
                                                  (lizzieLet0_4QVal_Bool_4QNone_Bool_d[0] && (! lizzieLet0_4QVal_Bool_4QNone_Bool_emitted[1]))};
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_3_d = {lizzieLet0_4QVal_Bool_4QNone_Bool_d[66:1],
                                                  (lizzieLet0_4QVal_Bool_4QNone_Bool_d[0] && (! lizzieLet0_4QVal_Bool_4QNone_Bool_emitted[2]))};
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_4_d = {lizzieLet0_4QVal_Bool_4QNone_Bool_d[66:1],
                                                  (lizzieLet0_4QVal_Bool_4QNone_Bool_d[0] && (! lizzieLet0_4QVal_Bool_4QNone_Bool_emitted[3]))};
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_5_d = {lizzieLet0_4QVal_Bool_4QNone_Bool_d[66:1],
                                                  (lizzieLet0_4QVal_Bool_4QNone_Bool_d[0] && (! lizzieLet0_4QVal_Bool_4QNone_Bool_emitted[4]))};
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_6_d = {lizzieLet0_4QVal_Bool_4QNone_Bool_d[66:1],
                                                  (lizzieLet0_4QVal_Bool_4QNone_Bool_d[0] && (! lizzieLet0_4QVal_Bool_4QNone_Bool_emitted[5]))};
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_done = (lizzieLet0_4QVal_Bool_4QNone_Bool_emitted | ({lizzieLet0_4QVal_Bool_4QNone_Bool_6_d[0],
                                                                                                 lizzieLet0_4QVal_Bool_4QNone_Bool_5_d[0],
                                                                                                 lizzieLet0_4QVal_Bool_4QNone_Bool_4_d[0],
                                                                                                 lizzieLet0_4QVal_Bool_4QNone_Bool_3_d[0],
                                                                                                 lizzieLet0_4QVal_Bool_4QNone_Bool_2_d[0],
                                                                                                 lizzieLet0_4QVal_Bool_4QNone_Bool_1_d[0]} & {lizzieLet0_4QVal_Bool_4QNone_Bool_6_r,
                                                                                                                                              lizzieLet0_4QVal_Bool_4QNone_Bool_5_r,
                                                                                                                                              lizzieLet0_4QVal_Bool_4QNone_Bool_4_r,
                                                                                                                                              lizzieLet0_4QVal_Bool_4QNone_Bool_3_r,
                                                                                                                                              lizzieLet0_4QVal_Bool_4QNone_Bool_2_r,
                                                                                                                                              lizzieLet0_4QVal_Bool_4QNone_Bool_1_r}));
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_r = (& lizzieLet0_4QVal_Bool_4QNone_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_4QNone_Bool_emitted <= 6'd0;
    else
      lizzieLet0_4QVal_Bool_4QNone_Bool_emitted <= (lizzieLet0_4QVal_Bool_4QNone_Bool_r ? 6'd0 :
                                                    lizzieLet0_4QVal_Bool_4QNone_Bool_done);
  
  /* destruct (Ty QTree_Bool,
          Dcon QVal_Bool) : (lizzieLet0_4QVal_Bool_4QNone_Bool_1QVal_Bool,QTree_Bool) > [(va8n_destruct,MyBool)] */
  assign va8n_destruct_d = {lizzieLet0_4QVal_Bool_4QNone_Bool_1QVal_Bool_d[3:3],
                            lizzieLet0_4QVal_Bool_4QNone_Bool_1QVal_Bool_d[0]};
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_1QVal_Bool_r = va8n_destruct_r;
  
  /* demux (Ty QTree_Bool,
       Ty QTree_Bool) : (lizzieLet0_4QVal_Bool_4QNone_Bool_2,QTree_Bool) (lizzieLet0_4QVal_Bool_4QNone_Bool_1,QTree_Bool) > [(_70,QTree_Bool),
                                                                                                                             (lizzieLet0_4QVal_Bool_4QNone_Bool_1QVal_Bool,QTree_Bool),
                                                                                                                             (_69,QTree_Bool),
                                                                                                                             (_68,QTree_Bool)] */
  logic [3:0] lizzieLet0_4QVal_Bool_4QNone_Bool_1_onehotd;
  always_comb
    if ((lizzieLet0_4QVal_Bool_4QNone_Bool_2_d[0] && lizzieLet0_4QVal_Bool_4QNone_Bool_1_d[0]))
      unique case (lizzieLet0_4QVal_Bool_4QNone_Bool_2_d[2:1])
        2'd0: lizzieLet0_4QVal_Bool_4QNone_Bool_1_onehotd = 4'd1;
        2'd1: lizzieLet0_4QVal_Bool_4QNone_Bool_1_onehotd = 4'd2;
        2'd2: lizzieLet0_4QVal_Bool_4QNone_Bool_1_onehotd = 4'd4;
        2'd3: lizzieLet0_4QVal_Bool_4QNone_Bool_1_onehotd = 4'd8;
        default: lizzieLet0_4QVal_Bool_4QNone_Bool_1_onehotd = 4'd0;
      endcase
    else lizzieLet0_4QVal_Bool_4QNone_Bool_1_onehotd = 4'd0;
  assign _70_d = {lizzieLet0_4QVal_Bool_4QNone_Bool_1_d[66:1],
                  lizzieLet0_4QVal_Bool_4QNone_Bool_1_onehotd[0]};
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_1QVal_Bool_d = {lizzieLet0_4QVal_Bool_4QNone_Bool_1_d[66:1],
                                                           lizzieLet0_4QVal_Bool_4QNone_Bool_1_onehotd[1]};
  assign _69_d = {lizzieLet0_4QVal_Bool_4QNone_Bool_1_d[66:1],
                  lizzieLet0_4QVal_Bool_4QNone_Bool_1_onehotd[2]};
  assign _68_d = {lizzieLet0_4QVal_Bool_4QNone_Bool_1_d[66:1],
                  lizzieLet0_4QVal_Bool_4QNone_Bool_1_onehotd[3]};
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_1_r = (| (lizzieLet0_4QVal_Bool_4QNone_Bool_1_onehotd & {_68_r,
                                                                                                    _69_r,
                                                                                                    lizzieLet0_4QVal_Bool_4QNone_Bool_1QVal_Bool_r,
                                                                                                    _70_r}));
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_2_r = lizzieLet0_4QVal_Bool_4QNone_Bool_1_r;
  
  /* demux (Ty QTree_Bool,
       Ty Go) : (lizzieLet0_4QVal_Bool_4QNone_Bool_3,QTree_Bool) (lizzieLet0_4QVal_Bool_3QNone_Bool,Go) > [(lizzieLet0_4QVal_Bool_4QNone_Bool_3QNone_Bool,Go),
                                                                                                           (lizzieLet0_4QVal_Bool_4QNone_Bool_3QVal_Bool,Go),
                                                                                                           (lizzieLet0_4QVal_Bool_4QNone_Bool_3QNode_Bool,Go),
                                                                                                           (lizzieLet0_4QVal_Bool_4QNone_Bool_3QError_Bool,Go)] */
  logic [3:0] lizzieLet0_4QVal_Bool_3QNone_Bool_onehotd;
  always_comb
    if ((lizzieLet0_4QVal_Bool_4QNone_Bool_3_d[0] && lizzieLet0_4QVal_Bool_3QNone_Bool_d[0]))
      unique case (lizzieLet0_4QVal_Bool_4QNone_Bool_3_d[2:1])
        2'd0: lizzieLet0_4QVal_Bool_3QNone_Bool_onehotd = 4'd1;
        2'd1: lizzieLet0_4QVal_Bool_3QNone_Bool_onehotd = 4'd2;
        2'd2: lizzieLet0_4QVal_Bool_3QNone_Bool_onehotd = 4'd4;
        2'd3: lizzieLet0_4QVal_Bool_3QNone_Bool_onehotd = 4'd8;
        default: lizzieLet0_4QVal_Bool_3QNone_Bool_onehotd = 4'd0;
      endcase
    else lizzieLet0_4QVal_Bool_3QNone_Bool_onehotd = 4'd0;
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_3QNone_Bool_d = lizzieLet0_4QVal_Bool_3QNone_Bool_onehotd[0];
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_3QVal_Bool_d = lizzieLet0_4QVal_Bool_3QNone_Bool_onehotd[1];
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_3QNode_Bool_d = lizzieLet0_4QVal_Bool_3QNone_Bool_onehotd[2];
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_3QError_Bool_d = lizzieLet0_4QVal_Bool_3QNone_Bool_onehotd[3];
  assign lizzieLet0_4QVal_Bool_3QNone_Bool_r = (| (lizzieLet0_4QVal_Bool_3QNone_Bool_onehotd & {lizzieLet0_4QVal_Bool_4QNone_Bool_3QError_Bool_r,
                                                                                                lizzieLet0_4QVal_Bool_4QNone_Bool_3QNode_Bool_r,
                                                                                                lizzieLet0_4QVal_Bool_4QNone_Bool_3QVal_Bool_r,
                                                                                                lizzieLet0_4QVal_Bool_4QNone_Bool_3QNone_Bool_r}));
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_3_r = lizzieLet0_4QVal_Bool_3QNone_Bool_r;
  
  /* fork (Ty Go) : (lizzieLet0_4QVal_Bool_4QNone_Bool_3QError_Bool,Go) > [(lizzieLet0_4QVal_Bool_4QNone_Bool_3QError_Bool_1,Go),
                                                                      (lizzieLet0_4QVal_Bool_4QNone_Bool_3QError_Bool_2,Go)] */
  logic [1:0] lizzieLet0_4QVal_Bool_4QNone_Bool_3QError_Bool_emitted;
  logic [1:0] lizzieLet0_4QVal_Bool_4QNone_Bool_3QError_Bool_done;
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_3QError_Bool_1_d = (lizzieLet0_4QVal_Bool_4QNone_Bool_3QError_Bool_d[0] && (! lizzieLet0_4QVal_Bool_4QNone_Bool_3QError_Bool_emitted[0]));
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_3QError_Bool_2_d = (lizzieLet0_4QVal_Bool_4QNone_Bool_3QError_Bool_d[0] && (! lizzieLet0_4QVal_Bool_4QNone_Bool_3QError_Bool_emitted[1]));
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_3QError_Bool_done = (lizzieLet0_4QVal_Bool_4QNone_Bool_3QError_Bool_emitted | ({lizzieLet0_4QVal_Bool_4QNone_Bool_3QError_Bool_2_d[0],
                                                                                                                           lizzieLet0_4QVal_Bool_4QNone_Bool_3QError_Bool_1_d[0]} & {lizzieLet0_4QVal_Bool_4QNone_Bool_3QError_Bool_2_r,
                                                                                                                                                                                     lizzieLet0_4QVal_Bool_4QNone_Bool_3QError_Bool_1_r}));
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_3QError_Bool_r = (& lizzieLet0_4QVal_Bool_4QNone_Bool_3QError_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_4QNone_Bool_3QError_Bool_emitted <= 2'd0;
    else
      lizzieLet0_4QVal_Bool_4QNone_Bool_3QError_Bool_emitted <= (lizzieLet0_4QVal_Bool_4QNone_Bool_3QError_Bool_r ? 2'd0 :
                                                                 lizzieLet0_4QVal_Bool_4QNone_Bool_3QError_Bool_done);
  
  /* dcon (Ty QTree_Bool,
      Dcon QError_Bool) : [(lizzieLet0_4QVal_Bool_4QNone_Bool_3QError_Bool_1,Go)] > (lizzieLet0_4QVal_Bool_4QNone_Bool_3QError_Bool_1QError_Bool,QTree_Bool) */
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_3QError_Bool_1QError_Bool_d = QError_Bool_dc((& {lizzieLet0_4QVal_Bool_4QNone_Bool_3QError_Bool_1_d[0]}), lizzieLet0_4QVal_Bool_4QNone_Bool_3QError_Bool_1_d);
  assign {lizzieLet0_4QVal_Bool_4QNone_Bool_3QError_Bool_1_r} = {1 {(lizzieLet0_4QVal_Bool_4QNone_Bool_3QError_Bool_1QError_Bool_r && lizzieLet0_4QVal_Bool_4QNone_Bool_3QError_Bool_1QError_Bool_d[0])}};
  
  /* buf (Ty QTree_Bool) : (lizzieLet0_4QVal_Bool_4QNone_Bool_3QError_Bool_1QError_Bool,QTree_Bool) > (lizzieLet19_1_argbuf,QTree_Bool) */
  QTree_Bool_t lizzieLet0_4QVal_Bool_4QNone_Bool_3QError_Bool_1QError_Bool_bufchan_d;
  logic lizzieLet0_4QVal_Bool_4QNone_Bool_3QError_Bool_1QError_Bool_bufchan_r;
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_3QError_Bool_1QError_Bool_r = ((! lizzieLet0_4QVal_Bool_4QNone_Bool_3QError_Bool_1QError_Bool_bufchan_d[0]) || lizzieLet0_4QVal_Bool_4QNone_Bool_3QError_Bool_1QError_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_4QNone_Bool_3QError_Bool_1QError_Bool_bufchan_d <= {66'd0,
                                                                                1'd0};
    else
      if (lizzieLet0_4QVal_Bool_4QNone_Bool_3QError_Bool_1QError_Bool_r)
        lizzieLet0_4QVal_Bool_4QNone_Bool_3QError_Bool_1QError_Bool_bufchan_d <= lizzieLet0_4QVal_Bool_4QNone_Bool_3QError_Bool_1QError_Bool_d;
  QTree_Bool_t lizzieLet0_4QVal_Bool_4QNone_Bool_3QError_Bool_1QError_Bool_bufchan_buf;
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_3QError_Bool_1QError_Bool_bufchan_r = (! lizzieLet0_4QVal_Bool_4QNone_Bool_3QError_Bool_1QError_Bool_bufchan_buf[0]);
  assign lizzieLet19_1_argbuf_d = (lizzieLet0_4QVal_Bool_4QNone_Bool_3QError_Bool_1QError_Bool_bufchan_buf[0] ? lizzieLet0_4QVal_Bool_4QNone_Bool_3QError_Bool_1QError_Bool_bufchan_buf :
                                   lizzieLet0_4QVal_Bool_4QNone_Bool_3QError_Bool_1QError_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_4QNone_Bool_3QError_Bool_1QError_Bool_bufchan_buf <= {66'd0,
                                                                                  1'd0};
    else
      if ((lizzieLet19_1_argbuf_r && lizzieLet0_4QVal_Bool_4QNone_Bool_3QError_Bool_1QError_Bool_bufchan_buf[0]))
        lizzieLet0_4QVal_Bool_4QNone_Bool_3QError_Bool_1QError_Bool_bufchan_buf <= {66'd0,
                                                                                    1'd0};
      else if (((! lizzieLet19_1_argbuf_r) && (! lizzieLet0_4QVal_Bool_4QNone_Bool_3QError_Bool_1QError_Bool_bufchan_buf[0])))
        lizzieLet0_4QVal_Bool_4QNone_Bool_3QError_Bool_1QError_Bool_bufchan_buf <= lizzieLet0_4QVal_Bool_4QNone_Bool_3QError_Bool_1QError_Bool_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet0_4QVal_Bool_4QNone_Bool_3QError_Bool_2,Go) > (lizzieLet0_4QVal_Bool_4QNone_Bool_3QError_Bool_2_argbuf,Go) */
  Go_t lizzieLet0_4QVal_Bool_4QNone_Bool_3QError_Bool_2_bufchan_d;
  logic lizzieLet0_4QVal_Bool_4QNone_Bool_3QError_Bool_2_bufchan_r;
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_3QError_Bool_2_r = ((! lizzieLet0_4QVal_Bool_4QNone_Bool_3QError_Bool_2_bufchan_d[0]) || lizzieLet0_4QVal_Bool_4QNone_Bool_3QError_Bool_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_4QNone_Bool_3QError_Bool_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet0_4QVal_Bool_4QNone_Bool_3QError_Bool_2_r)
        lizzieLet0_4QVal_Bool_4QNone_Bool_3QError_Bool_2_bufchan_d <= lizzieLet0_4QVal_Bool_4QNone_Bool_3QError_Bool_2_d;
  Go_t lizzieLet0_4QVal_Bool_4QNone_Bool_3QError_Bool_2_bufchan_buf;
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_3QError_Bool_2_bufchan_r = (! lizzieLet0_4QVal_Bool_4QNone_Bool_3QError_Bool_2_bufchan_buf[0]);
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_3QError_Bool_2_argbuf_d = (lizzieLet0_4QVal_Bool_4QNone_Bool_3QError_Bool_2_bufchan_buf[0] ? lizzieLet0_4QVal_Bool_4QNone_Bool_3QError_Bool_2_bufchan_buf :
                                                                      lizzieLet0_4QVal_Bool_4QNone_Bool_3QError_Bool_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_4QNone_Bool_3QError_Bool_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet0_4QVal_Bool_4QNone_Bool_3QError_Bool_2_argbuf_r && lizzieLet0_4QVal_Bool_4QNone_Bool_3QError_Bool_2_bufchan_buf[0]))
        lizzieLet0_4QVal_Bool_4QNone_Bool_3QError_Bool_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet0_4QVal_Bool_4QNone_Bool_3QError_Bool_2_argbuf_r) && (! lizzieLet0_4QVal_Bool_4QNone_Bool_3QError_Bool_2_bufchan_buf[0])))
        lizzieLet0_4QVal_Bool_4QNone_Bool_3QError_Bool_2_bufchan_buf <= lizzieLet0_4QVal_Bool_4QNone_Bool_3QError_Bool_2_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet0_4QVal_Bool_4QNone_Bool_3QNode_Bool,Go) > [(lizzieLet0_4QVal_Bool_4QNone_Bool_3QNode_Bool_1,Go),
                                                                     (lizzieLet0_4QVal_Bool_4QNone_Bool_3QNode_Bool_2,Go)] */
  logic [1:0] lizzieLet0_4QVal_Bool_4QNone_Bool_3QNode_Bool_emitted;
  logic [1:0] lizzieLet0_4QVal_Bool_4QNone_Bool_3QNode_Bool_done;
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_3QNode_Bool_1_d = (lizzieLet0_4QVal_Bool_4QNone_Bool_3QNode_Bool_d[0] && (! lizzieLet0_4QVal_Bool_4QNone_Bool_3QNode_Bool_emitted[0]));
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_3QNode_Bool_2_d = (lizzieLet0_4QVal_Bool_4QNone_Bool_3QNode_Bool_d[0] && (! lizzieLet0_4QVal_Bool_4QNone_Bool_3QNode_Bool_emitted[1]));
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_3QNode_Bool_done = (lizzieLet0_4QVal_Bool_4QNone_Bool_3QNode_Bool_emitted | ({lizzieLet0_4QVal_Bool_4QNone_Bool_3QNode_Bool_2_d[0],
                                                                                                                         lizzieLet0_4QVal_Bool_4QNone_Bool_3QNode_Bool_1_d[0]} & {lizzieLet0_4QVal_Bool_4QNone_Bool_3QNode_Bool_2_r,
                                                                                                                                                                                  lizzieLet0_4QVal_Bool_4QNone_Bool_3QNode_Bool_1_r}));
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_3QNode_Bool_r = (& lizzieLet0_4QVal_Bool_4QNone_Bool_3QNode_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_4QNone_Bool_3QNode_Bool_emitted <= 2'd0;
    else
      lizzieLet0_4QVal_Bool_4QNone_Bool_3QNode_Bool_emitted <= (lizzieLet0_4QVal_Bool_4QNone_Bool_3QNode_Bool_r ? 2'd0 :
                                                                lizzieLet0_4QVal_Bool_4QNone_Bool_3QNode_Bool_done);
  
  /* dcon (Ty QTree_Bool,
      Dcon QError_Bool) : [(lizzieLet0_4QVal_Bool_4QNone_Bool_3QNode_Bool_1,Go)] > (lizzieLet0_4QVal_Bool_4QNone_Bool_3QNode_Bool_1QError_Bool,QTree_Bool) */
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_3QNode_Bool_1QError_Bool_d = QError_Bool_dc((& {lizzieLet0_4QVal_Bool_4QNone_Bool_3QNode_Bool_1_d[0]}), lizzieLet0_4QVal_Bool_4QNone_Bool_3QNode_Bool_1_d);
  assign {lizzieLet0_4QVal_Bool_4QNone_Bool_3QNode_Bool_1_r} = {1 {(lizzieLet0_4QVal_Bool_4QNone_Bool_3QNode_Bool_1QError_Bool_r && lizzieLet0_4QVal_Bool_4QNone_Bool_3QNode_Bool_1QError_Bool_d[0])}};
  
  /* buf (Ty QTree_Bool) : (lizzieLet0_4QVal_Bool_4QNone_Bool_3QNode_Bool_1QError_Bool,QTree_Bool) > (lizzieLet18_1_argbuf,QTree_Bool) */
  QTree_Bool_t lizzieLet0_4QVal_Bool_4QNone_Bool_3QNode_Bool_1QError_Bool_bufchan_d;
  logic lizzieLet0_4QVal_Bool_4QNone_Bool_3QNode_Bool_1QError_Bool_bufchan_r;
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_3QNode_Bool_1QError_Bool_r = ((! lizzieLet0_4QVal_Bool_4QNone_Bool_3QNode_Bool_1QError_Bool_bufchan_d[0]) || lizzieLet0_4QVal_Bool_4QNone_Bool_3QNode_Bool_1QError_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_4QNone_Bool_3QNode_Bool_1QError_Bool_bufchan_d <= {66'd0,
                                                                               1'd0};
    else
      if (lizzieLet0_4QVal_Bool_4QNone_Bool_3QNode_Bool_1QError_Bool_r)
        lizzieLet0_4QVal_Bool_4QNone_Bool_3QNode_Bool_1QError_Bool_bufchan_d <= lizzieLet0_4QVal_Bool_4QNone_Bool_3QNode_Bool_1QError_Bool_d;
  QTree_Bool_t lizzieLet0_4QVal_Bool_4QNone_Bool_3QNode_Bool_1QError_Bool_bufchan_buf;
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_3QNode_Bool_1QError_Bool_bufchan_r = (! lizzieLet0_4QVal_Bool_4QNone_Bool_3QNode_Bool_1QError_Bool_bufchan_buf[0]);
  assign lizzieLet18_1_argbuf_d = (lizzieLet0_4QVal_Bool_4QNone_Bool_3QNode_Bool_1QError_Bool_bufchan_buf[0] ? lizzieLet0_4QVal_Bool_4QNone_Bool_3QNode_Bool_1QError_Bool_bufchan_buf :
                                   lizzieLet0_4QVal_Bool_4QNone_Bool_3QNode_Bool_1QError_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_4QNone_Bool_3QNode_Bool_1QError_Bool_bufchan_buf <= {66'd0,
                                                                                 1'd0};
    else
      if ((lizzieLet18_1_argbuf_r && lizzieLet0_4QVal_Bool_4QNone_Bool_3QNode_Bool_1QError_Bool_bufchan_buf[0]))
        lizzieLet0_4QVal_Bool_4QNone_Bool_3QNode_Bool_1QError_Bool_bufchan_buf <= {66'd0,
                                                                                   1'd0};
      else if (((! lizzieLet18_1_argbuf_r) && (! lizzieLet0_4QVal_Bool_4QNone_Bool_3QNode_Bool_1QError_Bool_bufchan_buf[0])))
        lizzieLet0_4QVal_Bool_4QNone_Bool_3QNode_Bool_1QError_Bool_bufchan_buf <= lizzieLet0_4QVal_Bool_4QNone_Bool_3QNode_Bool_1QError_Bool_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet0_4QVal_Bool_4QNone_Bool_3QNode_Bool_2,Go) > (lizzieLet0_4QVal_Bool_4QNone_Bool_3QNode_Bool_2_argbuf,Go) */
  Go_t lizzieLet0_4QVal_Bool_4QNone_Bool_3QNode_Bool_2_bufchan_d;
  logic lizzieLet0_4QVal_Bool_4QNone_Bool_3QNode_Bool_2_bufchan_r;
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_3QNode_Bool_2_r = ((! lizzieLet0_4QVal_Bool_4QNone_Bool_3QNode_Bool_2_bufchan_d[0]) || lizzieLet0_4QVal_Bool_4QNone_Bool_3QNode_Bool_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_4QNone_Bool_3QNode_Bool_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet0_4QVal_Bool_4QNone_Bool_3QNode_Bool_2_r)
        lizzieLet0_4QVal_Bool_4QNone_Bool_3QNode_Bool_2_bufchan_d <= lizzieLet0_4QVal_Bool_4QNone_Bool_3QNode_Bool_2_d;
  Go_t lizzieLet0_4QVal_Bool_4QNone_Bool_3QNode_Bool_2_bufchan_buf;
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_3QNode_Bool_2_bufchan_r = (! lizzieLet0_4QVal_Bool_4QNone_Bool_3QNode_Bool_2_bufchan_buf[0]);
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_3QNode_Bool_2_argbuf_d = (lizzieLet0_4QVal_Bool_4QNone_Bool_3QNode_Bool_2_bufchan_buf[0] ? lizzieLet0_4QVal_Bool_4QNone_Bool_3QNode_Bool_2_bufchan_buf :
                                                                     lizzieLet0_4QVal_Bool_4QNone_Bool_3QNode_Bool_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_4QNone_Bool_3QNode_Bool_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet0_4QVal_Bool_4QNone_Bool_3QNode_Bool_2_argbuf_r && lizzieLet0_4QVal_Bool_4QNone_Bool_3QNode_Bool_2_bufchan_buf[0]))
        lizzieLet0_4QVal_Bool_4QNone_Bool_3QNode_Bool_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet0_4QVal_Bool_4QNone_Bool_3QNode_Bool_2_argbuf_r) && (! lizzieLet0_4QVal_Bool_4QNone_Bool_3QNode_Bool_2_bufchan_buf[0])))
        lizzieLet0_4QVal_Bool_4QNone_Bool_3QNode_Bool_2_bufchan_buf <= lizzieLet0_4QVal_Bool_4QNone_Bool_3QNode_Bool_2_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet0_4QVal_Bool_4QNone_Bool_3QNone_Bool,Go) > (lizzieLet0_4QVal_Bool_4QNone_Bool_3QNone_Bool_1_argbuf,Go) */
  Go_t lizzieLet0_4QVal_Bool_4QNone_Bool_3QNone_Bool_bufchan_d;
  logic lizzieLet0_4QVal_Bool_4QNone_Bool_3QNone_Bool_bufchan_r;
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_3QNone_Bool_r = ((! lizzieLet0_4QVal_Bool_4QNone_Bool_3QNone_Bool_bufchan_d[0]) || lizzieLet0_4QVal_Bool_4QNone_Bool_3QNone_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_4QNone_Bool_3QNone_Bool_bufchan_d <= 1'd0;
    else
      if (lizzieLet0_4QVal_Bool_4QNone_Bool_3QNone_Bool_r)
        lizzieLet0_4QVal_Bool_4QNone_Bool_3QNone_Bool_bufchan_d <= lizzieLet0_4QVal_Bool_4QNone_Bool_3QNone_Bool_d;
  Go_t lizzieLet0_4QVal_Bool_4QNone_Bool_3QNone_Bool_bufchan_buf;
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_3QNone_Bool_bufchan_r = (! lizzieLet0_4QVal_Bool_4QNone_Bool_3QNone_Bool_bufchan_buf[0]);
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_3QNone_Bool_1_argbuf_d = (lizzieLet0_4QVal_Bool_4QNone_Bool_3QNone_Bool_bufchan_buf[0] ? lizzieLet0_4QVal_Bool_4QNone_Bool_3QNone_Bool_bufchan_buf :
                                                                     lizzieLet0_4QVal_Bool_4QNone_Bool_3QNone_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_4QNone_Bool_3QNone_Bool_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet0_4QVal_Bool_4QNone_Bool_3QNone_Bool_1_argbuf_r && lizzieLet0_4QVal_Bool_4QNone_Bool_3QNone_Bool_bufchan_buf[0]))
        lizzieLet0_4QVal_Bool_4QNone_Bool_3QNone_Bool_bufchan_buf <= 1'd0;
      else if (((! lizzieLet0_4QVal_Bool_4QNone_Bool_3QNone_Bool_1_argbuf_r) && (! lizzieLet0_4QVal_Bool_4QNone_Bool_3QNone_Bool_bufchan_buf[0])))
        lizzieLet0_4QVal_Bool_4QNone_Bool_3QNone_Bool_bufchan_buf <= lizzieLet0_4QVal_Bool_4QNone_Bool_3QNone_Bool_bufchan_d;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_QTree_Bool) : (lizzieLet0_4QVal_Bool_4QNone_Bool_4,QTree_Bool) (lizzieLet0_4QVal_Bool_5QNone_Bool,Pointer_QTree_Bool) > [(lizzieLet0_4QVal_Bool_4QNone_Bool_4QNone_Bool,Pointer_QTree_Bool),
                                                                                                                                           (_67,Pointer_QTree_Bool),
                                                                                                                                           (_66,Pointer_QTree_Bool),
                                                                                                                                           (_65,Pointer_QTree_Bool)] */
  logic [3:0] lizzieLet0_4QVal_Bool_5QNone_Bool_onehotd;
  always_comb
    if ((lizzieLet0_4QVal_Bool_4QNone_Bool_4_d[0] && lizzieLet0_4QVal_Bool_5QNone_Bool_d[0]))
      unique case (lizzieLet0_4QVal_Bool_4QNone_Bool_4_d[2:1])
        2'd0: lizzieLet0_4QVal_Bool_5QNone_Bool_onehotd = 4'd1;
        2'd1: lizzieLet0_4QVal_Bool_5QNone_Bool_onehotd = 4'd2;
        2'd2: lizzieLet0_4QVal_Bool_5QNone_Bool_onehotd = 4'd4;
        2'd3: lizzieLet0_4QVal_Bool_5QNone_Bool_onehotd = 4'd8;
        default: lizzieLet0_4QVal_Bool_5QNone_Bool_onehotd = 4'd0;
      endcase
    else lizzieLet0_4QVal_Bool_5QNone_Bool_onehotd = 4'd0;
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_4QNone_Bool_d = {lizzieLet0_4QVal_Bool_5QNone_Bool_d[16:1],
                                                            lizzieLet0_4QVal_Bool_5QNone_Bool_onehotd[0]};
  assign _67_d = {lizzieLet0_4QVal_Bool_5QNone_Bool_d[16:1],
                  lizzieLet0_4QVal_Bool_5QNone_Bool_onehotd[1]};
  assign _66_d = {lizzieLet0_4QVal_Bool_5QNone_Bool_d[16:1],
                  lizzieLet0_4QVal_Bool_5QNone_Bool_onehotd[2]};
  assign _65_d = {lizzieLet0_4QVal_Bool_5QNone_Bool_d[16:1],
                  lizzieLet0_4QVal_Bool_5QNone_Bool_onehotd[3]};
  assign lizzieLet0_4QVal_Bool_5QNone_Bool_r = (| (lizzieLet0_4QVal_Bool_5QNone_Bool_onehotd & {_65_r,
                                                                                                _66_r,
                                                                                                _67_r,
                                                                                                lizzieLet0_4QVal_Bool_4QNone_Bool_4QNone_Bool_r}));
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_4_r = lizzieLet0_4QVal_Bool_5QNone_Bool_r;
  
  /* buf (Ty Pointer_QTree_Bool) : (lizzieLet0_4QVal_Bool_4QNone_Bool_4QNone_Bool,Pointer_QTree_Bool) > (lizzieLet0_4QVal_Bool_4QNone_Bool_4QNone_Bool_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t lizzieLet0_4QVal_Bool_4QNone_Bool_4QNone_Bool_bufchan_d;
  logic lizzieLet0_4QVal_Bool_4QNone_Bool_4QNone_Bool_bufchan_r;
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_4QNone_Bool_r = ((! lizzieLet0_4QVal_Bool_4QNone_Bool_4QNone_Bool_bufchan_d[0]) || lizzieLet0_4QVal_Bool_4QNone_Bool_4QNone_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_4QNone_Bool_4QNone_Bool_bufchan_d <= {16'd0,
                                                                  1'd0};
    else
      if (lizzieLet0_4QVal_Bool_4QNone_Bool_4QNone_Bool_r)
        lizzieLet0_4QVal_Bool_4QNone_Bool_4QNone_Bool_bufchan_d <= lizzieLet0_4QVal_Bool_4QNone_Bool_4QNone_Bool_d;
  Pointer_QTree_Bool_t lizzieLet0_4QVal_Bool_4QNone_Bool_4QNone_Bool_bufchan_buf;
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_4QNone_Bool_bufchan_r = (! lizzieLet0_4QVal_Bool_4QNone_Bool_4QNone_Bool_bufchan_buf[0]);
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_4QNone_Bool_1_argbuf_d = (lizzieLet0_4QVal_Bool_4QNone_Bool_4QNone_Bool_bufchan_buf[0] ? lizzieLet0_4QVal_Bool_4QNone_Bool_4QNone_Bool_bufchan_buf :
                                                                     lizzieLet0_4QVal_Bool_4QNone_Bool_4QNone_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_4QNone_Bool_4QNone_Bool_bufchan_buf <= {16'd0,
                                                                    1'd0};
    else
      if ((lizzieLet0_4QVal_Bool_4QNone_Bool_4QNone_Bool_1_argbuf_r && lizzieLet0_4QVal_Bool_4QNone_Bool_4QNone_Bool_bufchan_buf[0]))
        lizzieLet0_4QVal_Bool_4QNone_Bool_4QNone_Bool_bufchan_buf <= {16'd0,
                                                                      1'd0};
      else if (((! lizzieLet0_4QVal_Bool_4QNone_Bool_4QNone_Bool_1_argbuf_r) && (! lizzieLet0_4QVal_Bool_4QNone_Bool_4QNone_Bool_bufchan_buf[0])))
        lizzieLet0_4QVal_Bool_4QNone_Bool_4QNone_Bool_bufchan_buf <= lizzieLet0_4QVal_Bool_4QNone_Bool_4QNone_Bool_bufchan_d;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_CTf) : (lizzieLet0_4QVal_Bool_4QNone_Bool_5,QTree_Bool) (lizzieLet0_4QVal_Bool_7QNone_Bool,Pointer_CTf) > [(lizzieLet0_4QVal_Bool_4QNone_Bool_5QNone_Bool,Pointer_CTf),
                                                                                                                             (lizzieLet0_4QVal_Bool_4QNone_Bool_5QVal_Bool,Pointer_CTf),
                                                                                                                             (lizzieLet0_4QVal_Bool_4QNone_Bool_5QNode_Bool,Pointer_CTf),
                                                                                                                             (lizzieLet0_4QVal_Bool_4QNone_Bool_5QError_Bool,Pointer_CTf)] */
  logic [3:0] lizzieLet0_4QVal_Bool_7QNone_Bool_onehotd;
  always_comb
    if ((lizzieLet0_4QVal_Bool_4QNone_Bool_5_d[0] && lizzieLet0_4QVal_Bool_7QNone_Bool_d[0]))
      unique case (lizzieLet0_4QVal_Bool_4QNone_Bool_5_d[2:1])
        2'd0: lizzieLet0_4QVal_Bool_7QNone_Bool_onehotd = 4'd1;
        2'd1: lizzieLet0_4QVal_Bool_7QNone_Bool_onehotd = 4'd2;
        2'd2: lizzieLet0_4QVal_Bool_7QNone_Bool_onehotd = 4'd4;
        2'd3: lizzieLet0_4QVal_Bool_7QNone_Bool_onehotd = 4'd8;
        default: lizzieLet0_4QVal_Bool_7QNone_Bool_onehotd = 4'd0;
      endcase
    else lizzieLet0_4QVal_Bool_7QNone_Bool_onehotd = 4'd0;
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_5QNone_Bool_d = {lizzieLet0_4QVal_Bool_7QNone_Bool_d[16:1],
                                                            lizzieLet0_4QVal_Bool_7QNone_Bool_onehotd[0]};
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_5QVal_Bool_d = {lizzieLet0_4QVal_Bool_7QNone_Bool_d[16:1],
                                                           lizzieLet0_4QVal_Bool_7QNone_Bool_onehotd[1]};
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_5QNode_Bool_d = {lizzieLet0_4QVal_Bool_7QNone_Bool_d[16:1],
                                                            lizzieLet0_4QVal_Bool_7QNone_Bool_onehotd[2]};
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_5QError_Bool_d = {lizzieLet0_4QVal_Bool_7QNone_Bool_d[16:1],
                                                             lizzieLet0_4QVal_Bool_7QNone_Bool_onehotd[3]};
  assign lizzieLet0_4QVal_Bool_7QNone_Bool_r = (| (lizzieLet0_4QVal_Bool_7QNone_Bool_onehotd & {lizzieLet0_4QVal_Bool_4QNone_Bool_5QError_Bool_r,
                                                                                                lizzieLet0_4QVal_Bool_4QNone_Bool_5QNode_Bool_r,
                                                                                                lizzieLet0_4QVal_Bool_4QNone_Bool_5QVal_Bool_r,
                                                                                                lizzieLet0_4QVal_Bool_4QNone_Bool_5QNone_Bool_r}));
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_5_r = lizzieLet0_4QVal_Bool_7QNone_Bool_r;
  
  /* buf (Ty Pointer_CTf) : (lizzieLet0_4QVal_Bool_4QNone_Bool_5QError_Bool,Pointer_CTf) > (lizzieLet0_4QVal_Bool_4QNone_Bool_5QError_Bool_1_argbuf,Pointer_CTf) */
  Pointer_CTf_t lizzieLet0_4QVal_Bool_4QNone_Bool_5QError_Bool_bufchan_d;
  logic lizzieLet0_4QVal_Bool_4QNone_Bool_5QError_Bool_bufchan_r;
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_5QError_Bool_r = ((! lizzieLet0_4QVal_Bool_4QNone_Bool_5QError_Bool_bufchan_d[0]) || lizzieLet0_4QVal_Bool_4QNone_Bool_5QError_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_4QNone_Bool_5QError_Bool_bufchan_d <= {16'd0,
                                                                   1'd0};
    else
      if (lizzieLet0_4QVal_Bool_4QNone_Bool_5QError_Bool_r)
        lizzieLet0_4QVal_Bool_4QNone_Bool_5QError_Bool_bufchan_d <= lizzieLet0_4QVal_Bool_4QNone_Bool_5QError_Bool_d;
  Pointer_CTf_t lizzieLet0_4QVal_Bool_4QNone_Bool_5QError_Bool_bufchan_buf;
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_5QError_Bool_bufchan_r = (! lizzieLet0_4QVal_Bool_4QNone_Bool_5QError_Bool_bufchan_buf[0]);
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_5QError_Bool_1_argbuf_d = (lizzieLet0_4QVal_Bool_4QNone_Bool_5QError_Bool_bufchan_buf[0] ? lizzieLet0_4QVal_Bool_4QNone_Bool_5QError_Bool_bufchan_buf :
                                                                      lizzieLet0_4QVal_Bool_4QNone_Bool_5QError_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_4QNone_Bool_5QError_Bool_bufchan_buf <= {16'd0,
                                                                     1'd0};
    else
      if ((lizzieLet0_4QVal_Bool_4QNone_Bool_5QError_Bool_1_argbuf_r && lizzieLet0_4QVal_Bool_4QNone_Bool_5QError_Bool_bufchan_buf[0]))
        lizzieLet0_4QVal_Bool_4QNone_Bool_5QError_Bool_bufchan_buf <= {16'd0,
                                                                       1'd0};
      else if (((! lizzieLet0_4QVal_Bool_4QNone_Bool_5QError_Bool_1_argbuf_r) && (! lizzieLet0_4QVal_Bool_4QNone_Bool_5QError_Bool_bufchan_buf[0])))
        lizzieLet0_4QVal_Bool_4QNone_Bool_5QError_Bool_bufchan_buf <= lizzieLet0_4QVal_Bool_4QNone_Bool_5QError_Bool_bufchan_d;
  
  /* buf (Ty Pointer_CTf) : (lizzieLet0_4QVal_Bool_4QNone_Bool_5QNode_Bool,Pointer_CTf) > (lizzieLet0_4QVal_Bool_4QNone_Bool_5QNode_Bool_1_argbuf,Pointer_CTf) */
  Pointer_CTf_t lizzieLet0_4QVal_Bool_4QNone_Bool_5QNode_Bool_bufchan_d;
  logic lizzieLet0_4QVal_Bool_4QNone_Bool_5QNode_Bool_bufchan_r;
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_5QNode_Bool_r = ((! lizzieLet0_4QVal_Bool_4QNone_Bool_5QNode_Bool_bufchan_d[0]) || lizzieLet0_4QVal_Bool_4QNone_Bool_5QNode_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_4QNone_Bool_5QNode_Bool_bufchan_d <= {16'd0,
                                                                  1'd0};
    else
      if (lizzieLet0_4QVal_Bool_4QNone_Bool_5QNode_Bool_r)
        lizzieLet0_4QVal_Bool_4QNone_Bool_5QNode_Bool_bufchan_d <= lizzieLet0_4QVal_Bool_4QNone_Bool_5QNode_Bool_d;
  Pointer_CTf_t lizzieLet0_4QVal_Bool_4QNone_Bool_5QNode_Bool_bufchan_buf;
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_5QNode_Bool_bufchan_r = (! lizzieLet0_4QVal_Bool_4QNone_Bool_5QNode_Bool_bufchan_buf[0]);
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_5QNode_Bool_1_argbuf_d = (lizzieLet0_4QVal_Bool_4QNone_Bool_5QNode_Bool_bufchan_buf[0] ? lizzieLet0_4QVal_Bool_4QNone_Bool_5QNode_Bool_bufchan_buf :
                                                                     lizzieLet0_4QVal_Bool_4QNone_Bool_5QNode_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_4QNone_Bool_5QNode_Bool_bufchan_buf <= {16'd0,
                                                                    1'd0};
    else
      if ((lizzieLet0_4QVal_Bool_4QNone_Bool_5QNode_Bool_1_argbuf_r && lizzieLet0_4QVal_Bool_4QNone_Bool_5QNode_Bool_bufchan_buf[0]))
        lizzieLet0_4QVal_Bool_4QNone_Bool_5QNode_Bool_bufchan_buf <= {16'd0,
                                                                      1'd0};
      else if (((! lizzieLet0_4QVal_Bool_4QNone_Bool_5QNode_Bool_1_argbuf_r) && (! lizzieLet0_4QVal_Bool_4QNone_Bool_5QNode_Bool_bufchan_buf[0])))
        lizzieLet0_4QVal_Bool_4QNone_Bool_5QNode_Bool_bufchan_buf <= lizzieLet0_4QVal_Bool_4QNone_Bool_5QNode_Bool_bufchan_d;
  
  /* buf (Ty Pointer_CTf) : (lizzieLet0_4QVal_Bool_4QNone_Bool_5QNone_Bool,Pointer_CTf) > (lizzieLet0_4QVal_Bool_4QNone_Bool_5QNone_Bool_1_argbuf,Pointer_CTf) */
  Pointer_CTf_t lizzieLet0_4QVal_Bool_4QNone_Bool_5QNone_Bool_bufchan_d;
  logic lizzieLet0_4QVal_Bool_4QNone_Bool_5QNone_Bool_bufchan_r;
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_5QNone_Bool_r = ((! lizzieLet0_4QVal_Bool_4QNone_Bool_5QNone_Bool_bufchan_d[0]) || lizzieLet0_4QVal_Bool_4QNone_Bool_5QNone_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_4QNone_Bool_5QNone_Bool_bufchan_d <= {16'd0,
                                                                  1'd0};
    else
      if (lizzieLet0_4QVal_Bool_4QNone_Bool_5QNone_Bool_r)
        lizzieLet0_4QVal_Bool_4QNone_Bool_5QNone_Bool_bufchan_d <= lizzieLet0_4QVal_Bool_4QNone_Bool_5QNone_Bool_d;
  Pointer_CTf_t lizzieLet0_4QVal_Bool_4QNone_Bool_5QNone_Bool_bufchan_buf;
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_5QNone_Bool_bufchan_r = (! lizzieLet0_4QVal_Bool_4QNone_Bool_5QNone_Bool_bufchan_buf[0]);
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_5QNone_Bool_1_argbuf_d = (lizzieLet0_4QVal_Bool_4QNone_Bool_5QNone_Bool_bufchan_buf[0] ? lizzieLet0_4QVal_Bool_4QNone_Bool_5QNone_Bool_bufchan_buf :
                                                                     lizzieLet0_4QVal_Bool_4QNone_Bool_5QNone_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_4QNone_Bool_5QNone_Bool_bufchan_buf <= {16'd0,
                                                                    1'd0};
    else
      if ((lizzieLet0_4QVal_Bool_4QNone_Bool_5QNone_Bool_1_argbuf_r && lizzieLet0_4QVal_Bool_4QNone_Bool_5QNone_Bool_bufchan_buf[0]))
        lizzieLet0_4QVal_Bool_4QNone_Bool_5QNone_Bool_bufchan_buf <= {16'd0,
                                                                      1'd0};
      else if (((! lizzieLet0_4QVal_Bool_4QNone_Bool_5QNone_Bool_1_argbuf_r) && (! lizzieLet0_4QVal_Bool_4QNone_Bool_5QNone_Bool_bufchan_buf[0])))
        lizzieLet0_4QVal_Bool_4QNone_Bool_5QNone_Bool_bufchan_buf <= lizzieLet0_4QVal_Bool_4QNone_Bool_5QNone_Bool_bufchan_d;
  
  /* demux (Ty QTree_Bool,
       Ty MyBool) : (lizzieLet0_4QVal_Bool_4QNone_Bool_6,QTree_Bool) (lizzieLet0_4QVal_Bool_8QNone_Bool,MyBool) > [(_64,MyBool),
                                                                                                                   (lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool,MyBool),
                                                                                                                   (_63,MyBool),
                                                                                                                   (_62,MyBool)] */
  logic [3:0] lizzieLet0_4QVal_Bool_8QNone_Bool_onehotd;
  always_comb
    if ((lizzieLet0_4QVal_Bool_4QNone_Bool_6_d[0] && lizzieLet0_4QVal_Bool_8QNone_Bool_d[0]))
      unique case (lizzieLet0_4QVal_Bool_4QNone_Bool_6_d[2:1])
        2'd0: lizzieLet0_4QVal_Bool_8QNone_Bool_onehotd = 4'd1;
        2'd1: lizzieLet0_4QVal_Bool_8QNone_Bool_onehotd = 4'd2;
        2'd2: lizzieLet0_4QVal_Bool_8QNone_Bool_onehotd = 4'd4;
        2'd3: lizzieLet0_4QVal_Bool_8QNone_Bool_onehotd = 4'd8;
        default: lizzieLet0_4QVal_Bool_8QNone_Bool_onehotd = 4'd0;
      endcase
    else lizzieLet0_4QVal_Bool_8QNone_Bool_onehotd = 4'd0;
  assign _64_d = {lizzieLet0_4QVal_Bool_8QNone_Bool_d[1:1],
                  lizzieLet0_4QVal_Bool_8QNone_Bool_onehotd[0]};
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_d = {lizzieLet0_4QVal_Bool_8QNone_Bool_d[1:1],
                                                           lizzieLet0_4QVal_Bool_8QNone_Bool_onehotd[1]};
  assign _63_d = {lizzieLet0_4QVal_Bool_8QNone_Bool_d[1:1],
                  lizzieLet0_4QVal_Bool_8QNone_Bool_onehotd[2]};
  assign _62_d = {lizzieLet0_4QVal_Bool_8QNone_Bool_d[1:1],
                  lizzieLet0_4QVal_Bool_8QNone_Bool_onehotd[3]};
  assign lizzieLet0_4QVal_Bool_8QNone_Bool_r = (| (lizzieLet0_4QVal_Bool_8QNone_Bool_onehotd & {_62_r,
                                                                                                _63_r,
                                                                                                lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_r,
                                                                                                _64_r}));
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_6_r = lizzieLet0_4QVal_Bool_8QNone_Bool_r;
  
  /* fork (Ty MyBool) : (lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool,MyBool) > [(lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1,MyBool),
                                                                            (lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_2,MyBool),
                                                                            (lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3,MyBool)] */
  logic [2:0] lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_emitted;
  logic [2:0] lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_done;
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1_d = {lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_d[1:1],
                                                             (lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_d[0] && (! lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_emitted[0]))};
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_2_d = {lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_d[1:1],
                                                             (lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_d[0] && (! lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_emitted[1]))};
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3_d = {lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_d[1:1],
                                                             (lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_d[0] && (! lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_emitted[2]))};
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_done = (lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_emitted | ({lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3_d[0],
                                                                                                                       lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_2_d[0],
                                                                                                                       lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1_d[0]} & {lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3_r,
                                                                                                                                                                               lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_2_r,
                                                                                                                                                                               lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1_r}));
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_r = (& lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_emitted <= 3'd0;
    else
      lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_emitted <= (lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_r ? 3'd0 :
                                                               lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_done);
  
  /* demux (Ty MyBool,
       Ty Go) : (lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1,MyBool) (lizzieLet0_4QVal_Bool_4QNone_Bool_3QVal_Bool,Go) > [(lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyFalse,Go),
                                                                                                                             (lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyTrue,Go)] */
  logic [1:0] lizzieLet0_4QVal_Bool_4QNone_Bool_3QVal_Bool_onehotd;
  always_comb
    if ((lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1_d[0] && lizzieLet0_4QVal_Bool_4QNone_Bool_3QVal_Bool_d[0]))
      unique case (lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1_d[1:1])
        1'd0: lizzieLet0_4QVal_Bool_4QNone_Bool_3QVal_Bool_onehotd = 2'd1;
        1'd1: lizzieLet0_4QVal_Bool_4QNone_Bool_3QVal_Bool_onehotd = 2'd2;
        default:
          lizzieLet0_4QVal_Bool_4QNone_Bool_3QVal_Bool_onehotd = 2'd0;
      endcase
    else lizzieLet0_4QVal_Bool_4QNone_Bool_3QVal_Bool_onehotd = 2'd0;
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyFalse_d = lizzieLet0_4QVal_Bool_4QNone_Bool_3QVal_Bool_onehotd[0];
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyTrue_d = lizzieLet0_4QVal_Bool_4QNone_Bool_3QVal_Bool_onehotd[1];
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_3QVal_Bool_r = (| (lizzieLet0_4QVal_Bool_4QNone_Bool_3QVal_Bool_onehotd & {lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyTrue_r,
                                                                                                                      lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyFalse_r}));
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1_r = lizzieLet0_4QVal_Bool_4QNone_Bool_3QVal_Bool_r;
  
  /* fork (Ty Go) : (lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyTrue,Go) > [(lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyTrue_1,Go),
                                                                            (lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyTrue_2,Go)] */
  logic [1:0] lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyTrue_emitted;
  logic [1:0] lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyTrue_done;
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyTrue_1_d = (lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyTrue_d[0] && (! lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyTrue_emitted[0]));
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyTrue_2_d = (lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyTrue_d[0] && (! lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyTrue_emitted[1]));
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyTrue_done = (lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyTrue_emitted | ({lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyTrue_2_d[0],
                                                                                                                                       lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyTrue_1_d[0]} & {lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyTrue_2_r,
                                                                                                                                                                                                       lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyTrue_1_r}));
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyTrue_r = (& lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyTrue_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyTrue_emitted <= 2'd0;
    else
      lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyTrue_emitted <= (lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyTrue_r ? 2'd0 :
                                                                       lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyTrue_done);
  
  /* buf (Ty Go) : (lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyTrue_1,Go) > (lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyTrue_1_argbuf,Go) */
  Go_t lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyTrue_1_bufchan_d;
  logic lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyTrue_1_bufchan_r;
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyTrue_1_r = ((! lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyTrue_1_bufchan_d[0]) || lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyTrue_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyTrue_1_bufchan_d <= 1'd0;
    else
      if (lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyTrue_1_r)
        lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyTrue_1_bufchan_d <= lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyTrue_1_d;
  Go_t lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyTrue_1_bufchan_buf;
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyTrue_1_bufchan_r = (! lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyTrue_1_bufchan_buf[0]);
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyTrue_1_argbuf_d = (lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyTrue_1_bufchan_buf[0] ? lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyTrue_1_bufchan_buf :
                                                                            lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyTrue_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyTrue_1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyTrue_1_argbuf_r && lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyTrue_1_bufchan_buf[0]))
        lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyTrue_1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyTrue_1_argbuf_r) && (! lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyTrue_1_bufchan_buf[0])))
        lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyTrue_1_bufchan_buf <= lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyTrue_1_bufchan_d;
  
  /* dcon (Ty TupGo,
      Dcon TupGo) : [(lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyTrue_1_argbuf,Go)] > (lvlrf2-0TupGo6,TupGo) */
  assign \lvlrf2-0TupGo6_d  = TupGo_dc((& {lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyTrue_1_argbuf_d[0]}), lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyTrue_1_argbuf_d);
  assign {lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyTrue_1_argbuf_r} = {1 {(\lvlrf2-0TupGo6_r  && \lvlrf2-0TupGo6_d [0])}};
  
  /* buf (Ty Go) : (lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyTrue_2,Go) > (lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyTrue_2_argbuf,Go) */
  Go_t lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyTrue_2_bufchan_d;
  logic lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyTrue_2_bufchan_r;
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyTrue_2_r = ((! lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyTrue_2_bufchan_d[0]) || lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyTrue_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyTrue_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyTrue_2_r)
        lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyTrue_2_bufchan_d <= lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyTrue_2_d;
  Go_t lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyTrue_2_bufchan_buf;
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyTrue_2_bufchan_r = (! lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyTrue_2_bufchan_buf[0]);
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyTrue_2_argbuf_d = (lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyTrue_2_bufchan_buf[0] ? lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyTrue_2_bufchan_buf :
                                                                            lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyTrue_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyTrue_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyTrue_2_argbuf_r && lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyTrue_2_bufchan_buf[0]))
        lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyTrue_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyTrue_2_argbuf_r) && (! lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyTrue_2_bufchan_buf[0])))
        lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyTrue_2_bufchan_buf <= lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyTrue_2_bufchan_d;
  
  /* demux (Ty MyBool,
       Ty Pointer_CTf) : (lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_2,MyBool) (lizzieLet0_4QVal_Bool_4QNone_Bool_5QVal_Bool,Pointer_CTf) > [(lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_2MyFalse,Pointer_CTf),
                                                                                                                                               (lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_2MyTrue,Pointer_CTf)] */
  logic [1:0] lizzieLet0_4QVal_Bool_4QNone_Bool_5QVal_Bool_onehotd;
  always_comb
    if ((lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_2_d[0] && lizzieLet0_4QVal_Bool_4QNone_Bool_5QVal_Bool_d[0]))
      unique case (lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_2_d[1:1])
        1'd0: lizzieLet0_4QVal_Bool_4QNone_Bool_5QVal_Bool_onehotd = 2'd1;
        1'd1: lizzieLet0_4QVal_Bool_4QNone_Bool_5QVal_Bool_onehotd = 2'd2;
        default:
          lizzieLet0_4QVal_Bool_4QNone_Bool_5QVal_Bool_onehotd = 2'd0;
      endcase
    else lizzieLet0_4QVal_Bool_4QNone_Bool_5QVal_Bool_onehotd = 2'd0;
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_2MyFalse_d = {lizzieLet0_4QVal_Bool_4QNone_Bool_5QVal_Bool_d[16:1],
                                                                    lizzieLet0_4QVal_Bool_4QNone_Bool_5QVal_Bool_onehotd[0]};
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_2MyTrue_d = {lizzieLet0_4QVal_Bool_4QNone_Bool_5QVal_Bool_d[16:1],
                                                                   lizzieLet0_4QVal_Bool_4QNone_Bool_5QVal_Bool_onehotd[1]};
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_5QVal_Bool_r = (| (lizzieLet0_4QVal_Bool_4QNone_Bool_5QVal_Bool_onehotd & {lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_2MyTrue_r,
                                                                                                                      lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_2MyFalse_r}));
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_2_r = lizzieLet0_4QVal_Bool_4QNone_Bool_5QVal_Bool_r;
  
  /* buf (Ty Pointer_CTf) : (lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_2MyTrue,Pointer_CTf) > (lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_2MyTrue_1_argbuf,Pointer_CTf) */
  Pointer_CTf_t lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_2MyTrue_bufchan_d;
  logic lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_2MyTrue_bufchan_r;
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_2MyTrue_r = ((! lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_2MyTrue_bufchan_d[0]) || lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_2MyTrue_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_2MyTrue_bufchan_d <= {16'd0,
                                                                         1'd0};
    else
      if (lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_2MyTrue_r)
        lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_2MyTrue_bufchan_d <= lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_2MyTrue_d;
  Pointer_CTf_t lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_2MyTrue_bufchan_buf;
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_2MyTrue_bufchan_r = (! lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_2MyTrue_bufchan_buf[0]);
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_2MyTrue_1_argbuf_d = (lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_2MyTrue_bufchan_buf[0] ? lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_2MyTrue_bufchan_buf :
                                                                            lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_2MyTrue_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_2MyTrue_bufchan_buf <= {16'd0,
                                                                           1'd0};
    else
      if ((lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_2MyTrue_1_argbuf_r && lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_2MyTrue_bufchan_buf[0]))
        lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_2MyTrue_bufchan_buf <= {16'd0,
                                                                             1'd0};
      else if (((! lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_2MyTrue_1_argbuf_r) && (! lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_2MyTrue_bufchan_buf[0])))
        lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_2MyTrue_bufchan_buf <= lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_2MyTrue_bufchan_d;
  
  /* demux (Ty MyBool,
       Ty MyBool) : (lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3,MyBool) (va8n_destruct,MyBool) > [(lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse,MyBool),
                                                                                                      (_61,MyBool)] */
  logic [1:0] va8n_destruct_onehotd;
  always_comb
    if ((lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3_d[0] && va8n_destruct_d[0]))
      unique case (lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3_d[1:1])
        1'd0: va8n_destruct_onehotd = 2'd1;
        1'd1: va8n_destruct_onehotd = 2'd2;
        default: va8n_destruct_onehotd = 2'd0;
      endcase
    else va8n_destruct_onehotd = 2'd0;
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_d = {va8n_destruct_d[1:1],
                                                                    va8n_destruct_onehotd[0]};
  assign _61_d = {va8n_destruct_d[1:1], va8n_destruct_onehotd[1]};
  assign va8n_destruct_r = (| (va8n_destruct_onehotd & {_61_r,
                                                        lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_r}));
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3_r = va8n_destruct_r;
  
  /* fork (Ty MyBool) : (lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse,MyBool) > [(lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1,MyBool),
                                                                                     (lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_2,MyBool)] */
  logic [1:0] lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_emitted;
  logic [1:0] lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_done;
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1_d = {lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_d[1:1],
                                                                      (lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_d[0] && (! lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_emitted[0]))};
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_2_d = {lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_d[1:1],
                                                                      (lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_d[0] && (! lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_emitted[1]))};
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_done = (lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_emitted | ({lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_2_d[0],
                                                                                                                                         lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1_d[0]} & {lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_2_r,
                                                                                                                                                                                                          lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1_r}));
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_r = (& lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_emitted <= 2'd0;
    else
      lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_emitted <= (lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_r ? 2'd0 :
                                                                        lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_done);
  
  /* demux (Ty MyBool,
       Ty Go) : (lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1,MyBool) (lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyFalse,Go) > [(lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyFalse,Go),
                                                                                                                                               (lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyTrue,Go)] */
  logic [1:0] lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyFalse_onehotd;
  always_comb
    if ((lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1_d[0] && lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyFalse_d[0]))
      unique case (lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1_d[1:1])
        1'd0:
          lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyFalse_onehotd = 2'd1;
        1'd1:
          lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyFalse_onehotd = 2'd2;
        default:
          lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyFalse_onehotd = 2'd0;
      endcase
    else
      lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyFalse_onehotd = 2'd0;
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyFalse_d = lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyFalse_onehotd[0];
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyTrue_d = lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyFalse_onehotd[1];
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyFalse_r = (| (lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyFalse_onehotd & {lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyTrue_r,
                                                                                                                                        lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyFalse_r}));
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1_r = lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_1MyFalse_r;
  
  /* fork (Ty Go) : (lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyFalse,Go) > [(lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyFalse_1,Go),
                                                                                      (lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyFalse_2,Go)] */
  logic [1:0] lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyFalse_emitted;
  logic [1:0] lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyFalse_done;
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyFalse_1_d = (lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyFalse_d[0] && (! lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyFalse_emitted[0]));
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_d = (lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyFalse_d[0] && (! lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyFalse_emitted[1]));
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyFalse_done = (lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyFalse_emitted | ({lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_d[0],
                                                                                                                                                           lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyFalse_1_d[0]} & {lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_r,
                                                                                                                                                                                                                                     lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyFalse_1_r}));
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyFalse_r = (& lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyFalse_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyFalse_emitted <= 2'd0;
    else
      lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyFalse_emitted <= (lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyFalse_r ? 2'd0 :
                                                                                 lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyFalse_done);
  
  /* dcon (Ty QTree_Bool,
      Dcon QNone_Bool) : [(lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyFalse_1,Go)] > (lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool,QTree_Bool) */
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_d = QNone_Bool_dc((& {lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyFalse_1_d[0]}), lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyFalse_1_d);
  assign {lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyFalse_1_r} = {1 {(lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_r && lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_d[0])}};
  
  /* buf (Ty QTree_Bool) : (lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool,QTree_Bool) > (lizzieLet15_1_1_argbuf,QTree_Bool) */
  QTree_Bool_t lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_bufchan_d;
  logic lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_bufchan_r;
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_r = ((! lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_bufchan_d[0]) || lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_bufchan_d <= {66'd0,
                                                                                               1'd0};
    else
      if (lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_r)
        lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_bufchan_d <= lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_d;
  QTree_Bool_t lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_bufchan_buf;
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_bufchan_r = (! lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_bufchan_buf[0]);
  assign lizzieLet15_1_1_argbuf_d = (lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_bufchan_buf[0] ? lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_bufchan_buf :
                                     lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_bufchan_buf <= {66'd0,
                                                                                                 1'd0};
    else
      if ((lizzieLet15_1_1_argbuf_r && lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_bufchan_buf[0]))
        lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_bufchan_buf <= {66'd0,
                                                                                                   1'd0};
      else if (((! lizzieLet15_1_1_argbuf_r) && (! lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_bufchan_buf[0])))
        lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_bufchan_buf <= lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyFalse_2,Go) > (lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_argbuf,Go) */
  Go_t lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_bufchan_d;
  logic lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_bufchan_r;
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_r = ((! lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_bufchan_d[0]) || lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_r)
        lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_bufchan_d <= lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_d;
  Go_t lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_bufchan_buf;
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_bufchan_r = (! lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_bufchan_buf[0]);
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_argbuf_d = (lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_bufchan_buf[0] ? lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_bufchan_buf :
                                                                                      lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_argbuf_r && lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_bufchan_buf[0]))
        lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_argbuf_r) && (! lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_bufchan_buf[0])))
        lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_bufchan_buf <= lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyTrue,Go) > [(lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyTrue_1,Go),
                                                                                     (lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyTrue_2,Go)] */
  logic [1:0] lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyTrue_emitted;
  logic [1:0] lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyTrue_done;
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_d = (lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyTrue_d[0] && (! lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyTrue_emitted[0]));
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_d = (lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyTrue_d[0] && (! lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyTrue_emitted[1]));
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyTrue_done = (lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyTrue_emitted | ({lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_d[0],
                                                                                                                                                         lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_d[0]} & {lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_r,
                                                                                                                                                                                                                                  lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_r}));
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyTrue_r = (& lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyTrue_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyTrue_emitted <= 2'd0;
    else
      lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyTrue_emitted <= (lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyTrue_r ? 2'd0 :
                                                                                lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyTrue_done);
  
  /* buf (Ty Go) : (lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyTrue_1,Go) > (lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_argbuf,Go) */
  Go_t lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_bufchan_d;
  logic lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_bufchan_r;
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_r = ((! lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_bufchan_d[0]) || lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_bufchan_d <= 1'd0;
    else
      if (lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_r)
        lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_bufchan_d <= lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_d;
  Go_t lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_bufchan_buf;
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_bufchan_r = (! lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_bufchan_buf[0]);
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_argbuf_d = (lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_bufchan_buf[0] ? lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_bufchan_buf :
                                                                                     lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_argbuf_r && lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_bufchan_buf[0]))
        lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_argbuf_r) && (! lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_bufchan_buf[0])))
        lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_bufchan_buf <= lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_bufchan_d;
  
  /* dcon (Ty TupGo,
      Dcon TupGo) : [(lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_argbuf,Go)] > (lvlrf2-0TupGo5,TupGo) */
  assign \lvlrf2-0TupGo5_d  = TupGo_dc((& {lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_argbuf_d[0]}), lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_argbuf_d);
  assign {lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_argbuf_r} = {1 {(\lvlrf2-0TupGo5_r  && \lvlrf2-0TupGo5_d [0])}};
  
  /* buf (Ty Go) : (lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyTrue_2,Go) > (lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_argbuf,Go) */
  Go_t lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_bufchan_d;
  logic lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_bufchan_r;
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_r = ((! lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_bufchan_d[0]) || lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_r)
        lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_bufchan_d <= lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_d;
  Go_t lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_bufchan_buf;
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_bufchan_r = (! lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_bufchan_buf[0]);
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_argbuf_d = (lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_bufchan_buf[0] ? lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_bufchan_buf :
                                                                                     lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_argbuf_r && lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_bufchan_buf[0]))
        lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_argbuf_r) && (! lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_bufchan_buf[0])))
        lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_bufchan_buf <= lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_bufchan_d;
  
  /* demux (Ty MyBool,
       Ty Pointer_CTf) : (lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_2,MyBool) (lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_2MyFalse,Pointer_CTf) > [(lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_2MyFalse,Pointer_CTf),
                                                                                                                                                                 (lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_2MyTrue,Pointer_CTf)] */
  logic [1:0] lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_2MyFalse_onehotd;
  always_comb
    if ((lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_2_d[0] && lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_2MyFalse_d[0]))
      unique case (lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_2_d[1:1])
        1'd0:
          lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_2MyFalse_onehotd = 2'd1;
        1'd1:
          lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_2MyFalse_onehotd = 2'd2;
        default:
          lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_2MyFalse_onehotd = 2'd0;
      endcase
    else
      lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_2MyFalse_onehotd = 2'd0;
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_2MyFalse_d = {lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_2MyFalse_d[16:1],
                                                                             lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_2MyFalse_onehotd[0]};
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_2MyTrue_d = {lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_2MyFalse_d[16:1],
                                                                            lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_2MyFalse_onehotd[1]};
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_2MyFalse_r = (| (lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_2MyFalse_onehotd & {lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_2MyTrue_r,
                                                                                                                                        lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_2MyFalse_r}));
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_2_r = lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_2MyFalse_r;
  
  /* buf (Ty Pointer_CTf) : (lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_2MyFalse,Pointer_CTf) > (lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_2MyFalse_1_argbuf,Pointer_CTf) */
  Pointer_CTf_t lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_2MyFalse_bufchan_d;
  logic lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_2MyFalse_bufchan_r;
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_2MyFalse_r = ((! lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_2MyFalse_bufchan_d[0]) || lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_2MyFalse_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_2MyFalse_bufchan_d <= {16'd0,
                                                                                   1'd0};
    else
      if (lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_2MyFalse_r)
        lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_2MyFalse_bufchan_d <= lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_2MyFalse_d;
  Pointer_CTf_t lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_2MyFalse_bufchan_buf;
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_2MyFalse_bufchan_r = (! lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_2MyFalse_bufchan_buf[0]);
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_2MyFalse_1_argbuf_d = (lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_2MyFalse_bufchan_buf[0] ? lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_2MyFalse_bufchan_buf :
                                                                                      lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_2MyFalse_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_2MyFalse_bufchan_buf <= {16'd0,
                                                                                     1'd0};
    else
      if ((lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_2MyFalse_1_argbuf_r && lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_2MyFalse_bufchan_buf[0]))
        lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_2MyFalse_bufchan_buf <= {16'd0,
                                                                                       1'd0};
      else if (((! lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_2MyFalse_1_argbuf_r) && (! lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_2MyFalse_bufchan_buf[0])))
        lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_2MyFalse_bufchan_buf <= lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_2MyFalse_bufchan_d;
  
  /* buf (Ty Pointer_CTf) : (lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_2MyTrue,Pointer_CTf) > (lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_2MyTrue_1_argbuf,Pointer_CTf) */
  Pointer_CTf_t lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_2MyTrue_bufchan_d;
  logic lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_2MyTrue_bufchan_r;
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_2MyTrue_r = ((! lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_2MyTrue_bufchan_d[0]) || lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_2MyTrue_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_2MyTrue_bufchan_d <= {16'd0,
                                                                                  1'd0};
    else
      if (lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_2MyTrue_r)
        lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_2MyTrue_bufchan_d <= lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_2MyTrue_d;
  Pointer_CTf_t lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_2MyTrue_bufchan_buf;
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_2MyTrue_bufchan_r = (! lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_2MyTrue_bufchan_buf[0]);
  assign lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_2MyTrue_1_argbuf_d = (lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_2MyTrue_bufchan_buf[0] ? lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_2MyTrue_bufchan_buf :
                                                                                     lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_2MyTrue_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_2MyTrue_bufchan_buf <= {16'd0,
                                                                                    1'd0};
    else
      if ((lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_2MyTrue_1_argbuf_r && lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_2MyTrue_bufchan_buf[0]))
        lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_2MyTrue_bufchan_buf <= {16'd0,
                                                                                      1'd0};
      else if (((! lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_2MyTrue_1_argbuf_r) && (! lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_2MyTrue_bufchan_buf[0])))
        lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_2MyTrue_bufchan_buf <= lizzieLet0_4QVal_Bool_4QNone_Bool_6QVal_Bool_3MyFalse_2MyTrue_bufchan_d;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_QTree_Bool) : (lizzieLet0_4QVal_Bool_5,QTree_Bool) (lizzieLet0_6QVal_Bool,Pointer_QTree_Bool) > [(lizzieLet0_4QVal_Bool_5QNone_Bool,Pointer_QTree_Bool),
                                                                                                                   (_60,Pointer_QTree_Bool),
                                                                                                                   (_59,Pointer_QTree_Bool),
                                                                                                                   (_58,Pointer_QTree_Bool)] */
  logic [3:0] lizzieLet0_6QVal_Bool_onehotd;
  always_comb
    if ((lizzieLet0_4QVal_Bool_5_d[0] && lizzieLet0_6QVal_Bool_d[0]))
      unique case (lizzieLet0_4QVal_Bool_5_d[2:1])
        2'd0: lizzieLet0_6QVal_Bool_onehotd = 4'd1;
        2'd1: lizzieLet0_6QVal_Bool_onehotd = 4'd2;
        2'd2: lizzieLet0_6QVal_Bool_onehotd = 4'd4;
        2'd3: lizzieLet0_6QVal_Bool_onehotd = 4'd8;
        default: lizzieLet0_6QVal_Bool_onehotd = 4'd0;
      endcase
    else lizzieLet0_6QVal_Bool_onehotd = 4'd0;
  assign lizzieLet0_4QVal_Bool_5QNone_Bool_d = {lizzieLet0_6QVal_Bool_d[16:1],
                                                lizzieLet0_6QVal_Bool_onehotd[0]};
  assign _60_d = {lizzieLet0_6QVal_Bool_d[16:1],
                  lizzieLet0_6QVal_Bool_onehotd[1]};
  assign _59_d = {lizzieLet0_6QVal_Bool_d[16:1],
                  lizzieLet0_6QVal_Bool_onehotd[2]};
  assign _58_d = {lizzieLet0_6QVal_Bool_d[16:1],
                  lizzieLet0_6QVal_Bool_onehotd[3]};
  assign lizzieLet0_6QVal_Bool_r = (| (lizzieLet0_6QVal_Bool_onehotd & {_58_r,
                                                                        _59_r,
                                                                        _60_r,
                                                                        lizzieLet0_4QVal_Bool_5QNone_Bool_r}));
  assign lizzieLet0_4QVal_Bool_5_r = lizzieLet0_6QVal_Bool_r;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_QTree_Bool) : (lizzieLet0_4QVal_Bool_6,QTree_Bool) (lizzieLet0_8QVal_Bool,Pointer_QTree_Bool) > [(_57,Pointer_QTree_Bool),
                                                                                                                   (lizzieLet0_4QVal_Bool_6QVal_Bool,Pointer_QTree_Bool),
                                                                                                                   (_56,Pointer_QTree_Bool),
                                                                                                                   (_55,Pointer_QTree_Bool)] */
  logic [3:0] lizzieLet0_8QVal_Bool_onehotd;
  always_comb
    if ((lizzieLet0_4QVal_Bool_6_d[0] && lizzieLet0_8QVal_Bool_d[0]))
      unique case (lizzieLet0_4QVal_Bool_6_d[2:1])
        2'd0: lizzieLet0_8QVal_Bool_onehotd = 4'd1;
        2'd1: lizzieLet0_8QVal_Bool_onehotd = 4'd2;
        2'd2: lizzieLet0_8QVal_Bool_onehotd = 4'd4;
        2'd3: lizzieLet0_8QVal_Bool_onehotd = 4'd8;
        default: lizzieLet0_8QVal_Bool_onehotd = 4'd0;
      endcase
    else lizzieLet0_8QVal_Bool_onehotd = 4'd0;
  assign _57_d = {lizzieLet0_8QVal_Bool_d[16:1],
                  lizzieLet0_8QVal_Bool_onehotd[0]};
  assign lizzieLet0_4QVal_Bool_6QVal_Bool_d = {lizzieLet0_8QVal_Bool_d[16:1],
                                               lizzieLet0_8QVal_Bool_onehotd[1]};
  assign _56_d = {lizzieLet0_8QVal_Bool_d[16:1],
                  lizzieLet0_8QVal_Bool_onehotd[2]};
  assign _55_d = {lizzieLet0_8QVal_Bool_d[16:1],
                  lizzieLet0_8QVal_Bool_onehotd[3]};
  assign lizzieLet0_8QVal_Bool_r = (| (lizzieLet0_8QVal_Bool_onehotd & {_55_r,
                                                                        _56_r,
                                                                        lizzieLet0_4QVal_Bool_6QVal_Bool_r,
                                                                        _57_r}));
  assign lizzieLet0_4QVal_Bool_6_r = lizzieLet0_8QVal_Bool_r;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_CTf) : (lizzieLet0_4QVal_Bool_7,QTree_Bool) (lizzieLet0_9QVal_Bool,Pointer_CTf) > [(lizzieLet0_4QVal_Bool_7QNone_Bool,Pointer_CTf),
                                                                                                     (lizzieLet0_4QVal_Bool_7QVal_Bool,Pointer_CTf),
                                                                                                     (lizzieLet0_4QVal_Bool_7QNode_Bool,Pointer_CTf),
                                                                                                     (lizzieLet0_4QVal_Bool_7QError_Bool,Pointer_CTf)] */
  logic [3:0] lizzieLet0_9QVal_Bool_onehotd;
  always_comb
    if ((lizzieLet0_4QVal_Bool_7_d[0] && lizzieLet0_9QVal_Bool_d[0]))
      unique case (lizzieLet0_4QVal_Bool_7_d[2:1])
        2'd0: lizzieLet0_9QVal_Bool_onehotd = 4'd1;
        2'd1: lizzieLet0_9QVal_Bool_onehotd = 4'd2;
        2'd2: lizzieLet0_9QVal_Bool_onehotd = 4'd4;
        2'd3: lizzieLet0_9QVal_Bool_onehotd = 4'd8;
        default: lizzieLet0_9QVal_Bool_onehotd = 4'd0;
      endcase
    else lizzieLet0_9QVal_Bool_onehotd = 4'd0;
  assign lizzieLet0_4QVal_Bool_7QNone_Bool_d = {lizzieLet0_9QVal_Bool_d[16:1],
                                                lizzieLet0_9QVal_Bool_onehotd[0]};
  assign lizzieLet0_4QVal_Bool_7QVal_Bool_d = {lizzieLet0_9QVal_Bool_d[16:1],
                                               lizzieLet0_9QVal_Bool_onehotd[1]};
  assign lizzieLet0_4QVal_Bool_7QNode_Bool_d = {lizzieLet0_9QVal_Bool_d[16:1],
                                                lizzieLet0_9QVal_Bool_onehotd[2]};
  assign lizzieLet0_4QVal_Bool_7QError_Bool_d = {lizzieLet0_9QVal_Bool_d[16:1],
                                                 lizzieLet0_9QVal_Bool_onehotd[3]};
  assign lizzieLet0_9QVal_Bool_r = (| (lizzieLet0_9QVal_Bool_onehotd & {lizzieLet0_4QVal_Bool_7QError_Bool_r,
                                                                        lizzieLet0_4QVal_Bool_7QNode_Bool_r,
                                                                        lizzieLet0_4QVal_Bool_7QVal_Bool_r,
                                                                        lizzieLet0_4QVal_Bool_7QNone_Bool_r}));
  assign lizzieLet0_4QVal_Bool_7_r = lizzieLet0_9QVal_Bool_r;
  
  /* buf (Ty Pointer_CTf) : (lizzieLet0_4QVal_Bool_7QError_Bool,Pointer_CTf) > (lizzieLet0_4QVal_Bool_7QError_Bool_1_argbuf,Pointer_CTf) */
  Pointer_CTf_t lizzieLet0_4QVal_Bool_7QError_Bool_bufchan_d;
  logic lizzieLet0_4QVal_Bool_7QError_Bool_bufchan_r;
  assign lizzieLet0_4QVal_Bool_7QError_Bool_r = ((! lizzieLet0_4QVal_Bool_7QError_Bool_bufchan_d[0]) || lizzieLet0_4QVal_Bool_7QError_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_7QError_Bool_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet0_4QVal_Bool_7QError_Bool_r)
        lizzieLet0_4QVal_Bool_7QError_Bool_bufchan_d <= lizzieLet0_4QVal_Bool_7QError_Bool_d;
  Pointer_CTf_t lizzieLet0_4QVal_Bool_7QError_Bool_bufchan_buf;
  assign lizzieLet0_4QVal_Bool_7QError_Bool_bufchan_r = (! lizzieLet0_4QVal_Bool_7QError_Bool_bufchan_buf[0]);
  assign lizzieLet0_4QVal_Bool_7QError_Bool_1_argbuf_d = (lizzieLet0_4QVal_Bool_7QError_Bool_bufchan_buf[0] ? lizzieLet0_4QVal_Bool_7QError_Bool_bufchan_buf :
                                                          lizzieLet0_4QVal_Bool_7QError_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_7QError_Bool_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet0_4QVal_Bool_7QError_Bool_1_argbuf_r && lizzieLet0_4QVal_Bool_7QError_Bool_bufchan_buf[0]))
        lizzieLet0_4QVal_Bool_7QError_Bool_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet0_4QVal_Bool_7QError_Bool_1_argbuf_r) && (! lizzieLet0_4QVal_Bool_7QError_Bool_bufchan_buf[0])))
        lizzieLet0_4QVal_Bool_7QError_Bool_bufchan_buf <= lizzieLet0_4QVal_Bool_7QError_Bool_bufchan_d;
  
  /* buf (Ty Pointer_CTf) : (lizzieLet0_4QVal_Bool_7QNode_Bool,Pointer_CTf) > (lizzieLet0_4QVal_Bool_7QNode_Bool_1_argbuf,Pointer_CTf) */
  Pointer_CTf_t lizzieLet0_4QVal_Bool_7QNode_Bool_bufchan_d;
  logic lizzieLet0_4QVal_Bool_7QNode_Bool_bufchan_r;
  assign lizzieLet0_4QVal_Bool_7QNode_Bool_r = ((! lizzieLet0_4QVal_Bool_7QNode_Bool_bufchan_d[0]) || lizzieLet0_4QVal_Bool_7QNode_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_7QNode_Bool_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet0_4QVal_Bool_7QNode_Bool_r)
        lizzieLet0_4QVal_Bool_7QNode_Bool_bufchan_d <= lizzieLet0_4QVal_Bool_7QNode_Bool_d;
  Pointer_CTf_t lizzieLet0_4QVal_Bool_7QNode_Bool_bufchan_buf;
  assign lizzieLet0_4QVal_Bool_7QNode_Bool_bufchan_r = (! lizzieLet0_4QVal_Bool_7QNode_Bool_bufchan_buf[0]);
  assign lizzieLet0_4QVal_Bool_7QNode_Bool_1_argbuf_d = (lizzieLet0_4QVal_Bool_7QNode_Bool_bufchan_buf[0] ? lizzieLet0_4QVal_Bool_7QNode_Bool_bufchan_buf :
                                                         lizzieLet0_4QVal_Bool_7QNode_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_7QNode_Bool_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet0_4QVal_Bool_7QNode_Bool_1_argbuf_r && lizzieLet0_4QVal_Bool_7QNode_Bool_bufchan_buf[0]))
        lizzieLet0_4QVal_Bool_7QNode_Bool_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet0_4QVal_Bool_7QNode_Bool_1_argbuf_r) && (! lizzieLet0_4QVal_Bool_7QNode_Bool_bufchan_buf[0])))
        lizzieLet0_4QVal_Bool_7QNode_Bool_bufchan_buf <= lizzieLet0_4QVal_Bool_7QNode_Bool_bufchan_d;
  
  /* demux (Ty QTree_Bool,
       Ty MyBool) : (lizzieLet0_4QVal_Bool_8,QTree_Bool) (v1a8m_destruct,MyBool) > [(lizzieLet0_4QVal_Bool_8QNone_Bool,MyBool),
                                                                                    (lizzieLet0_4QVal_Bool_8QVal_Bool,MyBool),
                                                                                    (_54,MyBool),
                                                                                    (_53,MyBool)] */
  logic [3:0] v1a8m_destruct_onehotd;
  always_comb
    if ((lizzieLet0_4QVal_Bool_8_d[0] && v1a8m_destruct_d[0]))
      unique case (lizzieLet0_4QVal_Bool_8_d[2:1])
        2'd0: v1a8m_destruct_onehotd = 4'd1;
        2'd1: v1a8m_destruct_onehotd = 4'd2;
        2'd2: v1a8m_destruct_onehotd = 4'd4;
        2'd3: v1a8m_destruct_onehotd = 4'd8;
        default: v1a8m_destruct_onehotd = 4'd0;
      endcase
    else v1a8m_destruct_onehotd = 4'd0;
  assign lizzieLet0_4QVal_Bool_8QNone_Bool_d = {v1a8m_destruct_d[1:1],
                                                v1a8m_destruct_onehotd[0]};
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_d = {v1a8m_destruct_d[1:1],
                                               v1a8m_destruct_onehotd[1]};
  assign _54_d = {v1a8m_destruct_d[1:1], v1a8m_destruct_onehotd[2]};
  assign _53_d = {v1a8m_destruct_d[1:1], v1a8m_destruct_onehotd[3]};
  assign v1a8m_destruct_r = (| (v1a8m_destruct_onehotd & {_53_r,
                                                          _54_r,
                                                          lizzieLet0_4QVal_Bool_8QVal_Bool_r,
                                                          lizzieLet0_4QVal_Bool_8QNone_Bool_r}));
  assign lizzieLet0_4QVal_Bool_8_r = v1a8m_destruct_r;
  
  /* fork (Ty MyBool) : (lizzieLet0_4QVal_Bool_8QVal_Bool,MyBool) > [(lizzieLet0_4QVal_Bool_8QVal_Bool_1,MyBool),
                                                                (lizzieLet0_4QVal_Bool_8QVal_Bool_2,MyBool),
                                                                (lizzieLet0_4QVal_Bool_8QVal_Bool_3,MyBool),
                                                                (lizzieLet0_4QVal_Bool_8QVal_Bool_4,MyBool),
                                                                (lizzieLet0_4QVal_Bool_8QVal_Bool_5,MyBool)] */
  logic [4:0] lizzieLet0_4QVal_Bool_8QVal_Bool_emitted;
  logic [4:0] lizzieLet0_4QVal_Bool_8QVal_Bool_done;
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_1_d = {lizzieLet0_4QVal_Bool_8QVal_Bool_d[1:1],
                                                 (lizzieLet0_4QVal_Bool_8QVal_Bool_d[0] && (! lizzieLet0_4QVal_Bool_8QVal_Bool_emitted[0]))};
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_2_d = {lizzieLet0_4QVal_Bool_8QVal_Bool_d[1:1],
                                                 (lizzieLet0_4QVal_Bool_8QVal_Bool_d[0] && (! lizzieLet0_4QVal_Bool_8QVal_Bool_emitted[1]))};
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_3_d = {lizzieLet0_4QVal_Bool_8QVal_Bool_d[1:1],
                                                 (lizzieLet0_4QVal_Bool_8QVal_Bool_d[0] && (! lizzieLet0_4QVal_Bool_8QVal_Bool_emitted[2]))};
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_4_d = {lizzieLet0_4QVal_Bool_8QVal_Bool_d[1:1],
                                                 (lizzieLet0_4QVal_Bool_8QVal_Bool_d[0] && (! lizzieLet0_4QVal_Bool_8QVal_Bool_emitted[3]))};
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_5_d = {lizzieLet0_4QVal_Bool_8QVal_Bool_d[1:1],
                                                 (lizzieLet0_4QVal_Bool_8QVal_Bool_d[0] && (! lizzieLet0_4QVal_Bool_8QVal_Bool_emitted[4]))};
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_done = (lizzieLet0_4QVal_Bool_8QVal_Bool_emitted | ({lizzieLet0_4QVal_Bool_8QVal_Bool_5_d[0],
                                                                                               lizzieLet0_4QVal_Bool_8QVal_Bool_4_d[0],
                                                                                               lizzieLet0_4QVal_Bool_8QVal_Bool_3_d[0],
                                                                                               lizzieLet0_4QVal_Bool_8QVal_Bool_2_d[0],
                                                                                               lizzieLet0_4QVal_Bool_8QVal_Bool_1_d[0]} & {lizzieLet0_4QVal_Bool_8QVal_Bool_5_r,
                                                                                                                                           lizzieLet0_4QVal_Bool_8QVal_Bool_4_r,
                                                                                                                                           lizzieLet0_4QVal_Bool_8QVal_Bool_3_r,
                                                                                                                                           lizzieLet0_4QVal_Bool_8QVal_Bool_2_r,
                                                                                                                                           lizzieLet0_4QVal_Bool_8QVal_Bool_1_r}));
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_r = (& lizzieLet0_4QVal_Bool_8QVal_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_8QVal_Bool_emitted <= 5'd0;
    else
      lizzieLet0_4QVal_Bool_8QVal_Bool_emitted <= (lizzieLet0_4QVal_Bool_8QVal_Bool_r ? 5'd0 :
                                                   lizzieLet0_4QVal_Bool_8QVal_Bool_done);
  
  /* demux (Ty MyBool,
       Ty Go) : (lizzieLet0_4QVal_Bool_8QVal_Bool_1,MyBool) (lizzieLet0_4QVal_Bool_3QVal_Bool,Go) > [(lizzieLet0_4QVal_Bool_8QVal_Bool_1MyFalse,Go),
                                                                                                     (lizzieLet0_4QVal_Bool_8QVal_Bool_1MyTrue,Go)] */
  logic [1:0] lizzieLet0_4QVal_Bool_3QVal_Bool_onehotd;
  always_comb
    if ((lizzieLet0_4QVal_Bool_8QVal_Bool_1_d[0] && lizzieLet0_4QVal_Bool_3QVal_Bool_d[0]))
      unique case (lizzieLet0_4QVal_Bool_8QVal_Bool_1_d[1:1])
        1'd0: lizzieLet0_4QVal_Bool_3QVal_Bool_onehotd = 2'd1;
        1'd1: lizzieLet0_4QVal_Bool_3QVal_Bool_onehotd = 2'd2;
        default: lizzieLet0_4QVal_Bool_3QVal_Bool_onehotd = 2'd0;
      endcase
    else lizzieLet0_4QVal_Bool_3QVal_Bool_onehotd = 2'd0;
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_1MyFalse_d = lizzieLet0_4QVal_Bool_3QVal_Bool_onehotd[0];
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_1MyTrue_d = lizzieLet0_4QVal_Bool_3QVal_Bool_onehotd[1];
  assign lizzieLet0_4QVal_Bool_3QVal_Bool_r = (| (lizzieLet0_4QVal_Bool_3QVal_Bool_onehotd & {lizzieLet0_4QVal_Bool_8QVal_Bool_1MyTrue_r,
                                                                                              lizzieLet0_4QVal_Bool_8QVal_Bool_1MyFalse_r}));
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_1_r = lizzieLet0_4QVal_Bool_3QVal_Bool_r;
  
  /* demux (Ty MyBool,
       Ty QTree_Bool) : (lizzieLet0_4QVal_Bool_8QVal_Bool_2,MyBool) (lizzieLet0_4QVal_Bool_4QVal_Bool,QTree_Bool) > [(lizzieLet0_4QVal_Bool_8QVal_Bool_2MyFalse,QTree_Bool),
                                                                                                                     (lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue,QTree_Bool)] */
  logic [1:0] lizzieLet0_4QVal_Bool_4QVal_Bool_onehotd;
  always_comb
    if ((lizzieLet0_4QVal_Bool_8QVal_Bool_2_d[0] && lizzieLet0_4QVal_Bool_4QVal_Bool_d[0]))
      unique case (lizzieLet0_4QVal_Bool_8QVal_Bool_2_d[1:1])
        1'd0: lizzieLet0_4QVal_Bool_4QVal_Bool_onehotd = 2'd1;
        1'd1: lizzieLet0_4QVal_Bool_4QVal_Bool_onehotd = 2'd2;
        default: lizzieLet0_4QVal_Bool_4QVal_Bool_onehotd = 2'd0;
      endcase
    else lizzieLet0_4QVal_Bool_4QVal_Bool_onehotd = 2'd0;
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_2MyFalse_d = {lizzieLet0_4QVal_Bool_4QVal_Bool_d[66:1],
                                                        lizzieLet0_4QVal_Bool_4QVal_Bool_onehotd[0]};
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_d = {lizzieLet0_4QVal_Bool_4QVal_Bool_d[66:1],
                                                       lizzieLet0_4QVal_Bool_4QVal_Bool_onehotd[1]};
  assign lizzieLet0_4QVal_Bool_4QVal_Bool_r = (| (lizzieLet0_4QVal_Bool_4QVal_Bool_onehotd & {lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_r,
                                                                                              lizzieLet0_4QVal_Bool_8QVal_Bool_2MyFalse_r}));
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_2_r = lizzieLet0_4QVal_Bool_4QVal_Bool_r;
  
  /* fork (Ty QTree_Bool) : (lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue,QTree_Bool) > [(lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1,QTree_Bool),
                                                                                (lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2,QTree_Bool)] */
  logic [1:0] lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_emitted;
  logic [1:0] lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_done;
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1_d = {lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_d[66:1],
                                                         (lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_d[0] && (! lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_emitted[0]))};
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2_d = {lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_d[66:1],
                                                         (lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_d[0] && (! lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_emitted[1]))};
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_done = (lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_emitted | ({lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2_d[0],
                                                                                                               lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1_d[0]} & {lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2_r,
                                                                                                                                                                   lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1_r}));
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_r = (& lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_emitted <= 2'd0;
    else
      lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_emitted <= (lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_r ? 2'd0 :
                                                           lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_done);
  
  /* demux (Ty QTree_Bool,
       Ty Go) : (lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1,QTree_Bool) (lizzieLet0_4QVal_Bool_8QVal_Bool_1MyTrue,Go) > [(lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNone_Bool,Go),
                                                                                                                         (lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QVal_Bool,Go),
                                                                                                                         (lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNode_Bool,Go),
                                                                                                                         (lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QError_Bool,Go)] */
  logic [3:0] lizzieLet0_4QVal_Bool_8QVal_Bool_1MyTrue_onehotd;
  always_comb
    if ((lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1_d[0] && lizzieLet0_4QVal_Bool_8QVal_Bool_1MyTrue_d[0]))
      unique case (lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1_d[2:1])
        2'd0: lizzieLet0_4QVal_Bool_8QVal_Bool_1MyTrue_onehotd = 4'd1;
        2'd1: lizzieLet0_4QVal_Bool_8QVal_Bool_1MyTrue_onehotd = 4'd2;
        2'd2: lizzieLet0_4QVal_Bool_8QVal_Bool_1MyTrue_onehotd = 4'd4;
        2'd3: lizzieLet0_4QVal_Bool_8QVal_Bool_1MyTrue_onehotd = 4'd8;
        default: lizzieLet0_4QVal_Bool_8QVal_Bool_1MyTrue_onehotd = 4'd0;
      endcase
    else lizzieLet0_4QVal_Bool_8QVal_Bool_1MyTrue_onehotd = 4'd0;
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNone_Bool_d = lizzieLet0_4QVal_Bool_8QVal_Bool_1MyTrue_onehotd[0];
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QVal_Bool_d = lizzieLet0_4QVal_Bool_8QVal_Bool_1MyTrue_onehotd[1];
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNode_Bool_d = lizzieLet0_4QVal_Bool_8QVal_Bool_1MyTrue_onehotd[2];
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QError_Bool_d = lizzieLet0_4QVal_Bool_8QVal_Bool_1MyTrue_onehotd[3];
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_1MyTrue_r = (| (lizzieLet0_4QVal_Bool_8QVal_Bool_1MyTrue_onehotd & {lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QError_Bool_r,
                                                                                                              lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNode_Bool_r,
                                                                                                              lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QVal_Bool_r,
                                                                                                              lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNone_Bool_r}));
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1_r = lizzieLet0_4QVal_Bool_8QVal_Bool_1MyTrue_r;
  
  /* fork (Ty Go) : (lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QError_Bool,Go) > [(lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QError_Bool_1,Go),
                                                                             (lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QError_Bool_2,Go)] */
  logic [1:0] lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QError_Bool_emitted;
  logic [1:0] lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QError_Bool_done;
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QError_Bool_1_d = (lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QError_Bool_d[0] && (! lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QError_Bool_emitted[0]));
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QError_Bool_2_d = (lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QError_Bool_d[0] && (! lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QError_Bool_emitted[1]));
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QError_Bool_done = (lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QError_Bool_emitted | ({lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QError_Bool_2_d[0],
                                                                                                                                         lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QError_Bool_1_d[0]} & {lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QError_Bool_2_r,
                                                                                                                                                                                                          lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QError_Bool_1_r}));
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QError_Bool_r = (& lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QError_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QError_Bool_emitted <= 2'd0;
    else
      lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QError_Bool_emitted <= (lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QError_Bool_r ? 2'd0 :
                                                                        lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QError_Bool_done);
  
  /* dcon (Ty QTree_Bool,
      Dcon QError_Bool) : [(lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QError_Bool_1,Go)] > (lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QError_Bool_1QError_Bool,QTree_Bool) */
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QError_Bool_1QError_Bool_d = QError_Bool_dc((& {lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QError_Bool_1_d[0]}), lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QError_Bool_1_d);
  assign {lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QError_Bool_1_r} = {1 {(lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QError_Bool_1QError_Bool_r && lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QError_Bool_1QError_Bool_d[0])}};
  
  /* buf (Ty QTree_Bool) : (lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QError_Bool_1QError_Bool,QTree_Bool) > (lizzieLet29_1_argbuf,QTree_Bool) */
  QTree_Bool_t lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QError_Bool_1QError_Bool_bufchan_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QError_Bool_1QError_Bool_bufchan_r;
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QError_Bool_1QError_Bool_r = ((! lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QError_Bool_1QError_Bool_bufchan_d[0]) || lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QError_Bool_1QError_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QError_Bool_1QError_Bool_bufchan_d <= {66'd0,
                                                                                       1'd0};
    else
      if (lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QError_Bool_1QError_Bool_r)
        lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QError_Bool_1QError_Bool_bufchan_d <= lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QError_Bool_1QError_Bool_d;
  QTree_Bool_t lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QError_Bool_1QError_Bool_bufchan_buf;
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QError_Bool_1QError_Bool_bufchan_r = (! lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QError_Bool_1QError_Bool_bufchan_buf[0]);
  assign lizzieLet29_1_argbuf_d = (lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QError_Bool_1QError_Bool_bufchan_buf[0] ? lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QError_Bool_1QError_Bool_bufchan_buf :
                                   lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QError_Bool_1QError_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QError_Bool_1QError_Bool_bufchan_buf <= {66'd0,
                                                                                         1'd0};
    else
      if ((lizzieLet29_1_argbuf_r && lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QError_Bool_1QError_Bool_bufchan_buf[0]))
        lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QError_Bool_1QError_Bool_bufchan_buf <= {66'd0,
                                                                                           1'd0};
      else if (((! lizzieLet29_1_argbuf_r) && (! lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QError_Bool_1QError_Bool_bufchan_buf[0])))
        lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QError_Bool_1QError_Bool_bufchan_buf <= lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QError_Bool_1QError_Bool_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QError_Bool_2,Go) > (lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QError_Bool_2_argbuf,Go) */
  Go_t lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QError_Bool_2_bufchan_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QError_Bool_2_bufchan_r;
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QError_Bool_2_r = ((! lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QError_Bool_2_bufchan_d[0]) || lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QError_Bool_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QError_Bool_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QError_Bool_2_r)
        lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QError_Bool_2_bufchan_d <= lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QError_Bool_2_d;
  Go_t lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QError_Bool_2_bufchan_buf;
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QError_Bool_2_bufchan_r = (! lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QError_Bool_2_bufchan_buf[0]);
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QError_Bool_2_argbuf_d = (lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QError_Bool_2_bufchan_buf[0] ? lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QError_Bool_2_bufchan_buf :
                                                                             lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QError_Bool_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QError_Bool_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QError_Bool_2_argbuf_r && lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QError_Bool_2_bufchan_buf[0]))
        lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QError_Bool_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QError_Bool_2_argbuf_r) && (! lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QError_Bool_2_bufchan_buf[0])))
        lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QError_Bool_2_bufchan_buf <= lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QError_Bool_2_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNode_Bool,Go) > [(lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNode_Bool_1,Go),
                                                                            (lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNode_Bool_2,Go)] */
  logic [1:0] lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNode_Bool_emitted;
  logic [1:0] lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNode_Bool_done;
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNode_Bool_1_d = (lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNode_Bool_d[0] && (! lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNode_Bool_emitted[0]));
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNode_Bool_2_d = (lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNode_Bool_d[0] && (! lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNode_Bool_emitted[1]));
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNode_Bool_done = (lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNode_Bool_emitted | ({lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNode_Bool_2_d[0],
                                                                                                                                       lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNode_Bool_1_d[0]} & {lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNode_Bool_2_r,
                                                                                                                                                                                                       lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNode_Bool_1_r}));
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNode_Bool_r = (& lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNode_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNode_Bool_emitted <= 2'd0;
    else
      lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNode_Bool_emitted <= (lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNode_Bool_r ? 2'd0 :
                                                                       lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNode_Bool_done);
  
  /* dcon (Ty QTree_Bool,
      Dcon QError_Bool) : [(lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNode_Bool_1,Go)] > (lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNode_Bool_1QError_Bool,QTree_Bool) */
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNode_Bool_1QError_Bool_d = QError_Bool_dc((& {lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNode_Bool_1_d[0]}), lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNode_Bool_1_d);
  assign {lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNode_Bool_1_r} = {1 {(lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNode_Bool_1QError_Bool_r && lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNode_Bool_1QError_Bool_d[0])}};
  
  /* buf (Ty QTree_Bool) : (lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNode_Bool_1QError_Bool,QTree_Bool) > (lizzieLet28_1_argbuf,QTree_Bool) */
  QTree_Bool_t lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNode_Bool_1QError_Bool_bufchan_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNode_Bool_1QError_Bool_bufchan_r;
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNode_Bool_1QError_Bool_r = ((! lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNode_Bool_1QError_Bool_bufchan_d[0]) || lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNode_Bool_1QError_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNode_Bool_1QError_Bool_bufchan_d <= {66'd0,
                                                                                      1'd0};
    else
      if (lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNode_Bool_1QError_Bool_r)
        lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNode_Bool_1QError_Bool_bufchan_d <= lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNode_Bool_1QError_Bool_d;
  QTree_Bool_t lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNode_Bool_1QError_Bool_bufchan_buf;
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNode_Bool_1QError_Bool_bufchan_r = (! lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNode_Bool_1QError_Bool_bufchan_buf[0]);
  assign lizzieLet28_1_argbuf_d = (lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNode_Bool_1QError_Bool_bufchan_buf[0] ? lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNode_Bool_1QError_Bool_bufchan_buf :
                                   lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNode_Bool_1QError_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNode_Bool_1QError_Bool_bufchan_buf <= {66'd0,
                                                                                        1'd0};
    else
      if ((lizzieLet28_1_argbuf_r && lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNode_Bool_1QError_Bool_bufchan_buf[0]))
        lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNode_Bool_1QError_Bool_bufchan_buf <= {66'd0,
                                                                                          1'd0};
      else if (((! lizzieLet28_1_argbuf_r) && (! lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNode_Bool_1QError_Bool_bufchan_buf[0])))
        lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNode_Bool_1QError_Bool_bufchan_buf <= lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNode_Bool_1QError_Bool_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNode_Bool_2,Go) > (lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNode_Bool_2_argbuf,Go) */
  Go_t lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNode_Bool_2_bufchan_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNode_Bool_2_bufchan_r;
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNode_Bool_2_r = ((! lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNode_Bool_2_bufchan_d[0]) || lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNode_Bool_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNode_Bool_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNode_Bool_2_r)
        lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNode_Bool_2_bufchan_d <= lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNode_Bool_2_d;
  Go_t lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNode_Bool_2_bufchan_buf;
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNode_Bool_2_bufchan_r = (! lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNode_Bool_2_bufchan_buf[0]);
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNode_Bool_2_argbuf_d = (lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNode_Bool_2_bufchan_buf[0] ? lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNode_Bool_2_bufchan_buf :
                                                                            lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNode_Bool_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNode_Bool_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNode_Bool_2_argbuf_r && lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNode_Bool_2_bufchan_buf[0]))
        lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNode_Bool_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNode_Bool_2_argbuf_r) && (! lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNode_Bool_2_bufchan_buf[0])))
        lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNode_Bool_2_bufchan_buf <= lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNode_Bool_2_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNone_Bool,Go) > [(lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNone_Bool_1,Go),
                                                                            (lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNone_Bool_2,Go)] */
  logic [1:0] lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNone_Bool_emitted;
  logic [1:0] lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNone_Bool_done;
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNone_Bool_1_d = (lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNone_Bool_d[0] && (! lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNone_Bool_emitted[0]));
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNone_Bool_2_d = (lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNone_Bool_d[0] && (! lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNone_Bool_emitted[1]));
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNone_Bool_done = (lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNone_Bool_emitted | ({lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNone_Bool_2_d[0],
                                                                                                                                       lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNone_Bool_1_d[0]} & {lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNone_Bool_2_r,
                                                                                                                                                                                                       lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNone_Bool_1_r}));
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNone_Bool_r = (& lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNone_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNone_Bool_emitted <= 2'd0;
    else
      lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNone_Bool_emitted <= (lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNone_Bool_r ? 2'd0 :
                                                                       lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNone_Bool_done);
  
  /* buf (Ty Go) : (lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNone_Bool_1,Go) > (lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNone_Bool_1_argbuf,Go) */
  Go_t lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNone_Bool_1_bufchan_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNone_Bool_1_bufchan_r;
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNone_Bool_1_r = ((! lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNone_Bool_1_bufchan_d[0]) || lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNone_Bool_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNone_Bool_1_bufchan_d <= 1'd0;
    else
      if (lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNone_Bool_1_r)
        lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNone_Bool_1_bufchan_d <= lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNone_Bool_1_d;
  Go_t lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNone_Bool_1_bufchan_buf;
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNone_Bool_1_bufchan_r = (! lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNone_Bool_1_bufchan_buf[0]);
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNone_Bool_1_argbuf_d = (lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNone_Bool_1_bufchan_buf[0] ? lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNone_Bool_1_bufchan_buf :
                                                                            lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNone_Bool_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNone_Bool_1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNone_Bool_1_argbuf_r && lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNone_Bool_1_bufchan_buf[0]))
        lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNone_Bool_1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNone_Bool_1_argbuf_r) && (! lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNone_Bool_1_bufchan_buf[0])))
        lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNone_Bool_1_bufchan_buf <= lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNone_Bool_1_bufchan_d;
  
  /* dcon (Ty TupGo,
      Dcon TupGo) : [(lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNone_Bool_1_argbuf,Go)] > (lvlrf2-0TupGo9,TupGo) */
  assign \lvlrf2-0TupGo9_d  = TupGo_dc((& {lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNone_Bool_1_argbuf_d[0]}), lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNone_Bool_1_argbuf_d);
  assign {lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNone_Bool_1_argbuf_r} = {1 {(\lvlrf2-0TupGo9_r  && \lvlrf2-0TupGo9_d [0])}};
  
  /* buf (Ty Go) : (lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNone_Bool_2,Go) > (lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNone_Bool_2_argbuf,Go) */
  Go_t lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNone_Bool_2_bufchan_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNone_Bool_2_bufchan_r;
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNone_Bool_2_r = ((! lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNone_Bool_2_bufchan_d[0]) || lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNone_Bool_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNone_Bool_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNone_Bool_2_r)
        lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNone_Bool_2_bufchan_d <= lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNone_Bool_2_d;
  Go_t lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNone_Bool_2_bufchan_buf;
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNone_Bool_2_bufchan_r = (! lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNone_Bool_2_bufchan_buf[0]);
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNone_Bool_2_argbuf_d = (lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNone_Bool_2_bufchan_buf[0] ? lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNone_Bool_2_bufchan_buf :
                                                                            lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNone_Bool_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNone_Bool_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNone_Bool_2_argbuf_r && lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNone_Bool_2_bufchan_buf[0]))
        lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNone_Bool_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNone_Bool_2_argbuf_r) && (! lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNone_Bool_2_bufchan_buf[0])))
        lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNone_Bool_2_bufchan_buf <= lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QNone_Bool_2_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QVal_Bool,Go) > [(lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QVal_Bool_1,Go),
                                                                           (lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QVal_Bool_2,Go)] */
  logic [1:0] lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QVal_Bool_emitted;
  logic [1:0] lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QVal_Bool_done;
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QVal_Bool_1_d = (lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QVal_Bool_d[0] && (! lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QVal_Bool_emitted[0]));
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QVal_Bool_2_d = (lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QVal_Bool_d[0] && (! lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QVal_Bool_emitted[1]));
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QVal_Bool_done = (lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QVal_Bool_emitted | ({lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QVal_Bool_2_d[0],
                                                                                                                                     lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QVal_Bool_1_d[0]} & {lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QVal_Bool_2_r,
                                                                                                                                                                                                    lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QVal_Bool_1_r}));
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QVal_Bool_r = (& lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QVal_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QVal_Bool_emitted <= 2'd0;
    else
      lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QVal_Bool_emitted <= (lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QVal_Bool_r ? 2'd0 :
                                                                      lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QVal_Bool_done);
  
  /* buf (Ty Go) : (lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QVal_Bool_1,Go) > (lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QVal_Bool_1_argbuf,Go) */
  Go_t lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QVal_Bool_1_bufchan_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QVal_Bool_1_bufchan_r;
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QVal_Bool_1_r = ((! lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QVal_Bool_1_bufchan_d[0]) || lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QVal_Bool_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QVal_Bool_1_bufchan_d <= 1'd0;
    else
      if (lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QVal_Bool_1_r)
        lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QVal_Bool_1_bufchan_d <= lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QVal_Bool_1_d;
  Go_t lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QVal_Bool_1_bufchan_buf;
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QVal_Bool_1_bufchan_r = (! lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QVal_Bool_1_bufchan_buf[0]);
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QVal_Bool_1_argbuf_d = (lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QVal_Bool_1_bufchan_buf[0] ? lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QVal_Bool_1_bufchan_buf :
                                                                           lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QVal_Bool_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QVal_Bool_1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QVal_Bool_1_argbuf_r && lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QVal_Bool_1_bufchan_buf[0]))
        lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QVal_Bool_1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QVal_Bool_1_argbuf_r) && (! lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QVal_Bool_1_bufchan_buf[0])))
        lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QVal_Bool_1_bufchan_buf <= lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QVal_Bool_1_bufchan_d;
  
  /* dcon (Ty TupGo,
      Dcon TupGo) : [(lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QVal_Bool_1_argbuf,Go)] > (lvlrf2-0TupGo10,TupGo) */
  assign \lvlrf2-0TupGo10_d  = TupGo_dc((& {lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QVal_Bool_1_argbuf_d[0]}), lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QVal_Bool_1_argbuf_d);
  assign {lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QVal_Bool_1_argbuf_r} = {1 {(\lvlrf2-0TupGo10_r  && \lvlrf2-0TupGo10_d [0])}};
  
  /* buf (Ty Go) : (lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QVal_Bool_2,Go) > (lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QVal_Bool_2_argbuf,Go) */
  Go_t lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QVal_Bool_2_bufchan_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QVal_Bool_2_bufchan_r;
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QVal_Bool_2_r = ((! lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QVal_Bool_2_bufchan_d[0]) || lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QVal_Bool_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QVal_Bool_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QVal_Bool_2_r)
        lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QVal_Bool_2_bufchan_d <= lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QVal_Bool_2_d;
  Go_t lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QVal_Bool_2_bufchan_buf;
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QVal_Bool_2_bufchan_r = (! lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QVal_Bool_2_bufchan_buf[0]);
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QVal_Bool_2_argbuf_d = (lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QVal_Bool_2_bufchan_buf[0] ? lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QVal_Bool_2_bufchan_buf :
                                                                           lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QVal_Bool_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QVal_Bool_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QVal_Bool_2_argbuf_r && lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QVal_Bool_2_bufchan_buf[0]))
        lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QVal_Bool_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QVal_Bool_2_argbuf_r) && (! lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QVal_Bool_2_bufchan_buf[0])))
        lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QVal_Bool_2_bufchan_buf <= lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_1QVal_Bool_2_bufchan_d;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_CTf) : (lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2,QTree_Bool) (lizzieLet0_4QVal_Bool_8QVal_Bool_4MyTrue,Pointer_CTf) > [(lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QNone_Bool,Pointer_CTf),
                                                                                                                                           (lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QVal_Bool,Pointer_CTf),
                                                                                                                                           (lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QNode_Bool,Pointer_CTf),
                                                                                                                                           (lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QError_Bool,Pointer_CTf)] */
  logic [3:0] lizzieLet0_4QVal_Bool_8QVal_Bool_4MyTrue_onehotd;
  always_comb
    if ((lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2_d[0] && lizzieLet0_4QVal_Bool_8QVal_Bool_4MyTrue_d[0]))
      unique case (lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2_d[2:1])
        2'd0: lizzieLet0_4QVal_Bool_8QVal_Bool_4MyTrue_onehotd = 4'd1;
        2'd1: lizzieLet0_4QVal_Bool_8QVal_Bool_4MyTrue_onehotd = 4'd2;
        2'd2: lizzieLet0_4QVal_Bool_8QVal_Bool_4MyTrue_onehotd = 4'd4;
        2'd3: lizzieLet0_4QVal_Bool_8QVal_Bool_4MyTrue_onehotd = 4'd8;
        default: lizzieLet0_4QVal_Bool_8QVal_Bool_4MyTrue_onehotd = 4'd0;
      endcase
    else lizzieLet0_4QVal_Bool_8QVal_Bool_4MyTrue_onehotd = 4'd0;
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QNone_Bool_d = {lizzieLet0_4QVal_Bool_8QVal_Bool_4MyTrue_d[16:1],
                                                                   lizzieLet0_4QVal_Bool_8QVal_Bool_4MyTrue_onehotd[0]};
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QVal_Bool_d = {lizzieLet0_4QVal_Bool_8QVal_Bool_4MyTrue_d[16:1],
                                                                  lizzieLet0_4QVal_Bool_8QVal_Bool_4MyTrue_onehotd[1]};
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QNode_Bool_d = {lizzieLet0_4QVal_Bool_8QVal_Bool_4MyTrue_d[16:1],
                                                                   lizzieLet0_4QVal_Bool_8QVal_Bool_4MyTrue_onehotd[2]};
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QError_Bool_d = {lizzieLet0_4QVal_Bool_8QVal_Bool_4MyTrue_d[16:1],
                                                                    lizzieLet0_4QVal_Bool_8QVal_Bool_4MyTrue_onehotd[3]};
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_4MyTrue_r = (| (lizzieLet0_4QVal_Bool_8QVal_Bool_4MyTrue_onehotd & {lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QError_Bool_r,
                                                                                                              lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QNode_Bool_r,
                                                                                                              lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QVal_Bool_r,
                                                                                                              lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QNone_Bool_r}));
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2_r = lizzieLet0_4QVal_Bool_8QVal_Bool_4MyTrue_r;
  
  /* buf (Ty Pointer_CTf) : (lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QError_Bool,Pointer_CTf) > (lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QError_Bool_1_argbuf,Pointer_CTf) */
  Pointer_CTf_t lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QError_Bool_bufchan_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QError_Bool_bufchan_r;
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QError_Bool_r = ((! lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QError_Bool_bufchan_d[0]) || lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QError_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QError_Bool_bufchan_d <= {16'd0,
                                                                          1'd0};
    else
      if (lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QError_Bool_r)
        lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QError_Bool_bufchan_d <= lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QError_Bool_d;
  Pointer_CTf_t lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QError_Bool_bufchan_buf;
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QError_Bool_bufchan_r = (! lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QError_Bool_bufchan_buf[0]);
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QError_Bool_1_argbuf_d = (lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QError_Bool_bufchan_buf[0] ? lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QError_Bool_bufchan_buf :
                                                                             lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QError_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QError_Bool_bufchan_buf <= {16'd0,
                                                                            1'd0};
    else
      if ((lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QError_Bool_1_argbuf_r && lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QError_Bool_bufchan_buf[0]))
        lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QError_Bool_bufchan_buf <= {16'd0,
                                                                              1'd0};
      else if (((! lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QError_Bool_1_argbuf_r) && (! lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QError_Bool_bufchan_buf[0])))
        lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QError_Bool_bufchan_buf <= lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QError_Bool_bufchan_d;
  
  /* buf (Ty Pointer_CTf) : (lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QNode_Bool,Pointer_CTf) > (lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QNode_Bool_1_argbuf,Pointer_CTf) */
  Pointer_CTf_t lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QNode_Bool_bufchan_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QNode_Bool_bufchan_r;
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QNode_Bool_r = ((! lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QNode_Bool_bufchan_d[0]) || lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QNode_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QNode_Bool_bufchan_d <= {16'd0,
                                                                         1'd0};
    else
      if (lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QNode_Bool_r)
        lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QNode_Bool_bufchan_d <= lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QNode_Bool_d;
  Pointer_CTf_t lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QNode_Bool_bufchan_buf;
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QNode_Bool_bufchan_r = (! lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QNode_Bool_bufchan_buf[0]);
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QNode_Bool_1_argbuf_d = (lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QNode_Bool_bufchan_buf[0] ? lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QNode_Bool_bufchan_buf :
                                                                            lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QNode_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QNode_Bool_bufchan_buf <= {16'd0,
                                                                           1'd0};
    else
      if ((lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QNode_Bool_1_argbuf_r && lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QNode_Bool_bufchan_buf[0]))
        lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QNode_Bool_bufchan_buf <= {16'd0,
                                                                             1'd0};
      else if (((! lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QNode_Bool_1_argbuf_r) && (! lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QNode_Bool_bufchan_buf[0])))
        lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QNode_Bool_bufchan_buf <= lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QNode_Bool_bufchan_d;
  
  /* buf (Ty Pointer_CTf) : (lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QNone_Bool,Pointer_CTf) > (lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QNone_Bool_1_argbuf,Pointer_CTf) */
  Pointer_CTf_t lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QNone_Bool_bufchan_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QNone_Bool_bufchan_r;
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QNone_Bool_r = ((! lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QNone_Bool_bufchan_d[0]) || lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QNone_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QNone_Bool_bufchan_d <= {16'd0,
                                                                         1'd0};
    else
      if (lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QNone_Bool_r)
        lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QNone_Bool_bufchan_d <= lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QNone_Bool_d;
  Pointer_CTf_t lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QNone_Bool_bufchan_buf;
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QNone_Bool_bufchan_r = (! lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QNone_Bool_bufchan_buf[0]);
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QNone_Bool_1_argbuf_d = (lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QNone_Bool_bufchan_buf[0] ? lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QNone_Bool_bufchan_buf :
                                                                            lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QNone_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QNone_Bool_bufchan_buf <= {16'd0,
                                                                           1'd0};
    else
      if ((lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QNone_Bool_1_argbuf_r && lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QNone_Bool_bufchan_buf[0]))
        lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QNone_Bool_bufchan_buf <= {16'd0,
                                                                             1'd0};
      else if (((! lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QNone_Bool_1_argbuf_r) && (! lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QNone_Bool_bufchan_buf[0])))
        lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QNone_Bool_bufchan_buf <= lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QNone_Bool_bufchan_d;
  
  /* buf (Ty Pointer_CTf) : (lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QVal_Bool,Pointer_CTf) > (lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QVal_Bool_1_argbuf,Pointer_CTf) */
  Pointer_CTf_t lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QVal_Bool_bufchan_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QVal_Bool_bufchan_r;
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QVal_Bool_r = ((! lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QVal_Bool_bufchan_d[0]) || lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QVal_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QVal_Bool_bufchan_d <= {16'd0,
                                                                        1'd0};
    else
      if (lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QVal_Bool_r)
        lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QVal_Bool_bufchan_d <= lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QVal_Bool_d;
  Pointer_CTf_t lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QVal_Bool_bufchan_buf;
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QVal_Bool_bufchan_r = (! lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QVal_Bool_bufchan_buf[0]);
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QVal_Bool_1_argbuf_d = (lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QVal_Bool_bufchan_buf[0] ? lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QVal_Bool_bufchan_buf :
                                                                           lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QVal_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QVal_Bool_bufchan_buf <= {16'd0,
                                                                          1'd0};
    else
      if ((lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QVal_Bool_1_argbuf_r && lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QVal_Bool_bufchan_buf[0]))
        lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QVal_Bool_bufchan_buf <= {16'd0,
                                                                            1'd0};
      else if (((! lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QVal_Bool_1_argbuf_r) && (! lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QVal_Bool_bufchan_buf[0])))
        lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QVal_Bool_bufchan_buf <= lizzieLet0_4QVal_Bool_8QVal_Bool_2MyTrue_2QVal_Bool_bufchan_d;
  
  /* demux (Ty MyBool,
       Ty Pointer_QTree_Bool) : (lizzieLet0_4QVal_Bool_8QVal_Bool_3,MyBool) (lizzieLet0_4QVal_Bool_6QVal_Bool,Pointer_QTree_Bool) > [(lizzieLet0_4QVal_Bool_8QVal_Bool_3MyFalse,Pointer_QTree_Bool),
                                                                                                                                     (_52,Pointer_QTree_Bool)] */
  logic [1:0] lizzieLet0_4QVal_Bool_6QVal_Bool_onehotd;
  always_comb
    if ((lizzieLet0_4QVal_Bool_8QVal_Bool_3_d[0] && lizzieLet0_4QVal_Bool_6QVal_Bool_d[0]))
      unique case (lizzieLet0_4QVal_Bool_8QVal_Bool_3_d[1:1])
        1'd0: lizzieLet0_4QVal_Bool_6QVal_Bool_onehotd = 2'd1;
        1'd1: lizzieLet0_4QVal_Bool_6QVal_Bool_onehotd = 2'd2;
        default: lizzieLet0_4QVal_Bool_6QVal_Bool_onehotd = 2'd0;
      endcase
    else lizzieLet0_4QVal_Bool_6QVal_Bool_onehotd = 2'd0;
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_3MyFalse_d = {lizzieLet0_4QVal_Bool_6QVal_Bool_d[16:1],
                                                        lizzieLet0_4QVal_Bool_6QVal_Bool_onehotd[0]};
  assign _52_d = {lizzieLet0_4QVal_Bool_6QVal_Bool_d[16:1],
                  lizzieLet0_4QVal_Bool_6QVal_Bool_onehotd[1]};
  assign lizzieLet0_4QVal_Bool_6QVal_Bool_r = (| (lizzieLet0_4QVal_Bool_6QVal_Bool_onehotd & {_52_r,
                                                                                              lizzieLet0_4QVal_Bool_8QVal_Bool_3MyFalse_r}));
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_3_r = lizzieLet0_4QVal_Bool_6QVal_Bool_r;
  
  /* demux (Ty MyBool,
       Ty Pointer_CTf) : (lizzieLet0_4QVal_Bool_8QVal_Bool_4,MyBool) (lizzieLet0_4QVal_Bool_7QVal_Bool,Pointer_CTf) > [(lizzieLet0_4QVal_Bool_8QVal_Bool_4MyFalse,Pointer_CTf),
                                                                                                                       (lizzieLet0_4QVal_Bool_8QVal_Bool_4MyTrue,Pointer_CTf)] */
  logic [1:0] lizzieLet0_4QVal_Bool_7QVal_Bool_onehotd;
  always_comb
    if ((lizzieLet0_4QVal_Bool_8QVal_Bool_4_d[0] && lizzieLet0_4QVal_Bool_7QVal_Bool_d[0]))
      unique case (lizzieLet0_4QVal_Bool_8QVal_Bool_4_d[1:1])
        1'd0: lizzieLet0_4QVal_Bool_7QVal_Bool_onehotd = 2'd1;
        1'd1: lizzieLet0_4QVal_Bool_7QVal_Bool_onehotd = 2'd2;
        default: lizzieLet0_4QVal_Bool_7QVal_Bool_onehotd = 2'd0;
      endcase
    else lizzieLet0_4QVal_Bool_7QVal_Bool_onehotd = 2'd0;
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_4MyFalse_d = {lizzieLet0_4QVal_Bool_7QVal_Bool_d[16:1],
                                                        lizzieLet0_4QVal_Bool_7QVal_Bool_onehotd[0]};
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_4MyTrue_d = {lizzieLet0_4QVal_Bool_7QVal_Bool_d[16:1],
                                                       lizzieLet0_4QVal_Bool_7QVal_Bool_onehotd[1]};
  assign lizzieLet0_4QVal_Bool_7QVal_Bool_r = (| (lizzieLet0_4QVal_Bool_7QVal_Bool_onehotd & {lizzieLet0_4QVal_Bool_8QVal_Bool_4MyTrue_r,
                                                                                              lizzieLet0_4QVal_Bool_8QVal_Bool_4MyFalse_r}));
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_4_r = lizzieLet0_4QVal_Bool_7QVal_Bool_r;
  
  /* demux (Ty MyBool,
       Ty MyBool) : (lizzieLet0_4QVal_Bool_8QVal_Bool_5,MyBool) (va8s_destruct,MyBool) > [(lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse,MyBool),
                                                                                          (_51,MyBool)] */
  logic [1:0] va8s_destruct_onehotd;
  always_comb
    if ((lizzieLet0_4QVal_Bool_8QVal_Bool_5_d[0] && va8s_destruct_d[0]))
      unique case (lizzieLet0_4QVal_Bool_8QVal_Bool_5_d[1:1])
        1'd0: va8s_destruct_onehotd = 2'd1;
        1'd1: va8s_destruct_onehotd = 2'd2;
        default: va8s_destruct_onehotd = 2'd0;
      endcase
    else va8s_destruct_onehotd = 2'd0;
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_d = {va8s_destruct_d[1:1],
                                                        va8s_destruct_onehotd[0]};
  assign _51_d = {va8s_destruct_d[1:1], va8s_destruct_onehotd[1]};
  assign va8s_destruct_r = (| (va8s_destruct_onehotd & {_51_r,
                                                        lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_r}));
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_5_r = va8s_destruct_r;
  
  /* fork (Ty MyBool) : (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse,MyBool) > [(lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_1,MyBool),
                                                                         (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2,MyBool),
                                                                         (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_3,MyBool),
                                                                         (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_4,MyBool)] */
  logic [3:0] lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_emitted;
  logic [3:0] lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_done;
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_1_d = {lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_d[1:1],
                                                          (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_d[0] && (! lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_emitted[0]))};
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2_d = {lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_d[1:1],
                                                          (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_d[0] && (! lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_emitted[1]))};
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_3_d = {lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_d[1:1],
                                                          (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_d[0] && (! lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_emitted[2]))};
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_4_d = {lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_d[1:1],
                                                          (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_d[0] && (! lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_emitted[3]))};
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_done = (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_emitted | ({lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_4_d[0],
                                                                                                                 lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_3_d[0],
                                                                                                                 lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2_d[0],
                                                                                                                 lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_1_d[0]} & {lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_4_r,
                                                                                                                                                                      lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_3_r,
                                                                                                                                                                      lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2_r,
                                                                                                                                                                      lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_1_r}));
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_r = (& lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_emitted <= 4'd0;
    else
      lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_emitted <= (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_r ? 4'd0 :
                                                            lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_done);
  
  /* demux (Ty MyBool,
       Ty Go) : (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_1,MyBool) (lizzieLet0_4QVal_Bool_8QVal_Bool_1MyFalse,Go) > [(lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_1MyFalse,Go),
                                                                                                                       (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_1MyTrue,Go)] */
  logic [1:0] lizzieLet0_4QVal_Bool_8QVal_Bool_1MyFalse_onehotd;
  always_comb
    if ((lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_1_d[0] && lizzieLet0_4QVal_Bool_8QVal_Bool_1MyFalse_d[0]))
      unique case (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_1_d[1:1])
        1'd0: lizzieLet0_4QVal_Bool_8QVal_Bool_1MyFalse_onehotd = 2'd1;
        1'd1: lizzieLet0_4QVal_Bool_8QVal_Bool_1MyFalse_onehotd = 2'd2;
        default: lizzieLet0_4QVal_Bool_8QVal_Bool_1MyFalse_onehotd = 2'd0;
      endcase
    else lizzieLet0_4QVal_Bool_8QVal_Bool_1MyFalse_onehotd = 2'd0;
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_1MyFalse_d = lizzieLet0_4QVal_Bool_8QVal_Bool_1MyFalse_onehotd[0];
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_1MyTrue_d = lizzieLet0_4QVal_Bool_8QVal_Bool_1MyFalse_onehotd[1];
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_1MyFalse_r = (| (lizzieLet0_4QVal_Bool_8QVal_Bool_1MyFalse_onehotd & {lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_1MyTrue_r,
                                                                                                                lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_1MyFalse_r}));
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_1_r = lizzieLet0_4QVal_Bool_8QVal_Bool_1MyFalse_r;
  
  /* buf (Ty Go) : (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_1MyFalse,Go) > (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_1MyFalse_1_argbuf,Go) */
  Go_t lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_1MyFalse_bufchan_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_1MyFalse_bufchan_r;
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_1MyFalse_r = ((! lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_1MyFalse_bufchan_d[0]) || lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_1MyFalse_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_1MyFalse_bufchan_d <= 1'd0;
    else
      if (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_1MyFalse_r)
        lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_1MyFalse_bufchan_d <= lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_1MyFalse_d;
  Go_t lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_1MyFalse_bufchan_buf;
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_1MyFalse_bufchan_r = (! lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_1MyFalse_bufchan_buf[0]);
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_1MyFalse_1_argbuf_d = (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_1MyFalse_bufchan_buf[0] ? lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_1MyFalse_bufchan_buf :
                                                                          lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_1MyFalse_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_1MyFalse_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_1MyFalse_1_argbuf_r && lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_1MyFalse_bufchan_buf[0]))
        lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_1MyFalse_bufchan_buf <= 1'd0;
      else if (((! lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_1MyFalse_1_argbuf_r) && (! lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_1MyFalse_bufchan_buf[0])))
        lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_1MyFalse_bufchan_buf <= lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_1MyFalse_bufchan_d;
  
  /* demux (Ty MyBool,
       Ty QTree_Bool) : (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2,MyBool) (lizzieLet0_4QVal_Bool_8QVal_Bool_2MyFalse,QTree_Bool) > [(_50,QTree_Bool),
                                                                                                                                       (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue,QTree_Bool)] */
  logic [1:0] lizzieLet0_4QVal_Bool_8QVal_Bool_2MyFalse_onehotd;
  always_comb
    if ((lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2_d[0] && lizzieLet0_4QVal_Bool_8QVal_Bool_2MyFalse_d[0]))
      unique case (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2_d[1:1])
        1'd0: lizzieLet0_4QVal_Bool_8QVal_Bool_2MyFalse_onehotd = 2'd1;
        1'd1: lizzieLet0_4QVal_Bool_8QVal_Bool_2MyFalse_onehotd = 2'd2;
        default: lizzieLet0_4QVal_Bool_8QVal_Bool_2MyFalse_onehotd = 2'd0;
      endcase
    else lizzieLet0_4QVal_Bool_8QVal_Bool_2MyFalse_onehotd = 2'd0;
  assign _50_d = {lizzieLet0_4QVal_Bool_8QVal_Bool_2MyFalse_d[66:1],
                  lizzieLet0_4QVal_Bool_8QVal_Bool_2MyFalse_onehotd[0]};
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_d = {lizzieLet0_4QVal_Bool_8QVal_Bool_2MyFalse_d[66:1],
                                                                lizzieLet0_4QVal_Bool_8QVal_Bool_2MyFalse_onehotd[1]};
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_2MyFalse_r = (| (lizzieLet0_4QVal_Bool_8QVal_Bool_2MyFalse_onehotd & {lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_r,
                                                                                                                _50_r}));
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2_r = lizzieLet0_4QVal_Bool_8QVal_Bool_2MyFalse_r;
  
  /* fork (Ty QTree_Bool) : (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue,QTree_Bool) > [(lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1,QTree_Bool),
                                                                                         (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2,QTree_Bool)] */
  logic [1:0] lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_emitted;
  logic [1:0] lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_done;
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1_d = {lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_d[66:1],
                                                                  (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_d[0] && (! lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_emitted[0]))};
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2_d = {lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_d[66:1],
                                                                  (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_d[0] && (! lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_emitted[1]))};
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_done = (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_emitted | ({lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2_d[0],
                                                                                                                                 lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1_d[0]} & {lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2_r,
                                                                                                                                                                                              lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1_r}));
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_r = (& lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_emitted <= 2'd0;
    else
      lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_emitted <= (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_r ? 2'd0 :
                                                                    lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_done);
  
  /* demux (Ty QTree_Bool,
       Ty Go) : (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1,QTree_Bool) (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_1MyTrue,Go) > [(lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNone_Bool,Go),
                                                                                                                                           (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QVal_Bool,Go),
                                                                                                                                           (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNode_Bool,Go),
                                                                                                                                           (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QError_Bool,Go)] */
  logic [3:0] lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_1MyTrue_onehotd;
  always_comb
    if ((lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1_d[0] && lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_1MyTrue_d[0]))
      unique case (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1_d[2:1])
        2'd0:
          lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_1MyTrue_onehotd = 4'd1;
        2'd1:
          lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_1MyTrue_onehotd = 4'd2;
        2'd2:
          lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_1MyTrue_onehotd = 4'd4;
        2'd3:
          lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_1MyTrue_onehotd = 4'd8;
        default:
          lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_1MyTrue_onehotd = 4'd0;
      endcase
    else
      lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_1MyTrue_onehotd = 4'd0;
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNone_Bool_d = lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_1MyTrue_onehotd[0];
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QVal_Bool_d = lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_1MyTrue_onehotd[1];
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNode_Bool_d = lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_1MyTrue_onehotd[2];
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QError_Bool_d = lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_1MyTrue_onehotd[3];
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_1MyTrue_r = (| (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_1MyTrue_onehotd & {lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QError_Bool_r,
                                                                                                                                lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNode_Bool_r,
                                                                                                                                lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QVal_Bool_r,
                                                                                                                                lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNone_Bool_r}));
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1_r = lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_1MyTrue_r;
  
  /* fork (Ty Go) : (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QError_Bool,Go) > [(lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QError_Bool_1,Go),
                                                                                      (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QError_Bool_2,Go)] */
  logic [1:0] lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QError_Bool_emitted;
  logic [1:0] lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QError_Bool_done;
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QError_Bool_1_d = (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QError_Bool_d[0] && (! lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QError_Bool_emitted[0]));
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QError_Bool_2_d = (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QError_Bool_d[0] && (! lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QError_Bool_emitted[1]));
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QError_Bool_done = (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QError_Bool_emitted | ({lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QError_Bool_2_d[0],
                                                                                                                                                           lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QError_Bool_1_d[0]} & {lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QError_Bool_2_r,
                                                                                                                                                                                                                                     lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QError_Bool_1_r}));
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QError_Bool_r = (& lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QError_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QError_Bool_emitted <= 2'd0;
    else
      lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QError_Bool_emitted <= (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QError_Bool_r ? 2'd0 :
                                                                                 lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QError_Bool_done);
  
  /* dcon (Ty QTree_Bool,
      Dcon QError_Bool) : [(lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QError_Bool_1,Go)] > (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QError_Bool_1QError_Bool,QTree_Bool) */
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QError_Bool_1QError_Bool_d = QError_Bool_dc((& {lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QError_Bool_1_d[0]}), lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QError_Bool_1_d);
  assign {lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QError_Bool_1_r} = {1 {(lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QError_Bool_1QError_Bool_r && lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QError_Bool_1QError_Bool_d[0])}};
  
  /* buf (Ty QTree_Bool) : (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QError_Bool_1QError_Bool,QTree_Bool) > (lizzieLet24_1_argbuf,QTree_Bool) */
  QTree_Bool_t lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QError_Bool_1QError_Bool_bufchan_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QError_Bool_1QError_Bool_bufchan_r;
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QError_Bool_1QError_Bool_r = ((! lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QError_Bool_1QError_Bool_bufchan_d[0]) || lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QError_Bool_1QError_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QError_Bool_1QError_Bool_bufchan_d <= {66'd0,
                                                                                                1'd0};
    else
      if (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QError_Bool_1QError_Bool_r)
        lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QError_Bool_1QError_Bool_bufchan_d <= lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QError_Bool_1QError_Bool_d;
  QTree_Bool_t lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QError_Bool_1QError_Bool_bufchan_buf;
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QError_Bool_1QError_Bool_bufchan_r = (! lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QError_Bool_1QError_Bool_bufchan_buf[0]);
  assign lizzieLet24_1_argbuf_d = (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QError_Bool_1QError_Bool_bufchan_buf[0] ? lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QError_Bool_1QError_Bool_bufchan_buf :
                                   lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QError_Bool_1QError_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QError_Bool_1QError_Bool_bufchan_buf <= {66'd0,
                                                                                                  1'd0};
    else
      if ((lizzieLet24_1_argbuf_r && lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QError_Bool_1QError_Bool_bufchan_buf[0]))
        lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QError_Bool_1QError_Bool_bufchan_buf <= {66'd0,
                                                                                                    1'd0};
      else if (((! lizzieLet24_1_argbuf_r) && (! lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QError_Bool_1QError_Bool_bufchan_buf[0])))
        lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QError_Bool_1QError_Bool_bufchan_buf <= lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QError_Bool_1QError_Bool_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QError_Bool_2,Go) > (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QError_Bool_2_argbuf,Go) */
  Go_t lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QError_Bool_2_bufchan_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QError_Bool_2_bufchan_r;
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QError_Bool_2_r = ((! lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QError_Bool_2_bufchan_d[0]) || lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QError_Bool_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QError_Bool_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QError_Bool_2_r)
        lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QError_Bool_2_bufchan_d <= lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QError_Bool_2_d;
  Go_t lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QError_Bool_2_bufchan_buf;
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QError_Bool_2_bufchan_r = (! lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QError_Bool_2_bufchan_buf[0]);
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QError_Bool_2_argbuf_d = (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QError_Bool_2_bufchan_buf[0] ? lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QError_Bool_2_bufchan_buf :
                                                                                      lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QError_Bool_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QError_Bool_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QError_Bool_2_argbuf_r && lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QError_Bool_2_bufchan_buf[0]))
        lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QError_Bool_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QError_Bool_2_argbuf_r) && (! lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QError_Bool_2_bufchan_buf[0])))
        lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QError_Bool_2_bufchan_buf <= lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QError_Bool_2_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNode_Bool,Go) > [(lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNode_Bool_1,Go),
                                                                                     (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNode_Bool_2,Go)] */
  logic [1:0] lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNode_Bool_emitted;
  logic [1:0] lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNode_Bool_done;
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNode_Bool_1_d = (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNode_Bool_d[0] && (! lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNode_Bool_emitted[0]));
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNode_Bool_2_d = (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNode_Bool_d[0] && (! lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNode_Bool_emitted[1]));
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNode_Bool_done = (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNode_Bool_emitted | ({lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNode_Bool_2_d[0],
                                                                                                                                                         lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNode_Bool_1_d[0]} & {lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNode_Bool_2_r,
                                                                                                                                                                                                                                  lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNode_Bool_1_r}));
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNode_Bool_r = (& lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNode_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNode_Bool_emitted <= 2'd0;
    else
      lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNode_Bool_emitted <= (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNode_Bool_r ? 2'd0 :
                                                                                lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNode_Bool_done);
  
  /* dcon (Ty QTree_Bool,
      Dcon QError_Bool) : [(lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNode_Bool_1,Go)] > (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNode_Bool_1QError_Bool,QTree_Bool) */
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNode_Bool_1QError_Bool_d = QError_Bool_dc((& {lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNode_Bool_1_d[0]}), lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNode_Bool_1_d);
  assign {lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNode_Bool_1_r} = {1 {(lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNode_Bool_1QError_Bool_r && lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNode_Bool_1QError_Bool_d[0])}};
  
  /* buf (Ty QTree_Bool) : (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNode_Bool_1QError_Bool,QTree_Bool) > (lizzieLet23_1_argbuf,QTree_Bool) */
  QTree_Bool_t lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNode_Bool_1QError_Bool_bufchan_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNode_Bool_1QError_Bool_bufchan_r;
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNode_Bool_1QError_Bool_r = ((! lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNode_Bool_1QError_Bool_bufchan_d[0]) || lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNode_Bool_1QError_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNode_Bool_1QError_Bool_bufchan_d <= {66'd0,
                                                                                               1'd0};
    else
      if (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNode_Bool_1QError_Bool_r)
        lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNode_Bool_1QError_Bool_bufchan_d <= lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNode_Bool_1QError_Bool_d;
  QTree_Bool_t lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNode_Bool_1QError_Bool_bufchan_buf;
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNode_Bool_1QError_Bool_bufchan_r = (! lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNode_Bool_1QError_Bool_bufchan_buf[0]);
  assign lizzieLet23_1_argbuf_d = (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNode_Bool_1QError_Bool_bufchan_buf[0] ? lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNode_Bool_1QError_Bool_bufchan_buf :
                                   lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNode_Bool_1QError_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNode_Bool_1QError_Bool_bufchan_buf <= {66'd0,
                                                                                                 1'd0};
    else
      if ((lizzieLet23_1_argbuf_r && lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNode_Bool_1QError_Bool_bufchan_buf[0]))
        lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNode_Bool_1QError_Bool_bufchan_buf <= {66'd0,
                                                                                                   1'd0};
      else if (((! lizzieLet23_1_argbuf_r) && (! lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNode_Bool_1QError_Bool_bufchan_buf[0])))
        lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNode_Bool_1QError_Bool_bufchan_buf <= lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNode_Bool_1QError_Bool_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNode_Bool_2,Go) > (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNode_Bool_2_argbuf,Go) */
  Go_t lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNode_Bool_2_bufchan_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNode_Bool_2_bufchan_r;
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNode_Bool_2_r = ((! lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNode_Bool_2_bufchan_d[0]) || lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNode_Bool_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNode_Bool_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNode_Bool_2_r)
        lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNode_Bool_2_bufchan_d <= lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNode_Bool_2_d;
  Go_t lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNode_Bool_2_bufchan_buf;
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNode_Bool_2_bufchan_r = (! lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNode_Bool_2_bufchan_buf[0]);
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNode_Bool_2_argbuf_d = (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNode_Bool_2_bufchan_buf[0] ? lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNode_Bool_2_bufchan_buf :
                                                                                     lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNode_Bool_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNode_Bool_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNode_Bool_2_argbuf_r && lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNode_Bool_2_bufchan_buf[0]))
        lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNode_Bool_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNode_Bool_2_argbuf_r) && (! lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNode_Bool_2_bufchan_buf[0])))
        lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNode_Bool_2_bufchan_buf <= lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNode_Bool_2_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNone_Bool,Go) > [(lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNone_Bool_1,Go),
                                                                                     (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNone_Bool_2,Go)] */
  logic [1:0] lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNone_Bool_emitted;
  logic [1:0] lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNone_Bool_done;
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNone_Bool_1_d = (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNone_Bool_d[0] && (! lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNone_Bool_emitted[0]));
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNone_Bool_2_d = (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNone_Bool_d[0] && (! lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNone_Bool_emitted[1]));
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNone_Bool_done = (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNone_Bool_emitted | ({lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNone_Bool_2_d[0],
                                                                                                                                                         lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNone_Bool_1_d[0]} & {lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNone_Bool_2_r,
                                                                                                                                                                                                                                  lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNone_Bool_1_r}));
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNone_Bool_r = (& lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNone_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNone_Bool_emitted <= 2'd0;
    else
      lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNone_Bool_emitted <= (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNone_Bool_r ? 2'd0 :
                                                                                lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNone_Bool_done);
  
  /* buf (Ty Go) : (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNone_Bool_1,Go) > (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNone_Bool_1_argbuf,Go) */
  Go_t lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNone_Bool_1_bufchan_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNone_Bool_1_bufchan_r;
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNone_Bool_1_r = ((! lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNone_Bool_1_bufchan_d[0]) || lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNone_Bool_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNone_Bool_1_bufchan_d <= 1'd0;
    else
      if (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNone_Bool_1_r)
        lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNone_Bool_1_bufchan_d <= lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNone_Bool_1_d;
  Go_t lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNone_Bool_1_bufchan_buf;
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNone_Bool_1_bufchan_r = (! lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNone_Bool_1_bufchan_buf[0]);
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNone_Bool_1_argbuf_d = (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNone_Bool_1_bufchan_buf[0] ? lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNone_Bool_1_bufchan_buf :
                                                                                     lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNone_Bool_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNone_Bool_1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNone_Bool_1_argbuf_r && lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNone_Bool_1_bufchan_buf[0]))
        lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNone_Bool_1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNone_Bool_1_argbuf_r) && (! lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNone_Bool_1_bufchan_buf[0])))
        lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNone_Bool_1_bufchan_buf <= lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNone_Bool_1_bufchan_d;
  
  /* dcon (Ty TupGo,
      Dcon TupGo) : [(lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNone_Bool_1_argbuf,Go)] > (lvlrf2-0TupGo7,TupGo) */
  assign \lvlrf2-0TupGo7_d  = TupGo_dc((& {lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNone_Bool_1_argbuf_d[0]}), lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNone_Bool_1_argbuf_d);
  assign {lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNone_Bool_1_argbuf_r} = {1 {(\lvlrf2-0TupGo7_r  && \lvlrf2-0TupGo7_d [0])}};
  
  /* buf (Ty Go) : (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNone_Bool_2,Go) > (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNone_Bool_2_argbuf,Go) */
  Go_t lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNone_Bool_2_bufchan_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNone_Bool_2_bufchan_r;
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNone_Bool_2_r = ((! lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNone_Bool_2_bufchan_d[0]) || lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNone_Bool_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNone_Bool_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNone_Bool_2_r)
        lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNone_Bool_2_bufchan_d <= lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNone_Bool_2_d;
  Go_t lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNone_Bool_2_bufchan_buf;
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNone_Bool_2_bufchan_r = (! lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNone_Bool_2_bufchan_buf[0]);
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNone_Bool_2_argbuf_d = (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNone_Bool_2_bufchan_buf[0] ? lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNone_Bool_2_bufchan_buf :
                                                                                     lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNone_Bool_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNone_Bool_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNone_Bool_2_argbuf_r && lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNone_Bool_2_bufchan_buf[0]))
        lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNone_Bool_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNone_Bool_2_argbuf_r) && (! lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNone_Bool_2_bufchan_buf[0])))
        lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNone_Bool_2_bufchan_buf <= lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QNone_Bool_2_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QVal_Bool,Go) > [(lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QVal_Bool_1,Go),
                                                                                    (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QVal_Bool_2,Go)] */
  logic [1:0] lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QVal_Bool_emitted;
  logic [1:0] lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QVal_Bool_done;
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QVal_Bool_1_d = (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QVal_Bool_d[0] && (! lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QVal_Bool_emitted[0]));
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QVal_Bool_2_d = (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QVal_Bool_d[0] && (! lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QVal_Bool_emitted[1]));
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QVal_Bool_done = (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QVal_Bool_emitted | ({lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QVal_Bool_2_d[0],
                                                                                                                                                       lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QVal_Bool_1_d[0]} & {lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QVal_Bool_2_r,
                                                                                                                                                                                                                               lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QVal_Bool_1_r}));
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QVal_Bool_r = (& lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QVal_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QVal_Bool_emitted <= 2'd0;
    else
      lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QVal_Bool_emitted <= (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QVal_Bool_r ? 2'd0 :
                                                                               lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QVal_Bool_done);
  
  /* buf (Ty Go) : (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QVal_Bool_1,Go) > (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QVal_Bool_1_argbuf,Go) */
  Go_t lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QVal_Bool_1_bufchan_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QVal_Bool_1_bufchan_r;
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QVal_Bool_1_r = ((! lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QVal_Bool_1_bufchan_d[0]) || lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QVal_Bool_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QVal_Bool_1_bufchan_d <= 1'd0;
    else
      if (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QVal_Bool_1_r)
        lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QVal_Bool_1_bufchan_d <= lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QVal_Bool_1_d;
  Go_t lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QVal_Bool_1_bufchan_buf;
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QVal_Bool_1_bufchan_r = (! lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QVal_Bool_1_bufchan_buf[0]);
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QVal_Bool_1_argbuf_d = (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QVal_Bool_1_bufchan_buf[0] ? lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QVal_Bool_1_bufchan_buf :
                                                                                    lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QVal_Bool_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QVal_Bool_1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QVal_Bool_1_argbuf_r && lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QVal_Bool_1_bufchan_buf[0]))
        lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QVal_Bool_1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QVal_Bool_1_argbuf_r) && (! lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QVal_Bool_1_bufchan_buf[0])))
        lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QVal_Bool_1_bufchan_buf <= lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QVal_Bool_1_bufchan_d;
  
  /* dcon (Ty TupGo,
      Dcon TupGo) : [(lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QVal_Bool_1_argbuf,Go)] > (lvlrf2-0TupGo8,TupGo) */
  assign \lvlrf2-0TupGo8_d  = TupGo_dc((& {lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QVal_Bool_1_argbuf_d[0]}), lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QVal_Bool_1_argbuf_d);
  assign {lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QVal_Bool_1_argbuf_r} = {1 {(\lvlrf2-0TupGo8_r  && \lvlrf2-0TupGo8_d [0])}};
  
  /* buf (Ty Go) : (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QVal_Bool_2,Go) > (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QVal_Bool_2_argbuf,Go) */
  Go_t lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QVal_Bool_2_bufchan_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QVal_Bool_2_bufchan_r;
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QVal_Bool_2_r = ((! lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QVal_Bool_2_bufchan_d[0]) || lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QVal_Bool_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QVal_Bool_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QVal_Bool_2_r)
        lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QVal_Bool_2_bufchan_d <= lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QVal_Bool_2_d;
  Go_t lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QVal_Bool_2_bufchan_buf;
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QVal_Bool_2_bufchan_r = (! lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QVal_Bool_2_bufchan_buf[0]);
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QVal_Bool_2_argbuf_d = (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QVal_Bool_2_bufchan_buf[0] ? lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QVal_Bool_2_bufchan_buf :
                                                                                    lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QVal_Bool_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QVal_Bool_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QVal_Bool_2_argbuf_r && lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QVal_Bool_2_bufchan_buf[0]))
        lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QVal_Bool_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QVal_Bool_2_argbuf_r) && (! lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QVal_Bool_2_bufchan_buf[0])))
        lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QVal_Bool_2_bufchan_buf <= lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_1QVal_Bool_2_bufchan_d;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_CTf) : (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2,QTree_Bool) (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_4MyTrue,Pointer_CTf) > [(lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QNone_Bool,Pointer_CTf),
                                                                                                                                                             (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QVal_Bool,Pointer_CTf),
                                                                                                                                                             (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QNode_Bool,Pointer_CTf),
                                                                                                                                                             (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QError_Bool,Pointer_CTf)] */
  logic [3:0] lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_4MyTrue_onehotd;
  always_comb
    if ((lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2_d[0] && lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_4MyTrue_d[0]))
      unique case (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2_d[2:1])
        2'd0:
          lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_4MyTrue_onehotd = 4'd1;
        2'd1:
          lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_4MyTrue_onehotd = 4'd2;
        2'd2:
          lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_4MyTrue_onehotd = 4'd4;
        2'd3:
          lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_4MyTrue_onehotd = 4'd8;
        default:
          lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_4MyTrue_onehotd = 4'd0;
      endcase
    else
      lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_4MyTrue_onehotd = 4'd0;
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QNone_Bool_d = {lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_4MyTrue_d[16:1],
                                                                            lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_4MyTrue_onehotd[0]};
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QVal_Bool_d = {lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_4MyTrue_d[16:1],
                                                                           lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_4MyTrue_onehotd[1]};
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QNode_Bool_d = {lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_4MyTrue_d[16:1],
                                                                            lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_4MyTrue_onehotd[2]};
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QError_Bool_d = {lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_4MyTrue_d[16:1],
                                                                             lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_4MyTrue_onehotd[3]};
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_4MyTrue_r = (| (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_4MyTrue_onehotd & {lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QError_Bool_r,
                                                                                                                                lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QNode_Bool_r,
                                                                                                                                lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QVal_Bool_r,
                                                                                                                                lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QNone_Bool_r}));
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2_r = lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_4MyTrue_r;
  
  /* buf (Ty Pointer_CTf) : (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QError_Bool,Pointer_CTf) > (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QError_Bool_1_argbuf,Pointer_CTf) */
  Pointer_CTf_t lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QError_Bool_bufchan_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QError_Bool_bufchan_r;
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QError_Bool_r = ((! lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QError_Bool_bufchan_d[0]) || lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QError_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QError_Bool_bufchan_d <= {16'd0,
                                                                                   1'd0};
    else
      if (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QError_Bool_r)
        lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QError_Bool_bufchan_d <= lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QError_Bool_d;
  Pointer_CTf_t lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QError_Bool_bufchan_buf;
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QError_Bool_bufchan_r = (! lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QError_Bool_bufchan_buf[0]);
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QError_Bool_1_argbuf_d = (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QError_Bool_bufchan_buf[0] ? lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QError_Bool_bufchan_buf :
                                                                                      lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QError_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QError_Bool_bufchan_buf <= {16'd0,
                                                                                     1'd0};
    else
      if ((lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QError_Bool_1_argbuf_r && lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QError_Bool_bufchan_buf[0]))
        lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QError_Bool_bufchan_buf <= {16'd0,
                                                                                       1'd0};
      else if (((! lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QError_Bool_1_argbuf_r) && (! lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QError_Bool_bufchan_buf[0])))
        lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QError_Bool_bufchan_buf <= lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QError_Bool_bufchan_d;
  
  /* buf (Ty Pointer_CTf) : (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QNode_Bool,Pointer_CTf) > (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QNode_Bool_1_argbuf,Pointer_CTf) */
  Pointer_CTf_t lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QNode_Bool_bufchan_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QNode_Bool_bufchan_r;
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QNode_Bool_r = ((! lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QNode_Bool_bufchan_d[0]) || lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QNode_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QNode_Bool_bufchan_d <= {16'd0,
                                                                                  1'd0};
    else
      if (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QNode_Bool_r)
        lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QNode_Bool_bufchan_d <= lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QNode_Bool_d;
  Pointer_CTf_t lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QNode_Bool_bufchan_buf;
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QNode_Bool_bufchan_r = (! lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QNode_Bool_bufchan_buf[0]);
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QNode_Bool_1_argbuf_d = (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QNode_Bool_bufchan_buf[0] ? lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QNode_Bool_bufchan_buf :
                                                                                     lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QNode_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QNode_Bool_bufchan_buf <= {16'd0,
                                                                                    1'd0};
    else
      if ((lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QNode_Bool_1_argbuf_r && lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QNode_Bool_bufchan_buf[0]))
        lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QNode_Bool_bufchan_buf <= {16'd0,
                                                                                      1'd0};
      else if (((! lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QNode_Bool_1_argbuf_r) && (! lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QNode_Bool_bufchan_buf[0])))
        lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QNode_Bool_bufchan_buf <= lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QNode_Bool_bufchan_d;
  
  /* buf (Ty Pointer_CTf) : (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QNone_Bool,Pointer_CTf) > (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QNone_Bool_1_argbuf,Pointer_CTf) */
  Pointer_CTf_t lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QNone_Bool_bufchan_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QNone_Bool_bufchan_r;
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QNone_Bool_r = ((! lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QNone_Bool_bufchan_d[0]) || lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QNone_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QNone_Bool_bufchan_d <= {16'd0,
                                                                                  1'd0};
    else
      if (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QNone_Bool_r)
        lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QNone_Bool_bufchan_d <= lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QNone_Bool_d;
  Pointer_CTf_t lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QNone_Bool_bufchan_buf;
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QNone_Bool_bufchan_r = (! lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QNone_Bool_bufchan_buf[0]);
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QNone_Bool_1_argbuf_d = (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QNone_Bool_bufchan_buf[0] ? lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QNone_Bool_bufchan_buf :
                                                                                     lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QNone_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QNone_Bool_bufchan_buf <= {16'd0,
                                                                                    1'd0};
    else
      if ((lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QNone_Bool_1_argbuf_r && lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QNone_Bool_bufchan_buf[0]))
        lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QNone_Bool_bufchan_buf <= {16'd0,
                                                                                      1'd0};
      else if (((! lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QNone_Bool_1_argbuf_r) && (! lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QNone_Bool_bufchan_buf[0])))
        lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QNone_Bool_bufchan_buf <= lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QNone_Bool_bufchan_d;
  
  /* buf (Ty Pointer_CTf) : (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QVal_Bool,Pointer_CTf) > (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QVal_Bool_1_argbuf,Pointer_CTf) */
  Pointer_CTf_t lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QVal_Bool_bufchan_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QVal_Bool_bufchan_r;
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QVal_Bool_r = ((! lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QVal_Bool_bufchan_d[0]) || lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QVal_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QVal_Bool_bufchan_d <= {16'd0,
                                                                                 1'd0};
    else
      if (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QVal_Bool_r)
        lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QVal_Bool_bufchan_d <= lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QVal_Bool_d;
  Pointer_CTf_t lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QVal_Bool_bufchan_buf;
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QVal_Bool_bufchan_r = (! lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QVal_Bool_bufchan_buf[0]);
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QVal_Bool_1_argbuf_d = (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QVal_Bool_bufchan_buf[0] ? lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QVal_Bool_bufchan_buf :
                                                                                    lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QVal_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QVal_Bool_bufchan_buf <= {16'd0,
                                                                                   1'd0};
    else
      if ((lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QVal_Bool_1_argbuf_r && lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QVal_Bool_bufchan_buf[0]))
        lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QVal_Bool_bufchan_buf <= {16'd0,
                                                                                     1'd0};
      else if (((! lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QVal_Bool_1_argbuf_r) && (! lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QVal_Bool_bufchan_buf[0])))
        lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QVal_Bool_bufchan_buf <= lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_2MyTrue_2QVal_Bool_bufchan_d;
  
  /* demux (Ty MyBool,
       Ty Pointer_QTree_Bool) : (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_3,MyBool) (lizzieLet0_4QVal_Bool_8QVal_Bool_3MyFalse,Pointer_QTree_Bool) > [(lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_3MyFalse,Pointer_QTree_Bool),
                                                                                                                                                       (_49,Pointer_QTree_Bool)] */
  logic [1:0] lizzieLet0_4QVal_Bool_8QVal_Bool_3MyFalse_onehotd;
  always_comb
    if ((lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_3_d[0] && lizzieLet0_4QVal_Bool_8QVal_Bool_3MyFalse_d[0]))
      unique case (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_3_d[1:1])
        1'd0: lizzieLet0_4QVal_Bool_8QVal_Bool_3MyFalse_onehotd = 2'd1;
        1'd1: lizzieLet0_4QVal_Bool_8QVal_Bool_3MyFalse_onehotd = 2'd2;
        default: lizzieLet0_4QVal_Bool_8QVal_Bool_3MyFalse_onehotd = 2'd0;
      endcase
    else lizzieLet0_4QVal_Bool_8QVal_Bool_3MyFalse_onehotd = 2'd0;
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_3MyFalse_d = {lizzieLet0_4QVal_Bool_8QVal_Bool_3MyFalse_d[16:1],
                                                                 lizzieLet0_4QVal_Bool_8QVal_Bool_3MyFalse_onehotd[0]};
  assign _49_d = {lizzieLet0_4QVal_Bool_8QVal_Bool_3MyFalse_d[16:1],
                  lizzieLet0_4QVal_Bool_8QVal_Bool_3MyFalse_onehotd[1]};
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_3MyFalse_r = (| (lizzieLet0_4QVal_Bool_8QVal_Bool_3MyFalse_onehotd & {_49_r,
                                                                                                                lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_3MyFalse_r}));
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_3_r = lizzieLet0_4QVal_Bool_8QVal_Bool_3MyFalse_r;
  
  /* buf (Ty Pointer_QTree_Bool) : (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_3MyFalse,Pointer_QTree_Bool) > (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_3MyFalse_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_3MyFalse_bufchan_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_3MyFalse_bufchan_r;
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_3MyFalse_r = ((! lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_3MyFalse_bufchan_d[0]) || lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_3MyFalse_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_3MyFalse_bufchan_d <= {16'd0,
                                                                       1'd0};
    else
      if (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_3MyFalse_r)
        lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_3MyFalse_bufchan_d <= lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_3MyFalse_d;
  Pointer_QTree_Bool_t lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_3MyFalse_bufchan_buf;
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_3MyFalse_bufchan_r = (! lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_3MyFalse_bufchan_buf[0]);
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_3MyFalse_1_argbuf_d = (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_3MyFalse_bufchan_buf[0] ? lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_3MyFalse_bufchan_buf :
                                                                          lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_3MyFalse_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_3MyFalse_bufchan_buf <= {16'd0,
                                                                         1'd0};
    else
      if ((lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_3MyFalse_1_argbuf_r && lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_3MyFalse_bufchan_buf[0]))
        lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_3MyFalse_bufchan_buf <= {16'd0,
                                                                           1'd0};
      else if (((! lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_3MyFalse_1_argbuf_r) && (! lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_3MyFalse_bufchan_buf[0])))
        lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_3MyFalse_bufchan_buf <= lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_3MyFalse_bufchan_d;
  
  /* demux (Ty MyBool,
       Ty Pointer_CTf) : (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_4,MyBool) (lizzieLet0_4QVal_Bool_8QVal_Bool_4MyFalse,Pointer_CTf) > [(lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_4MyFalse,Pointer_CTf),
                                                                                                                                         (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_4MyTrue,Pointer_CTf)] */
  logic [1:0] lizzieLet0_4QVal_Bool_8QVal_Bool_4MyFalse_onehotd;
  always_comb
    if ((lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_4_d[0] && lizzieLet0_4QVal_Bool_8QVal_Bool_4MyFalse_d[0]))
      unique case (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_4_d[1:1])
        1'd0: lizzieLet0_4QVal_Bool_8QVal_Bool_4MyFalse_onehotd = 2'd1;
        1'd1: lizzieLet0_4QVal_Bool_8QVal_Bool_4MyFalse_onehotd = 2'd2;
        default: lizzieLet0_4QVal_Bool_8QVal_Bool_4MyFalse_onehotd = 2'd0;
      endcase
    else lizzieLet0_4QVal_Bool_8QVal_Bool_4MyFalse_onehotd = 2'd0;
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_4MyFalse_d = {lizzieLet0_4QVal_Bool_8QVal_Bool_4MyFalse_d[16:1],
                                                                 lizzieLet0_4QVal_Bool_8QVal_Bool_4MyFalse_onehotd[0]};
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_4MyTrue_d = {lizzieLet0_4QVal_Bool_8QVal_Bool_4MyFalse_d[16:1],
                                                                lizzieLet0_4QVal_Bool_8QVal_Bool_4MyFalse_onehotd[1]};
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_4MyFalse_r = (| (lizzieLet0_4QVal_Bool_8QVal_Bool_4MyFalse_onehotd & {lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_4MyTrue_r,
                                                                                                                lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_4MyFalse_r}));
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_4_r = lizzieLet0_4QVal_Bool_8QVal_Bool_4MyFalse_r;
  
  /* buf (Ty Pointer_CTf) : (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_4MyFalse,Pointer_CTf) > (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_4MyFalse_1_argbuf,Pointer_CTf) */
  Pointer_CTf_t lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_4MyFalse_bufchan_d;
  logic lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_4MyFalse_bufchan_r;
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_4MyFalse_r = ((! lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_4MyFalse_bufchan_d[0]) || lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_4MyFalse_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_4MyFalse_bufchan_d <= {16'd0,
                                                                       1'd0};
    else
      if (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_4MyFalse_r)
        lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_4MyFalse_bufchan_d <= lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_4MyFalse_d;
  Pointer_CTf_t lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_4MyFalse_bufchan_buf;
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_4MyFalse_bufchan_r = (! lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_4MyFalse_bufchan_buf[0]);
  assign lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_4MyFalse_1_argbuf_d = (lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_4MyFalse_bufchan_buf[0] ? lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_4MyFalse_bufchan_buf :
                                                                          lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_4MyFalse_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_4MyFalse_bufchan_buf <= {16'd0,
                                                                         1'd0};
    else
      if ((lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_4MyFalse_1_argbuf_r && lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_4MyFalse_bufchan_buf[0]))
        lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_4MyFalse_bufchan_buf <= {16'd0,
                                                                           1'd0};
      else if (((! lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_4MyFalse_1_argbuf_r) && (! lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_4MyFalse_bufchan_buf[0])))
        lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_4MyFalse_bufchan_buf <= lizzieLet0_4QVal_Bool_8QVal_Bool_5MyFalse_4MyFalse_bufchan_d;
  
  /* demux (Ty QTree_Bool,
       Ty QTree_Bool) : (lizzieLet0_5,QTree_Bool) (readPointer_QTree_Boolm3a86_1_argbuf_rwb,QTree_Bool) > [(lizzieLet0_5QNone_Bool,QTree_Bool),
                                                                                                           (lizzieLet0_5QVal_Bool,QTree_Bool),
                                                                                                           (lizzieLet0_5QNode_Bool,QTree_Bool),
                                                                                                           (_48,QTree_Bool)] */
  logic [3:0] readPointer_QTree_Boolm3a86_1_argbuf_rwb_onehotd;
  always_comb
    if ((lizzieLet0_5_d[0] && readPointer_QTree_Boolm3a86_1_argbuf_rwb_d[0]))
      unique case (lizzieLet0_5_d[2:1])
        2'd0: readPointer_QTree_Boolm3a86_1_argbuf_rwb_onehotd = 4'd1;
        2'd1: readPointer_QTree_Boolm3a86_1_argbuf_rwb_onehotd = 4'd2;
        2'd2: readPointer_QTree_Boolm3a86_1_argbuf_rwb_onehotd = 4'd4;
        2'd3: readPointer_QTree_Boolm3a86_1_argbuf_rwb_onehotd = 4'd8;
        default: readPointer_QTree_Boolm3a86_1_argbuf_rwb_onehotd = 4'd0;
      endcase
    else readPointer_QTree_Boolm3a86_1_argbuf_rwb_onehotd = 4'd0;
  assign lizzieLet0_5QNone_Bool_d = {readPointer_QTree_Boolm3a86_1_argbuf_rwb_d[66:1],
                                     readPointer_QTree_Boolm3a86_1_argbuf_rwb_onehotd[0]};
  assign lizzieLet0_5QVal_Bool_d = {readPointer_QTree_Boolm3a86_1_argbuf_rwb_d[66:1],
                                    readPointer_QTree_Boolm3a86_1_argbuf_rwb_onehotd[1]};
  assign lizzieLet0_5QNode_Bool_d = {readPointer_QTree_Boolm3a86_1_argbuf_rwb_d[66:1],
                                     readPointer_QTree_Boolm3a86_1_argbuf_rwb_onehotd[2]};
  assign _48_d = {readPointer_QTree_Boolm3a86_1_argbuf_rwb_d[66:1],
                  readPointer_QTree_Boolm3a86_1_argbuf_rwb_onehotd[3]};
  assign readPointer_QTree_Boolm3a86_1_argbuf_rwb_r = (| (readPointer_QTree_Boolm3a86_1_argbuf_rwb_onehotd & {_48_r,
                                                                                                              lizzieLet0_5QNode_Bool_r,
                                                                                                              lizzieLet0_5QVal_Bool_r,
                                                                                                              lizzieLet0_5QNone_Bool_r}));
  assign lizzieLet0_5_r = readPointer_QTree_Boolm3a86_1_argbuf_rwb_r;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_QTree_Bool) : (lizzieLet0_6,QTree_Bool) (m1a84_2,Pointer_QTree_Bool) > [(_47,Pointer_QTree_Bool),
                                                                                          (lizzieLet0_6QVal_Bool,Pointer_QTree_Bool),
                                                                                          (lizzieLet0_6QNode_Bool,Pointer_QTree_Bool),
                                                                                          (_46,Pointer_QTree_Bool)] */
  logic [3:0] m1a84_2_onehotd;
  always_comb
    if ((lizzieLet0_6_d[0] && m1a84_2_d[0]))
      unique case (lizzieLet0_6_d[2:1])
        2'd0: m1a84_2_onehotd = 4'd1;
        2'd1: m1a84_2_onehotd = 4'd2;
        2'd2: m1a84_2_onehotd = 4'd4;
        2'd3: m1a84_2_onehotd = 4'd8;
        default: m1a84_2_onehotd = 4'd0;
      endcase
    else m1a84_2_onehotd = 4'd0;
  assign _47_d = {m1a84_2_d[16:1], m1a84_2_onehotd[0]};
  assign lizzieLet0_6QVal_Bool_d = {m1a84_2_d[16:1],
                                    m1a84_2_onehotd[1]};
  assign lizzieLet0_6QNode_Bool_d = {m1a84_2_d[16:1],
                                     m1a84_2_onehotd[2]};
  assign _46_d = {m1a84_2_d[16:1], m1a84_2_onehotd[3]};
  assign m1a84_2_r = (| (m1a84_2_onehotd & {_46_r,
                                            lizzieLet0_6QNode_Bool_r,
                                            lizzieLet0_6QVal_Bool_r,
                                            _47_r}));
  assign lizzieLet0_6_r = m1a84_2_r;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_QTree_Bool) : (lizzieLet0_7,QTree_Bool) (m2a85_2,Pointer_QTree_Bool) > [(lizzieLet0_7QNone_Bool,Pointer_QTree_Bool),
                                                                                          (_45,Pointer_QTree_Bool),
                                                                                          (_44,Pointer_QTree_Bool),
                                                                                          (_43,Pointer_QTree_Bool)] */
  logic [3:0] m2a85_2_onehotd;
  always_comb
    if ((lizzieLet0_7_d[0] && m2a85_2_d[0]))
      unique case (lizzieLet0_7_d[2:1])
        2'd0: m2a85_2_onehotd = 4'd1;
        2'd1: m2a85_2_onehotd = 4'd2;
        2'd2: m2a85_2_onehotd = 4'd4;
        2'd3: m2a85_2_onehotd = 4'd8;
        default: m2a85_2_onehotd = 4'd0;
      endcase
    else m2a85_2_onehotd = 4'd0;
  assign lizzieLet0_7QNone_Bool_d = {m2a85_2_d[16:1],
                                     m2a85_2_onehotd[0]};
  assign _45_d = {m2a85_2_d[16:1], m2a85_2_onehotd[1]};
  assign _44_d = {m2a85_2_d[16:1], m2a85_2_onehotd[2]};
  assign _43_d = {m2a85_2_d[16:1], m2a85_2_onehotd[3]};
  assign m2a85_2_r = (| (m2a85_2_onehotd & {_43_r,
                                            _44_r,
                                            _45_r,
                                            lizzieLet0_7QNone_Bool_r}));
  assign lizzieLet0_7_r = m2a85_2_r;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_QTree_Bool) : (lizzieLet0_8,QTree_Bool) (m3a86_2,Pointer_QTree_Bool) > [(lizzieLet0_8QNone_Bool,Pointer_QTree_Bool),
                                                                                          (lizzieLet0_8QVal_Bool,Pointer_QTree_Bool),
                                                                                          (_42,Pointer_QTree_Bool),
                                                                                          (_41,Pointer_QTree_Bool)] */
  logic [3:0] m3a86_2_onehotd;
  always_comb
    if ((lizzieLet0_8_d[0] && m3a86_2_d[0]))
      unique case (lizzieLet0_8_d[2:1])
        2'd0: m3a86_2_onehotd = 4'd1;
        2'd1: m3a86_2_onehotd = 4'd2;
        2'd2: m3a86_2_onehotd = 4'd4;
        2'd3: m3a86_2_onehotd = 4'd8;
        default: m3a86_2_onehotd = 4'd0;
      endcase
    else m3a86_2_onehotd = 4'd0;
  assign lizzieLet0_8QNone_Bool_d = {m3a86_2_d[16:1],
                                     m3a86_2_onehotd[0]};
  assign lizzieLet0_8QVal_Bool_d = {m3a86_2_d[16:1],
                                    m3a86_2_onehotd[1]};
  assign _42_d = {m3a86_2_d[16:1], m3a86_2_onehotd[2]};
  assign _41_d = {m3a86_2_d[16:1], m3a86_2_onehotd[3]};
  assign m3a86_2_r = (| (m3a86_2_onehotd & {_41_r,
                                            _42_r,
                                            lizzieLet0_8QVal_Bool_r,
                                            lizzieLet0_8QNone_Bool_r}));
  assign lizzieLet0_8_r = m3a86_2_r;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_CTf) : (lizzieLet0_9,QTree_Bool) (sc_0_goMux_mux,Pointer_CTf) > [(lizzieLet0_9QNone_Bool,Pointer_CTf),
                                                                                   (lizzieLet0_9QVal_Bool,Pointer_CTf),
                                                                                   (lizzieLet0_9QNode_Bool,Pointer_CTf),
                                                                                   (lizzieLet0_9QError_Bool,Pointer_CTf)] */
  logic [3:0] sc_0_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet0_9_d[0] && sc_0_goMux_mux_d[0]))
      unique case (lizzieLet0_9_d[2:1])
        2'd0: sc_0_goMux_mux_onehotd = 4'd1;
        2'd1: sc_0_goMux_mux_onehotd = 4'd2;
        2'd2: sc_0_goMux_mux_onehotd = 4'd4;
        2'd3: sc_0_goMux_mux_onehotd = 4'd8;
        default: sc_0_goMux_mux_onehotd = 4'd0;
      endcase
    else sc_0_goMux_mux_onehotd = 4'd0;
  assign lizzieLet0_9QNone_Bool_d = {sc_0_goMux_mux_d[16:1],
                                     sc_0_goMux_mux_onehotd[0]};
  assign lizzieLet0_9QVal_Bool_d = {sc_0_goMux_mux_d[16:1],
                                    sc_0_goMux_mux_onehotd[1]};
  assign lizzieLet0_9QNode_Bool_d = {sc_0_goMux_mux_d[16:1],
                                     sc_0_goMux_mux_onehotd[2]};
  assign lizzieLet0_9QError_Bool_d = {sc_0_goMux_mux_d[16:1],
                                      sc_0_goMux_mux_onehotd[3]};
  assign sc_0_goMux_mux_r = (| (sc_0_goMux_mux_onehotd & {lizzieLet0_9QError_Bool_r,
                                                          lizzieLet0_9QNode_Bool_r,
                                                          lizzieLet0_9QVal_Bool_r,
                                                          lizzieLet0_9QNone_Bool_r}));
  assign lizzieLet0_9_r = sc_0_goMux_mux_r;
  
  /* buf (Ty Pointer_CTf) : (lizzieLet0_9QError_Bool,Pointer_CTf) > (lizzieLet0_9QError_Bool_1_argbuf,Pointer_CTf) */
  Pointer_CTf_t lizzieLet0_9QError_Bool_bufchan_d;
  logic lizzieLet0_9QError_Bool_bufchan_r;
  assign lizzieLet0_9QError_Bool_r = ((! lizzieLet0_9QError_Bool_bufchan_d[0]) || lizzieLet0_9QError_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_9QError_Bool_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet0_9QError_Bool_r)
        lizzieLet0_9QError_Bool_bufchan_d <= lizzieLet0_9QError_Bool_d;
  Pointer_CTf_t lizzieLet0_9QError_Bool_bufchan_buf;
  assign lizzieLet0_9QError_Bool_bufchan_r = (! lizzieLet0_9QError_Bool_bufchan_buf[0]);
  assign lizzieLet0_9QError_Bool_1_argbuf_d = (lizzieLet0_9QError_Bool_bufchan_buf[0] ? lizzieLet0_9QError_Bool_bufchan_buf :
                                               lizzieLet0_9QError_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_9QError_Bool_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet0_9QError_Bool_1_argbuf_r && lizzieLet0_9QError_Bool_bufchan_buf[0]))
        lizzieLet0_9QError_Bool_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet0_9QError_Bool_1_argbuf_r) && (! lizzieLet0_9QError_Bool_bufchan_buf[0])))
        lizzieLet0_9QError_Bool_bufchan_buf <= lizzieLet0_9QError_Bool_bufchan_d;
  
  /* destruct (Ty QTree_Bool,
          Dcon QNode_Bool) : (lizzieLet45_1QNode_Bool,QTree_Bool) > [(q1a98_destruct,Pointer_QTree_Bool),
                                                                     (q2a99_destruct,Pointer_QTree_Bool),
                                                                     (q3a9a_destruct,Pointer_QTree_Bool),
                                                                     (q5a9b_destruct,Pointer_QTree_Bool)] */
  logic [3:0] lizzieLet45_1QNode_Bool_emitted;
  logic [3:0] lizzieLet45_1QNode_Bool_done;
  assign q1a98_destruct_d = {lizzieLet45_1QNode_Bool_d[18:3],
                             (lizzieLet45_1QNode_Bool_d[0] && (! lizzieLet45_1QNode_Bool_emitted[0]))};
  assign q2a99_destruct_d = {lizzieLet45_1QNode_Bool_d[34:19],
                             (lizzieLet45_1QNode_Bool_d[0] && (! lizzieLet45_1QNode_Bool_emitted[1]))};
  assign q3a9a_destruct_d = {lizzieLet45_1QNode_Bool_d[50:35],
                             (lizzieLet45_1QNode_Bool_d[0] && (! lizzieLet45_1QNode_Bool_emitted[2]))};
  assign q5a9b_destruct_d = {lizzieLet45_1QNode_Bool_d[66:51],
                             (lizzieLet45_1QNode_Bool_d[0] && (! lizzieLet45_1QNode_Bool_emitted[3]))};
  assign lizzieLet45_1QNode_Bool_done = (lizzieLet45_1QNode_Bool_emitted | ({q5a9b_destruct_d[0],
                                                                             q3a9a_destruct_d[0],
                                                                             q2a99_destruct_d[0],
                                                                             q1a98_destruct_d[0]} & {q5a9b_destruct_r,
                                                                                                     q3a9a_destruct_r,
                                                                                                     q2a99_destruct_r,
                                                                                                     q1a98_destruct_r}));
  assign lizzieLet45_1QNode_Bool_r = (& lizzieLet45_1QNode_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet45_1QNode_Bool_emitted <= 4'd0;
    else
      lizzieLet45_1QNode_Bool_emitted <= (lizzieLet45_1QNode_Bool_r ? 4'd0 :
                                          lizzieLet45_1QNode_Bool_done);
  
  /* destruct (Ty QTree_Bool,
          Dcon QVal_Bool) : (lizzieLet45_1QVal_Bool,QTree_Bool) > [(v1a92_destruct,MyBool)] */
  assign v1a92_destruct_d = {lizzieLet45_1QVal_Bool_d[3:3],
                             lizzieLet45_1QVal_Bool_d[0]};
  assign lizzieLet45_1QVal_Bool_r = v1a92_destruct_r;
  
  /* demux (Ty QTree_Bool,
       Ty QTree_Bool) : (lizzieLet45_2,QTree_Bool) (lizzieLet45_1,QTree_Bool) > [(_40,QTree_Bool),
                                                                                 (lizzieLet45_1QVal_Bool,QTree_Bool),
                                                                                 (lizzieLet45_1QNode_Bool,QTree_Bool),
                                                                                 (_39,QTree_Bool)] */
  logic [3:0] lizzieLet45_1_onehotd;
  always_comb
    if ((lizzieLet45_2_d[0] && lizzieLet45_1_d[0]))
      unique case (lizzieLet45_2_d[2:1])
        2'd0: lizzieLet45_1_onehotd = 4'd1;
        2'd1: lizzieLet45_1_onehotd = 4'd2;
        2'd2: lizzieLet45_1_onehotd = 4'd4;
        2'd3: lizzieLet45_1_onehotd = 4'd8;
        default: lizzieLet45_1_onehotd = 4'd0;
      endcase
    else lizzieLet45_1_onehotd = 4'd0;
  assign _40_d = {lizzieLet45_1_d[66:1], lizzieLet45_1_onehotd[0]};
  assign lizzieLet45_1QVal_Bool_d = {lizzieLet45_1_d[66:1],
                                     lizzieLet45_1_onehotd[1]};
  assign lizzieLet45_1QNode_Bool_d = {lizzieLet45_1_d[66:1],
                                      lizzieLet45_1_onehotd[2]};
  assign _39_d = {lizzieLet45_1_d[66:1], lizzieLet45_1_onehotd[3]};
  assign lizzieLet45_1_r = (| (lizzieLet45_1_onehotd & {_39_r,
                                                        lizzieLet45_1QNode_Bool_r,
                                                        lizzieLet45_1QVal_Bool_r,
                                                        _40_r}));
  assign lizzieLet45_2_r = lizzieLet45_1_r;
  
  /* demux (Ty QTree_Bool,
       Ty Go) : (lizzieLet45_3,QTree_Bool) (go_3_goMux_data,Go) > [(lizzieLet45_3QNone_Bool,Go),
                                                                   (lizzieLet45_3QVal_Bool,Go),
                                                                   (lizzieLet45_3QNode_Bool,Go),
                                                                   (lizzieLet45_3QError_Bool,Go)] */
  logic [3:0] go_3_goMux_data_onehotd;
  always_comb
    if ((lizzieLet45_3_d[0] && go_3_goMux_data_d[0]))
      unique case (lizzieLet45_3_d[2:1])
        2'd0: go_3_goMux_data_onehotd = 4'd1;
        2'd1: go_3_goMux_data_onehotd = 4'd2;
        2'd2: go_3_goMux_data_onehotd = 4'd4;
        2'd3: go_3_goMux_data_onehotd = 4'd8;
        default: go_3_goMux_data_onehotd = 4'd0;
      endcase
    else go_3_goMux_data_onehotd = 4'd0;
  assign lizzieLet45_3QNone_Bool_d = go_3_goMux_data_onehotd[0];
  assign lizzieLet45_3QVal_Bool_d = go_3_goMux_data_onehotd[1];
  assign lizzieLet45_3QNode_Bool_d = go_3_goMux_data_onehotd[2];
  assign lizzieLet45_3QError_Bool_d = go_3_goMux_data_onehotd[3];
  assign go_3_goMux_data_r = (| (go_3_goMux_data_onehotd & {lizzieLet45_3QError_Bool_r,
                                                            lizzieLet45_3QNode_Bool_r,
                                                            lizzieLet45_3QVal_Bool_r,
                                                            lizzieLet45_3QNone_Bool_r}));
  assign lizzieLet45_3_r = go_3_goMux_data_r;
  
  /* fork (Ty Go) : (lizzieLet45_3QError_Bool,Go) > [(lizzieLet45_3QError_Bool_1,Go),
                                                (lizzieLet45_3QError_Bool_2,Go)] */
  logic [1:0] lizzieLet45_3QError_Bool_emitted;
  logic [1:0] lizzieLet45_3QError_Bool_done;
  assign lizzieLet45_3QError_Bool_1_d = (lizzieLet45_3QError_Bool_d[0] && (! lizzieLet45_3QError_Bool_emitted[0]));
  assign lizzieLet45_3QError_Bool_2_d = (lizzieLet45_3QError_Bool_d[0] && (! lizzieLet45_3QError_Bool_emitted[1]));
  assign lizzieLet45_3QError_Bool_done = (lizzieLet45_3QError_Bool_emitted | ({lizzieLet45_3QError_Bool_2_d[0],
                                                                               lizzieLet45_3QError_Bool_1_d[0]} & {lizzieLet45_3QError_Bool_2_r,
                                                                                                                   lizzieLet45_3QError_Bool_1_r}));
  assign lizzieLet45_3QError_Bool_r = (& lizzieLet45_3QError_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet45_3QError_Bool_emitted <= 2'd0;
    else
      lizzieLet45_3QError_Bool_emitted <= (lizzieLet45_3QError_Bool_r ? 2'd0 :
                                           lizzieLet45_3QError_Bool_done);
  
  /* dcon (Ty QTree_Bool,
      Dcon QError_Bool) : [(lizzieLet45_3QError_Bool_1,Go)] > (lizzieLet45_3QError_Bool_1QError_Bool,QTree_Bool) */
  assign lizzieLet45_3QError_Bool_1QError_Bool_d = QError_Bool_dc((& {lizzieLet45_3QError_Bool_1_d[0]}), lizzieLet45_3QError_Bool_1_d);
  assign {lizzieLet45_3QError_Bool_1_r} = {1 {(lizzieLet45_3QError_Bool_1QError_Bool_r && lizzieLet45_3QError_Bool_1QError_Bool_d[0])}};
  
  /* buf (Ty QTree_Bool) : (lizzieLet45_3QError_Bool_1QError_Bool,QTree_Bool) > (lizzieLet56_1_argbuf,QTree_Bool) */
  QTree_Bool_t lizzieLet45_3QError_Bool_1QError_Bool_bufchan_d;
  logic lizzieLet45_3QError_Bool_1QError_Bool_bufchan_r;
  assign lizzieLet45_3QError_Bool_1QError_Bool_r = ((! lizzieLet45_3QError_Bool_1QError_Bool_bufchan_d[0]) || lizzieLet45_3QError_Bool_1QError_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet45_3QError_Bool_1QError_Bool_bufchan_d <= {66'd0, 1'd0};
    else
      if (lizzieLet45_3QError_Bool_1QError_Bool_r)
        lizzieLet45_3QError_Bool_1QError_Bool_bufchan_d <= lizzieLet45_3QError_Bool_1QError_Bool_d;
  QTree_Bool_t lizzieLet45_3QError_Bool_1QError_Bool_bufchan_buf;
  assign lizzieLet45_3QError_Bool_1QError_Bool_bufchan_r = (! lizzieLet45_3QError_Bool_1QError_Bool_bufchan_buf[0]);
  assign lizzieLet56_1_argbuf_d = (lizzieLet45_3QError_Bool_1QError_Bool_bufchan_buf[0] ? lizzieLet45_3QError_Bool_1QError_Bool_bufchan_buf :
                                   lizzieLet45_3QError_Bool_1QError_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet45_3QError_Bool_1QError_Bool_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((lizzieLet56_1_argbuf_r && lizzieLet45_3QError_Bool_1QError_Bool_bufchan_buf[0]))
        lizzieLet45_3QError_Bool_1QError_Bool_bufchan_buf <= {66'd0, 1'd0};
      else if (((! lizzieLet56_1_argbuf_r) && (! lizzieLet45_3QError_Bool_1QError_Bool_bufchan_buf[0])))
        lizzieLet45_3QError_Bool_1QError_Bool_bufchan_buf <= lizzieLet45_3QError_Bool_1QError_Bool_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet45_3QError_Bool_2,Go) > (lizzieLet45_3QError_Bool_2_argbuf,Go) */
  Go_t lizzieLet45_3QError_Bool_2_bufchan_d;
  logic lizzieLet45_3QError_Bool_2_bufchan_r;
  assign lizzieLet45_3QError_Bool_2_r = ((! lizzieLet45_3QError_Bool_2_bufchan_d[0]) || lizzieLet45_3QError_Bool_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet45_3QError_Bool_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet45_3QError_Bool_2_r)
        lizzieLet45_3QError_Bool_2_bufchan_d <= lizzieLet45_3QError_Bool_2_d;
  Go_t lizzieLet45_3QError_Bool_2_bufchan_buf;
  assign lizzieLet45_3QError_Bool_2_bufchan_r = (! lizzieLet45_3QError_Bool_2_bufchan_buf[0]);
  assign lizzieLet45_3QError_Bool_2_argbuf_d = (lizzieLet45_3QError_Bool_2_bufchan_buf[0] ? lizzieLet45_3QError_Bool_2_bufchan_buf :
                                                lizzieLet45_3QError_Bool_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet45_3QError_Bool_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet45_3QError_Bool_2_argbuf_r && lizzieLet45_3QError_Bool_2_bufchan_buf[0]))
        lizzieLet45_3QError_Bool_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet45_3QError_Bool_2_argbuf_r) && (! lizzieLet45_3QError_Bool_2_bufchan_buf[0])))
        lizzieLet45_3QError_Bool_2_bufchan_buf <= lizzieLet45_3QError_Bool_2_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet45_3QNone_Bool,Go) > (lizzieLet45_3QNone_Bool_1_argbuf,Go) */
  Go_t lizzieLet45_3QNone_Bool_bufchan_d;
  logic lizzieLet45_3QNone_Bool_bufchan_r;
  assign lizzieLet45_3QNone_Bool_r = ((! lizzieLet45_3QNone_Bool_bufchan_d[0]) || lizzieLet45_3QNone_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet45_3QNone_Bool_bufchan_d <= 1'd0;
    else
      if (lizzieLet45_3QNone_Bool_r)
        lizzieLet45_3QNone_Bool_bufchan_d <= lizzieLet45_3QNone_Bool_d;
  Go_t lizzieLet45_3QNone_Bool_bufchan_buf;
  assign lizzieLet45_3QNone_Bool_bufchan_r = (! lizzieLet45_3QNone_Bool_bufchan_buf[0]);
  assign lizzieLet45_3QNone_Bool_1_argbuf_d = (lizzieLet45_3QNone_Bool_bufchan_buf[0] ? lizzieLet45_3QNone_Bool_bufchan_buf :
                                               lizzieLet45_3QNone_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet45_3QNone_Bool_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet45_3QNone_Bool_1_argbuf_r && lizzieLet45_3QNone_Bool_bufchan_buf[0]))
        lizzieLet45_3QNone_Bool_bufchan_buf <= 1'd0;
      else if (((! lizzieLet45_3QNone_Bool_1_argbuf_r) && (! lizzieLet45_3QNone_Bool_bufchan_buf[0])))
        lizzieLet45_3QNone_Bool_bufchan_buf <= lizzieLet45_3QNone_Bool_bufchan_d;
  
  /* mergectrl (Ty C12,Ty Go) : [(lizzieLet45_3QNone_Bool_1_argbuf,Go),
                            (lizzieLet65_3Lcall_f''''''''''''0_1_argbuf,Go),
                            (lizzieLet45_4QVal_Bool_3QNone_Bool_1_argbuf,Go),
                            (lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_argbuf,Go),
                            (lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_argbuf,Go),
                            (lizzieLet45_4QVal_Bool_6QVal_Bool_1MyTrue_2_argbuf,Go),
                            (lizzieLet45_4QVal_Bool_3QNode_Bool_2_argbuf,Go),
                            (lizzieLet45_4QVal_Bool_3QError_Bool_2_argbuf,Go),
                            (lizzieLet45_4QNode_Bool_3QNone_Bool_1_argbuf,Go),
                            (lizzieLet45_4QNode_Bool_3QVal_Bool_2_argbuf,Go),
                            (lizzieLet45_4QNode_Bool_3QError_Bool_2_argbuf,Go),
                            (lizzieLet45_3QError_Bool_2_argbuf,Go)] > (go_8_goMux_choice,C12) (go_8_goMux_data,Go) */
  logic [11:0] lizzieLet45_3QNone_Bool_1_argbuf_select_d;
  assign lizzieLet45_3QNone_Bool_1_argbuf_select_d = ((| lizzieLet45_3QNone_Bool_1_argbuf_select_q) ? lizzieLet45_3QNone_Bool_1_argbuf_select_q :
                                                      (lizzieLet45_3QNone_Bool_1_argbuf_d[0] ? 12'd1 :
                                                       (\lizzieLet65_3Lcall_f''''''''''''0_1_argbuf_d [0] ? 12'd2 :
                                                        (lizzieLet45_4QVal_Bool_3QNone_Bool_1_argbuf_d[0] ? 12'd4 :
                                                         (lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_argbuf_d[0] ? 12'd8 :
                                                          (lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_argbuf_d[0] ? 12'd16 :
                                                           (lizzieLet45_4QVal_Bool_6QVal_Bool_1MyTrue_2_argbuf_d[0] ? 12'd32 :
                                                            (lizzieLet45_4QVal_Bool_3QNode_Bool_2_argbuf_d[0] ? 12'd64 :
                                                             (lizzieLet45_4QVal_Bool_3QError_Bool_2_argbuf_d[0] ? 12'd128 :
                                                              (lizzieLet45_4QNode_Bool_3QNone_Bool_1_argbuf_d[0] ? 12'd256 :
                                                               (lizzieLet45_4QNode_Bool_3QVal_Bool_2_argbuf_d[0] ? 12'd512 :
                                                                (lizzieLet45_4QNode_Bool_3QError_Bool_2_argbuf_d[0] ? 12'd1024 :
                                                                 (lizzieLet45_3QError_Bool_2_argbuf_d[0] ? 12'd2048 :
                                                                  12'd0)))))))))))));
  logic [11:0] lizzieLet45_3QNone_Bool_1_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet45_3QNone_Bool_1_argbuf_select_q <= 12'd0;
    else
      lizzieLet45_3QNone_Bool_1_argbuf_select_q <= (lizzieLet45_3QNone_Bool_1_argbuf_done ? 12'd0 :
                                                    lizzieLet45_3QNone_Bool_1_argbuf_select_d);
  logic [1:0] lizzieLet45_3QNone_Bool_1_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet45_3QNone_Bool_1_argbuf_emit_q <= 2'd0;
    else
      lizzieLet45_3QNone_Bool_1_argbuf_emit_q <= (lizzieLet45_3QNone_Bool_1_argbuf_done ? 2'd0 :
                                                  lizzieLet45_3QNone_Bool_1_argbuf_emit_d);
  logic [1:0] lizzieLet45_3QNone_Bool_1_argbuf_emit_d;
  assign lizzieLet45_3QNone_Bool_1_argbuf_emit_d = (lizzieLet45_3QNone_Bool_1_argbuf_emit_q | ({go_8_goMux_choice_d[0],
                                                                                                go_8_goMux_data_d[0]} & {go_8_goMux_choice_r,
                                                                                                                         go_8_goMux_data_r}));
  logic lizzieLet45_3QNone_Bool_1_argbuf_done;
  assign lizzieLet45_3QNone_Bool_1_argbuf_done = (& lizzieLet45_3QNone_Bool_1_argbuf_emit_d);
  assign {lizzieLet45_3QError_Bool_2_argbuf_r,
          lizzieLet45_4QNode_Bool_3QError_Bool_2_argbuf_r,
          lizzieLet45_4QNode_Bool_3QVal_Bool_2_argbuf_r,
          lizzieLet45_4QNode_Bool_3QNone_Bool_1_argbuf_r,
          lizzieLet45_4QVal_Bool_3QError_Bool_2_argbuf_r,
          lizzieLet45_4QVal_Bool_3QNode_Bool_2_argbuf_r,
          lizzieLet45_4QVal_Bool_6QVal_Bool_1MyTrue_2_argbuf_r,
          lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_argbuf_r,
          lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_argbuf_r,
          lizzieLet45_4QVal_Bool_3QNone_Bool_1_argbuf_r,
          \lizzieLet65_3Lcall_f''''''''''''0_1_argbuf_r ,
          lizzieLet45_3QNone_Bool_1_argbuf_r} = (lizzieLet45_3QNone_Bool_1_argbuf_done ? lizzieLet45_3QNone_Bool_1_argbuf_select_d :
                                                 12'd0);
  assign go_8_goMux_data_d = ((lizzieLet45_3QNone_Bool_1_argbuf_select_d[0] && (! lizzieLet45_3QNone_Bool_1_argbuf_emit_q[0])) ? lizzieLet45_3QNone_Bool_1_argbuf_d :
                              ((lizzieLet45_3QNone_Bool_1_argbuf_select_d[1] && (! lizzieLet45_3QNone_Bool_1_argbuf_emit_q[0])) ? \lizzieLet65_3Lcall_f''''''''''''0_1_argbuf_d  :
                               ((lizzieLet45_3QNone_Bool_1_argbuf_select_d[2] && (! lizzieLet45_3QNone_Bool_1_argbuf_emit_q[0])) ? lizzieLet45_4QVal_Bool_3QNone_Bool_1_argbuf_d :
                                ((lizzieLet45_3QNone_Bool_1_argbuf_select_d[3] && (! lizzieLet45_3QNone_Bool_1_argbuf_emit_q[0])) ? lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_argbuf_d :
                                 ((lizzieLet45_3QNone_Bool_1_argbuf_select_d[4] && (! lizzieLet45_3QNone_Bool_1_argbuf_emit_q[0])) ? lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_argbuf_d :
                                  ((lizzieLet45_3QNone_Bool_1_argbuf_select_d[5] && (! lizzieLet45_3QNone_Bool_1_argbuf_emit_q[0])) ? lizzieLet45_4QVal_Bool_6QVal_Bool_1MyTrue_2_argbuf_d :
                                   ((lizzieLet45_3QNone_Bool_1_argbuf_select_d[6] && (! lizzieLet45_3QNone_Bool_1_argbuf_emit_q[0])) ? lizzieLet45_4QVal_Bool_3QNode_Bool_2_argbuf_d :
                                    ((lizzieLet45_3QNone_Bool_1_argbuf_select_d[7] && (! lizzieLet45_3QNone_Bool_1_argbuf_emit_q[0])) ? lizzieLet45_4QVal_Bool_3QError_Bool_2_argbuf_d :
                                     ((lizzieLet45_3QNone_Bool_1_argbuf_select_d[8] && (! lizzieLet45_3QNone_Bool_1_argbuf_emit_q[0])) ? lizzieLet45_4QNode_Bool_3QNone_Bool_1_argbuf_d :
                                      ((lizzieLet45_3QNone_Bool_1_argbuf_select_d[9] && (! lizzieLet45_3QNone_Bool_1_argbuf_emit_q[0])) ? lizzieLet45_4QNode_Bool_3QVal_Bool_2_argbuf_d :
                                       ((lizzieLet45_3QNone_Bool_1_argbuf_select_d[10] && (! lizzieLet45_3QNone_Bool_1_argbuf_emit_q[0])) ? lizzieLet45_4QNode_Bool_3QError_Bool_2_argbuf_d :
                                        ((lizzieLet45_3QNone_Bool_1_argbuf_select_d[11] && (! lizzieLet45_3QNone_Bool_1_argbuf_emit_q[0])) ? lizzieLet45_3QError_Bool_2_argbuf_d :
                                         1'd0))))))))))));
  assign go_8_goMux_choice_d = ((lizzieLet45_3QNone_Bool_1_argbuf_select_d[0] && (! lizzieLet45_3QNone_Bool_1_argbuf_emit_q[1])) ? C1_12_dc(1'd1) :
                                ((lizzieLet45_3QNone_Bool_1_argbuf_select_d[1] && (! lizzieLet45_3QNone_Bool_1_argbuf_emit_q[1])) ? C2_12_dc(1'd1) :
                                 ((lizzieLet45_3QNone_Bool_1_argbuf_select_d[2] && (! lizzieLet45_3QNone_Bool_1_argbuf_emit_q[1])) ? C3_12_dc(1'd1) :
                                  ((lizzieLet45_3QNone_Bool_1_argbuf_select_d[3] && (! lizzieLet45_3QNone_Bool_1_argbuf_emit_q[1])) ? C4_12_dc(1'd1) :
                                   ((lizzieLet45_3QNone_Bool_1_argbuf_select_d[4] && (! lizzieLet45_3QNone_Bool_1_argbuf_emit_q[1])) ? C5_12_dc(1'd1) :
                                    ((lizzieLet45_3QNone_Bool_1_argbuf_select_d[5] && (! lizzieLet45_3QNone_Bool_1_argbuf_emit_q[1])) ? C6_12_dc(1'd1) :
                                     ((lizzieLet45_3QNone_Bool_1_argbuf_select_d[6] && (! lizzieLet45_3QNone_Bool_1_argbuf_emit_q[1])) ? C7_12_dc(1'd1) :
                                      ((lizzieLet45_3QNone_Bool_1_argbuf_select_d[7] && (! lizzieLet45_3QNone_Bool_1_argbuf_emit_q[1])) ? C8_12_dc(1'd1) :
                                       ((lizzieLet45_3QNone_Bool_1_argbuf_select_d[8] && (! lizzieLet45_3QNone_Bool_1_argbuf_emit_q[1])) ? C9_12_dc(1'd1) :
                                        ((lizzieLet45_3QNone_Bool_1_argbuf_select_d[9] && (! lizzieLet45_3QNone_Bool_1_argbuf_emit_q[1])) ? C10_12_dc(1'd1) :
                                         ((lizzieLet45_3QNone_Bool_1_argbuf_select_d[10] && (! lizzieLet45_3QNone_Bool_1_argbuf_emit_q[1])) ? C11_12_dc(1'd1) :
                                          ((lizzieLet45_3QNone_Bool_1_argbuf_select_d[11] && (! lizzieLet45_3QNone_Bool_1_argbuf_emit_q[1])) ? C12_12_dc(1'd1) :
                                           {4'd0, 1'd0}))))))))))));
  
  /* demux (Ty QTree_Bool,
       Ty QTree_Bool) : (lizzieLet45_4,QTree_Bool) (readPointer_QTree_Boolt4a91_1_argbuf_rwb,QTree_Bool) > [(_38,QTree_Bool),
                                                                                                            (lizzieLet45_4QVal_Bool,QTree_Bool),
                                                                                                            (lizzieLet45_4QNode_Bool,QTree_Bool),
                                                                                                            (_37,QTree_Bool)] */
  logic [3:0] readPointer_QTree_Boolt4a91_1_argbuf_rwb_onehotd;
  always_comb
    if ((lizzieLet45_4_d[0] && readPointer_QTree_Boolt4a91_1_argbuf_rwb_d[0]))
      unique case (lizzieLet45_4_d[2:1])
        2'd0: readPointer_QTree_Boolt4a91_1_argbuf_rwb_onehotd = 4'd1;
        2'd1: readPointer_QTree_Boolt4a91_1_argbuf_rwb_onehotd = 4'd2;
        2'd2: readPointer_QTree_Boolt4a91_1_argbuf_rwb_onehotd = 4'd4;
        2'd3: readPointer_QTree_Boolt4a91_1_argbuf_rwb_onehotd = 4'd8;
        default: readPointer_QTree_Boolt4a91_1_argbuf_rwb_onehotd = 4'd0;
      endcase
    else readPointer_QTree_Boolt4a91_1_argbuf_rwb_onehotd = 4'd0;
  assign _38_d = {readPointer_QTree_Boolt4a91_1_argbuf_rwb_d[66:1],
                  readPointer_QTree_Boolt4a91_1_argbuf_rwb_onehotd[0]};
  assign lizzieLet45_4QVal_Bool_d = {readPointer_QTree_Boolt4a91_1_argbuf_rwb_d[66:1],
                                     readPointer_QTree_Boolt4a91_1_argbuf_rwb_onehotd[1]};
  assign lizzieLet45_4QNode_Bool_d = {readPointer_QTree_Boolt4a91_1_argbuf_rwb_d[66:1],
                                      readPointer_QTree_Boolt4a91_1_argbuf_rwb_onehotd[2]};
  assign _37_d = {readPointer_QTree_Boolt4a91_1_argbuf_rwb_d[66:1],
                  readPointer_QTree_Boolt4a91_1_argbuf_rwb_onehotd[3]};
  assign readPointer_QTree_Boolt4a91_1_argbuf_rwb_r = (| (readPointer_QTree_Boolt4a91_1_argbuf_rwb_onehotd & {_37_r,
                                                                                                              lizzieLet45_4QNode_Bool_r,
                                                                                                              lizzieLet45_4QVal_Bool_r,
                                                                                                              _38_r}));
  assign lizzieLet45_4_r = readPointer_QTree_Boolt4a91_1_argbuf_rwb_r;
  
  /* fork (Ty QTree_Bool) : (lizzieLet45_4QNode_Bool,QTree_Bool) > [(lizzieLet45_4QNode_Bool_1,QTree_Bool),
                                                               (lizzieLet45_4QNode_Bool_2,QTree_Bool),
                                                               (lizzieLet45_4QNode_Bool_3,QTree_Bool),
                                                               (lizzieLet45_4QNode_Bool_4,QTree_Bool),
                                                               (lizzieLet45_4QNode_Bool_5,QTree_Bool),
                                                               (lizzieLet45_4QNode_Bool_6,QTree_Bool),
                                                               (lizzieLet45_4QNode_Bool_7,QTree_Bool),
                                                               (lizzieLet45_4QNode_Bool_8,QTree_Bool),
                                                               (lizzieLet45_4QNode_Bool_9,QTree_Bool)] */
  logic [8:0] lizzieLet45_4QNode_Bool_emitted;
  logic [8:0] lizzieLet45_4QNode_Bool_done;
  assign lizzieLet45_4QNode_Bool_1_d = {lizzieLet45_4QNode_Bool_d[66:1],
                                        (lizzieLet45_4QNode_Bool_d[0] && (! lizzieLet45_4QNode_Bool_emitted[0]))};
  assign lizzieLet45_4QNode_Bool_2_d = {lizzieLet45_4QNode_Bool_d[66:1],
                                        (lizzieLet45_4QNode_Bool_d[0] && (! lizzieLet45_4QNode_Bool_emitted[1]))};
  assign lizzieLet45_4QNode_Bool_3_d = {lizzieLet45_4QNode_Bool_d[66:1],
                                        (lizzieLet45_4QNode_Bool_d[0] && (! lizzieLet45_4QNode_Bool_emitted[2]))};
  assign lizzieLet45_4QNode_Bool_4_d = {lizzieLet45_4QNode_Bool_d[66:1],
                                        (lizzieLet45_4QNode_Bool_d[0] && (! lizzieLet45_4QNode_Bool_emitted[3]))};
  assign lizzieLet45_4QNode_Bool_5_d = {lizzieLet45_4QNode_Bool_d[66:1],
                                        (lizzieLet45_4QNode_Bool_d[0] && (! lizzieLet45_4QNode_Bool_emitted[4]))};
  assign lizzieLet45_4QNode_Bool_6_d = {lizzieLet45_4QNode_Bool_d[66:1],
                                        (lizzieLet45_4QNode_Bool_d[0] && (! lizzieLet45_4QNode_Bool_emitted[5]))};
  assign lizzieLet45_4QNode_Bool_7_d = {lizzieLet45_4QNode_Bool_d[66:1],
                                        (lizzieLet45_4QNode_Bool_d[0] && (! lizzieLet45_4QNode_Bool_emitted[6]))};
  assign lizzieLet45_4QNode_Bool_8_d = {lizzieLet45_4QNode_Bool_d[66:1],
                                        (lizzieLet45_4QNode_Bool_d[0] && (! lizzieLet45_4QNode_Bool_emitted[7]))};
  assign lizzieLet45_4QNode_Bool_9_d = {lizzieLet45_4QNode_Bool_d[66:1],
                                        (lizzieLet45_4QNode_Bool_d[0] && (! lizzieLet45_4QNode_Bool_emitted[8]))};
  assign lizzieLet45_4QNode_Bool_done = (lizzieLet45_4QNode_Bool_emitted | ({lizzieLet45_4QNode_Bool_9_d[0],
                                                                             lizzieLet45_4QNode_Bool_8_d[0],
                                                                             lizzieLet45_4QNode_Bool_7_d[0],
                                                                             lizzieLet45_4QNode_Bool_6_d[0],
                                                                             lizzieLet45_4QNode_Bool_5_d[0],
                                                                             lizzieLet45_4QNode_Bool_4_d[0],
                                                                             lizzieLet45_4QNode_Bool_3_d[0],
                                                                             lizzieLet45_4QNode_Bool_2_d[0],
                                                                             lizzieLet45_4QNode_Bool_1_d[0]} & {lizzieLet45_4QNode_Bool_9_r,
                                                                                                                lizzieLet45_4QNode_Bool_8_r,
                                                                                                                lizzieLet45_4QNode_Bool_7_r,
                                                                                                                lizzieLet45_4QNode_Bool_6_r,
                                                                                                                lizzieLet45_4QNode_Bool_5_r,
                                                                                                                lizzieLet45_4QNode_Bool_4_r,
                                                                                                                lizzieLet45_4QNode_Bool_3_r,
                                                                                                                lizzieLet45_4QNode_Bool_2_r,
                                                                                                                lizzieLet45_4QNode_Bool_1_r}));
  assign lizzieLet45_4QNode_Bool_r = (& lizzieLet45_4QNode_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet45_4QNode_Bool_emitted <= 9'd0;
    else
      lizzieLet45_4QNode_Bool_emitted <= (lizzieLet45_4QNode_Bool_r ? 9'd0 :
                                          lizzieLet45_4QNode_Bool_done);
  
  /* destruct (Ty QTree_Bool,
          Dcon QNode_Bool) : (lizzieLet45_4QNode_Bool_1QNode_Bool,QTree_Bool) > [(t1a9d_destruct,Pointer_QTree_Bool),
                                                                                 (t2a9e_destruct,Pointer_QTree_Bool),
                                                                                 (t3a9f_destruct,Pointer_QTree_Bool),
                                                                                 (t5a9g_destruct,Pointer_QTree_Bool)] */
  logic [3:0] lizzieLet45_4QNode_Bool_1QNode_Bool_emitted;
  logic [3:0] lizzieLet45_4QNode_Bool_1QNode_Bool_done;
  assign t1a9d_destruct_d = {lizzieLet45_4QNode_Bool_1QNode_Bool_d[18:3],
                             (lizzieLet45_4QNode_Bool_1QNode_Bool_d[0] && (! lizzieLet45_4QNode_Bool_1QNode_Bool_emitted[0]))};
  assign t2a9e_destruct_d = {lizzieLet45_4QNode_Bool_1QNode_Bool_d[34:19],
                             (lizzieLet45_4QNode_Bool_1QNode_Bool_d[0] && (! lizzieLet45_4QNode_Bool_1QNode_Bool_emitted[1]))};
  assign t3a9f_destruct_d = {lizzieLet45_4QNode_Bool_1QNode_Bool_d[50:35],
                             (lizzieLet45_4QNode_Bool_1QNode_Bool_d[0] && (! lizzieLet45_4QNode_Bool_1QNode_Bool_emitted[2]))};
  assign t5a9g_destruct_d = {lizzieLet45_4QNode_Bool_1QNode_Bool_d[66:51],
                             (lizzieLet45_4QNode_Bool_1QNode_Bool_d[0] && (! lizzieLet45_4QNode_Bool_1QNode_Bool_emitted[3]))};
  assign lizzieLet45_4QNode_Bool_1QNode_Bool_done = (lizzieLet45_4QNode_Bool_1QNode_Bool_emitted | ({t5a9g_destruct_d[0],
                                                                                                     t3a9f_destruct_d[0],
                                                                                                     t2a9e_destruct_d[0],
                                                                                                     t1a9d_destruct_d[0]} & {t5a9g_destruct_r,
                                                                                                                             t3a9f_destruct_r,
                                                                                                                             t2a9e_destruct_r,
                                                                                                                             t1a9d_destruct_r}));
  assign lizzieLet45_4QNode_Bool_1QNode_Bool_r = (& lizzieLet45_4QNode_Bool_1QNode_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet45_4QNode_Bool_1QNode_Bool_emitted <= 4'd0;
    else
      lizzieLet45_4QNode_Bool_1QNode_Bool_emitted <= (lizzieLet45_4QNode_Bool_1QNode_Bool_r ? 4'd0 :
                                                      lizzieLet45_4QNode_Bool_1QNode_Bool_done);
  
  /* demux (Ty QTree_Bool,
       Ty QTree_Bool) : (lizzieLet45_4QNode_Bool_2,QTree_Bool) (lizzieLet45_4QNode_Bool_1,QTree_Bool) > [(_36,QTree_Bool),
                                                                                                         (_35,QTree_Bool),
                                                                                                         (lizzieLet45_4QNode_Bool_1QNode_Bool,QTree_Bool),
                                                                                                         (_34,QTree_Bool)] */
  logic [3:0] lizzieLet45_4QNode_Bool_1_onehotd;
  always_comb
    if ((lizzieLet45_4QNode_Bool_2_d[0] && lizzieLet45_4QNode_Bool_1_d[0]))
      unique case (lizzieLet45_4QNode_Bool_2_d[2:1])
        2'd0: lizzieLet45_4QNode_Bool_1_onehotd = 4'd1;
        2'd1: lizzieLet45_4QNode_Bool_1_onehotd = 4'd2;
        2'd2: lizzieLet45_4QNode_Bool_1_onehotd = 4'd4;
        2'd3: lizzieLet45_4QNode_Bool_1_onehotd = 4'd8;
        default: lizzieLet45_4QNode_Bool_1_onehotd = 4'd0;
      endcase
    else lizzieLet45_4QNode_Bool_1_onehotd = 4'd0;
  assign _36_d = {lizzieLet45_4QNode_Bool_1_d[66:1],
                  lizzieLet45_4QNode_Bool_1_onehotd[0]};
  assign _35_d = {lizzieLet45_4QNode_Bool_1_d[66:1],
                  lizzieLet45_4QNode_Bool_1_onehotd[1]};
  assign lizzieLet45_4QNode_Bool_1QNode_Bool_d = {lizzieLet45_4QNode_Bool_1_d[66:1],
                                                  lizzieLet45_4QNode_Bool_1_onehotd[2]};
  assign _34_d = {lizzieLet45_4QNode_Bool_1_d[66:1],
                  lizzieLet45_4QNode_Bool_1_onehotd[3]};
  assign lizzieLet45_4QNode_Bool_1_r = (| (lizzieLet45_4QNode_Bool_1_onehotd & {_34_r,
                                                                                lizzieLet45_4QNode_Bool_1QNode_Bool_r,
                                                                                _35_r,
                                                                                _36_r}));
  assign lizzieLet45_4QNode_Bool_2_r = lizzieLet45_4QNode_Bool_1_r;
  
  /* demux (Ty QTree_Bool,
       Ty Go) : (lizzieLet45_4QNode_Bool_3,QTree_Bool) (lizzieLet45_3QNode_Bool,Go) > [(lizzieLet45_4QNode_Bool_3QNone_Bool,Go),
                                                                                       (lizzieLet45_4QNode_Bool_3QVal_Bool,Go),
                                                                                       (lizzieLet45_4QNode_Bool_3QNode_Bool,Go),
                                                                                       (lizzieLet45_4QNode_Bool_3QError_Bool,Go)] */
  logic [3:0] lizzieLet45_3QNode_Bool_onehotd;
  always_comb
    if ((lizzieLet45_4QNode_Bool_3_d[0] && lizzieLet45_3QNode_Bool_d[0]))
      unique case (lizzieLet45_4QNode_Bool_3_d[2:1])
        2'd0: lizzieLet45_3QNode_Bool_onehotd = 4'd1;
        2'd1: lizzieLet45_3QNode_Bool_onehotd = 4'd2;
        2'd2: lizzieLet45_3QNode_Bool_onehotd = 4'd4;
        2'd3: lizzieLet45_3QNode_Bool_onehotd = 4'd8;
        default: lizzieLet45_3QNode_Bool_onehotd = 4'd0;
      endcase
    else lizzieLet45_3QNode_Bool_onehotd = 4'd0;
  assign lizzieLet45_4QNode_Bool_3QNone_Bool_d = lizzieLet45_3QNode_Bool_onehotd[0];
  assign lizzieLet45_4QNode_Bool_3QVal_Bool_d = lizzieLet45_3QNode_Bool_onehotd[1];
  assign lizzieLet45_4QNode_Bool_3QNode_Bool_d = lizzieLet45_3QNode_Bool_onehotd[2];
  assign lizzieLet45_4QNode_Bool_3QError_Bool_d = lizzieLet45_3QNode_Bool_onehotd[3];
  assign lizzieLet45_3QNode_Bool_r = (| (lizzieLet45_3QNode_Bool_onehotd & {lizzieLet45_4QNode_Bool_3QError_Bool_r,
                                                                            lizzieLet45_4QNode_Bool_3QNode_Bool_r,
                                                                            lizzieLet45_4QNode_Bool_3QVal_Bool_r,
                                                                            lizzieLet45_4QNode_Bool_3QNone_Bool_r}));
  assign lizzieLet45_4QNode_Bool_3_r = lizzieLet45_3QNode_Bool_r;
  
  /* fork (Ty Go) : (lizzieLet45_4QNode_Bool_3QError_Bool,Go) > [(lizzieLet45_4QNode_Bool_3QError_Bool_1,Go),
                                                            (lizzieLet45_4QNode_Bool_3QError_Bool_2,Go)] */
  logic [1:0] lizzieLet45_4QNode_Bool_3QError_Bool_emitted;
  logic [1:0] lizzieLet45_4QNode_Bool_3QError_Bool_done;
  assign lizzieLet45_4QNode_Bool_3QError_Bool_1_d = (lizzieLet45_4QNode_Bool_3QError_Bool_d[0] && (! lizzieLet45_4QNode_Bool_3QError_Bool_emitted[0]));
  assign lizzieLet45_4QNode_Bool_3QError_Bool_2_d = (lizzieLet45_4QNode_Bool_3QError_Bool_d[0] && (! lizzieLet45_4QNode_Bool_3QError_Bool_emitted[1]));
  assign lizzieLet45_4QNode_Bool_3QError_Bool_done = (lizzieLet45_4QNode_Bool_3QError_Bool_emitted | ({lizzieLet45_4QNode_Bool_3QError_Bool_2_d[0],
                                                                                                       lizzieLet45_4QNode_Bool_3QError_Bool_1_d[0]} & {lizzieLet45_4QNode_Bool_3QError_Bool_2_r,
                                                                                                                                                       lizzieLet45_4QNode_Bool_3QError_Bool_1_r}));
  assign lizzieLet45_4QNode_Bool_3QError_Bool_r = (& lizzieLet45_4QNode_Bool_3QError_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet45_4QNode_Bool_3QError_Bool_emitted <= 2'd0;
    else
      lizzieLet45_4QNode_Bool_3QError_Bool_emitted <= (lizzieLet45_4QNode_Bool_3QError_Bool_r ? 2'd0 :
                                                       lizzieLet45_4QNode_Bool_3QError_Bool_done);
  
  /* dcon (Ty QTree_Bool,
      Dcon QError_Bool) : [(lizzieLet45_4QNode_Bool_3QError_Bool_1,Go)] > (lizzieLet45_4QNode_Bool_3QError_Bool_1QError_Bool,QTree_Bool) */
  assign lizzieLet45_4QNode_Bool_3QError_Bool_1QError_Bool_d = QError_Bool_dc((& {lizzieLet45_4QNode_Bool_3QError_Bool_1_d[0]}), lizzieLet45_4QNode_Bool_3QError_Bool_1_d);
  assign {lizzieLet45_4QNode_Bool_3QError_Bool_1_r} = {1 {(lizzieLet45_4QNode_Bool_3QError_Bool_1QError_Bool_r && lizzieLet45_4QNode_Bool_3QError_Bool_1QError_Bool_d[0])}};
  
  /* buf (Ty QTree_Bool) : (lizzieLet45_4QNode_Bool_3QError_Bool_1QError_Bool,QTree_Bool) > (lizzieLet55_1_argbuf,QTree_Bool) */
  QTree_Bool_t lizzieLet45_4QNode_Bool_3QError_Bool_1QError_Bool_bufchan_d;
  logic lizzieLet45_4QNode_Bool_3QError_Bool_1QError_Bool_bufchan_r;
  assign lizzieLet45_4QNode_Bool_3QError_Bool_1QError_Bool_r = ((! lizzieLet45_4QNode_Bool_3QError_Bool_1QError_Bool_bufchan_d[0]) || lizzieLet45_4QNode_Bool_3QError_Bool_1QError_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet45_4QNode_Bool_3QError_Bool_1QError_Bool_bufchan_d <= {66'd0,
                                                                      1'd0};
    else
      if (lizzieLet45_4QNode_Bool_3QError_Bool_1QError_Bool_r)
        lizzieLet45_4QNode_Bool_3QError_Bool_1QError_Bool_bufchan_d <= lizzieLet45_4QNode_Bool_3QError_Bool_1QError_Bool_d;
  QTree_Bool_t lizzieLet45_4QNode_Bool_3QError_Bool_1QError_Bool_bufchan_buf;
  assign lizzieLet45_4QNode_Bool_3QError_Bool_1QError_Bool_bufchan_r = (! lizzieLet45_4QNode_Bool_3QError_Bool_1QError_Bool_bufchan_buf[0]);
  assign lizzieLet55_1_argbuf_d = (lizzieLet45_4QNode_Bool_3QError_Bool_1QError_Bool_bufchan_buf[0] ? lizzieLet45_4QNode_Bool_3QError_Bool_1QError_Bool_bufchan_buf :
                                   lizzieLet45_4QNode_Bool_3QError_Bool_1QError_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet45_4QNode_Bool_3QError_Bool_1QError_Bool_bufchan_buf <= {66'd0,
                                                                        1'd0};
    else
      if ((lizzieLet55_1_argbuf_r && lizzieLet45_4QNode_Bool_3QError_Bool_1QError_Bool_bufchan_buf[0]))
        lizzieLet45_4QNode_Bool_3QError_Bool_1QError_Bool_bufchan_buf <= {66'd0,
                                                                          1'd0};
      else if (((! lizzieLet55_1_argbuf_r) && (! lizzieLet45_4QNode_Bool_3QError_Bool_1QError_Bool_bufchan_buf[0])))
        lizzieLet45_4QNode_Bool_3QError_Bool_1QError_Bool_bufchan_buf <= lizzieLet45_4QNode_Bool_3QError_Bool_1QError_Bool_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet45_4QNode_Bool_3QError_Bool_2,Go) > (lizzieLet45_4QNode_Bool_3QError_Bool_2_argbuf,Go) */
  Go_t lizzieLet45_4QNode_Bool_3QError_Bool_2_bufchan_d;
  logic lizzieLet45_4QNode_Bool_3QError_Bool_2_bufchan_r;
  assign lizzieLet45_4QNode_Bool_3QError_Bool_2_r = ((! lizzieLet45_4QNode_Bool_3QError_Bool_2_bufchan_d[0]) || lizzieLet45_4QNode_Bool_3QError_Bool_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet45_4QNode_Bool_3QError_Bool_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet45_4QNode_Bool_3QError_Bool_2_r)
        lizzieLet45_4QNode_Bool_3QError_Bool_2_bufchan_d <= lizzieLet45_4QNode_Bool_3QError_Bool_2_d;
  Go_t lizzieLet45_4QNode_Bool_3QError_Bool_2_bufchan_buf;
  assign lizzieLet45_4QNode_Bool_3QError_Bool_2_bufchan_r = (! lizzieLet45_4QNode_Bool_3QError_Bool_2_bufchan_buf[0]);
  assign lizzieLet45_4QNode_Bool_3QError_Bool_2_argbuf_d = (lizzieLet45_4QNode_Bool_3QError_Bool_2_bufchan_buf[0] ? lizzieLet45_4QNode_Bool_3QError_Bool_2_bufchan_buf :
                                                            lizzieLet45_4QNode_Bool_3QError_Bool_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet45_4QNode_Bool_3QError_Bool_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet45_4QNode_Bool_3QError_Bool_2_argbuf_r && lizzieLet45_4QNode_Bool_3QError_Bool_2_bufchan_buf[0]))
        lizzieLet45_4QNode_Bool_3QError_Bool_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet45_4QNode_Bool_3QError_Bool_2_argbuf_r) && (! lizzieLet45_4QNode_Bool_3QError_Bool_2_bufchan_buf[0])))
        lizzieLet45_4QNode_Bool_3QError_Bool_2_bufchan_buf <= lizzieLet45_4QNode_Bool_3QError_Bool_2_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet45_4QNode_Bool_3QNode_Bool,Go) > (lizzieLet45_4QNode_Bool_3QNode_Bool_1_argbuf,Go) */
  Go_t lizzieLet45_4QNode_Bool_3QNode_Bool_bufchan_d;
  logic lizzieLet45_4QNode_Bool_3QNode_Bool_bufchan_r;
  assign lizzieLet45_4QNode_Bool_3QNode_Bool_r = ((! lizzieLet45_4QNode_Bool_3QNode_Bool_bufchan_d[0]) || lizzieLet45_4QNode_Bool_3QNode_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet45_4QNode_Bool_3QNode_Bool_bufchan_d <= 1'd0;
    else
      if (lizzieLet45_4QNode_Bool_3QNode_Bool_r)
        lizzieLet45_4QNode_Bool_3QNode_Bool_bufchan_d <= lizzieLet45_4QNode_Bool_3QNode_Bool_d;
  Go_t lizzieLet45_4QNode_Bool_3QNode_Bool_bufchan_buf;
  assign lizzieLet45_4QNode_Bool_3QNode_Bool_bufchan_r = (! lizzieLet45_4QNode_Bool_3QNode_Bool_bufchan_buf[0]);
  assign lizzieLet45_4QNode_Bool_3QNode_Bool_1_argbuf_d = (lizzieLet45_4QNode_Bool_3QNode_Bool_bufchan_buf[0] ? lizzieLet45_4QNode_Bool_3QNode_Bool_bufchan_buf :
                                                           lizzieLet45_4QNode_Bool_3QNode_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet45_4QNode_Bool_3QNode_Bool_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet45_4QNode_Bool_3QNode_Bool_1_argbuf_r && lizzieLet45_4QNode_Bool_3QNode_Bool_bufchan_buf[0]))
        lizzieLet45_4QNode_Bool_3QNode_Bool_bufchan_buf <= 1'd0;
      else if (((! lizzieLet45_4QNode_Bool_3QNode_Bool_1_argbuf_r) && (! lizzieLet45_4QNode_Bool_3QNode_Bool_bufchan_buf[0])))
        lizzieLet45_4QNode_Bool_3QNode_Bool_bufchan_buf <= lizzieLet45_4QNode_Bool_3QNode_Bool_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet45_4QNode_Bool_3QNone_Bool,Go) > (lizzieLet45_4QNode_Bool_3QNone_Bool_1_argbuf,Go) */
  Go_t lizzieLet45_4QNode_Bool_3QNone_Bool_bufchan_d;
  logic lizzieLet45_4QNode_Bool_3QNone_Bool_bufchan_r;
  assign lizzieLet45_4QNode_Bool_3QNone_Bool_r = ((! lizzieLet45_4QNode_Bool_3QNone_Bool_bufchan_d[0]) || lizzieLet45_4QNode_Bool_3QNone_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet45_4QNode_Bool_3QNone_Bool_bufchan_d <= 1'd0;
    else
      if (lizzieLet45_4QNode_Bool_3QNone_Bool_r)
        lizzieLet45_4QNode_Bool_3QNone_Bool_bufchan_d <= lizzieLet45_4QNode_Bool_3QNone_Bool_d;
  Go_t lizzieLet45_4QNode_Bool_3QNone_Bool_bufchan_buf;
  assign lizzieLet45_4QNode_Bool_3QNone_Bool_bufchan_r = (! lizzieLet45_4QNode_Bool_3QNone_Bool_bufchan_buf[0]);
  assign lizzieLet45_4QNode_Bool_3QNone_Bool_1_argbuf_d = (lizzieLet45_4QNode_Bool_3QNone_Bool_bufchan_buf[0] ? lizzieLet45_4QNode_Bool_3QNone_Bool_bufchan_buf :
                                                           lizzieLet45_4QNode_Bool_3QNone_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet45_4QNode_Bool_3QNone_Bool_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet45_4QNode_Bool_3QNone_Bool_1_argbuf_r && lizzieLet45_4QNode_Bool_3QNone_Bool_bufchan_buf[0]))
        lizzieLet45_4QNode_Bool_3QNone_Bool_bufchan_buf <= 1'd0;
      else if (((! lizzieLet45_4QNode_Bool_3QNone_Bool_1_argbuf_r) && (! lizzieLet45_4QNode_Bool_3QNone_Bool_bufchan_buf[0])))
        lizzieLet45_4QNode_Bool_3QNone_Bool_bufchan_buf <= lizzieLet45_4QNode_Bool_3QNone_Bool_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet45_4QNode_Bool_3QVal_Bool,Go) > [(lizzieLet45_4QNode_Bool_3QVal_Bool_1,Go),
                                                          (lizzieLet45_4QNode_Bool_3QVal_Bool_2,Go)] */
  logic [1:0] lizzieLet45_4QNode_Bool_3QVal_Bool_emitted;
  logic [1:0] lizzieLet45_4QNode_Bool_3QVal_Bool_done;
  assign lizzieLet45_4QNode_Bool_3QVal_Bool_1_d = (lizzieLet45_4QNode_Bool_3QVal_Bool_d[0] && (! lizzieLet45_4QNode_Bool_3QVal_Bool_emitted[0]));
  assign lizzieLet45_4QNode_Bool_3QVal_Bool_2_d = (lizzieLet45_4QNode_Bool_3QVal_Bool_d[0] && (! lizzieLet45_4QNode_Bool_3QVal_Bool_emitted[1]));
  assign lizzieLet45_4QNode_Bool_3QVal_Bool_done = (lizzieLet45_4QNode_Bool_3QVal_Bool_emitted | ({lizzieLet45_4QNode_Bool_3QVal_Bool_2_d[0],
                                                                                                   lizzieLet45_4QNode_Bool_3QVal_Bool_1_d[0]} & {lizzieLet45_4QNode_Bool_3QVal_Bool_2_r,
                                                                                                                                                 lizzieLet45_4QNode_Bool_3QVal_Bool_1_r}));
  assign lizzieLet45_4QNode_Bool_3QVal_Bool_r = (& lizzieLet45_4QNode_Bool_3QVal_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet45_4QNode_Bool_3QVal_Bool_emitted <= 2'd0;
    else
      lizzieLet45_4QNode_Bool_3QVal_Bool_emitted <= (lizzieLet45_4QNode_Bool_3QVal_Bool_r ? 2'd0 :
                                                     lizzieLet45_4QNode_Bool_3QVal_Bool_done);
  
  /* dcon (Ty QTree_Bool,
      Dcon QError_Bool) : [(lizzieLet45_4QNode_Bool_3QVal_Bool_1,Go)] > (lizzieLet45_4QNode_Bool_3QVal_Bool_1QError_Bool,QTree_Bool) */
  assign lizzieLet45_4QNode_Bool_3QVal_Bool_1QError_Bool_d = QError_Bool_dc((& {lizzieLet45_4QNode_Bool_3QVal_Bool_1_d[0]}), lizzieLet45_4QNode_Bool_3QVal_Bool_1_d);
  assign {lizzieLet45_4QNode_Bool_3QVal_Bool_1_r} = {1 {(lizzieLet45_4QNode_Bool_3QVal_Bool_1QError_Bool_r && lizzieLet45_4QNode_Bool_3QVal_Bool_1QError_Bool_d[0])}};
  
  /* buf (Ty QTree_Bool) : (lizzieLet45_4QNode_Bool_3QVal_Bool_1QError_Bool,QTree_Bool) > (lizzieLet53_1_argbuf,QTree_Bool) */
  QTree_Bool_t lizzieLet45_4QNode_Bool_3QVal_Bool_1QError_Bool_bufchan_d;
  logic lizzieLet45_4QNode_Bool_3QVal_Bool_1QError_Bool_bufchan_r;
  assign lizzieLet45_4QNode_Bool_3QVal_Bool_1QError_Bool_r = ((! lizzieLet45_4QNode_Bool_3QVal_Bool_1QError_Bool_bufchan_d[0]) || lizzieLet45_4QNode_Bool_3QVal_Bool_1QError_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet45_4QNode_Bool_3QVal_Bool_1QError_Bool_bufchan_d <= {66'd0,
                                                                    1'd0};
    else
      if (lizzieLet45_4QNode_Bool_3QVal_Bool_1QError_Bool_r)
        lizzieLet45_4QNode_Bool_3QVal_Bool_1QError_Bool_bufchan_d <= lizzieLet45_4QNode_Bool_3QVal_Bool_1QError_Bool_d;
  QTree_Bool_t lizzieLet45_4QNode_Bool_3QVal_Bool_1QError_Bool_bufchan_buf;
  assign lizzieLet45_4QNode_Bool_3QVal_Bool_1QError_Bool_bufchan_r = (! lizzieLet45_4QNode_Bool_3QVal_Bool_1QError_Bool_bufchan_buf[0]);
  assign lizzieLet53_1_argbuf_d = (lizzieLet45_4QNode_Bool_3QVal_Bool_1QError_Bool_bufchan_buf[0] ? lizzieLet45_4QNode_Bool_3QVal_Bool_1QError_Bool_bufchan_buf :
                                   lizzieLet45_4QNode_Bool_3QVal_Bool_1QError_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet45_4QNode_Bool_3QVal_Bool_1QError_Bool_bufchan_buf <= {66'd0,
                                                                      1'd0};
    else
      if ((lizzieLet53_1_argbuf_r && lizzieLet45_4QNode_Bool_3QVal_Bool_1QError_Bool_bufchan_buf[0]))
        lizzieLet45_4QNode_Bool_3QVal_Bool_1QError_Bool_bufchan_buf <= {66'd0,
                                                                        1'd0};
      else if (((! lizzieLet53_1_argbuf_r) && (! lizzieLet45_4QNode_Bool_3QVal_Bool_1QError_Bool_bufchan_buf[0])))
        lizzieLet45_4QNode_Bool_3QVal_Bool_1QError_Bool_bufchan_buf <= lizzieLet45_4QNode_Bool_3QVal_Bool_1QError_Bool_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet45_4QNode_Bool_3QVal_Bool_2,Go) > (lizzieLet45_4QNode_Bool_3QVal_Bool_2_argbuf,Go) */
  Go_t lizzieLet45_4QNode_Bool_3QVal_Bool_2_bufchan_d;
  logic lizzieLet45_4QNode_Bool_3QVal_Bool_2_bufchan_r;
  assign lizzieLet45_4QNode_Bool_3QVal_Bool_2_r = ((! lizzieLet45_4QNode_Bool_3QVal_Bool_2_bufchan_d[0]) || lizzieLet45_4QNode_Bool_3QVal_Bool_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet45_4QNode_Bool_3QVal_Bool_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet45_4QNode_Bool_3QVal_Bool_2_r)
        lizzieLet45_4QNode_Bool_3QVal_Bool_2_bufchan_d <= lizzieLet45_4QNode_Bool_3QVal_Bool_2_d;
  Go_t lizzieLet45_4QNode_Bool_3QVal_Bool_2_bufchan_buf;
  assign lizzieLet45_4QNode_Bool_3QVal_Bool_2_bufchan_r = (! lizzieLet45_4QNode_Bool_3QVal_Bool_2_bufchan_buf[0]);
  assign lizzieLet45_4QNode_Bool_3QVal_Bool_2_argbuf_d = (lizzieLet45_4QNode_Bool_3QVal_Bool_2_bufchan_buf[0] ? lizzieLet45_4QNode_Bool_3QVal_Bool_2_bufchan_buf :
                                                          lizzieLet45_4QNode_Bool_3QVal_Bool_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet45_4QNode_Bool_3QVal_Bool_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet45_4QNode_Bool_3QVal_Bool_2_argbuf_r && lizzieLet45_4QNode_Bool_3QVal_Bool_2_bufchan_buf[0]))
        lizzieLet45_4QNode_Bool_3QVal_Bool_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet45_4QNode_Bool_3QVal_Bool_2_argbuf_r) && (! lizzieLet45_4QNode_Bool_3QVal_Bool_2_bufchan_buf[0])))
        lizzieLet45_4QNode_Bool_3QVal_Bool_2_bufchan_buf <= lizzieLet45_4QNode_Bool_3QVal_Bool_2_bufchan_d;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_QTree_Bool) : (lizzieLet45_4QNode_Bool_4,QTree_Bool) (lizzieLet45_5QNode_Bool,Pointer_QTree_Bool) > [(lizzieLet45_4QNode_Bool_4QNone_Bool,Pointer_QTree_Bool),
                                                                                                                       (_33,Pointer_QTree_Bool),
                                                                                                                       (_32,Pointer_QTree_Bool),
                                                                                                                       (_31,Pointer_QTree_Bool)] */
  logic [3:0] lizzieLet45_5QNode_Bool_onehotd;
  always_comb
    if ((lizzieLet45_4QNode_Bool_4_d[0] && lizzieLet45_5QNode_Bool_d[0]))
      unique case (lizzieLet45_4QNode_Bool_4_d[2:1])
        2'd0: lizzieLet45_5QNode_Bool_onehotd = 4'd1;
        2'd1: lizzieLet45_5QNode_Bool_onehotd = 4'd2;
        2'd2: lizzieLet45_5QNode_Bool_onehotd = 4'd4;
        2'd3: lizzieLet45_5QNode_Bool_onehotd = 4'd8;
        default: lizzieLet45_5QNode_Bool_onehotd = 4'd0;
      endcase
    else lizzieLet45_5QNode_Bool_onehotd = 4'd0;
  assign lizzieLet45_4QNode_Bool_4QNone_Bool_d = {lizzieLet45_5QNode_Bool_d[16:1],
                                                  lizzieLet45_5QNode_Bool_onehotd[0]};
  assign _33_d = {lizzieLet45_5QNode_Bool_d[16:1],
                  lizzieLet45_5QNode_Bool_onehotd[1]};
  assign _32_d = {lizzieLet45_5QNode_Bool_d[16:1],
                  lizzieLet45_5QNode_Bool_onehotd[2]};
  assign _31_d = {lizzieLet45_5QNode_Bool_d[16:1],
                  lizzieLet45_5QNode_Bool_onehotd[3]};
  assign lizzieLet45_5QNode_Bool_r = (| (lizzieLet45_5QNode_Bool_onehotd & {_31_r,
                                                                            _32_r,
                                                                            _33_r,
                                                                            lizzieLet45_4QNode_Bool_4QNone_Bool_r}));
  assign lizzieLet45_4QNode_Bool_4_r = lizzieLet45_5QNode_Bool_r;
  
  /* buf (Ty Pointer_QTree_Bool) : (lizzieLet45_4QNode_Bool_4QNone_Bool,Pointer_QTree_Bool) > (lizzieLet45_4QNode_Bool_4QNone_Bool_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t lizzieLet45_4QNode_Bool_4QNone_Bool_bufchan_d;
  logic lizzieLet45_4QNode_Bool_4QNone_Bool_bufchan_r;
  assign lizzieLet45_4QNode_Bool_4QNone_Bool_r = ((! lizzieLet45_4QNode_Bool_4QNone_Bool_bufchan_d[0]) || lizzieLet45_4QNode_Bool_4QNone_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet45_4QNode_Bool_4QNone_Bool_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet45_4QNode_Bool_4QNone_Bool_r)
        lizzieLet45_4QNode_Bool_4QNone_Bool_bufchan_d <= lizzieLet45_4QNode_Bool_4QNone_Bool_d;
  Pointer_QTree_Bool_t lizzieLet45_4QNode_Bool_4QNone_Bool_bufchan_buf;
  assign lizzieLet45_4QNode_Bool_4QNone_Bool_bufchan_r = (! lizzieLet45_4QNode_Bool_4QNone_Bool_bufchan_buf[0]);
  assign lizzieLet45_4QNode_Bool_4QNone_Bool_1_argbuf_d = (lizzieLet45_4QNode_Bool_4QNone_Bool_bufchan_buf[0] ? lizzieLet45_4QNode_Bool_4QNone_Bool_bufchan_buf :
                                                           lizzieLet45_4QNode_Bool_4QNone_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet45_4QNode_Bool_4QNone_Bool_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet45_4QNode_Bool_4QNone_Bool_1_argbuf_r && lizzieLet45_4QNode_Bool_4QNone_Bool_bufchan_buf[0]))
        lizzieLet45_4QNode_Bool_4QNone_Bool_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet45_4QNode_Bool_4QNone_Bool_1_argbuf_r) && (! lizzieLet45_4QNode_Bool_4QNone_Bool_bufchan_buf[0])))
        lizzieLet45_4QNode_Bool_4QNone_Bool_bufchan_buf <= lizzieLet45_4QNode_Bool_4QNone_Bool_bufchan_d;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_CTf'''''''''''') : (lizzieLet45_4QNode_Bool_5,QTree_Bool) (lizzieLet45_6QNode_Bool,Pointer_CTf'''''''''''') > [(lizzieLet45_4QNode_Bool_5QNone_Bool,Pointer_CTf''''''''''''),
                                                                                                                                 (lizzieLet45_4QNode_Bool_5QVal_Bool,Pointer_CTf''''''''''''),
                                                                                                                                 (lizzieLet45_4QNode_Bool_5QNode_Bool,Pointer_CTf''''''''''''),
                                                                                                                                 (lizzieLet45_4QNode_Bool_5QError_Bool,Pointer_CTf'''''''''''')] */
  logic [3:0] lizzieLet45_6QNode_Bool_onehotd;
  always_comb
    if ((lizzieLet45_4QNode_Bool_5_d[0] && lizzieLet45_6QNode_Bool_d[0]))
      unique case (lizzieLet45_4QNode_Bool_5_d[2:1])
        2'd0: lizzieLet45_6QNode_Bool_onehotd = 4'd1;
        2'd1: lizzieLet45_6QNode_Bool_onehotd = 4'd2;
        2'd2: lizzieLet45_6QNode_Bool_onehotd = 4'd4;
        2'd3: lizzieLet45_6QNode_Bool_onehotd = 4'd8;
        default: lizzieLet45_6QNode_Bool_onehotd = 4'd0;
      endcase
    else lizzieLet45_6QNode_Bool_onehotd = 4'd0;
  assign lizzieLet45_4QNode_Bool_5QNone_Bool_d = {lizzieLet45_6QNode_Bool_d[16:1],
                                                  lizzieLet45_6QNode_Bool_onehotd[0]};
  assign lizzieLet45_4QNode_Bool_5QVal_Bool_d = {lizzieLet45_6QNode_Bool_d[16:1],
                                                 lizzieLet45_6QNode_Bool_onehotd[1]};
  assign lizzieLet45_4QNode_Bool_5QNode_Bool_d = {lizzieLet45_6QNode_Bool_d[16:1],
                                                  lizzieLet45_6QNode_Bool_onehotd[2]};
  assign lizzieLet45_4QNode_Bool_5QError_Bool_d = {lizzieLet45_6QNode_Bool_d[16:1],
                                                   lizzieLet45_6QNode_Bool_onehotd[3]};
  assign lizzieLet45_6QNode_Bool_r = (| (lizzieLet45_6QNode_Bool_onehotd & {lizzieLet45_4QNode_Bool_5QError_Bool_r,
                                                                            lizzieLet45_4QNode_Bool_5QNode_Bool_r,
                                                                            lizzieLet45_4QNode_Bool_5QVal_Bool_r,
                                                                            lizzieLet45_4QNode_Bool_5QNone_Bool_r}));
  assign lizzieLet45_4QNode_Bool_5_r = lizzieLet45_6QNode_Bool_r;
  
  /* buf (Ty Pointer_CTf'''''''''''') : (lizzieLet45_4QNode_Bool_5QError_Bool,Pointer_CTf'''''''''''') > (lizzieLet45_4QNode_Bool_5QError_Bool_1_argbuf,Pointer_CTf'''''''''''') */
  \Pointer_CTf''''''''''''_t  lizzieLet45_4QNode_Bool_5QError_Bool_bufchan_d;
  logic lizzieLet45_4QNode_Bool_5QError_Bool_bufchan_r;
  assign lizzieLet45_4QNode_Bool_5QError_Bool_r = ((! lizzieLet45_4QNode_Bool_5QError_Bool_bufchan_d[0]) || lizzieLet45_4QNode_Bool_5QError_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet45_4QNode_Bool_5QError_Bool_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet45_4QNode_Bool_5QError_Bool_r)
        lizzieLet45_4QNode_Bool_5QError_Bool_bufchan_d <= lizzieLet45_4QNode_Bool_5QError_Bool_d;
  \Pointer_CTf''''''''''''_t  lizzieLet45_4QNode_Bool_5QError_Bool_bufchan_buf;
  assign lizzieLet45_4QNode_Bool_5QError_Bool_bufchan_r = (! lizzieLet45_4QNode_Bool_5QError_Bool_bufchan_buf[0]);
  assign lizzieLet45_4QNode_Bool_5QError_Bool_1_argbuf_d = (lizzieLet45_4QNode_Bool_5QError_Bool_bufchan_buf[0] ? lizzieLet45_4QNode_Bool_5QError_Bool_bufchan_buf :
                                                            lizzieLet45_4QNode_Bool_5QError_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet45_4QNode_Bool_5QError_Bool_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet45_4QNode_Bool_5QError_Bool_1_argbuf_r && lizzieLet45_4QNode_Bool_5QError_Bool_bufchan_buf[0]))
        lizzieLet45_4QNode_Bool_5QError_Bool_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet45_4QNode_Bool_5QError_Bool_1_argbuf_r) && (! lizzieLet45_4QNode_Bool_5QError_Bool_bufchan_buf[0])))
        lizzieLet45_4QNode_Bool_5QError_Bool_bufchan_buf <= lizzieLet45_4QNode_Bool_5QError_Bool_bufchan_d;
  
  /* dcon (Ty CTf'''''''''''',
      Dcon Lcall_f''''''''''''3) : [(lizzieLet45_4QNode_Bool_5QNode_Bool,Pointer_CTf''''''''''''),
                                    (lizzieLet45_4QNode_Bool_6QNode_Bool,Pointer_QTree_Bool),
                                    (t1a9d_destruct,Pointer_QTree_Bool),
                                    (lizzieLet45_4QNode_Bool_7QNode_Bool,Pointer_QTree_Bool),
                                    (t2a9e_destruct,Pointer_QTree_Bool),
                                    (lizzieLet45_4QNode_Bool_8QNode_Bool,Pointer_QTree_Bool),
                                    (t3a9f_destruct,Pointer_QTree_Bool)] > (lizzieLet45_4QNode_Bool_5QNode_Bool_1lizzieLet45_4QNode_Bool_6QNode_Bool_1t1a9d_1lizzieLet45_4QNode_Bool_7QNode_Bool_1t2a9e_1lizzieLet45_4QNode_Bool_8QNode_Bool_1t3a9f_1Lcall_f''''''''''''3,CTf'''''''''''') */
  assign \lizzieLet45_4QNode_Bool_5QNode_Bool_1lizzieLet45_4QNode_Bool_6QNode_Bool_1t1a9d_1lizzieLet45_4QNode_Bool_7QNode_Bool_1t2a9e_1lizzieLet45_4QNode_Bool_8QNode_Bool_1t3a9f_1Lcall_f''''''''''''3_d  = \Lcall_f''''''''''''3_dc ((& {lizzieLet45_4QNode_Bool_5QNode_Bool_d[0],
                                                                                                                                                                                                                                           lizzieLet45_4QNode_Bool_6QNode_Bool_d[0],
                                                                                                                                                                                                                                           t1a9d_destruct_d[0],
                                                                                                                                                                                                                                           lizzieLet45_4QNode_Bool_7QNode_Bool_d[0],
                                                                                                                                                                                                                                           t2a9e_destruct_d[0],
                                                                                                                                                                                                                                           lizzieLet45_4QNode_Bool_8QNode_Bool_d[0],
                                                                                                                                                                                                                                           t3a9f_destruct_d[0]}), lizzieLet45_4QNode_Bool_5QNode_Bool_d, lizzieLet45_4QNode_Bool_6QNode_Bool_d, t1a9d_destruct_d, lizzieLet45_4QNode_Bool_7QNode_Bool_d, t2a9e_destruct_d, lizzieLet45_4QNode_Bool_8QNode_Bool_d, t3a9f_destruct_d);
  assign {lizzieLet45_4QNode_Bool_5QNode_Bool_r,
          lizzieLet45_4QNode_Bool_6QNode_Bool_r,
          t1a9d_destruct_r,
          lizzieLet45_4QNode_Bool_7QNode_Bool_r,
          t2a9e_destruct_r,
          lizzieLet45_4QNode_Bool_8QNode_Bool_r,
          t3a9f_destruct_r} = {7 {(\lizzieLet45_4QNode_Bool_5QNode_Bool_1lizzieLet45_4QNode_Bool_6QNode_Bool_1t1a9d_1lizzieLet45_4QNode_Bool_7QNode_Bool_1t2a9e_1lizzieLet45_4QNode_Bool_8QNode_Bool_1t3a9f_1Lcall_f''''''''''''3_r  && \lizzieLet45_4QNode_Bool_5QNode_Bool_1lizzieLet45_4QNode_Bool_6QNode_Bool_1t1a9d_1lizzieLet45_4QNode_Bool_7QNode_Bool_1t2a9e_1lizzieLet45_4QNode_Bool_8QNode_Bool_1t3a9f_1Lcall_f''''''''''''3_d [0])}};
  
  /* buf (Ty CTf'''''''''''') : (lizzieLet45_4QNode_Bool_5QNode_Bool_1lizzieLet45_4QNode_Bool_6QNode_Bool_1t1a9d_1lizzieLet45_4QNode_Bool_7QNode_Bool_1t2a9e_1lizzieLet45_4QNode_Bool_8QNode_Bool_1t3a9f_1Lcall_f''''''''''''3,CTf'''''''''''') > (lizzieLet54_1_argbuf,CTf'''''''''''') */
  \CTf''''''''''''_t  \lizzieLet45_4QNode_Bool_5QNode_Bool_1lizzieLet45_4QNode_Bool_6QNode_Bool_1t1a9d_1lizzieLet45_4QNode_Bool_7QNode_Bool_1t2a9e_1lizzieLet45_4QNode_Bool_8QNode_Bool_1t3a9f_1Lcall_f''''''''''''3_bufchan_d ;
  logic \lizzieLet45_4QNode_Bool_5QNode_Bool_1lizzieLet45_4QNode_Bool_6QNode_Bool_1t1a9d_1lizzieLet45_4QNode_Bool_7QNode_Bool_1t2a9e_1lizzieLet45_4QNode_Bool_8QNode_Bool_1t3a9f_1Lcall_f''''''''''''3_bufchan_r ;
  assign \lizzieLet45_4QNode_Bool_5QNode_Bool_1lizzieLet45_4QNode_Bool_6QNode_Bool_1t1a9d_1lizzieLet45_4QNode_Bool_7QNode_Bool_1t2a9e_1lizzieLet45_4QNode_Bool_8QNode_Bool_1t3a9f_1Lcall_f''''''''''''3_r  = ((! \lizzieLet45_4QNode_Bool_5QNode_Bool_1lizzieLet45_4QNode_Bool_6QNode_Bool_1t1a9d_1lizzieLet45_4QNode_Bool_7QNode_Bool_1t2a9e_1lizzieLet45_4QNode_Bool_8QNode_Bool_1t3a9f_1Lcall_f''''''''''''3_bufchan_d [0]) || \lizzieLet45_4QNode_Bool_5QNode_Bool_1lizzieLet45_4QNode_Bool_6QNode_Bool_1t1a9d_1lizzieLet45_4QNode_Bool_7QNode_Bool_1t2a9e_1lizzieLet45_4QNode_Bool_8QNode_Bool_1t3a9f_1Lcall_f''''''''''''3_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet45_4QNode_Bool_5QNode_Bool_1lizzieLet45_4QNode_Bool_6QNode_Bool_1t1a9d_1lizzieLet45_4QNode_Bool_7QNode_Bool_1t2a9e_1lizzieLet45_4QNode_Bool_8QNode_Bool_1t3a9f_1Lcall_f''''''''''''3_bufchan_d  <= {115'd0,
                                                                                                                                                                                                                    1'd0};
    else
      if (\lizzieLet45_4QNode_Bool_5QNode_Bool_1lizzieLet45_4QNode_Bool_6QNode_Bool_1t1a9d_1lizzieLet45_4QNode_Bool_7QNode_Bool_1t2a9e_1lizzieLet45_4QNode_Bool_8QNode_Bool_1t3a9f_1Lcall_f''''''''''''3_r )
        \lizzieLet45_4QNode_Bool_5QNode_Bool_1lizzieLet45_4QNode_Bool_6QNode_Bool_1t1a9d_1lizzieLet45_4QNode_Bool_7QNode_Bool_1t2a9e_1lizzieLet45_4QNode_Bool_8QNode_Bool_1t3a9f_1Lcall_f''''''''''''3_bufchan_d  <= \lizzieLet45_4QNode_Bool_5QNode_Bool_1lizzieLet45_4QNode_Bool_6QNode_Bool_1t1a9d_1lizzieLet45_4QNode_Bool_7QNode_Bool_1t2a9e_1lizzieLet45_4QNode_Bool_8QNode_Bool_1t3a9f_1Lcall_f''''''''''''3_d ;
  \CTf''''''''''''_t  \lizzieLet45_4QNode_Bool_5QNode_Bool_1lizzieLet45_4QNode_Bool_6QNode_Bool_1t1a9d_1lizzieLet45_4QNode_Bool_7QNode_Bool_1t2a9e_1lizzieLet45_4QNode_Bool_8QNode_Bool_1t3a9f_1Lcall_f''''''''''''3_bufchan_buf ;
  assign \lizzieLet45_4QNode_Bool_5QNode_Bool_1lizzieLet45_4QNode_Bool_6QNode_Bool_1t1a9d_1lizzieLet45_4QNode_Bool_7QNode_Bool_1t2a9e_1lizzieLet45_4QNode_Bool_8QNode_Bool_1t3a9f_1Lcall_f''''''''''''3_bufchan_r  = (! \lizzieLet45_4QNode_Bool_5QNode_Bool_1lizzieLet45_4QNode_Bool_6QNode_Bool_1t1a9d_1lizzieLet45_4QNode_Bool_7QNode_Bool_1t2a9e_1lizzieLet45_4QNode_Bool_8QNode_Bool_1t3a9f_1Lcall_f''''''''''''3_bufchan_buf [0]);
  assign lizzieLet54_1_argbuf_d = (\lizzieLet45_4QNode_Bool_5QNode_Bool_1lizzieLet45_4QNode_Bool_6QNode_Bool_1t1a9d_1lizzieLet45_4QNode_Bool_7QNode_Bool_1t2a9e_1lizzieLet45_4QNode_Bool_8QNode_Bool_1t3a9f_1Lcall_f''''''''''''3_bufchan_buf [0] ? \lizzieLet45_4QNode_Bool_5QNode_Bool_1lizzieLet45_4QNode_Bool_6QNode_Bool_1t1a9d_1lizzieLet45_4QNode_Bool_7QNode_Bool_1t2a9e_1lizzieLet45_4QNode_Bool_8QNode_Bool_1t3a9f_1Lcall_f''''''''''''3_bufchan_buf  :
                                   \lizzieLet45_4QNode_Bool_5QNode_Bool_1lizzieLet45_4QNode_Bool_6QNode_Bool_1t1a9d_1lizzieLet45_4QNode_Bool_7QNode_Bool_1t2a9e_1lizzieLet45_4QNode_Bool_8QNode_Bool_1t3a9f_1Lcall_f''''''''''''3_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet45_4QNode_Bool_5QNode_Bool_1lizzieLet45_4QNode_Bool_6QNode_Bool_1t1a9d_1lizzieLet45_4QNode_Bool_7QNode_Bool_1t2a9e_1lizzieLet45_4QNode_Bool_8QNode_Bool_1t3a9f_1Lcall_f''''''''''''3_bufchan_buf  <= {115'd0,
                                                                                                                                                                                                                      1'd0};
    else
      if ((lizzieLet54_1_argbuf_r && \lizzieLet45_4QNode_Bool_5QNode_Bool_1lizzieLet45_4QNode_Bool_6QNode_Bool_1t1a9d_1lizzieLet45_4QNode_Bool_7QNode_Bool_1t2a9e_1lizzieLet45_4QNode_Bool_8QNode_Bool_1t3a9f_1Lcall_f''''''''''''3_bufchan_buf [0]))
        \lizzieLet45_4QNode_Bool_5QNode_Bool_1lizzieLet45_4QNode_Bool_6QNode_Bool_1t1a9d_1lizzieLet45_4QNode_Bool_7QNode_Bool_1t2a9e_1lizzieLet45_4QNode_Bool_8QNode_Bool_1t3a9f_1Lcall_f''''''''''''3_bufchan_buf  <= {115'd0,
                                                                                                                                                                                                                        1'd0};
      else if (((! lizzieLet54_1_argbuf_r) && (! \lizzieLet45_4QNode_Bool_5QNode_Bool_1lizzieLet45_4QNode_Bool_6QNode_Bool_1t1a9d_1lizzieLet45_4QNode_Bool_7QNode_Bool_1t2a9e_1lizzieLet45_4QNode_Bool_8QNode_Bool_1t3a9f_1Lcall_f''''''''''''3_bufchan_buf [0])))
        \lizzieLet45_4QNode_Bool_5QNode_Bool_1lizzieLet45_4QNode_Bool_6QNode_Bool_1t1a9d_1lizzieLet45_4QNode_Bool_7QNode_Bool_1t2a9e_1lizzieLet45_4QNode_Bool_8QNode_Bool_1t3a9f_1Lcall_f''''''''''''3_bufchan_buf  <= \lizzieLet45_4QNode_Bool_5QNode_Bool_1lizzieLet45_4QNode_Bool_6QNode_Bool_1t1a9d_1lizzieLet45_4QNode_Bool_7QNode_Bool_1t2a9e_1lizzieLet45_4QNode_Bool_8QNode_Bool_1t3a9f_1Lcall_f''''''''''''3_bufchan_d ;
  
  /* buf (Ty Pointer_CTf'''''''''''') : (lizzieLet45_4QNode_Bool_5QNone_Bool,Pointer_CTf'''''''''''') > (lizzieLet45_4QNode_Bool_5QNone_Bool_1_argbuf,Pointer_CTf'''''''''''') */
  \Pointer_CTf''''''''''''_t  lizzieLet45_4QNode_Bool_5QNone_Bool_bufchan_d;
  logic lizzieLet45_4QNode_Bool_5QNone_Bool_bufchan_r;
  assign lizzieLet45_4QNode_Bool_5QNone_Bool_r = ((! lizzieLet45_4QNode_Bool_5QNone_Bool_bufchan_d[0]) || lizzieLet45_4QNode_Bool_5QNone_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet45_4QNode_Bool_5QNone_Bool_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet45_4QNode_Bool_5QNone_Bool_r)
        lizzieLet45_4QNode_Bool_5QNone_Bool_bufchan_d <= lizzieLet45_4QNode_Bool_5QNone_Bool_d;
  \Pointer_CTf''''''''''''_t  lizzieLet45_4QNode_Bool_5QNone_Bool_bufchan_buf;
  assign lizzieLet45_4QNode_Bool_5QNone_Bool_bufchan_r = (! lizzieLet45_4QNode_Bool_5QNone_Bool_bufchan_buf[0]);
  assign lizzieLet45_4QNode_Bool_5QNone_Bool_1_argbuf_d = (lizzieLet45_4QNode_Bool_5QNone_Bool_bufchan_buf[0] ? lizzieLet45_4QNode_Bool_5QNone_Bool_bufchan_buf :
                                                           lizzieLet45_4QNode_Bool_5QNone_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet45_4QNode_Bool_5QNone_Bool_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet45_4QNode_Bool_5QNone_Bool_1_argbuf_r && lizzieLet45_4QNode_Bool_5QNone_Bool_bufchan_buf[0]))
        lizzieLet45_4QNode_Bool_5QNone_Bool_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet45_4QNode_Bool_5QNone_Bool_1_argbuf_r) && (! lizzieLet45_4QNode_Bool_5QNone_Bool_bufchan_buf[0])))
        lizzieLet45_4QNode_Bool_5QNone_Bool_bufchan_buf <= lizzieLet45_4QNode_Bool_5QNone_Bool_bufchan_d;
  
  /* buf (Ty Pointer_CTf'''''''''''') : (lizzieLet45_4QNode_Bool_5QVal_Bool,Pointer_CTf'''''''''''') > (lizzieLet45_4QNode_Bool_5QVal_Bool_1_argbuf,Pointer_CTf'''''''''''') */
  \Pointer_CTf''''''''''''_t  lizzieLet45_4QNode_Bool_5QVal_Bool_bufchan_d;
  logic lizzieLet45_4QNode_Bool_5QVal_Bool_bufchan_r;
  assign lizzieLet45_4QNode_Bool_5QVal_Bool_r = ((! lizzieLet45_4QNode_Bool_5QVal_Bool_bufchan_d[0]) || lizzieLet45_4QNode_Bool_5QVal_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet45_4QNode_Bool_5QVal_Bool_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet45_4QNode_Bool_5QVal_Bool_r)
        lizzieLet45_4QNode_Bool_5QVal_Bool_bufchan_d <= lizzieLet45_4QNode_Bool_5QVal_Bool_d;
  \Pointer_CTf''''''''''''_t  lizzieLet45_4QNode_Bool_5QVal_Bool_bufchan_buf;
  assign lizzieLet45_4QNode_Bool_5QVal_Bool_bufchan_r = (! lizzieLet45_4QNode_Bool_5QVal_Bool_bufchan_buf[0]);
  assign lizzieLet45_4QNode_Bool_5QVal_Bool_1_argbuf_d = (lizzieLet45_4QNode_Bool_5QVal_Bool_bufchan_buf[0] ? lizzieLet45_4QNode_Bool_5QVal_Bool_bufchan_buf :
                                                          lizzieLet45_4QNode_Bool_5QVal_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet45_4QNode_Bool_5QVal_Bool_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet45_4QNode_Bool_5QVal_Bool_1_argbuf_r && lizzieLet45_4QNode_Bool_5QVal_Bool_bufchan_buf[0]))
        lizzieLet45_4QNode_Bool_5QVal_Bool_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet45_4QNode_Bool_5QVal_Bool_1_argbuf_r) && (! lizzieLet45_4QNode_Bool_5QVal_Bool_bufchan_buf[0])))
        lizzieLet45_4QNode_Bool_5QVal_Bool_bufchan_buf <= lizzieLet45_4QNode_Bool_5QVal_Bool_bufchan_d;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_QTree_Bool) : (lizzieLet45_4QNode_Bool_6,QTree_Bool) (q1a98_destruct,Pointer_QTree_Bool) > [(_30,Pointer_QTree_Bool),
                                                                                                              (_29,Pointer_QTree_Bool),
                                                                                                              (lizzieLet45_4QNode_Bool_6QNode_Bool,Pointer_QTree_Bool),
                                                                                                              (_28,Pointer_QTree_Bool)] */
  logic [3:0] q1a98_destruct_onehotd;
  always_comb
    if ((lizzieLet45_4QNode_Bool_6_d[0] && q1a98_destruct_d[0]))
      unique case (lizzieLet45_4QNode_Bool_6_d[2:1])
        2'd0: q1a98_destruct_onehotd = 4'd1;
        2'd1: q1a98_destruct_onehotd = 4'd2;
        2'd2: q1a98_destruct_onehotd = 4'd4;
        2'd3: q1a98_destruct_onehotd = 4'd8;
        default: q1a98_destruct_onehotd = 4'd0;
      endcase
    else q1a98_destruct_onehotd = 4'd0;
  assign _30_d = {q1a98_destruct_d[16:1], q1a98_destruct_onehotd[0]};
  assign _29_d = {q1a98_destruct_d[16:1], q1a98_destruct_onehotd[1]};
  assign lizzieLet45_4QNode_Bool_6QNode_Bool_d = {q1a98_destruct_d[16:1],
                                                  q1a98_destruct_onehotd[2]};
  assign _28_d = {q1a98_destruct_d[16:1], q1a98_destruct_onehotd[3]};
  assign q1a98_destruct_r = (| (q1a98_destruct_onehotd & {_28_r,
                                                          lizzieLet45_4QNode_Bool_6QNode_Bool_r,
                                                          _29_r,
                                                          _30_r}));
  assign lizzieLet45_4QNode_Bool_6_r = q1a98_destruct_r;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_QTree_Bool) : (lizzieLet45_4QNode_Bool_7,QTree_Bool) (q2a99_destruct,Pointer_QTree_Bool) > [(_27,Pointer_QTree_Bool),
                                                                                                              (_26,Pointer_QTree_Bool),
                                                                                                              (lizzieLet45_4QNode_Bool_7QNode_Bool,Pointer_QTree_Bool),
                                                                                                              (_25,Pointer_QTree_Bool)] */
  logic [3:0] q2a99_destruct_onehotd;
  always_comb
    if ((lizzieLet45_4QNode_Bool_7_d[0] && q2a99_destruct_d[0]))
      unique case (lizzieLet45_4QNode_Bool_7_d[2:1])
        2'd0: q2a99_destruct_onehotd = 4'd1;
        2'd1: q2a99_destruct_onehotd = 4'd2;
        2'd2: q2a99_destruct_onehotd = 4'd4;
        2'd3: q2a99_destruct_onehotd = 4'd8;
        default: q2a99_destruct_onehotd = 4'd0;
      endcase
    else q2a99_destruct_onehotd = 4'd0;
  assign _27_d = {q2a99_destruct_d[16:1], q2a99_destruct_onehotd[0]};
  assign _26_d = {q2a99_destruct_d[16:1], q2a99_destruct_onehotd[1]};
  assign lizzieLet45_4QNode_Bool_7QNode_Bool_d = {q2a99_destruct_d[16:1],
                                                  q2a99_destruct_onehotd[2]};
  assign _25_d = {q2a99_destruct_d[16:1], q2a99_destruct_onehotd[3]};
  assign q2a99_destruct_r = (| (q2a99_destruct_onehotd & {_25_r,
                                                          lizzieLet45_4QNode_Bool_7QNode_Bool_r,
                                                          _26_r,
                                                          _27_r}));
  assign lizzieLet45_4QNode_Bool_7_r = q2a99_destruct_r;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_QTree_Bool) : (lizzieLet45_4QNode_Bool_8,QTree_Bool) (q3a9a_destruct,Pointer_QTree_Bool) > [(_24,Pointer_QTree_Bool),
                                                                                                              (_23,Pointer_QTree_Bool),
                                                                                                              (lizzieLet45_4QNode_Bool_8QNode_Bool,Pointer_QTree_Bool),
                                                                                                              (_22,Pointer_QTree_Bool)] */
  logic [3:0] q3a9a_destruct_onehotd;
  always_comb
    if ((lizzieLet45_4QNode_Bool_8_d[0] && q3a9a_destruct_d[0]))
      unique case (lizzieLet45_4QNode_Bool_8_d[2:1])
        2'd0: q3a9a_destruct_onehotd = 4'd1;
        2'd1: q3a9a_destruct_onehotd = 4'd2;
        2'd2: q3a9a_destruct_onehotd = 4'd4;
        2'd3: q3a9a_destruct_onehotd = 4'd8;
        default: q3a9a_destruct_onehotd = 4'd0;
      endcase
    else q3a9a_destruct_onehotd = 4'd0;
  assign _24_d = {q3a9a_destruct_d[16:1], q3a9a_destruct_onehotd[0]};
  assign _23_d = {q3a9a_destruct_d[16:1], q3a9a_destruct_onehotd[1]};
  assign lizzieLet45_4QNode_Bool_8QNode_Bool_d = {q3a9a_destruct_d[16:1],
                                                  q3a9a_destruct_onehotd[2]};
  assign _22_d = {q3a9a_destruct_d[16:1], q3a9a_destruct_onehotd[3]};
  assign q3a9a_destruct_r = (| (q3a9a_destruct_onehotd & {_22_r,
                                                          lizzieLet45_4QNode_Bool_8QNode_Bool_r,
                                                          _23_r,
                                                          _24_r}));
  assign lizzieLet45_4QNode_Bool_8_r = q3a9a_destruct_r;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_QTree_Bool) : (lizzieLet45_4QNode_Bool_9,QTree_Bool) (q5a9b_destruct,Pointer_QTree_Bool) > [(_21,Pointer_QTree_Bool),
                                                                                                              (_20,Pointer_QTree_Bool),
                                                                                                              (lizzieLet45_4QNode_Bool_9QNode_Bool,Pointer_QTree_Bool),
                                                                                                              (_19,Pointer_QTree_Bool)] */
  logic [3:0] q5a9b_destruct_onehotd;
  always_comb
    if ((lizzieLet45_4QNode_Bool_9_d[0] && q5a9b_destruct_d[0]))
      unique case (lizzieLet45_4QNode_Bool_9_d[2:1])
        2'd0: q5a9b_destruct_onehotd = 4'd1;
        2'd1: q5a9b_destruct_onehotd = 4'd2;
        2'd2: q5a9b_destruct_onehotd = 4'd4;
        2'd3: q5a9b_destruct_onehotd = 4'd8;
        default: q5a9b_destruct_onehotd = 4'd0;
      endcase
    else q5a9b_destruct_onehotd = 4'd0;
  assign _21_d = {q5a9b_destruct_d[16:1], q5a9b_destruct_onehotd[0]};
  assign _20_d = {q5a9b_destruct_d[16:1], q5a9b_destruct_onehotd[1]};
  assign lizzieLet45_4QNode_Bool_9QNode_Bool_d = {q5a9b_destruct_d[16:1],
                                                  q5a9b_destruct_onehotd[2]};
  assign _19_d = {q5a9b_destruct_d[16:1], q5a9b_destruct_onehotd[3]};
  assign q5a9b_destruct_r = (| (q5a9b_destruct_onehotd & {_19_r,
                                                          lizzieLet45_4QNode_Bool_9QNode_Bool_r,
                                                          _20_r,
                                                          _21_r}));
  assign lizzieLet45_4QNode_Bool_9_r = q5a9b_destruct_r;
  
  /* buf (Ty Pointer_QTree_Bool) : (lizzieLet45_4QNode_Bool_9QNode_Bool,Pointer_QTree_Bool) > (lizzieLet45_4QNode_Bool_9QNode_Bool_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t lizzieLet45_4QNode_Bool_9QNode_Bool_bufchan_d;
  logic lizzieLet45_4QNode_Bool_9QNode_Bool_bufchan_r;
  assign lizzieLet45_4QNode_Bool_9QNode_Bool_r = ((! lizzieLet45_4QNode_Bool_9QNode_Bool_bufchan_d[0]) || lizzieLet45_4QNode_Bool_9QNode_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet45_4QNode_Bool_9QNode_Bool_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet45_4QNode_Bool_9QNode_Bool_r)
        lizzieLet45_4QNode_Bool_9QNode_Bool_bufchan_d <= lizzieLet45_4QNode_Bool_9QNode_Bool_d;
  Pointer_QTree_Bool_t lizzieLet45_4QNode_Bool_9QNode_Bool_bufchan_buf;
  assign lizzieLet45_4QNode_Bool_9QNode_Bool_bufchan_r = (! lizzieLet45_4QNode_Bool_9QNode_Bool_bufchan_buf[0]);
  assign lizzieLet45_4QNode_Bool_9QNode_Bool_1_argbuf_d = (lizzieLet45_4QNode_Bool_9QNode_Bool_bufchan_buf[0] ? lizzieLet45_4QNode_Bool_9QNode_Bool_bufchan_buf :
                                                           lizzieLet45_4QNode_Bool_9QNode_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet45_4QNode_Bool_9QNode_Bool_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet45_4QNode_Bool_9QNode_Bool_1_argbuf_r && lizzieLet45_4QNode_Bool_9QNode_Bool_bufchan_buf[0]))
        lizzieLet45_4QNode_Bool_9QNode_Bool_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet45_4QNode_Bool_9QNode_Bool_1_argbuf_r) && (! lizzieLet45_4QNode_Bool_9QNode_Bool_bufchan_buf[0])))
        lizzieLet45_4QNode_Bool_9QNode_Bool_bufchan_buf <= lizzieLet45_4QNode_Bool_9QNode_Bool_bufchan_d;
  
  /* fork (Ty QTree_Bool) : (lizzieLet45_4QVal_Bool,QTree_Bool) > [(lizzieLet45_4QVal_Bool_1,QTree_Bool),
                                                              (lizzieLet45_4QVal_Bool_2,QTree_Bool),
                                                              (lizzieLet45_4QVal_Bool_3,QTree_Bool),
                                                              (lizzieLet45_4QVal_Bool_4,QTree_Bool),
                                                              (lizzieLet45_4QVal_Bool_5,QTree_Bool),
                                                              (lizzieLet45_4QVal_Bool_6,QTree_Bool)] */
  logic [5:0] lizzieLet45_4QVal_Bool_emitted;
  logic [5:0] lizzieLet45_4QVal_Bool_done;
  assign lizzieLet45_4QVal_Bool_1_d = {lizzieLet45_4QVal_Bool_d[66:1],
                                       (lizzieLet45_4QVal_Bool_d[0] && (! lizzieLet45_4QVal_Bool_emitted[0]))};
  assign lizzieLet45_4QVal_Bool_2_d = {lizzieLet45_4QVal_Bool_d[66:1],
                                       (lizzieLet45_4QVal_Bool_d[0] && (! lizzieLet45_4QVal_Bool_emitted[1]))};
  assign lizzieLet45_4QVal_Bool_3_d = {lizzieLet45_4QVal_Bool_d[66:1],
                                       (lizzieLet45_4QVal_Bool_d[0] && (! lizzieLet45_4QVal_Bool_emitted[2]))};
  assign lizzieLet45_4QVal_Bool_4_d = {lizzieLet45_4QVal_Bool_d[66:1],
                                       (lizzieLet45_4QVal_Bool_d[0] && (! lizzieLet45_4QVal_Bool_emitted[3]))};
  assign lizzieLet45_4QVal_Bool_5_d = {lizzieLet45_4QVal_Bool_d[66:1],
                                       (lizzieLet45_4QVal_Bool_d[0] && (! lizzieLet45_4QVal_Bool_emitted[4]))};
  assign lizzieLet45_4QVal_Bool_6_d = {lizzieLet45_4QVal_Bool_d[66:1],
                                       (lizzieLet45_4QVal_Bool_d[0] && (! lizzieLet45_4QVal_Bool_emitted[5]))};
  assign lizzieLet45_4QVal_Bool_done = (lizzieLet45_4QVal_Bool_emitted | ({lizzieLet45_4QVal_Bool_6_d[0],
                                                                           lizzieLet45_4QVal_Bool_5_d[0],
                                                                           lizzieLet45_4QVal_Bool_4_d[0],
                                                                           lizzieLet45_4QVal_Bool_3_d[0],
                                                                           lizzieLet45_4QVal_Bool_2_d[0],
                                                                           lizzieLet45_4QVal_Bool_1_d[0]} & {lizzieLet45_4QVal_Bool_6_r,
                                                                                                             lizzieLet45_4QVal_Bool_5_r,
                                                                                                             lizzieLet45_4QVal_Bool_4_r,
                                                                                                             lizzieLet45_4QVal_Bool_3_r,
                                                                                                             lizzieLet45_4QVal_Bool_2_r,
                                                                                                             lizzieLet45_4QVal_Bool_1_r}));
  assign lizzieLet45_4QVal_Bool_r = (& lizzieLet45_4QVal_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet45_4QVal_Bool_emitted <= 6'd0;
    else
      lizzieLet45_4QVal_Bool_emitted <= (lizzieLet45_4QVal_Bool_r ? 6'd0 :
                                         lizzieLet45_4QVal_Bool_done);
  
  /* destruct (Ty QTree_Bool,
          Dcon QVal_Bool) : (lizzieLet45_4QVal_Bool_1QVal_Bool,QTree_Bool) > [(va93_destruct,MyBool)] */
  assign va93_destruct_d = {lizzieLet45_4QVal_Bool_1QVal_Bool_d[3:3],
                            lizzieLet45_4QVal_Bool_1QVal_Bool_d[0]};
  assign lizzieLet45_4QVal_Bool_1QVal_Bool_r = va93_destruct_r;
  
  /* demux (Ty QTree_Bool,
       Ty QTree_Bool) : (lizzieLet45_4QVal_Bool_2,QTree_Bool) (lizzieLet45_4QVal_Bool_1,QTree_Bool) > [(_18,QTree_Bool),
                                                                                                       (lizzieLet45_4QVal_Bool_1QVal_Bool,QTree_Bool),
                                                                                                       (_17,QTree_Bool),
                                                                                                       (_16,QTree_Bool)] */
  logic [3:0] lizzieLet45_4QVal_Bool_1_onehotd;
  always_comb
    if ((lizzieLet45_4QVal_Bool_2_d[0] && lizzieLet45_4QVal_Bool_1_d[0]))
      unique case (lizzieLet45_4QVal_Bool_2_d[2:1])
        2'd0: lizzieLet45_4QVal_Bool_1_onehotd = 4'd1;
        2'd1: lizzieLet45_4QVal_Bool_1_onehotd = 4'd2;
        2'd2: lizzieLet45_4QVal_Bool_1_onehotd = 4'd4;
        2'd3: lizzieLet45_4QVal_Bool_1_onehotd = 4'd8;
        default: lizzieLet45_4QVal_Bool_1_onehotd = 4'd0;
      endcase
    else lizzieLet45_4QVal_Bool_1_onehotd = 4'd0;
  assign _18_d = {lizzieLet45_4QVal_Bool_1_d[66:1],
                  lizzieLet45_4QVal_Bool_1_onehotd[0]};
  assign lizzieLet45_4QVal_Bool_1QVal_Bool_d = {lizzieLet45_4QVal_Bool_1_d[66:1],
                                                lizzieLet45_4QVal_Bool_1_onehotd[1]};
  assign _17_d = {lizzieLet45_4QVal_Bool_1_d[66:1],
                  lizzieLet45_4QVal_Bool_1_onehotd[2]};
  assign _16_d = {lizzieLet45_4QVal_Bool_1_d[66:1],
                  lizzieLet45_4QVal_Bool_1_onehotd[3]};
  assign lizzieLet45_4QVal_Bool_1_r = (| (lizzieLet45_4QVal_Bool_1_onehotd & {_16_r,
                                                                              _17_r,
                                                                              lizzieLet45_4QVal_Bool_1QVal_Bool_r,
                                                                              _18_r}));
  assign lizzieLet45_4QVal_Bool_2_r = lizzieLet45_4QVal_Bool_1_r;
  
  /* demux (Ty QTree_Bool,
       Ty Go) : (lizzieLet45_4QVal_Bool_3,QTree_Bool) (lizzieLet45_3QVal_Bool,Go) > [(lizzieLet45_4QVal_Bool_3QNone_Bool,Go),
                                                                                     (lizzieLet45_4QVal_Bool_3QVal_Bool,Go),
                                                                                     (lizzieLet45_4QVal_Bool_3QNode_Bool,Go),
                                                                                     (lizzieLet45_4QVal_Bool_3QError_Bool,Go)] */
  logic [3:0] lizzieLet45_3QVal_Bool_onehotd;
  always_comb
    if ((lizzieLet45_4QVal_Bool_3_d[0] && lizzieLet45_3QVal_Bool_d[0]))
      unique case (lizzieLet45_4QVal_Bool_3_d[2:1])
        2'd0: lizzieLet45_3QVal_Bool_onehotd = 4'd1;
        2'd1: lizzieLet45_3QVal_Bool_onehotd = 4'd2;
        2'd2: lizzieLet45_3QVal_Bool_onehotd = 4'd4;
        2'd3: lizzieLet45_3QVal_Bool_onehotd = 4'd8;
        default: lizzieLet45_3QVal_Bool_onehotd = 4'd0;
      endcase
    else lizzieLet45_3QVal_Bool_onehotd = 4'd0;
  assign lizzieLet45_4QVal_Bool_3QNone_Bool_d = lizzieLet45_3QVal_Bool_onehotd[0];
  assign lizzieLet45_4QVal_Bool_3QVal_Bool_d = lizzieLet45_3QVal_Bool_onehotd[1];
  assign lizzieLet45_4QVal_Bool_3QNode_Bool_d = lizzieLet45_3QVal_Bool_onehotd[2];
  assign lizzieLet45_4QVal_Bool_3QError_Bool_d = lizzieLet45_3QVal_Bool_onehotd[3];
  assign lizzieLet45_3QVal_Bool_r = (| (lizzieLet45_3QVal_Bool_onehotd & {lizzieLet45_4QVal_Bool_3QError_Bool_r,
                                                                          lizzieLet45_4QVal_Bool_3QNode_Bool_r,
                                                                          lizzieLet45_4QVal_Bool_3QVal_Bool_r,
                                                                          lizzieLet45_4QVal_Bool_3QNone_Bool_r}));
  assign lizzieLet45_4QVal_Bool_3_r = lizzieLet45_3QVal_Bool_r;
  
  /* fork (Ty Go) : (lizzieLet45_4QVal_Bool_3QError_Bool,Go) > [(lizzieLet45_4QVal_Bool_3QError_Bool_1,Go),
                                                           (lizzieLet45_4QVal_Bool_3QError_Bool_2,Go)] */
  logic [1:0] lizzieLet45_4QVal_Bool_3QError_Bool_emitted;
  logic [1:0] lizzieLet45_4QVal_Bool_3QError_Bool_done;
  assign lizzieLet45_4QVal_Bool_3QError_Bool_1_d = (lizzieLet45_4QVal_Bool_3QError_Bool_d[0] && (! lizzieLet45_4QVal_Bool_3QError_Bool_emitted[0]));
  assign lizzieLet45_4QVal_Bool_3QError_Bool_2_d = (lizzieLet45_4QVal_Bool_3QError_Bool_d[0] && (! lizzieLet45_4QVal_Bool_3QError_Bool_emitted[1]));
  assign lizzieLet45_4QVal_Bool_3QError_Bool_done = (lizzieLet45_4QVal_Bool_3QError_Bool_emitted | ({lizzieLet45_4QVal_Bool_3QError_Bool_2_d[0],
                                                                                                     lizzieLet45_4QVal_Bool_3QError_Bool_1_d[0]} & {lizzieLet45_4QVal_Bool_3QError_Bool_2_r,
                                                                                                                                                    lizzieLet45_4QVal_Bool_3QError_Bool_1_r}));
  assign lizzieLet45_4QVal_Bool_3QError_Bool_r = (& lizzieLet45_4QVal_Bool_3QError_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet45_4QVal_Bool_3QError_Bool_emitted <= 2'd0;
    else
      lizzieLet45_4QVal_Bool_3QError_Bool_emitted <= (lizzieLet45_4QVal_Bool_3QError_Bool_r ? 2'd0 :
                                                      lizzieLet45_4QVal_Bool_3QError_Bool_done);
  
  /* dcon (Ty QTree_Bool,
      Dcon QError_Bool) : [(lizzieLet45_4QVal_Bool_3QError_Bool_1,Go)] > (lizzieLet45_4QVal_Bool_3QError_Bool_1QError_Bool,QTree_Bool) */
  assign lizzieLet45_4QVal_Bool_3QError_Bool_1QError_Bool_d = QError_Bool_dc((& {lizzieLet45_4QVal_Bool_3QError_Bool_1_d[0]}), lizzieLet45_4QVal_Bool_3QError_Bool_1_d);
  assign {lizzieLet45_4QVal_Bool_3QError_Bool_1_r} = {1 {(lizzieLet45_4QVal_Bool_3QError_Bool_1QError_Bool_r && lizzieLet45_4QVal_Bool_3QError_Bool_1QError_Bool_d[0])}};
  
  /* buf (Ty QTree_Bool) : (lizzieLet45_4QVal_Bool_3QError_Bool_1QError_Bool,QTree_Bool) > (lizzieLet51_1_argbuf,QTree_Bool) */
  QTree_Bool_t lizzieLet45_4QVal_Bool_3QError_Bool_1QError_Bool_bufchan_d;
  logic lizzieLet45_4QVal_Bool_3QError_Bool_1QError_Bool_bufchan_r;
  assign lizzieLet45_4QVal_Bool_3QError_Bool_1QError_Bool_r = ((! lizzieLet45_4QVal_Bool_3QError_Bool_1QError_Bool_bufchan_d[0]) || lizzieLet45_4QVal_Bool_3QError_Bool_1QError_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet45_4QVal_Bool_3QError_Bool_1QError_Bool_bufchan_d <= {66'd0,
                                                                     1'd0};
    else
      if (lizzieLet45_4QVal_Bool_3QError_Bool_1QError_Bool_r)
        lizzieLet45_4QVal_Bool_3QError_Bool_1QError_Bool_bufchan_d <= lizzieLet45_4QVal_Bool_3QError_Bool_1QError_Bool_d;
  QTree_Bool_t lizzieLet45_4QVal_Bool_3QError_Bool_1QError_Bool_bufchan_buf;
  assign lizzieLet45_4QVal_Bool_3QError_Bool_1QError_Bool_bufchan_r = (! lizzieLet45_4QVal_Bool_3QError_Bool_1QError_Bool_bufchan_buf[0]);
  assign lizzieLet51_1_argbuf_d = (lizzieLet45_4QVal_Bool_3QError_Bool_1QError_Bool_bufchan_buf[0] ? lizzieLet45_4QVal_Bool_3QError_Bool_1QError_Bool_bufchan_buf :
                                   lizzieLet45_4QVal_Bool_3QError_Bool_1QError_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet45_4QVal_Bool_3QError_Bool_1QError_Bool_bufchan_buf <= {66'd0,
                                                                       1'd0};
    else
      if ((lizzieLet51_1_argbuf_r && lizzieLet45_4QVal_Bool_3QError_Bool_1QError_Bool_bufchan_buf[0]))
        lizzieLet45_4QVal_Bool_3QError_Bool_1QError_Bool_bufchan_buf <= {66'd0,
                                                                         1'd0};
      else if (((! lizzieLet51_1_argbuf_r) && (! lizzieLet45_4QVal_Bool_3QError_Bool_1QError_Bool_bufchan_buf[0])))
        lizzieLet45_4QVal_Bool_3QError_Bool_1QError_Bool_bufchan_buf <= lizzieLet45_4QVal_Bool_3QError_Bool_1QError_Bool_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet45_4QVal_Bool_3QError_Bool_2,Go) > (lizzieLet45_4QVal_Bool_3QError_Bool_2_argbuf,Go) */
  Go_t lizzieLet45_4QVal_Bool_3QError_Bool_2_bufchan_d;
  logic lizzieLet45_4QVal_Bool_3QError_Bool_2_bufchan_r;
  assign lizzieLet45_4QVal_Bool_3QError_Bool_2_r = ((! lizzieLet45_4QVal_Bool_3QError_Bool_2_bufchan_d[0]) || lizzieLet45_4QVal_Bool_3QError_Bool_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet45_4QVal_Bool_3QError_Bool_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet45_4QVal_Bool_3QError_Bool_2_r)
        lizzieLet45_4QVal_Bool_3QError_Bool_2_bufchan_d <= lizzieLet45_4QVal_Bool_3QError_Bool_2_d;
  Go_t lizzieLet45_4QVal_Bool_3QError_Bool_2_bufchan_buf;
  assign lizzieLet45_4QVal_Bool_3QError_Bool_2_bufchan_r = (! lizzieLet45_4QVal_Bool_3QError_Bool_2_bufchan_buf[0]);
  assign lizzieLet45_4QVal_Bool_3QError_Bool_2_argbuf_d = (lizzieLet45_4QVal_Bool_3QError_Bool_2_bufchan_buf[0] ? lizzieLet45_4QVal_Bool_3QError_Bool_2_bufchan_buf :
                                                           lizzieLet45_4QVal_Bool_3QError_Bool_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet45_4QVal_Bool_3QError_Bool_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet45_4QVal_Bool_3QError_Bool_2_argbuf_r && lizzieLet45_4QVal_Bool_3QError_Bool_2_bufchan_buf[0]))
        lizzieLet45_4QVal_Bool_3QError_Bool_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet45_4QVal_Bool_3QError_Bool_2_argbuf_r) && (! lizzieLet45_4QVal_Bool_3QError_Bool_2_bufchan_buf[0])))
        lizzieLet45_4QVal_Bool_3QError_Bool_2_bufchan_buf <= lizzieLet45_4QVal_Bool_3QError_Bool_2_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet45_4QVal_Bool_3QNode_Bool,Go) > [(lizzieLet45_4QVal_Bool_3QNode_Bool_1,Go),
                                                          (lizzieLet45_4QVal_Bool_3QNode_Bool_2,Go)] */
  logic [1:0] lizzieLet45_4QVal_Bool_3QNode_Bool_emitted;
  logic [1:0] lizzieLet45_4QVal_Bool_3QNode_Bool_done;
  assign lizzieLet45_4QVal_Bool_3QNode_Bool_1_d = (lizzieLet45_4QVal_Bool_3QNode_Bool_d[0] && (! lizzieLet45_4QVal_Bool_3QNode_Bool_emitted[0]));
  assign lizzieLet45_4QVal_Bool_3QNode_Bool_2_d = (lizzieLet45_4QVal_Bool_3QNode_Bool_d[0] && (! lizzieLet45_4QVal_Bool_3QNode_Bool_emitted[1]));
  assign lizzieLet45_4QVal_Bool_3QNode_Bool_done = (lizzieLet45_4QVal_Bool_3QNode_Bool_emitted | ({lizzieLet45_4QVal_Bool_3QNode_Bool_2_d[0],
                                                                                                   lizzieLet45_4QVal_Bool_3QNode_Bool_1_d[0]} & {lizzieLet45_4QVal_Bool_3QNode_Bool_2_r,
                                                                                                                                                 lizzieLet45_4QVal_Bool_3QNode_Bool_1_r}));
  assign lizzieLet45_4QVal_Bool_3QNode_Bool_r = (& lizzieLet45_4QVal_Bool_3QNode_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet45_4QVal_Bool_3QNode_Bool_emitted <= 2'd0;
    else
      lizzieLet45_4QVal_Bool_3QNode_Bool_emitted <= (lizzieLet45_4QVal_Bool_3QNode_Bool_r ? 2'd0 :
                                                     lizzieLet45_4QVal_Bool_3QNode_Bool_done);
  
  /* dcon (Ty QTree_Bool,
      Dcon QError_Bool) : [(lizzieLet45_4QVal_Bool_3QNode_Bool_1,Go)] > (lizzieLet45_4QVal_Bool_3QNode_Bool_1QError_Bool,QTree_Bool) */
  assign lizzieLet45_4QVal_Bool_3QNode_Bool_1QError_Bool_d = QError_Bool_dc((& {lizzieLet45_4QVal_Bool_3QNode_Bool_1_d[0]}), lizzieLet45_4QVal_Bool_3QNode_Bool_1_d);
  assign {lizzieLet45_4QVal_Bool_3QNode_Bool_1_r} = {1 {(lizzieLet45_4QVal_Bool_3QNode_Bool_1QError_Bool_r && lizzieLet45_4QVal_Bool_3QNode_Bool_1QError_Bool_d[0])}};
  
  /* buf (Ty QTree_Bool) : (lizzieLet45_4QVal_Bool_3QNode_Bool_1QError_Bool,QTree_Bool) > (lizzieLet50_1_argbuf,QTree_Bool) */
  QTree_Bool_t lizzieLet45_4QVal_Bool_3QNode_Bool_1QError_Bool_bufchan_d;
  logic lizzieLet45_4QVal_Bool_3QNode_Bool_1QError_Bool_bufchan_r;
  assign lizzieLet45_4QVal_Bool_3QNode_Bool_1QError_Bool_r = ((! lizzieLet45_4QVal_Bool_3QNode_Bool_1QError_Bool_bufchan_d[0]) || lizzieLet45_4QVal_Bool_3QNode_Bool_1QError_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet45_4QVal_Bool_3QNode_Bool_1QError_Bool_bufchan_d <= {66'd0,
                                                                    1'd0};
    else
      if (lizzieLet45_4QVal_Bool_3QNode_Bool_1QError_Bool_r)
        lizzieLet45_4QVal_Bool_3QNode_Bool_1QError_Bool_bufchan_d <= lizzieLet45_4QVal_Bool_3QNode_Bool_1QError_Bool_d;
  QTree_Bool_t lizzieLet45_4QVal_Bool_3QNode_Bool_1QError_Bool_bufchan_buf;
  assign lizzieLet45_4QVal_Bool_3QNode_Bool_1QError_Bool_bufchan_r = (! lizzieLet45_4QVal_Bool_3QNode_Bool_1QError_Bool_bufchan_buf[0]);
  assign lizzieLet50_1_argbuf_d = (lizzieLet45_4QVal_Bool_3QNode_Bool_1QError_Bool_bufchan_buf[0] ? lizzieLet45_4QVal_Bool_3QNode_Bool_1QError_Bool_bufchan_buf :
                                   lizzieLet45_4QVal_Bool_3QNode_Bool_1QError_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet45_4QVal_Bool_3QNode_Bool_1QError_Bool_bufchan_buf <= {66'd0,
                                                                      1'd0};
    else
      if ((lizzieLet50_1_argbuf_r && lizzieLet45_4QVal_Bool_3QNode_Bool_1QError_Bool_bufchan_buf[0]))
        lizzieLet45_4QVal_Bool_3QNode_Bool_1QError_Bool_bufchan_buf <= {66'd0,
                                                                        1'd0};
      else if (((! lizzieLet50_1_argbuf_r) && (! lizzieLet45_4QVal_Bool_3QNode_Bool_1QError_Bool_bufchan_buf[0])))
        lizzieLet45_4QVal_Bool_3QNode_Bool_1QError_Bool_bufchan_buf <= lizzieLet45_4QVal_Bool_3QNode_Bool_1QError_Bool_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet45_4QVal_Bool_3QNode_Bool_2,Go) > (lizzieLet45_4QVal_Bool_3QNode_Bool_2_argbuf,Go) */
  Go_t lizzieLet45_4QVal_Bool_3QNode_Bool_2_bufchan_d;
  logic lizzieLet45_4QVal_Bool_3QNode_Bool_2_bufchan_r;
  assign lizzieLet45_4QVal_Bool_3QNode_Bool_2_r = ((! lizzieLet45_4QVal_Bool_3QNode_Bool_2_bufchan_d[0]) || lizzieLet45_4QVal_Bool_3QNode_Bool_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet45_4QVal_Bool_3QNode_Bool_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet45_4QVal_Bool_3QNode_Bool_2_r)
        lizzieLet45_4QVal_Bool_3QNode_Bool_2_bufchan_d <= lizzieLet45_4QVal_Bool_3QNode_Bool_2_d;
  Go_t lizzieLet45_4QVal_Bool_3QNode_Bool_2_bufchan_buf;
  assign lizzieLet45_4QVal_Bool_3QNode_Bool_2_bufchan_r = (! lizzieLet45_4QVal_Bool_3QNode_Bool_2_bufchan_buf[0]);
  assign lizzieLet45_4QVal_Bool_3QNode_Bool_2_argbuf_d = (lizzieLet45_4QVal_Bool_3QNode_Bool_2_bufchan_buf[0] ? lizzieLet45_4QVal_Bool_3QNode_Bool_2_bufchan_buf :
                                                          lizzieLet45_4QVal_Bool_3QNode_Bool_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet45_4QVal_Bool_3QNode_Bool_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet45_4QVal_Bool_3QNode_Bool_2_argbuf_r && lizzieLet45_4QVal_Bool_3QNode_Bool_2_bufchan_buf[0]))
        lizzieLet45_4QVal_Bool_3QNode_Bool_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet45_4QVal_Bool_3QNode_Bool_2_argbuf_r) && (! lizzieLet45_4QVal_Bool_3QNode_Bool_2_bufchan_buf[0])))
        lizzieLet45_4QVal_Bool_3QNode_Bool_2_bufchan_buf <= lizzieLet45_4QVal_Bool_3QNode_Bool_2_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet45_4QVal_Bool_3QNone_Bool,Go) > (lizzieLet45_4QVal_Bool_3QNone_Bool_1_argbuf,Go) */
  Go_t lizzieLet45_4QVal_Bool_3QNone_Bool_bufchan_d;
  logic lizzieLet45_4QVal_Bool_3QNone_Bool_bufchan_r;
  assign lizzieLet45_4QVal_Bool_3QNone_Bool_r = ((! lizzieLet45_4QVal_Bool_3QNone_Bool_bufchan_d[0]) || lizzieLet45_4QVal_Bool_3QNone_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet45_4QVal_Bool_3QNone_Bool_bufchan_d <= 1'd0;
    else
      if (lizzieLet45_4QVal_Bool_3QNone_Bool_r)
        lizzieLet45_4QVal_Bool_3QNone_Bool_bufchan_d <= lizzieLet45_4QVal_Bool_3QNone_Bool_d;
  Go_t lizzieLet45_4QVal_Bool_3QNone_Bool_bufchan_buf;
  assign lizzieLet45_4QVal_Bool_3QNone_Bool_bufchan_r = (! lizzieLet45_4QVal_Bool_3QNone_Bool_bufchan_buf[0]);
  assign lizzieLet45_4QVal_Bool_3QNone_Bool_1_argbuf_d = (lizzieLet45_4QVal_Bool_3QNone_Bool_bufchan_buf[0] ? lizzieLet45_4QVal_Bool_3QNone_Bool_bufchan_buf :
                                                          lizzieLet45_4QVal_Bool_3QNone_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet45_4QVal_Bool_3QNone_Bool_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet45_4QVal_Bool_3QNone_Bool_1_argbuf_r && lizzieLet45_4QVal_Bool_3QNone_Bool_bufchan_buf[0]))
        lizzieLet45_4QVal_Bool_3QNone_Bool_bufchan_buf <= 1'd0;
      else if (((! lizzieLet45_4QVal_Bool_3QNone_Bool_1_argbuf_r) && (! lizzieLet45_4QVal_Bool_3QNone_Bool_bufchan_buf[0])))
        lizzieLet45_4QVal_Bool_3QNone_Bool_bufchan_buf <= lizzieLet45_4QVal_Bool_3QNone_Bool_bufchan_d;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_QTree_Bool) : (lizzieLet45_4QVal_Bool_4,QTree_Bool) (lizzieLet45_5QVal_Bool,Pointer_QTree_Bool) > [(lizzieLet45_4QVal_Bool_4QNone_Bool,Pointer_QTree_Bool),
                                                                                                                     (_15,Pointer_QTree_Bool),
                                                                                                                     (_14,Pointer_QTree_Bool),
                                                                                                                     (_13,Pointer_QTree_Bool)] */
  logic [3:0] lizzieLet45_5QVal_Bool_onehotd;
  always_comb
    if ((lizzieLet45_4QVal_Bool_4_d[0] && lizzieLet45_5QVal_Bool_d[0]))
      unique case (lizzieLet45_4QVal_Bool_4_d[2:1])
        2'd0: lizzieLet45_5QVal_Bool_onehotd = 4'd1;
        2'd1: lizzieLet45_5QVal_Bool_onehotd = 4'd2;
        2'd2: lizzieLet45_5QVal_Bool_onehotd = 4'd4;
        2'd3: lizzieLet45_5QVal_Bool_onehotd = 4'd8;
        default: lizzieLet45_5QVal_Bool_onehotd = 4'd0;
      endcase
    else lizzieLet45_5QVal_Bool_onehotd = 4'd0;
  assign lizzieLet45_4QVal_Bool_4QNone_Bool_d = {lizzieLet45_5QVal_Bool_d[16:1],
                                                 lizzieLet45_5QVal_Bool_onehotd[0]};
  assign _15_d = {lizzieLet45_5QVal_Bool_d[16:1],
                  lizzieLet45_5QVal_Bool_onehotd[1]};
  assign _14_d = {lizzieLet45_5QVal_Bool_d[16:1],
                  lizzieLet45_5QVal_Bool_onehotd[2]};
  assign _13_d = {lizzieLet45_5QVal_Bool_d[16:1],
                  lizzieLet45_5QVal_Bool_onehotd[3]};
  assign lizzieLet45_5QVal_Bool_r = (| (lizzieLet45_5QVal_Bool_onehotd & {_13_r,
                                                                          _14_r,
                                                                          _15_r,
                                                                          lizzieLet45_4QVal_Bool_4QNone_Bool_r}));
  assign lizzieLet45_4QVal_Bool_4_r = lizzieLet45_5QVal_Bool_r;
  
  /* buf (Ty Pointer_QTree_Bool) : (lizzieLet45_4QVal_Bool_4QNone_Bool,Pointer_QTree_Bool) > (lizzieLet45_4QVal_Bool_4QNone_Bool_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t lizzieLet45_4QVal_Bool_4QNone_Bool_bufchan_d;
  logic lizzieLet45_4QVal_Bool_4QNone_Bool_bufchan_r;
  assign lizzieLet45_4QVal_Bool_4QNone_Bool_r = ((! lizzieLet45_4QVal_Bool_4QNone_Bool_bufchan_d[0]) || lizzieLet45_4QVal_Bool_4QNone_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet45_4QVal_Bool_4QNone_Bool_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet45_4QVal_Bool_4QNone_Bool_r)
        lizzieLet45_4QVal_Bool_4QNone_Bool_bufchan_d <= lizzieLet45_4QVal_Bool_4QNone_Bool_d;
  Pointer_QTree_Bool_t lizzieLet45_4QVal_Bool_4QNone_Bool_bufchan_buf;
  assign lizzieLet45_4QVal_Bool_4QNone_Bool_bufchan_r = (! lizzieLet45_4QVal_Bool_4QNone_Bool_bufchan_buf[0]);
  assign lizzieLet45_4QVal_Bool_4QNone_Bool_1_argbuf_d = (lizzieLet45_4QVal_Bool_4QNone_Bool_bufchan_buf[0] ? lizzieLet45_4QVal_Bool_4QNone_Bool_bufchan_buf :
                                                          lizzieLet45_4QVal_Bool_4QNone_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet45_4QVal_Bool_4QNone_Bool_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet45_4QVal_Bool_4QNone_Bool_1_argbuf_r && lizzieLet45_4QVal_Bool_4QNone_Bool_bufchan_buf[0]))
        lizzieLet45_4QVal_Bool_4QNone_Bool_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet45_4QVal_Bool_4QNone_Bool_1_argbuf_r) && (! lizzieLet45_4QVal_Bool_4QNone_Bool_bufchan_buf[0])))
        lizzieLet45_4QVal_Bool_4QNone_Bool_bufchan_buf <= lizzieLet45_4QVal_Bool_4QNone_Bool_bufchan_d;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_CTf'''''''''''') : (lizzieLet45_4QVal_Bool_5,QTree_Bool) (lizzieLet45_6QVal_Bool,Pointer_CTf'''''''''''') > [(lizzieLet45_4QVal_Bool_5QNone_Bool,Pointer_CTf''''''''''''),
                                                                                                                               (lizzieLet45_4QVal_Bool_5QVal_Bool,Pointer_CTf''''''''''''),
                                                                                                                               (lizzieLet45_4QVal_Bool_5QNode_Bool,Pointer_CTf''''''''''''),
                                                                                                                               (lizzieLet45_4QVal_Bool_5QError_Bool,Pointer_CTf'''''''''''')] */
  logic [3:0] lizzieLet45_6QVal_Bool_onehotd;
  always_comb
    if ((lizzieLet45_4QVal_Bool_5_d[0] && lizzieLet45_6QVal_Bool_d[0]))
      unique case (lizzieLet45_4QVal_Bool_5_d[2:1])
        2'd0: lizzieLet45_6QVal_Bool_onehotd = 4'd1;
        2'd1: lizzieLet45_6QVal_Bool_onehotd = 4'd2;
        2'd2: lizzieLet45_6QVal_Bool_onehotd = 4'd4;
        2'd3: lizzieLet45_6QVal_Bool_onehotd = 4'd8;
        default: lizzieLet45_6QVal_Bool_onehotd = 4'd0;
      endcase
    else lizzieLet45_6QVal_Bool_onehotd = 4'd0;
  assign lizzieLet45_4QVal_Bool_5QNone_Bool_d = {lizzieLet45_6QVal_Bool_d[16:1],
                                                 lizzieLet45_6QVal_Bool_onehotd[0]};
  assign lizzieLet45_4QVal_Bool_5QVal_Bool_d = {lizzieLet45_6QVal_Bool_d[16:1],
                                                lizzieLet45_6QVal_Bool_onehotd[1]};
  assign lizzieLet45_4QVal_Bool_5QNode_Bool_d = {lizzieLet45_6QVal_Bool_d[16:1],
                                                 lizzieLet45_6QVal_Bool_onehotd[2]};
  assign lizzieLet45_4QVal_Bool_5QError_Bool_d = {lizzieLet45_6QVal_Bool_d[16:1],
                                                  lizzieLet45_6QVal_Bool_onehotd[3]};
  assign lizzieLet45_6QVal_Bool_r = (| (lizzieLet45_6QVal_Bool_onehotd & {lizzieLet45_4QVal_Bool_5QError_Bool_r,
                                                                          lizzieLet45_4QVal_Bool_5QNode_Bool_r,
                                                                          lizzieLet45_4QVal_Bool_5QVal_Bool_r,
                                                                          lizzieLet45_4QVal_Bool_5QNone_Bool_r}));
  assign lizzieLet45_4QVal_Bool_5_r = lizzieLet45_6QVal_Bool_r;
  
  /* buf (Ty Pointer_CTf'''''''''''') : (lizzieLet45_4QVal_Bool_5QError_Bool,Pointer_CTf'''''''''''') > (lizzieLet45_4QVal_Bool_5QError_Bool_1_argbuf,Pointer_CTf'''''''''''') */
  \Pointer_CTf''''''''''''_t  lizzieLet45_4QVal_Bool_5QError_Bool_bufchan_d;
  logic lizzieLet45_4QVal_Bool_5QError_Bool_bufchan_r;
  assign lizzieLet45_4QVal_Bool_5QError_Bool_r = ((! lizzieLet45_4QVal_Bool_5QError_Bool_bufchan_d[0]) || lizzieLet45_4QVal_Bool_5QError_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet45_4QVal_Bool_5QError_Bool_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet45_4QVal_Bool_5QError_Bool_r)
        lizzieLet45_4QVal_Bool_5QError_Bool_bufchan_d <= lizzieLet45_4QVal_Bool_5QError_Bool_d;
  \Pointer_CTf''''''''''''_t  lizzieLet45_4QVal_Bool_5QError_Bool_bufchan_buf;
  assign lizzieLet45_4QVal_Bool_5QError_Bool_bufchan_r = (! lizzieLet45_4QVal_Bool_5QError_Bool_bufchan_buf[0]);
  assign lizzieLet45_4QVal_Bool_5QError_Bool_1_argbuf_d = (lizzieLet45_4QVal_Bool_5QError_Bool_bufchan_buf[0] ? lizzieLet45_4QVal_Bool_5QError_Bool_bufchan_buf :
                                                           lizzieLet45_4QVal_Bool_5QError_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet45_4QVal_Bool_5QError_Bool_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet45_4QVal_Bool_5QError_Bool_1_argbuf_r && lizzieLet45_4QVal_Bool_5QError_Bool_bufchan_buf[0]))
        lizzieLet45_4QVal_Bool_5QError_Bool_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet45_4QVal_Bool_5QError_Bool_1_argbuf_r) && (! lizzieLet45_4QVal_Bool_5QError_Bool_bufchan_buf[0])))
        lizzieLet45_4QVal_Bool_5QError_Bool_bufchan_buf <= lizzieLet45_4QVal_Bool_5QError_Bool_bufchan_d;
  
  /* buf (Ty Pointer_CTf'''''''''''') : (lizzieLet45_4QVal_Bool_5QNode_Bool,Pointer_CTf'''''''''''') > (lizzieLet45_4QVal_Bool_5QNode_Bool_1_argbuf,Pointer_CTf'''''''''''') */
  \Pointer_CTf''''''''''''_t  lizzieLet45_4QVal_Bool_5QNode_Bool_bufchan_d;
  logic lizzieLet45_4QVal_Bool_5QNode_Bool_bufchan_r;
  assign lizzieLet45_4QVal_Bool_5QNode_Bool_r = ((! lizzieLet45_4QVal_Bool_5QNode_Bool_bufchan_d[0]) || lizzieLet45_4QVal_Bool_5QNode_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet45_4QVal_Bool_5QNode_Bool_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet45_4QVal_Bool_5QNode_Bool_r)
        lizzieLet45_4QVal_Bool_5QNode_Bool_bufchan_d <= lizzieLet45_4QVal_Bool_5QNode_Bool_d;
  \Pointer_CTf''''''''''''_t  lizzieLet45_4QVal_Bool_5QNode_Bool_bufchan_buf;
  assign lizzieLet45_4QVal_Bool_5QNode_Bool_bufchan_r = (! lizzieLet45_4QVal_Bool_5QNode_Bool_bufchan_buf[0]);
  assign lizzieLet45_4QVal_Bool_5QNode_Bool_1_argbuf_d = (lizzieLet45_4QVal_Bool_5QNode_Bool_bufchan_buf[0] ? lizzieLet45_4QVal_Bool_5QNode_Bool_bufchan_buf :
                                                          lizzieLet45_4QVal_Bool_5QNode_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet45_4QVal_Bool_5QNode_Bool_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet45_4QVal_Bool_5QNode_Bool_1_argbuf_r && lizzieLet45_4QVal_Bool_5QNode_Bool_bufchan_buf[0]))
        lizzieLet45_4QVal_Bool_5QNode_Bool_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet45_4QVal_Bool_5QNode_Bool_1_argbuf_r) && (! lizzieLet45_4QVal_Bool_5QNode_Bool_bufchan_buf[0])))
        lizzieLet45_4QVal_Bool_5QNode_Bool_bufchan_buf <= lizzieLet45_4QVal_Bool_5QNode_Bool_bufchan_d;
  
  /* buf (Ty Pointer_CTf'''''''''''') : (lizzieLet45_4QVal_Bool_5QNone_Bool,Pointer_CTf'''''''''''') > (lizzieLet45_4QVal_Bool_5QNone_Bool_1_argbuf,Pointer_CTf'''''''''''') */
  \Pointer_CTf''''''''''''_t  lizzieLet45_4QVal_Bool_5QNone_Bool_bufchan_d;
  logic lizzieLet45_4QVal_Bool_5QNone_Bool_bufchan_r;
  assign lizzieLet45_4QVal_Bool_5QNone_Bool_r = ((! lizzieLet45_4QVal_Bool_5QNone_Bool_bufchan_d[0]) || lizzieLet45_4QVal_Bool_5QNone_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet45_4QVal_Bool_5QNone_Bool_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet45_4QVal_Bool_5QNone_Bool_r)
        lizzieLet45_4QVal_Bool_5QNone_Bool_bufchan_d <= lizzieLet45_4QVal_Bool_5QNone_Bool_d;
  \Pointer_CTf''''''''''''_t  lizzieLet45_4QVal_Bool_5QNone_Bool_bufchan_buf;
  assign lizzieLet45_4QVal_Bool_5QNone_Bool_bufchan_r = (! lizzieLet45_4QVal_Bool_5QNone_Bool_bufchan_buf[0]);
  assign lizzieLet45_4QVal_Bool_5QNone_Bool_1_argbuf_d = (lizzieLet45_4QVal_Bool_5QNone_Bool_bufchan_buf[0] ? lizzieLet45_4QVal_Bool_5QNone_Bool_bufchan_buf :
                                                          lizzieLet45_4QVal_Bool_5QNone_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet45_4QVal_Bool_5QNone_Bool_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet45_4QVal_Bool_5QNone_Bool_1_argbuf_r && lizzieLet45_4QVal_Bool_5QNone_Bool_bufchan_buf[0]))
        lizzieLet45_4QVal_Bool_5QNone_Bool_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet45_4QVal_Bool_5QNone_Bool_1_argbuf_r) && (! lizzieLet45_4QVal_Bool_5QNone_Bool_bufchan_buf[0])))
        lizzieLet45_4QVal_Bool_5QNone_Bool_bufchan_buf <= lizzieLet45_4QVal_Bool_5QNone_Bool_bufchan_d;
  
  /* demux (Ty QTree_Bool,
       Ty MyBool) : (lizzieLet45_4QVal_Bool_6,QTree_Bool) (v1a92_destruct,MyBool) > [(_12,MyBool),
                                                                                     (lizzieLet45_4QVal_Bool_6QVal_Bool,MyBool),
                                                                                     (_11,MyBool),
                                                                                     (_10,MyBool)] */
  logic [3:0] v1a92_destruct_onehotd;
  always_comb
    if ((lizzieLet45_4QVal_Bool_6_d[0] && v1a92_destruct_d[0]))
      unique case (lizzieLet45_4QVal_Bool_6_d[2:1])
        2'd0: v1a92_destruct_onehotd = 4'd1;
        2'd1: v1a92_destruct_onehotd = 4'd2;
        2'd2: v1a92_destruct_onehotd = 4'd4;
        2'd3: v1a92_destruct_onehotd = 4'd8;
        default: v1a92_destruct_onehotd = 4'd0;
      endcase
    else v1a92_destruct_onehotd = 4'd0;
  assign _12_d = {v1a92_destruct_d[1:1], v1a92_destruct_onehotd[0]};
  assign lizzieLet45_4QVal_Bool_6QVal_Bool_d = {v1a92_destruct_d[1:1],
                                                v1a92_destruct_onehotd[1]};
  assign _11_d = {v1a92_destruct_d[1:1], v1a92_destruct_onehotd[2]};
  assign _10_d = {v1a92_destruct_d[1:1], v1a92_destruct_onehotd[3]};
  assign v1a92_destruct_r = (| (v1a92_destruct_onehotd & {_10_r,
                                                          _11_r,
                                                          lizzieLet45_4QVal_Bool_6QVal_Bool_r,
                                                          _12_r}));
  assign lizzieLet45_4QVal_Bool_6_r = v1a92_destruct_r;
  
  /* fork (Ty MyBool) : (lizzieLet45_4QVal_Bool_6QVal_Bool,MyBool) > [(lizzieLet45_4QVal_Bool_6QVal_Bool_1,MyBool),
                                                                 (lizzieLet45_4QVal_Bool_6QVal_Bool_2,MyBool),
                                                                 (lizzieLet45_4QVal_Bool_6QVal_Bool_3,MyBool)] */
  logic [2:0] lizzieLet45_4QVal_Bool_6QVal_Bool_emitted;
  logic [2:0] lizzieLet45_4QVal_Bool_6QVal_Bool_done;
  assign lizzieLet45_4QVal_Bool_6QVal_Bool_1_d = {lizzieLet45_4QVal_Bool_6QVal_Bool_d[1:1],
                                                  (lizzieLet45_4QVal_Bool_6QVal_Bool_d[0] && (! lizzieLet45_4QVal_Bool_6QVal_Bool_emitted[0]))};
  assign lizzieLet45_4QVal_Bool_6QVal_Bool_2_d = {lizzieLet45_4QVal_Bool_6QVal_Bool_d[1:1],
                                                  (lizzieLet45_4QVal_Bool_6QVal_Bool_d[0] && (! lizzieLet45_4QVal_Bool_6QVal_Bool_emitted[1]))};
  assign lizzieLet45_4QVal_Bool_6QVal_Bool_3_d = {lizzieLet45_4QVal_Bool_6QVal_Bool_d[1:1],
                                                  (lizzieLet45_4QVal_Bool_6QVal_Bool_d[0] && (! lizzieLet45_4QVal_Bool_6QVal_Bool_emitted[2]))};
  assign lizzieLet45_4QVal_Bool_6QVal_Bool_done = (lizzieLet45_4QVal_Bool_6QVal_Bool_emitted | ({lizzieLet45_4QVal_Bool_6QVal_Bool_3_d[0],
                                                                                                 lizzieLet45_4QVal_Bool_6QVal_Bool_2_d[0],
                                                                                                 lizzieLet45_4QVal_Bool_6QVal_Bool_1_d[0]} & {lizzieLet45_4QVal_Bool_6QVal_Bool_3_r,
                                                                                                                                              lizzieLet45_4QVal_Bool_6QVal_Bool_2_r,
                                                                                                                                              lizzieLet45_4QVal_Bool_6QVal_Bool_1_r}));
  assign lizzieLet45_4QVal_Bool_6QVal_Bool_r = (& lizzieLet45_4QVal_Bool_6QVal_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet45_4QVal_Bool_6QVal_Bool_emitted <= 3'd0;
    else
      lizzieLet45_4QVal_Bool_6QVal_Bool_emitted <= (lizzieLet45_4QVal_Bool_6QVal_Bool_r ? 3'd0 :
                                                    lizzieLet45_4QVal_Bool_6QVal_Bool_done);
  
  /* demux (Ty MyBool,
       Ty Go) : (lizzieLet45_4QVal_Bool_6QVal_Bool_1,MyBool) (lizzieLet45_4QVal_Bool_3QVal_Bool,Go) > [(lizzieLet45_4QVal_Bool_6QVal_Bool_1MyFalse,Go),
                                                                                                       (lizzieLet45_4QVal_Bool_6QVal_Bool_1MyTrue,Go)] */
  logic [1:0] lizzieLet45_4QVal_Bool_3QVal_Bool_onehotd;
  always_comb
    if ((lizzieLet45_4QVal_Bool_6QVal_Bool_1_d[0] && lizzieLet45_4QVal_Bool_3QVal_Bool_d[0]))
      unique case (lizzieLet45_4QVal_Bool_6QVal_Bool_1_d[1:1])
        1'd0: lizzieLet45_4QVal_Bool_3QVal_Bool_onehotd = 2'd1;
        1'd1: lizzieLet45_4QVal_Bool_3QVal_Bool_onehotd = 2'd2;
        default: lizzieLet45_4QVal_Bool_3QVal_Bool_onehotd = 2'd0;
      endcase
    else lizzieLet45_4QVal_Bool_3QVal_Bool_onehotd = 2'd0;
  assign lizzieLet45_4QVal_Bool_6QVal_Bool_1MyFalse_d = lizzieLet45_4QVal_Bool_3QVal_Bool_onehotd[0];
  assign lizzieLet45_4QVal_Bool_6QVal_Bool_1MyTrue_d = lizzieLet45_4QVal_Bool_3QVal_Bool_onehotd[1];
  assign lizzieLet45_4QVal_Bool_3QVal_Bool_r = (| (lizzieLet45_4QVal_Bool_3QVal_Bool_onehotd & {lizzieLet45_4QVal_Bool_6QVal_Bool_1MyTrue_r,
                                                                                                lizzieLet45_4QVal_Bool_6QVal_Bool_1MyFalse_r}));
  assign lizzieLet45_4QVal_Bool_6QVal_Bool_1_r = lizzieLet45_4QVal_Bool_3QVal_Bool_r;
  
  /* fork (Ty Go) : (lizzieLet45_4QVal_Bool_6QVal_Bool_1MyTrue,Go) > [(lizzieLet45_4QVal_Bool_6QVal_Bool_1MyTrue_1,Go),
                                                                 (lizzieLet45_4QVal_Bool_6QVal_Bool_1MyTrue_2,Go)] */
  logic [1:0] lizzieLet45_4QVal_Bool_6QVal_Bool_1MyTrue_emitted;
  logic [1:0] lizzieLet45_4QVal_Bool_6QVal_Bool_1MyTrue_done;
  assign lizzieLet45_4QVal_Bool_6QVal_Bool_1MyTrue_1_d = (lizzieLet45_4QVal_Bool_6QVal_Bool_1MyTrue_d[0] && (! lizzieLet45_4QVal_Bool_6QVal_Bool_1MyTrue_emitted[0]));
  assign lizzieLet45_4QVal_Bool_6QVal_Bool_1MyTrue_2_d = (lizzieLet45_4QVal_Bool_6QVal_Bool_1MyTrue_d[0] && (! lizzieLet45_4QVal_Bool_6QVal_Bool_1MyTrue_emitted[1]));
  assign lizzieLet45_4QVal_Bool_6QVal_Bool_1MyTrue_done = (lizzieLet45_4QVal_Bool_6QVal_Bool_1MyTrue_emitted | ({lizzieLet45_4QVal_Bool_6QVal_Bool_1MyTrue_2_d[0],
                                                                                                                 lizzieLet45_4QVal_Bool_6QVal_Bool_1MyTrue_1_d[0]} & {lizzieLet45_4QVal_Bool_6QVal_Bool_1MyTrue_2_r,
                                                                                                                                                                      lizzieLet45_4QVal_Bool_6QVal_Bool_1MyTrue_1_r}));
  assign lizzieLet45_4QVal_Bool_6QVal_Bool_1MyTrue_r = (& lizzieLet45_4QVal_Bool_6QVal_Bool_1MyTrue_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet45_4QVal_Bool_6QVal_Bool_1MyTrue_emitted <= 2'd0;
    else
      lizzieLet45_4QVal_Bool_6QVal_Bool_1MyTrue_emitted <= (lizzieLet45_4QVal_Bool_6QVal_Bool_1MyTrue_r ? 2'd0 :
                                                            lizzieLet45_4QVal_Bool_6QVal_Bool_1MyTrue_done);
  
  /* buf (Ty Go) : (lizzieLet45_4QVal_Bool_6QVal_Bool_1MyTrue_1,Go) > (lizzieLet45_4QVal_Bool_6QVal_Bool_1MyTrue_1_argbuf,Go) */
  Go_t lizzieLet45_4QVal_Bool_6QVal_Bool_1MyTrue_1_bufchan_d;
  logic lizzieLet45_4QVal_Bool_6QVal_Bool_1MyTrue_1_bufchan_r;
  assign lizzieLet45_4QVal_Bool_6QVal_Bool_1MyTrue_1_r = ((! lizzieLet45_4QVal_Bool_6QVal_Bool_1MyTrue_1_bufchan_d[0]) || lizzieLet45_4QVal_Bool_6QVal_Bool_1MyTrue_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet45_4QVal_Bool_6QVal_Bool_1MyTrue_1_bufchan_d <= 1'd0;
    else
      if (lizzieLet45_4QVal_Bool_6QVal_Bool_1MyTrue_1_r)
        lizzieLet45_4QVal_Bool_6QVal_Bool_1MyTrue_1_bufchan_d <= lizzieLet45_4QVal_Bool_6QVal_Bool_1MyTrue_1_d;
  Go_t lizzieLet45_4QVal_Bool_6QVal_Bool_1MyTrue_1_bufchan_buf;
  assign lizzieLet45_4QVal_Bool_6QVal_Bool_1MyTrue_1_bufchan_r = (! lizzieLet45_4QVal_Bool_6QVal_Bool_1MyTrue_1_bufchan_buf[0]);
  assign lizzieLet45_4QVal_Bool_6QVal_Bool_1MyTrue_1_argbuf_d = (lizzieLet45_4QVal_Bool_6QVal_Bool_1MyTrue_1_bufchan_buf[0] ? lizzieLet45_4QVal_Bool_6QVal_Bool_1MyTrue_1_bufchan_buf :
                                                                 lizzieLet45_4QVal_Bool_6QVal_Bool_1MyTrue_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet45_4QVal_Bool_6QVal_Bool_1MyTrue_1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet45_4QVal_Bool_6QVal_Bool_1MyTrue_1_argbuf_r && lizzieLet45_4QVal_Bool_6QVal_Bool_1MyTrue_1_bufchan_buf[0]))
        lizzieLet45_4QVal_Bool_6QVal_Bool_1MyTrue_1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet45_4QVal_Bool_6QVal_Bool_1MyTrue_1_argbuf_r) && (! lizzieLet45_4QVal_Bool_6QVal_Bool_1MyTrue_1_bufchan_buf[0])))
        lizzieLet45_4QVal_Bool_6QVal_Bool_1MyTrue_1_bufchan_buf <= lizzieLet45_4QVal_Bool_6QVal_Bool_1MyTrue_1_bufchan_d;
  
  /* dcon (Ty TupGo,
      Dcon TupGo) : [(lizzieLet45_4QVal_Bool_6QVal_Bool_1MyTrue_1_argbuf,Go)] > (lvlrf2-0TupGo4,TupGo) */
  assign \lvlrf2-0TupGo4_d  = TupGo_dc((& {lizzieLet45_4QVal_Bool_6QVal_Bool_1MyTrue_1_argbuf_d[0]}), lizzieLet45_4QVal_Bool_6QVal_Bool_1MyTrue_1_argbuf_d);
  assign {lizzieLet45_4QVal_Bool_6QVal_Bool_1MyTrue_1_argbuf_r} = {1 {(\lvlrf2-0TupGo4_r  && \lvlrf2-0TupGo4_d [0])}};
  
  /* buf (Ty Go) : (lizzieLet45_4QVal_Bool_6QVal_Bool_1MyTrue_2,Go) > (lizzieLet45_4QVal_Bool_6QVal_Bool_1MyTrue_2_argbuf,Go) */
  Go_t lizzieLet45_4QVal_Bool_6QVal_Bool_1MyTrue_2_bufchan_d;
  logic lizzieLet45_4QVal_Bool_6QVal_Bool_1MyTrue_2_bufchan_r;
  assign lizzieLet45_4QVal_Bool_6QVal_Bool_1MyTrue_2_r = ((! lizzieLet45_4QVal_Bool_6QVal_Bool_1MyTrue_2_bufchan_d[0]) || lizzieLet45_4QVal_Bool_6QVal_Bool_1MyTrue_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet45_4QVal_Bool_6QVal_Bool_1MyTrue_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet45_4QVal_Bool_6QVal_Bool_1MyTrue_2_r)
        lizzieLet45_4QVal_Bool_6QVal_Bool_1MyTrue_2_bufchan_d <= lizzieLet45_4QVal_Bool_6QVal_Bool_1MyTrue_2_d;
  Go_t lizzieLet45_4QVal_Bool_6QVal_Bool_1MyTrue_2_bufchan_buf;
  assign lizzieLet45_4QVal_Bool_6QVal_Bool_1MyTrue_2_bufchan_r = (! lizzieLet45_4QVal_Bool_6QVal_Bool_1MyTrue_2_bufchan_buf[0]);
  assign lizzieLet45_4QVal_Bool_6QVal_Bool_1MyTrue_2_argbuf_d = (lizzieLet45_4QVal_Bool_6QVal_Bool_1MyTrue_2_bufchan_buf[0] ? lizzieLet45_4QVal_Bool_6QVal_Bool_1MyTrue_2_bufchan_buf :
                                                                 lizzieLet45_4QVal_Bool_6QVal_Bool_1MyTrue_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet45_4QVal_Bool_6QVal_Bool_1MyTrue_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet45_4QVal_Bool_6QVal_Bool_1MyTrue_2_argbuf_r && lizzieLet45_4QVal_Bool_6QVal_Bool_1MyTrue_2_bufchan_buf[0]))
        lizzieLet45_4QVal_Bool_6QVal_Bool_1MyTrue_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet45_4QVal_Bool_6QVal_Bool_1MyTrue_2_argbuf_r) && (! lizzieLet45_4QVal_Bool_6QVal_Bool_1MyTrue_2_bufchan_buf[0])))
        lizzieLet45_4QVal_Bool_6QVal_Bool_1MyTrue_2_bufchan_buf <= lizzieLet45_4QVal_Bool_6QVal_Bool_1MyTrue_2_bufchan_d;
  
  /* demux (Ty MyBool,
       Ty Pointer_CTf'''''''''''') : (lizzieLet45_4QVal_Bool_6QVal_Bool_2,MyBool) (lizzieLet45_4QVal_Bool_5QVal_Bool,Pointer_CTf'''''''''''') > [(lizzieLet45_4QVal_Bool_6QVal_Bool_2MyFalse,Pointer_CTf''''''''''''),
                                                                                                                                                 (lizzieLet45_4QVal_Bool_6QVal_Bool_2MyTrue,Pointer_CTf'''''''''''')] */
  logic [1:0] lizzieLet45_4QVal_Bool_5QVal_Bool_onehotd;
  always_comb
    if ((lizzieLet45_4QVal_Bool_6QVal_Bool_2_d[0] && lizzieLet45_4QVal_Bool_5QVal_Bool_d[0]))
      unique case (lizzieLet45_4QVal_Bool_6QVal_Bool_2_d[1:1])
        1'd0: lizzieLet45_4QVal_Bool_5QVal_Bool_onehotd = 2'd1;
        1'd1: lizzieLet45_4QVal_Bool_5QVal_Bool_onehotd = 2'd2;
        default: lizzieLet45_4QVal_Bool_5QVal_Bool_onehotd = 2'd0;
      endcase
    else lizzieLet45_4QVal_Bool_5QVal_Bool_onehotd = 2'd0;
  assign lizzieLet45_4QVal_Bool_6QVal_Bool_2MyFalse_d = {lizzieLet45_4QVal_Bool_5QVal_Bool_d[16:1],
                                                         lizzieLet45_4QVal_Bool_5QVal_Bool_onehotd[0]};
  assign lizzieLet45_4QVal_Bool_6QVal_Bool_2MyTrue_d = {lizzieLet45_4QVal_Bool_5QVal_Bool_d[16:1],
                                                        lizzieLet45_4QVal_Bool_5QVal_Bool_onehotd[1]};
  assign lizzieLet45_4QVal_Bool_5QVal_Bool_r = (| (lizzieLet45_4QVal_Bool_5QVal_Bool_onehotd & {lizzieLet45_4QVal_Bool_6QVal_Bool_2MyTrue_r,
                                                                                                lizzieLet45_4QVal_Bool_6QVal_Bool_2MyFalse_r}));
  assign lizzieLet45_4QVal_Bool_6QVal_Bool_2_r = lizzieLet45_4QVal_Bool_5QVal_Bool_r;
  
  /* buf (Ty Pointer_CTf'''''''''''') : (lizzieLet45_4QVal_Bool_6QVal_Bool_2MyTrue,Pointer_CTf'''''''''''') > (lizzieLet45_4QVal_Bool_6QVal_Bool_2MyTrue_1_argbuf,Pointer_CTf'''''''''''') */
  \Pointer_CTf''''''''''''_t  lizzieLet45_4QVal_Bool_6QVal_Bool_2MyTrue_bufchan_d;
  logic lizzieLet45_4QVal_Bool_6QVal_Bool_2MyTrue_bufchan_r;
  assign lizzieLet45_4QVal_Bool_6QVal_Bool_2MyTrue_r = ((! lizzieLet45_4QVal_Bool_6QVal_Bool_2MyTrue_bufchan_d[0]) || lizzieLet45_4QVal_Bool_6QVal_Bool_2MyTrue_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet45_4QVal_Bool_6QVal_Bool_2MyTrue_bufchan_d <= {16'd0,
                                                              1'd0};
    else
      if (lizzieLet45_4QVal_Bool_6QVal_Bool_2MyTrue_r)
        lizzieLet45_4QVal_Bool_6QVal_Bool_2MyTrue_bufchan_d <= lizzieLet45_4QVal_Bool_6QVal_Bool_2MyTrue_d;
  \Pointer_CTf''''''''''''_t  lizzieLet45_4QVal_Bool_6QVal_Bool_2MyTrue_bufchan_buf;
  assign lizzieLet45_4QVal_Bool_6QVal_Bool_2MyTrue_bufchan_r = (! lizzieLet45_4QVal_Bool_6QVal_Bool_2MyTrue_bufchan_buf[0]);
  assign lizzieLet45_4QVal_Bool_6QVal_Bool_2MyTrue_1_argbuf_d = (lizzieLet45_4QVal_Bool_6QVal_Bool_2MyTrue_bufchan_buf[0] ? lizzieLet45_4QVal_Bool_6QVal_Bool_2MyTrue_bufchan_buf :
                                                                 lizzieLet45_4QVal_Bool_6QVal_Bool_2MyTrue_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet45_4QVal_Bool_6QVal_Bool_2MyTrue_bufchan_buf <= {16'd0,
                                                                1'd0};
    else
      if ((lizzieLet45_4QVal_Bool_6QVal_Bool_2MyTrue_1_argbuf_r && lizzieLet45_4QVal_Bool_6QVal_Bool_2MyTrue_bufchan_buf[0]))
        lizzieLet45_4QVal_Bool_6QVal_Bool_2MyTrue_bufchan_buf <= {16'd0,
                                                                  1'd0};
      else if (((! lizzieLet45_4QVal_Bool_6QVal_Bool_2MyTrue_1_argbuf_r) && (! lizzieLet45_4QVal_Bool_6QVal_Bool_2MyTrue_bufchan_buf[0])))
        lizzieLet45_4QVal_Bool_6QVal_Bool_2MyTrue_bufchan_buf <= lizzieLet45_4QVal_Bool_6QVal_Bool_2MyTrue_bufchan_d;
  
  /* demux (Ty MyBool,
       Ty MyBool) : (lizzieLet45_4QVal_Bool_6QVal_Bool_3,MyBool) (va93_destruct,MyBool) > [(lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse,MyBool),
                                                                                           (_9,MyBool)] */
  logic [1:0] va93_destruct_onehotd;
  always_comb
    if ((lizzieLet45_4QVal_Bool_6QVal_Bool_3_d[0] && va93_destruct_d[0]))
      unique case (lizzieLet45_4QVal_Bool_6QVal_Bool_3_d[1:1])
        1'd0: va93_destruct_onehotd = 2'd1;
        1'd1: va93_destruct_onehotd = 2'd2;
        default: va93_destruct_onehotd = 2'd0;
      endcase
    else va93_destruct_onehotd = 2'd0;
  assign lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_d = {va93_destruct_d[1:1],
                                                         va93_destruct_onehotd[0]};
  assign _9_d = {va93_destruct_d[1:1], va93_destruct_onehotd[1]};
  assign va93_destruct_r = (| (va93_destruct_onehotd & {_9_r,
                                                        lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_r}));
  assign lizzieLet45_4QVal_Bool_6QVal_Bool_3_r = va93_destruct_r;
  
  /* fork (Ty MyBool) : (lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse,MyBool) > [(lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1,MyBool),
                                                                          (lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_2,MyBool)] */
  logic [1:0] lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_emitted;
  logic [1:0] lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_done;
  assign lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1_d = {lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_d[1:1],
                                                           (lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_d[0] && (! lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_emitted[0]))};
  assign lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_2_d = {lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_d[1:1],
                                                           (lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_d[0] && (! lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_emitted[1]))};
  assign lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_done = (lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_emitted | ({lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_2_d[0],
                                                                                                                   lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1_d[0]} & {lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_2_r,
                                                                                                                                                                         lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1_r}));
  assign lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_r = (& lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_emitted <= 2'd0;
    else
      lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_emitted <= (lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_r ? 2'd0 :
                                                             lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_done);
  
  /* demux (Ty MyBool,
       Ty Go) : (lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1,MyBool) (lizzieLet45_4QVal_Bool_6QVal_Bool_1MyFalse,Go) > [(lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse,Go),
                                                                                                                         (lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue,Go)] */
  logic [1:0] lizzieLet45_4QVal_Bool_6QVal_Bool_1MyFalse_onehotd;
  always_comb
    if ((lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1_d[0] && lizzieLet45_4QVal_Bool_6QVal_Bool_1MyFalse_d[0]))
      unique case (lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1_d[1:1])
        1'd0: lizzieLet45_4QVal_Bool_6QVal_Bool_1MyFalse_onehotd = 2'd1;
        1'd1: lizzieLet45_4QVal_Bool_6QVal_Bool_1MyFalse_onehotd = 2'd2;
        default: lizzieLet45_4QVal_Bool_6QVal_Bool_1MyFalse_onehotd = 2'd0;
      endcase
    else lizzieLet45_4QVal_Bool_6QVal_Bool_1MyFalse_onehotd = 2'd0;
  assign lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_d = lizzieLet45_4QVal_Bool_6QVal_Bool_1MyFalse_onehotd[0];
  assign lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_d = lizzieLet45_4QVal_Bool_6QVal_Bool_1MyFalse_onehotd[1];
  assign lizzieLet45_4QVal_Bool_6QVal_Bool_1MyFalse_r = (| (lizzieLet45_4QVal_Bool_6QVal_Bool_1MyFalse_onehotd & {lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_r,
                                                                                                                  lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_r}));
  assign lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1_r = lizzieLet45_4QVal_Bool_6QVal_Bool_1MyFalse_r;
  
  /* fork (Ty Go) : (lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse,Go) > [(lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1,Go),
                                                                           (lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2,Go)] */
  logic [1:0] lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_emitted;
  logic [1:0] lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_done;
  assign lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1_d = (lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_d[0] && (! lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_emitted[0]));
  assign lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_d = (lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_d[0] && (! lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_emitted[1]));
  assign lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_done = (lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_emitted | ({lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_d[0],
                                                                                                                                     lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1_d[0]} & {lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_r,
                                                                                                                                                                                                    lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1_r}));
  assign lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_r = (& lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_emitted <= 2'd0;
    else
      lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_emitted <= (lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_r ? 2'd0 :
                                                                      lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_done);
  
  /* dcon (Ty QTree_Bool,
      Dcon QNone_Bool) : [(lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1,Go)] > (lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool,QTree_Bool) */
  assign lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_d = QNone_Bool_dc((& {lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1_d[0]}), lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1_d);
  assign {lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1_r} = {1 {(lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_r && lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_d[0])}};
  
  /* buf (Ty QTree_Bool) : (lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool,QTree_Bool) > (lizzieLet47_1_argbuf,QTree_Bool) */
  QTree_Bool_t lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_bufchan_d;
  logic lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_bufchan_r;
  assign lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_r = ((! lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_bufchan_d[0]) || lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_bufchan_d <= {66'd0,
                                                                                    1'd0};
    else
      if (lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_r)
        lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_bufchan_d <= lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_d;
  QTree_Bool_t lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_bufchan_buf;
  assign lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_bufchan_r = (! lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_bufchan_buf[0]);
  assign lizzieLet47_1_argbuf_d = (lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_bufchan_buf[0] ? lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_bufchan_buf :
                                   lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_bufchan_buf <= {66'd0,
                                                                                      1'd0};
    else
      if ((lizzieLet47_1_argbuf_r && lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_bufchan_buf[0]))
        lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_bufchan_buf <= {66'd0,
                                                                                        1'd0};
      else if (((! lizzieLet47_1_argbuf_r) && (! lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_bufchan_buf[0])))
        lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_bufchan_buf <= lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2,Go) > (lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_argbuf,Go) */
  Go_t lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_bufchan_d;
  logic lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_bufchan_r;
  assign lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_r = ((! lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_bufchan_d[0]) || lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_r)
        lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_bufchan_d <= lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_d;
  Go_t lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_bufchan_buf;
  assign lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_bufchan_r = (! lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_bufchan_buf[0]);
  assign lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_argbuf_d = (lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_bufchan_buf[0] ? lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_bufchan_buf :
                                                                           lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_argbuf_r && lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_bufchan_buf[0]))
        lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_argbuf_r) && (! lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_bufchan_buf[0])))
        lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_bufchan_buf <= lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue,Go) > [(lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1,Go),
                                                                          (lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2,Go)] */
  logic [1:0] lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_emitted;
  logic [1:0] lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_done;
  assign lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_d = (lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_d[0] && (! lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_emitted[0]));
  assign lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_d = (lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_d[0] && (! lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_emitted[1]));
  assign lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_done = (lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_emitted | ({lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_d[0],
                                                                                                                                   lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_d[0]} & {lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_r,
                                                                                                                                                                                                 lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_r}));
  assign lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_r = (& lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_emitted <= 2'd0;
    else
      lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_emitted <= (lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_r ? 2'd0 :
                                                                     lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_done);
  
  /* buf (Ty Go) : (lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1,Go) > (lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_argbuf,Go) */
  Go_t lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_bufchan_d;
  logic lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_bufchan_r;
  assign lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_r = ((! lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_bufchan_d[0]) || lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_bufchan_d <= 1'd0;
    else
      if (lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_r)
        lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_bufchan_d <= lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_d;
  Go_t lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_bufchan_buf;
  assign lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_bufchan_r = (! lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_bufchan_buf[0]);
  assign lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_argbuf_d = (lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_bufchan_buf[0] ? lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_bufchan_buf :
                                                                          lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_argbuf_r && lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_bufchan_buf[0]))
        lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_argbuf_r) && (! lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_bufchan_buf[0])))
        lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_bufchan_buf <= lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_bufchan_d;
  
  /* dcon (Ty TupGo,
      Dcon TupGo) : [(lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_argbuf,Go)] > (lvlrf2-0TupGo3,TupGo) */
  assign \lvlrf2-0TupGo3_d  = TupGo_dc((& {lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_argbuf_d[0]}), lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_argbuf_d);
  assign {lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_argbuf_r} = {1 {(\lvlrf2-0TupGo3_r  && \lvlrf2-0TupGo3_d [0])}};
  
  /* buf (Ty Go) : (lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2,Go) > (lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_argbuf,Go) */
  Go_t lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_bufchan_d;
  logic lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_bufchan_r;
  assign lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_r = ((! lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_bufchan_d[0]) || lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_r)
        lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_bufchan_d <= lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_d;
  Go_t lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_bufchan_buf;
  assign lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_bufchan_r = (! lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_bufchan_buf[0]);
  assign lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_argbuf_d = (lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_bufchan_buf[0] ? lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_bufchan_buf :
                                                                          lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_argbuf_r && lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_bufchan_buf[0]))
        lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_argbuf_r) && (! lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_bufchan_buf[0])))
        lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_bufchan_buf <= lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_bufchan_d;
  
  /* demux (Ty MyBool,
       Ty Pointer_CTf'''''''''''') : (lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_2,MyBool) (lizzieLet45_4QVal_Bool_6QVal_Bool_2MyFalse,Pointer_CTf'''''''''''') > [(lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_2MyFalse,Pointer_CTf''''''''''''),
                                                                                                                                                                   (lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_2MyTrue,Pointer_CTf'''''''''''')] */
  logic [1:0] lizzieLet45_4QVal_Bool_6QVal_Bool_2MyFalse_onehotd;
  always_comb
    if ((lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_2_d[0] && lizzieLet45_4QVal_Bool_6QVal_Bool_2MyFalse_d[0]))
      unique case (lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_2_d[1:1])
        1'd0: lizzieLet45_4QVal_Bool_6QVal_Bool_2MyFalse_onehotd = 2'd1;
        1'd1: lizzieLet45_4QVal_Bool_6QVal_Bool_2MyFalse_onehotd = 2'd2;
        default: lizzieLet45_4QVal_Bool_6QVal_Bool_2MyFalse_onehotd = 2'd0;
      endcase
    else lizzieLet45_4QVal_Bool_6QVal_Bool_2MyFalse_onehotd = 2'd0;
  assign lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_2MyFalse_d = {lizzieLet45_4QVal_Bool_6QVal_Bool_2MyFalse_d[16:1],
                                                                  lizzieLet45_4QVal_Bool_6QVal_Bool_2MyFalse_onehotd[0]};
  assign lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_2MyTrue_d = {lizzieLet45_4QVal_Bool_6QVal_Bool_2MyFalse_d[16:1],
                                                                 lizzieLet45_4QVal_Bool_6QVal_Bool_2MyFalse_onehotd[1]};
  assign lizzieLet45_4QVal_Bool_6QVal_Bool_2MyFalse_r = (| (lizzieLet45_4QVal_Bool_6QVal_Bool_2MyFalse_onehotd & {lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_2MyTrue_r,
                                                                                                                  lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_2MyFalse_r}));
  assign lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_2_r = lizzieLet45_4QVal_Bool_6QVal_Bool_2MyFalse_r;
  
  /* buf (Ty Pointer_CTf'''''''''''') : (lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_2MyFalse,Pointer_CTf'''''''''''') > (lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_2MyFalse_1_argbuf,Pointer_CTf'''''''''''') */
  \Pointer_CTf''''''''''''_t  lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_2MyFalse_bufchan_d;
  logic lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_2MyFalse_bufchan_r;
  assign lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_2MyFalse_r = ((! lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_2MyFalse_bufchan_d[0]) || lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_2MyFalse_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_2MyFalse_bufchan_d <= {16'd0,
                                                                        1'd0};
    else
      if (lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_2MyFalse_r)
        lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_2MyFalse_bufchan_d <= lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_2MyFalse_d;
  \Pointer_CTf''''''''''''_t  lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_2MyFalse_bufchan_buf;
  assign lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_2MyFalse_bufchan_r = (! lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_2MyFalse_bufchan_buf[0]);
  assign lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_2MyFalse_1_argbuf_d = (lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_2MyFalse_bufchan_buf[0] ? lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_2MyFalse_bufchan_buf :
                                                                           lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_2MyFalse_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_2MyFalse_bufchan_buf <= {16'd0,
                                                                          1'd0};
    else
      if ((lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_2MyFalse_1_argbuf_r && lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_2MyFalse_bufchan_buf[0]))
        lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_2MyFalse_bufchan_buf <= {16'd0,
                                                                            1'd0};
      else if (((! lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_2MyFalse_1_argbuf_r) && (! lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_2MyFalse_bufchan_buf[0])))
        lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_2MyFalse_bufchan_buf <= lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_2MyFalse_bufchan_d;
  
  /* buf (Ty Pointer_CTf'''''''''''') : (lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_2MyTrue,Pointer_CTf'''''''''''') > (lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_2MyTrue_1_argbuf,Pointer_CTf'''''''''''') */
  \Pointer_CTf''''''''''''_t  lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_2MyTrue_bufchan_d;
  logic lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_2MyTrue_bufchan_r;
  assign lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_2MyTrue_r = ((! lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_2MyTrue_bufchan_d[0]) || lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_2MyTrue_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_2MyTrue_bufchan_d <= {16'd0,
                                                                       1'd0};
    else
      if (lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_2MyTrue_r)
        lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_2MyTrue_bufchan_d <= lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_2MyTrue_d;
  \Pointer_CTf''''''''''''_t  lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_2MyTrue_bufchan_buf;
  assign lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_2MyTrue_bufchan_r = (! lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_2MyTrue_bufchan_buf[0]);
  assign lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_2MyTrue_1_argbuf_d = (lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_2MyTrue_bufchan_buf[0] ? lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_2MyTrue_bufchan_buf :
                                                                          lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_2MyTrue_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_2MyTrue_bufchan_buf <= {16'd0,
                                                                         1'd0};
    else
      if ((lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_2MyTrue_1_argbuf_r && lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_2MyTrue_bufchan_buf[0]))
        lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_2MyTrue_bufchan_buf <= {16'd0,
                                                                           1'd0};
      else if (((! lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_2MyTrue_1_argbuf_r) && (! lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_2MyTrue_bufchan_buf[0])))
        lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_2MyTrue_bufchan_buf <= lizzieLet45_4QVal_Bool_6QVal_Bool_3MyFalse_2MyTrue_bufchan_d;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_QTree_Bool) : (lizzieLet45_5,QTree_Bool) (q4a90_2,Pointer_QTree_Bool) > [(_8,Pointer_QTree_Bool),
                                                                                           (lizzieLet45_5QVal_Bool,Pointer_QTree_Bool),
                                                                                           (lizzieLet45_5QNode_Bool,Pointer_QTree_Bool),
                                                                                           (_7,Pointer_QTree_Bool)] */
  logic [3:0] q4a90_2_onehotd;
  always_comb
    if ((lizzieLet45_5_d[0] && q4a90_2_d[0]))
      unique case (lizzieLet45_5_d[2:1])
        2'd0: q4a90_2_onehotd = 4'd1;
        2'd1: q4a90_2_onehotd = 4'd2;
        2'd2: q4a90_2_onehotd = 4'd4;
        2'd3: q4a90_2_onehotd = 4'd8;
        default: q4a90_2_onehotd = 4'd0;
      endcase
    else q4a90_2_onehotd = 4'd0;
  assign _8_d = {q4a90_2_d[16:1], q4a90_2_onehotd[0]};
  assign lizzieLet45_5QVal_Bool_d = {q4a90_2_d[16:1],
                                     q4a90_2_onehotd[1]};
  assign lizzieLet45_5QNode_Bool_d = {q4a90_2_d[16:1],
                                      q4a90_2_onehotd[2]};
  assign _7_d = {q4a90_2_d[16:1], q4a90_2_onehotd[3]};
  assign q4a90_2_r = (| (q4a90_2_onehotd & {_7_r,
                                            lizzieLet45_5QNode_Bool_r,
                                            lizzieLet45_5QVal_Bool_r,
                                            _8_r}));
  assign lizzieLet45_5_r = q4a90_2_r;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_CTf'''''''''''') : (lizzieLet45_6,QTree_Bool) (sc_0_1_goMux_mux,Pointer_CTf'''''''''''') > [(lizzieLet45_6QNone_Bool,Pointer_CTf''''''''''''),
                                                                                                              (lizzieLet45_6QVal_Bool,Pointer_CTf''''''''''''),
                                                                                                              (lizzieLet45_6QNode_Bool,Pointer_CTf''''''''''''),
                                                                                                              (lizzieLet45_6QError_Bool,Pointer_CTf'''''''''''')] */
  logic [3:0] sc_0_1_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet45_6_d[0] && sc_0_1_goMux_mux_d[0]))
      unique case (lizzieLet45_6_d[2:1])
        2'd0: sc_0_1_goMux_mux_onehotd = 4'd1;
        2'd1: sc_0_1_goMux_mux_onehotd = 4'd2;
        2'd2: sc_0_1_goMux_mux_onehotd = 4'd4;
        2'd3: sc_0_1_goMux_mux_onehotd = 4'd8;
        default: sc_0_1_goMux_mux_onehotd = 4'd0;
      endcase
    else sc_0_1_goMux_mux_onehotd = 4'd0;
  assign lizzieLet45_6QNone_Bool_d = {sc_0_1_goMux_mux_d[16:1],
                                      sc_0_1_goMux_mux_onehotd[0]};
  assign lizzieLet45_6QVal_Bool_d = {sc_0_1_goMux_mux_d[16:1],
                                     sc_0_1_goMux_mux_onehotd[1]};
  assign lizzieLet45_6QNode_Bool_d = {sc_0_1_goMux_mux_d[16:1],
                                      sc_0_1_goMux_mux_onehotd[2]};
  assign lizzieLet45_6QError_Bool_d = {sc_0_1_goMux_mux_d[16:1],
                                       sc_0_1_goMux_mux_onehotd[3]};
  assign sc_0_1_goMux_mux_r = (| (sc_0_1_goMux_mux_onehotd & {lizzieLet45_6QError_Bool_r,
                                                              lizzieLet45_6QNode_Bool_r,
                                                              lizzieLet45_6QVal_Bool_r,
                                                              lizzieLet45_6QNone_Bool_r}));
  assign lizzieLet45_6_r = sc_0_1_goMux_mux_r;
  
  /* buf (Ty Pointer_CTf'''''''''''') : (lizzieLet45_6QError_Bool,Pointer_CTf'''''''''''') > (lizzieLet45_6QError_Bool_1_argbuf,Pointer_CTf'''''''''''') */
  \Pointer_CTf''''''''''''_t  lizzieLet45_6QError_Bool_bufchan_d;
  logic lizzieLet45_6QError_Bool_bufchan_r;
  assign lizzieLet45_6QError_Bool_r = ((! lizzieLet45_6QError_Bool_bufchan_d[0]) || lizzieLet45_6QError_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet45_6QError_Bool_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet45_6QError_Bool_r)
        lizzieLet45_6QError_Bool_bufchan_d <= lizzieLet45_6QError_Bool_d;
  \Pointer_CTf''''''''''''_t  lizzieLet45_6QError_Bool_bufchan_buf;
  assign lizzieLet45_6QError_Bool_bufchan_r = (! lizzieLet45_6QError_Bool_bufchan_buf[0]);
  assign lizzieLet45_6QError_Bool_1_argbuf_d = (lizzieLet45_6QError_Bool_bufchan_buf[0] ? lizzieLet45_6QError_Bool_bufchan_buf :
                                                lizzieLet45_6QError_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet45_6QError_Bool_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet45_6QError_Bool_1_argbuf_r && lizzieLet45_6QError_Bool_bufchan_buf[0]))
        lizzieLet45_6QError_Bool_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet45_6QError_Bool_1_argbuf_r) && (! lizzieLet45_6QError_Bool_bufchan_buf[0])))
        lizzieLet45_6QError_Bool_bufchan_buf <= lizzieLet45_6QError_Bool_bufchan_d;
  
  /* buf (Ty Pointer_CTf'''''''''''') : (lizzieLet45_6QNone_Bool,Pointer_CTf'''''''''''') > (lizzieLet45_6QNone_Bool_1_argbuf,Pointer_CTf'''''''''''') */
  \Pointer_CTf''''''''''''_t  lizzieLet45_6QNone_Bool_bufchan_d;
  logic lizzieLet45_6QNone_Bool_bufchan_r;
  assign lizzieLet45_6QNone_Bool_r = ((! lizzieLet45_6QNone_Bool_bufchan_d[0]) || lizzieLet45_6QNone_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet45_6QNone_Bool_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet45_6QNone_Bool_r)
        lizzieLet45_6QNone_Bool_bufchan_d <= lizzieLet45_6QNone_Bool_d;
  \Pointer_CTf''''''''''''_t  lizzieLet45_6QNone_Bool_bufchan_buf;
  assign lizzieLet45_6QNone_Bool_bufchan_r = (! lizzieLet45_6QNone_Bool_bufchan_buf[0]);
  assign lizzieLet45_6QNone_Bool_1_argbuf_d = (lizzieLet45_6QNone_Bool_bufchan_buf[0] ? lizzieLet45_6QNone_Bool_bufchan_buf :
                                               lizzieLet45_6QNone_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet45_6QNone_Bool_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet45_6QNone_Bool_1_argbuf_r && lizzieLet45_6QNone_Bool_bufchan_buf[0]))
        lizzieLet45_6QNone_Bool_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet45_6QNone_Bool_1_argbuf_r) && (! lizzieLet45_6QNone_Bool_bufchan_buf[0])))
        lizzieLet45_6QNone_Bool_bufchan_buf <= lizzieLet45_6QNone_Bool_bufchan_d;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_QTree_Bool) : (lizzieLet45_7,QTree_Bool) (t4a91_2,Pointer_QTree_Bool) > [(lizzieLet45_7QNone_Bool,Pointer_QTree_Bool),
                                                                                           (_6,Pointer_QTree_Bool),
                                                                                           (_5,Pointer_QTree_Bool),
                                                                                           (_4,Pointer_QTree_Bool)] */
  logic [3:0] t4a91_2_onehotd;
  always_comb
    if ((lizzieLet45_7_d[0] && t4a91_2_d[0]))
      unique case (lizzieLet45_7_d[2:1])
        2'd0: t4a91_2_onehotd = 4'd1;
        2'd1: t4a91_2_onehotd = 4'd2;
        2'd2: t4a91_2_onehotd = 4'd4;
        2'd3: t4a91_2_onehotd = 4'd8;
        default: t4a91_2_onehotd = 4'd0;
      endcase
    else t4a91_2_onehotd = 4'd0;
  assign lizzieLet45_7QNone_Bool_d = {t4a91_2_d[16:1],
                                      t4a91_2_onehotd[0]};
  assign _6_d = {t4a91_2_d[16:1], t4a91_2_onehotd[1]};
  assign _5_d = {t4a91_2_d[16:1], t4a91_2_onehotd[2]};
  assign _4_d = {t4a91_2_d[16:1], t4a91_2_onehotd[3]};
  assign t4a91_2_r = (| (t4a91_2_onehotd & {_4_r,
                                            _5_r,
                                            _6_r,
                                            lizzieLet45_7QNone_Bool_r}));
  assign lizzieLet45_7_r = t4a91_2_r;
  
  /* buf (Ty Pointer_QTree_Bool) : (lizzieLet45_7QNone_Bool,Pointer_QTree_Bool) > (lizzieLet45_7QNone_Bool_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t lizzieLet45_7QNone_Bool_bufchan_d;
  logic lizzieLet45_7QNone_Bool_bufchan_r;
  assign lizzieLet45_7QNone_Bool_r = ((! lizzieLet45_7QNone_Bool_bufchan_d[0]) || lizzieLet45_7QNone_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet45_7QNone_Bool_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet45_7QNone_Bool_r)
        lizzieLet45_7QNone_Bool_bufchan_d <= lizzieLet45_7QNone_Bool_d;
  Pointer_QTree_Bool_t lizzieLet45_7QNone_Bool_bufchan_buf;
  assign lizzieLet45_7QNone_Bool_bufchan_r = (! lizzieLet45_7QNone_Bool_bufchan_buf[0]);
  assign lizzieLet45_7QNone_Bool_1_argbuf_d = (lizzieLet45_7QNone_Bool_bufchan_buf[0] ? lizzieLet45_7QNone_Bool_bufchan_buf :
                                               lizzieLet45_7QNone_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet45_7QNone_Bool_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet45_7QNone_Bool_1_argbuf_r && lizzieLet45_7QNone_Bool_bufchan_buf[0]))
        lizzieLet45_7QNone_Bool_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet45_7QNone_Bool_1_argbuf_r) && (! lizzieLet45_7QNone_Bool_bufchan_buf[0])))
        lizzieLet45_7QNone_Bool_bufchan_buf <= lizzieLet45_7QNone_Bool_bufchan_d;
  
  /* destruct (Ty CTf,
          Dcon Lcall_f0) : (lizzieLet60_1Lcall_f0,CTf) > [(es_13_destruct,Pointer_QTree_Bool),
                                                          (es_14_1_destruct,Pointer_QTree_Bool),
                                                          (es_15_2_destruct,Pointer_QTree_Bool),
                                                          (sc_0_5_destruct,Pointer_CTf)] */
  logic [3:0] lizzieLet60_1Lcall_f0_emitted;
  logic [3:0] lizzieLet60_1Lcall_f0_done;
  assign es_13_destruct_d = {lizzieLet60_1Lcall_f0_d[19:4],
                             (lizzieLet60_1Lcall_f0_d[0] && (! lizzieLet60_1Lcall_f0_emitted[0]))};
  assign es_14_1_destruct_d = {lizzieLet60_1Lcall_f0_d[35:20],
                               (lizzieLet60_1Lcall_f0_d[0] && (! lizzieLet60_1Lcall_f0_emitted[1]))};
  assign es_15_2_destruct_d = {lizzieLet60_1Lcall_f0_d[51:36],
                               (lizzieLet60_1Lcall_f0_d[0] && (! lizzieLet60_1Lcall_f0_emitted[2]))};
  assign sc_0_5_destruct_d = {lizzieLet60_1Lcall_f0_d[67:52],
                              (lizzieLet60_1Lcall_f0_d[0] && (! lizzieLet60_1Lcall_f0_emitted[3]))};
  assign lizzieLet60_1Lcall_f0_done = (lizzieLet60_1Lcall_f0_emitted | ({sc_0_5_destruct_d[0],
                                                                         es_15_2_destruct_d[0],
                                                                         es_14_1_destruct_d[0],
                                                                         es_13_destruct_d[0]} & {sc_0_5_destruct_r,
                                                                                                 es_15_2_destruct_r,
                                                                                                 es_14_1_destruct_r,
                                                                                                 es_13_destruct_r}));
  assign lizzieLet60_1Lcall_f0_r = (& lizzieLet60_1Lcall_f0_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet60_1Lcall_f0_emitted <= 4'd0;
    else
      lizzieLet60_1Lcall_f0_emitted <= (lizzieLet60_1Lcall_f0_r ? 4'd0 :
                                        lizzieLet60_1Lcall_f0_done);
  
  /* destruct (Ty CTf,
          Dcon Lcall_f1) : (lizzieLet60_1Lcall_f1,CTf) > [(es_14_destruct,Pointer_QTree_Bool),
                                                          (es_15_1_destruct,Pointer_QTree_Bool),
                                                          (sc_0_4_destruct,Pointer_CTf),
                                                          (q1a8H_3_destruct,Pointer_QTree_Bool),
                                                          (t1a8R_3_destruct,Pointer_QTree_Bool),
                                                          (t1'a8W_3_destruct,Pointer_QTree_Bool)] */
  logic [5:0] lizzieLet60_1Lcall_f1_emitted;
  logic [5:0] lizzieLet60_1Lcall_f1_done;
  assign es_14_destruct_d = {lizzieLet60_1Lcall_f1_d[19:4],
                             (lizzieLet60_1Lcall_f1_d[0] && (! lizzieLet60_1Lcall_f1_emitted[0]))};
  assign es_15_1_destruct_d = {lizzieLet60_1Lcall_f1_d[35:20],
                               (lizzieLet60_1Lcall_f1_d[0] && (! lizzieLet60_1Lcall_f1_emitted[1]))};
  assign sc_0_4_destruct_d = {lizzieLet60_1Lcall_f1_d[51:36],
                              (lizzieLet60_1Lcall_f1_d[0] && (! lizzieLet60_1Lcall_f1_emitted[2]))};
  assign q1a8H_3_destruct_d = {lizzieLet60_1Lcall_f1_d[67:52],
                               (lizzieLet60_1Lcall_f1_d[0] && (! lizzieLet60_1Lcall_f1_emitted[3]))};
  assign t1a8R_3_destruct_d = {lizzieLet60_1Lcall_f1_d[83:68],
                               (lizzieLet60_1Lcall_f1_d[0] && (! lizzieLet60_1Lcall_f1_emitted[4]))};
  assign \t1'a8W_3_destruct_d  = {lizzieLet60_1Lcall_f1_d[99:84],
                                  (lizzieLet60_1Lcall_f1_d[0] && (! lizzieLet60_1Lcall_f1_emitted[5]))};
  assign lizzieLet60_1Lcall_f1_done = (lizzieLet60_1Lcall_f1_emitted | ({\t1'a8W_3_destruct_d [0],
                                                                         t1a8R_3_destruct_d[0],
                                                                         q1a8H_3_destruct_d[0],
                                                                         sc_0_4_destruct_d[0],
                                                                         es_15_1_destruct_d[0],
                                                                         es_14_destruct_d[0]} & {\t1'a8W_3_destruct_r ,
                                                                                                 t1a8R_3_destruct_r,
                                                                                                 q1a8H_3_destruct_r,
                                                                                                 sc_0_4_destruct_r,
                                                                                                 es_15_1_destruct_r,
                                                                                                 es_14_destruct_r}));
  assign lizzieLet60_1Lcall_f1_r = (& lizzieLet60_1Lcall_f1_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet60_1Lcall_f1_emitted <= 6'd0;
    else
      lizzieLet60_1Lcall_f1_emitted <= (lizzieLet60_1Lcall_f1_r ? 6'd0 :
                                        lizzieLet60_1Lcall_f1_done);
  
  /* destruct (Ty CTf,
          Dcon Lcall_f2) : (lizzieLet60_1Lcall_f2,CTf) > [(es_15_destruct,Pointer_QTree_Bool),
                                                          (sc_0_3_destruct,Pointer_CTf),
                                                          (q1a8H_2_destruct,Pointer_QTree_Bool),
                                                          (t1a8R_2_destruct,Pointer_QTree_Bool),
                                                          (t1'a8W_2_destruct,Pointer_QTree_Bool),
                                                          (q2a8I_2_destruct,Pointer_QTree_Bool),
                                                          (t2a8S_2_destruct,Pointer_QTree_Bool),
                                                          (t2'a8X_2_destruct,Pointer_QTree_Bool)] */
  logic [7:0] lizzieLet60_1Lcall_f2_emitted;
  logic [7:0] lizzieLet60_1Lcall_f2_done;
  assign es_15_destruct_d = {lizzieLet60_1Lcall_f2_d[19:4],
                             (lizzieLet60_1Lcall_f2_d[0] && (! lizzieLet60_1Lcall_f2_emitted[0]))};
  assign sc_0_3_destruct_d = {lizzieLet60_1Lcall_f2_d[35:20],
                              (lizzieLet60_1Lcall_f2_d[0] && (! lizzieLet60_1Lcall_f2_emitted[1]))};
  assign q1a8H_2_destruct_d = {lizzieLet60_1Lcall_f2_d[51:36],
                               (lizzieLet60_1Lcall_f2_d[0] && (! lizzieLet60_1Lcall_f2_emitted[2]))};
  assign t1a8R_2_destruct_d = {lizzieLet60_1Lcall_f2_d[67:52],
                               (lizzieLet60_1Lcall_f2_d[0] && (! lizzieLet60_1Lcall_f2_emitted[3]))};
  assign \t1'a8W_2_destruct_d  = {lizzieLet60_1Lcall_f2_d[83:68],
                                  (lizzieLet60_1Lcall_f2_d[0] && (! lizzieLet60_1Lcall_f2_emitted[4]))};
  assign q2a8I_2_destruct_d = {lizzieLet60_1Lcall_f2_d[99:84],
                               (lizzieLet60_1Lcall_f2_d[0] && (! lizzieLet60_1Lcall_f2_emitted[5]))};
  assign t2a8S_2_destruct_d = {lizzieLet60_1Lcall_f2_d[115:100],
                               (lizzieLet60_1Lcall_f2_d[0] && (! lizzieLet60_1Lcall_f2_emitted[6]))};
  assign \t2'a8X_2_destruct_d  = {lizzieLet60_1Lcall_f2_d[131:116],
                                  (lizzieLet60_1Lcall_f2_d[0] && (! lizzieLet60_1Lcall_f2_emitted[7]))};
  assign lizzieLet60_1Lcall_f2_done = (lizzieLet60_1Lcall_f2_emitted | ({\t2'a8X_2_destruct_d [0],
                                                                         t2a8S_2_destruct_d[0],
                                                                         q2a8I_2_destruct_d[0],
                                                                         \t1'a8W_2_destruct_d [0],
                                                                         t1a8R_2_destruct_d[0],
                                                                         q1a8H_2_destruct_d[0],
                                                                         sc_0_3_destruct_d[0],
                                                                         es_15_destruct_d[0]} & {\t2'a8X_2_destruct_r ,
                                                                                                 t2a8S_2_destruct_r,
                                                                                                 q2a8I_2_destruct_r,
                                                                                                 \t1'a8W_2_destruct_r ,
                                                                                                 t1a8R_2_destruct_r,
                                                                                                 q1a8H_2_destruct_r,
                                                                                                 sc_0_3_destruct_r,
                                                                                                 es_15_destruct_r}));
  assign lizzieLet60_1Lcall_f2_r = (& lizzieLet60_1Lcall_f2_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet60_1Lcall_f2_emitted <= 8'd0;
    else
      lizzieLet60_1Lcall_f2_emitted <= (lizzieLet60_1Lcall_f2_r ? 8'd0 :
                                        lizzieLet60_1Lcall_f2_done);
  
  /* destruct (Ty CTf,
          Dcon Lcall_f3) : (lizzieLet60_1Lcall_f3,CTf) > [(sc_0_2_destruct,Pointer_CTf),
                                                          (q1a8H_1_destruct,Pointer_QTree_Bool),
                                                          (t1a8R_1_destruct,Pointer_QTree_Bool),
                                                          (t1'a8W_1_destruct,Pointer_QTree_Bool),
                                                          (q2a8I_1_destruct,Pointer_QTree_Bool),
                                                          (t2a8S_1_destruct,Pointer_QTree_Bool),
                                                          (t2'a8X_1_destruct,Pointer_QTree_Bool),
                                                          (q3a8J_1_destruct,Pointer_QTree_Bool),
                                                          (t3a8T_1_destruct,Pointer_QTree_Bool),
                                                          (t3'a8Y_1_destruct,Pointer_QTree_Bool)] */
  logic [9:0] lizzieLet60_1Lcall_f3_emitted;
  logic [9:0] lizzieLet60_1Lcall_f3_done;
  assign sc_0_2_destruct_d = {lizzieLet60_1Lcall_f3_d[19:4],
                              (lizzieLet60_1Lcall_f3_d[0] && (! lizzieLet60_1Lcall_f3_emitted[0]))};
  assign q1a8H_1_destruct_d = {lizzieLet60_1Lcall_f3_d[35:20],
                               (lizzieLet60_1Lcall_f3_d[0] && (! lizzieLet60_1Lcall_f3_emitted[1]))};
  assign t1a8R_1_destruct_d = {lizzieLet60_1Lcall_f3_d[51:36],
                               (lizzieLet60_1Lcall_f3_d[0] && (! lizzieLet60_1Lcall_f3_emitted[2]))};
  assign \t1'a8W_1_destruct_d  = {lizzieLet60_1Lcall_f3_d[67:52],
                                  (lizzieLet60_1Lcall_f3_d[0] && (! lizzieLet60_1Lcall_f3_emitted[3]))};
  assign q2a8I_1_destruct_d = {lizzieLet60_1Lcall_f3_d[83:68],
                               (lizzieLet60_1Lcall_f3_d[0] && (! lizzieLet60_1Lcall_f3_emitted[4]))};
  assign t2a8S_1_destruct_d = {lizzieLet60_1Lcall_f3_d[99:84],
                               (lizzieLet60_1Lcall_f3_d[0] && (! lizzieLet60_1Lcall_f3_emitted[5]))};
  assign \t2'a8X_1_destruct_d  = {lizzieLet60_1Lcall_f3_d[115:100],
                                  (lizzieLet60_1Lcall_f3_d[0] && (! lizzieLet60_1Lcall_f3_emitted[6]))};
  assign q3a8J_1_destruct_d = {lizzieLet60_1Lcall_f3_d[131:116],
                               (lizzieLet60_1Lcall_f3_d[0] && (! lizzieLet60_1Lcall_f3_emitted[7]))};
  assign t3a8T_1_destruct_d = {lizzieLet60_1Lcall_f3_d[147:132],
                               (lizzieLet60_1Lcall_f3_d[0] && (! lizzieLet60_1Lcall_f3_emitted[8]))};
  assign \t3'a8Y_1_destruct_d  = {lizzieLet60_1Lcall_f3_d[163:148],
                                  (lizzieLet60_1Lcall_f3_d[0] && (! lizzieLet60_1Lcall_f3_emitted[9]))};
  assign lizzieLet60_1Lcall_f3_done = (lizzieLet60_1Lcall_f3_emitted | ({\t3'a8Y_1_destruct_d [0],
                                                                         t3a8T_1_destruct_d[0],
                                                                         q3a8J_1_destruct_d[0],
                                                                         \t2'a8X_1_destruct_d [0],
                                                                         t2a8S_1_destruct_d[0],
                                                                         q2a8I_1_destruct_d[0],
                                                                         \t1'a8W_1_destruct_d [0],
                                                                         t1a8R_1_destruct_d[0],
                                                                         q1a8H_1_destruct_d[0],
                                                                         sc_0_2_destruct_d[0]} & {\t3'a8Y_1_destruct_r ,
                                                                                                  t3a8T_1_destruct_r,
                                                                                                  q3a8J_1_destruct_r,
                                                                                                  \t2'a8X_1_destruct_r ,
                                                                                                  t2a8S_1_destruct_r,
                                                                                                  q2a8I_1_destruct_r,
                                                                                                  \t1'a8W_1_destruct_r ,
                                                                                                  t1a8R_1_destruct_r,
                                                                                                  q1a8H_1_destruct_r,
                                                                                                  sc_0_2_destruct_r}));
  assign lizzieLet60_1Lcall_f3_r = (& lizzieLet60_1Lcall_f3_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet60_1Lcall_f3_emitted <= 10'd0;
    else
      lizzieLet60_1Lcall_f3_emitted <= (lizzieLet60_1Lcall_f3_r ? 10'd0 :
                                        lizzieLet60_1Lcall_f3_done);
  
  /* demux (Ty CTf,
       Ty CTf) : (lizzieLet60_2,CTf) (lizzieLet60_1,CTf) > [(_3,CTf),
                                                            (lizzieLet60_1Lcall_f3,CTf),
                                                            (lizzieLet60_1Lcall_f2,CTf),
                                                            (lizzieLet60_1Lcall_f1,CTf),
                                                            (lizzieLet60_1Lcall_f0,CTf)] */
  logic [4:0] lizzieLet60_1_onehotd;
  always_comb
    if ((lizzieLet60_2_d[0] && lizzieLet60_1_d[0]))
      unique case (lizzieLet60_2_d[3:1])
        3'd0: lizzieLet60_1_onehotd = 5'd1;
        3'd1: lizzieLet60_1_onehotd = 5'd2;
        3'd2: lizzieLet60_1_onehotd = 5'd4;
        3'd3: lizzieLet60_1_onehotd = 5'd8;
        3'd4: lizzieLet60_1_onehotd = 5'd16;
        default: lizzieLet60_1_onehotd = 5'd0;
      endcase
    else lizzieLet60_1_onehotd = 5'd0;
  assign _3_d = {lizzieLet60_1_d[163:1], lizzieLet60_1_onehotd[0]};
  assign lizzieLet60_1Lcall_f3_d = {lizzieLet60_1_d[163:1],
                                    lizzieLet60_1_onehotd[1]};
  assign lizzieLet60_1Lcall_f2_d = {lizzieLet60_1_d[163:1],
                                    lizzieLet60_1_onehotd[2]};
  assign lizzieLet60_1Lcall_f1_d = {lizzieLet60_1_d[163:1],
                                    lizzieLet60_1_onehotd[3]};
  assign lizzieLet60_1Lcall_f0_d = {lizzieLet60_1_d[163:1],
                                    lizzieLet60_1_onehotd[4]};
  assign lizzieLet60_1_r = (| (lizzieLet60_1_onehotd & {lizzieLet60_1Lcall_f0_r,
                                                        lizzieLet60_1Lcall_f1_r,
                                                        lizzieLet60_1Lcall_f2_r,
                                                        lizzieLet60_1Lcall_f3_r,
                                                        _3_r}));
  assign lizzieLet60_2_r = lizzieLet60_1_r;
  
  /* demux (Ty CTf,
       Ty Go) : (lizzieLet60_3,CTf) (go_7_goMux_data,Go) > [(_2,Go),
                                                            (lizzieLet60_3Lcall_f3,Go),
                                                            (lizzieLet60_3Lcall_f2,Go),
                                                            (lizzieLet60_3Lcall_f1,Go),
                                                            (lizzieLet60_3Lcall_f0,Go)] */
  logic [4:0] go_7_goMux_data_onehotd;
  always_comb
    if ((lizzieLet60_3_d[0] && go_7_goMux_data_d[0]))
      unique case (lizzieLet60_3_d[3:1])
        3'd0: go_7_goMux_data_onehotd = 5'd1;
        3'd1: go_7_goMux_data_onehotd = 5'd2;
        3'd2: go_7_goMux_data_onehotd = 5'd4;
        3'd3: go_7_goMux_data_onehotd = 5'd8;
        3'd4: go_7_goMux_data_onehotd = 5'd16;
        default: go_7_goMux_data_onehotd = 5'd0;
      endcase
    else go_7_goMux_data_onehotd = 5'd0;
  assign _2_d = go_7_goMux_data_onehotd[0];
  assign lizzieLet60_3Lcall_f3_d = go_7_goMux_data_onehotd[1];
  assign lizzieLet60_3Lcall_f2_d = go_7_goMux_data_onehotd[2];
  assign lizzieLet60_3Lcall_f1_d = go_7_goMux_data_onehotd[3];
  assign lizzieLet60_3Lcall_f0_d = go_7_goMux_data_onehotd[4];
  assign go_7_goMux_data_r = (| (go_7_goMux_data_onehotd & {lizzieLet60_3Lcall_f0_r,
                                                            lizzieLet60_3Lcall_f1_r,
                                                            lizzieLet60_3Lcall_f2_r,
                                                            lizzieLet60_3Lcall_f3_r,
                                                            _2_r}));
  assign lizzieLet60_3_r = go_7_goMux_data_r;
  
  /* buf (Ty Go) : (lizzieLet60_3Lcall_f0,Go) > (lizzieLet60_3Lcall_f0_1_argbuf,Go) */
  Go_t lizzieLet60_3Lcall_f0_bufchan_d;
  logic lizzieLet60_3Lcall_f0_bufchan_r;
  assign lizzieLet60_3Lcall_f0_r = ((! lizzieLet60_3Lcall_f0_bufchan_d[0]) || lizzieLet60_3Lcall_f0_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet60_3Lcall_f0_bufchan_d <= 1'd0;
    else
      if (lizzieLet60_3Lcall_f0_r)
        lizzieLet60_3Lcall_f0_bufchan_d <= lizzieLet60_3Lcall_f0_d;
  Go_t lizzieLet60_3Lcall_f0_bufchan_buf;
  assign lizzieLet60_3Lcall_f0_bufchan_r = (! lizzieLet60_3Lcall_f0_bufchan_buf[0]);
  assign lizzieLet60_3Lcall_f0_1_argbuf_d = (lizzieLet60_3Lcall_f0_bufchan_buf[0] ? lizzieLet60_3Lcall_f0_bufchan_buf :
                                             lizzieLet60_3Lcall_f0_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet60_3Lcall_f0_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet60_3Lcall_f0_1_argbuf_r && lizzieLet60_3Lcall_f0_bufchan_buf[0]))
        lizzieLet60_3Lcall_f0_bufchan_buf <= 1'd0;
      else if (((! lizzieLet60_3Lcall_f0_1_argbuf_r) && (! lizzieLet60_3Lcall_f0_bufchan_buf[0])))
        lizzieLet60_3Lcall_f0_bufchan_buf <= lizzieLet60_3Lcall_f0_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet60_3Lcall_f1,Go) > (lizzieLet60_3Lcall_f1_1_argbuf,Go) */
  Go_t lizzieLet60_3Lcall_f1_bufchan_d;
  logic lizzieLet60_3Lcall_f1_bufchan_r;
  assign lizzieLet60_3Lcall_f1_r = ((! lizzieLet60_3Lcall_f1_bufchan_d[0]) || lizzieLet60_3Lcall_f1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet60_3Lcall_f1_bufchan_d <= 1'd0;
    else
      if (lizzieLet60_3Lcall_f1_r)
        lizzieLet60_3Lcall_f1_bufchan_d <= lizzieLet60_3Lcall_f1_d;
  Go_t lizzieLet60_3Lcall_f1_bufchan_buf;
  assign lizzieLet60_3Lcall_f1_bufchan_r = (! lizzieLet60_3Lcall_f1_bufchan_buf[0]);
  assign lizzieLet60_3Lcall_f1_1_argbuf_d = (lizzieLet60_3Lcall_f1_bufchan_buf[0] ? lizzieLet60_3Lcall_f1_bufchan_buf :
                                             lizzieLet60_3Lcall_f1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet60_3Lcall_f1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet60_3Lcall_f1_1_argbuf_r && lizzieLet60_3Lcall_f1_bufchan_buf[0]))
        lizzieLet60_3Lcall_f1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet60_3Lcall_f1_1_argbuf_r) && (! lizzieLet60_3Lcall_f1_bufchan_buf[0])))
        lizzieLet60_3Lcall_f1_bufchan_buf <= lizzieLet60_3Lcall_f1_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet60_3Lcall_f2,Go) > (lizzieLet60_3Lcall_f2_1_argbuf,Go) */
  Go_t lizzieLet60_3Lcall_f2_bufchan_d;
  logic lizzieLet60_3Lcall_f2_bufchan_r;
  assign lizzieLet60_3Lcall_f2_r = ((! lizzieLet60_3Lcall_f2_bufchan_d[0]) || lizzieLet60_3Lcall_f2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet60_3Lcall_f2_bufchan_d <= 1'd0;
    else
      if (lizzieLet60_3Lcall_f2_r)
        lizzieLet60_3Lcall_f2_bufchan_d <= lizzieLet60_3Lcall_f2_d;
  Go_t lizzieLet60_3Lcall_f2_bufchan_buf;
  assign lizzieLet60_3Lcall_f2_bufchan_r = (! lizzieLet60_3Lcall_f2_bufchan_buf[0]);
  assign lizzieLet60_3Lcall_f2_1_argbuf_d = (lizzieLet60_3Lcall_f2_bufchan_buf[0] ? lizzieLet60_3Lcall_f2_bufchan_buf :
                                             lizzieLet60_3Lcall_f2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet60_3Lcall_f2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet60_3Lcall_f2_1_argbuf_r && lizzieLet60_3Lcall_f2_bufchan_buf[0]))
        lizzieLet60_3Lcall_f2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet60_3Lcall_f2_1_argbuf_r) && (! lizzieLet60_3Lcall_f2_bufchan_buf[0])))
        lizzieLet60_3Lcall_f2_bufchan_buf <= lizzieLet60_3Lcall_f2_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet60_3Lcall_f3,Go) > (lizzieLet60_3Lcall_f3_1_argbuf,Go) */
  Go_t lizzieLet60_3Lcall_f3_bufchan_d;
  logic lizzieLet60_3Lcall_f3_bufchan_r;
  assign lizzieLet60_3Lcall_f3_r = ((! lizzieLet60_3Lcall_f3_bufchan_d[0]) || lizzieLet60_3Lcall_f3_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet60_3Lcall_f3_bufchan_d <= 1'd0;
    else
      if (lizzieLet60_3Lcall_f3_r)
        lizzieLet60_3Lcall_f3_bufchan_d <= lizzieLet60_3Lcall_f3_d;
  Go_t lizzieLet60_3Lcall_f3_bufchan_buf;
  assign lizzieLet60_3Lcall_f3_bufchan_r = (! lizzieLet60_3Lcall_f3_bufchan_buf[0]);
  assign lizzieLet60_3Lcall_f3_1_argbuf_d = (lizzieLet60_3Lcall_f3_bufchan_buf[0] ? lizzieLet60_3Lcall_f3_bufchan_buf :
                                             lizzieLet60_3Lcall_f3_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet60_3Lcall_f3_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet60_3Lcall_f3_1_argbuf_r && lizzieLet60_3Lcall_f3_bufchan_buf[0]))
        lizzieLet60_3Lcall_f3_bufchan_buf <= 1'd0;
      else if (((! lizzieLet60_3Lcall_f3_1_argbuf_r) && (! lizzieLet60_3Lcall_f3_bufchan_buf[0])))
        lizzieLet60_3Lcall_f3_bufchan_buf <= lizzieLet60_3Lcall_f3_bufchan_d;
  
  /* demux (Ty CTf,
       Ty Pointer_QTree_Bool) : (lizzieLet60_4,CTf) (srtarg_0_goMux_mux,Pointer_QTree_Bool) > [(lizzieLet60_4Lfsbos,Pointer_QTree_Bool),
                                                                                               (lizzieLet60_4Lcall_f3,Pointer_QTree_Bool),
                                                                                               (lizzieLet60_4Lcall_f2,Pointer_QTree_Bool),
                                                                                               (lizzieLet60_4Lcall_f1,Pointer_QTree_Bool),
                                                                                               (lizzieLet60_4Lcall_f0,Pointer_QTree_Bool)] */
  logic [4:0] srtarg_0_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet60_4_d[0] && srtarg_0_goMux_mux_d[0]))
      unique case (lizzieLet60_4_d[3:1])
        3'd0: srtarg_0_goMux_mux_onehotd = 5'd1;
        3'd1: srtarg_0_goMux_mux_onehotd = 5'd2;
        3'd2: srtarg_0_goMux_mux_onehotd = 5'd4;
        3'd3: srtarg_0_goMux_mux_onehotd = 5'd8;
        3'd4: srtarg_0_goMux_mux_onehotd = 5'd16;
        default: srtarg_0_goMux_mux_onehotd = 5'd0;
      endcase
    else srtarg_0_goMux_mux_onehotd = 5'd0;
  assign lizzieLet60_4Lfsbos_d = {srtarg_0_goMux_mux_d[16:1],
                                  srtarg_0_goMux_mux_onehotd[0]};
  assign lizzieLet60_4Lcall_f3_d = {srtarg_0_goMux_mux_d[16:1],
                                    srtarg_0_goMux_mux_onehotd[1]};
  assign lizzieLet60_4Lcall_f2_d = {srtarg_0_goMux_mux_d[16:1],
                                    srtarg_0_goMux_mux_onehotd[2]};
  assign lizzieLet60_4Lcall_f1_d = {srtarg_0_goMux_mux_d[16:1],
                                    srtarg_0_goMux_mux_onehotd[3]};
  assign lizzieLet60_4Lcall_f0_d = {srtarg_0_goMux_mux_d[16:1],
                                    srtarg_0_goMux_mux_onehotd[4]};
  assign srtarg_0_goMux_mux_r = (| (srtarg_0_goMux_mux_onehotd & {lizzieLet60_4Lcall_f0_r,
                                                                  lizzieLet60_4Lcall_f1_r,
                                                                  lizzieLet60_4Lcall_f2_r,
                                                                  lizzieLet60_4Lcall_f3_r,
                                                                  lizzieLet60_4Lfsbos_r}));
  assign lizzieLet60_4_r = srtarg_0_goMux_mux_r;
  
  /* dcon (Ty QTree_Bool,
      Dcon QNode_Bool) : [(lizzieLet60_4Lcall_f0,Pointer_QTree_Bool),
                          (es_13_destruct,Pointer_QTree_Bool),
                          (es_14_1_destruct,Pointer_QTree_Bool),
                          (es_15_2_destruct,Pointer_QTree_Bool)] > (lizzieLet60_4Lcall_f0_1es_13_1es_14_1_1es_15_2_1QNode_Bool,QTree_Bool) */
  assign lizzieLet60_4Lcall_f0_1es_13_1es_14_1_1es_15_2_1QNode_Bool_d = QNode_Bool_dc((& {lizzieLet60_4Lcall_f0_d[0],
                                                                                          es_13_destruct_d[0],
                                                                                          es_14_1_destruct_d[0],
                                                                                          es_15_2_destruct_d[0]}), lizzieLet60_4Lcall_f0_d, es_13_destruct_d, es_14_1_destruct_d, es_15_2_destruct_d);
  assign {lizzieLet60_4Lcall_f0_r,
          es_13_destruct_r,
          es_14_1_destruct_r,
          es_15_2_destruct_r} = {4 {(lizzieLet60_4Lcall_f0_1es_13_1es_14_1_1es_15_2_1QNode_Bool_r && lizzieLet60_4Lcall_f0_1es_13_1es_14_1_1es_15_2_1QNode_Bool_d[0])}};
  
  /* buf (Ty QTree_Bool) : (lizzieLet60_4Lcall_f0_1es_13_1es_14_1_1es_15_2_1QNode_Bool,QTree_Bool) > (lizzieLet64_1_argbuf,QTree_Bool) */
  QTree_Bool_t lizzieLet60_4Lcall_f0_1es_13_1es_14_1_1es_15_2_1QNode_Bool_bufchan_d;
  logic lizzieLet60_4Lcall_f0_1es_13_1es_14_1_1es_15_2_1QNode_Bool_bufchan_r;
  assign lizzieLet60_4Lcall_f0_1es_13_1es_14_1_1es_15_2_1QNode_Bool_r = ((! lizzieLet60_4Lcall_f0_1es_13_1es_14_1_1es_15_2_1QNode_Bool_bufchan_d[0]) || lizzieLet60_4Lcall_f0_1es_13_1es_14_1_1es_15_2_1QNode_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet60_4Lcall_f0_1es_13_1es_14_1_1es_15_2_1QNode_Bool_bufchan_d <= {66'd0,
                                                                               1'd0};
    else
      if (lizzieLet60_4Lcall_f0_1es_13_1es_14_1_1es_15_2_1QNode_Bool_r)
        lizzieLet60_4Lcall_f0_1es_13_1es_14_1_1es_15_2_1QNode_Bool_bufchan_d <= lizzieLet60_4Lcall_f0_1es_13_1es_14_1_1es_15_2_1QNode_Bool_d;
  QTree_Bool_t lizzieLet60_4Lcall_f0_1es_13_1es_14_1_1es_15_2_1QNode_Bool_bufchan_buf;
  assign lizzieLet60_4Lcall_f0_1es_13_1es_14_1_1es_15_2_1QNode_Bool_bufchan_r = (! lizzieLet60_4Lcall_f0_1es_13_1es_14_1_1es_15_2_1QNode_Bool_bufchan_buf[0]);
  assign lizzieLet64_1_argbuf_d = (lizzieLet60_4Lcall_f0_1es_13_1es_14_1_1es_15_2_1QNode_Bool_bufchan_buf[0] ? lizzieLet60_4Lcall_f0_1es_13_1es_14_1_1es_15_2_1QNode_Bool_bufchan_buf :
                                   lizzieLet60_4Lcall_f0_1es_13_1es_14_1_1es_15_2_1QNode_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet60_4Lcall_f0_1es_13_1es_14_1_1es_15_2_1QNode_Bool_bufchan_buf <= {66'd0,
                                                                                 1'd0};
    else
      if ((lizzieLet64_1_argbuf_r && lizzieLet60_4Lcall_f0_1es_13_1es_14_1_1es_15_2_1QNode_Bool_bufchan_buf[0]))
        lizzieLet60_4Lcall_f0_1es_13_1es_14_1_1es_15_2_1QNode_Bool_bufchan_buf <= {66'd0,
                                                                                   1'd0};
      else if (((! lizzieLet64_1_argbuf_r) && (! lizzieLet60_4Lcall_f0_1es_13_1es_14_1_1es_15_2_1QNode_Bool_bufchan_buf[0])))
        lizzieLet60_4Lcall_f0_1es_13_1es_14_1_1es_15_2_1QNode_Bool_bufchan_buf <= lizzieLet60_4Lcall_f0_1es_13_1es_14_1_1es_15_2_1QNode_Bool_bufchan_d;
  
  /* dcon (Ty CTf,
      Dcon Lcall_f0) : [(lizzieLet60_4Lcall_f1,Pointer_QTree_Bool),
                        (es_14_destruct,Pointer_QTree_Bool),
                        (es_15_1_destruct,Pointer_QTree_Bool),
                        (sc_0_4_destruct,Pointer_CTf)] > (lizzieLet60_4Lcall_f1_1es_14_1es_15_1_1sc_0_4_1Lcall_f0,CTf) */
  assign lizzieLet60_4Lcall_f1_1es_14_1es_15_1_1sc_0_4_1Lcall_f0_d = Lcall_f0_dc((& {lizzieLet60_4Lcall_f1_d[0],
                                                                                     es_14_destruct_d[0],
                                                                                     es_15_1_destruct_d[0],
                                                                                     sc_0_4_destruct_d[0]}), lizzieLet60_4Lcall_f1_d, es_14_destruct_d, es_15_1_destruct_d, sc_0_4_destruct_d);
  assign {lizzieLet60_4Lcall_f1_r,
          es_14_destruct_r,
          es_15_1_destruct_r,
          sc_0_4_destruct_r} = {4 {(lizzieLet60_4Lcall_f1_1es_14_1es_15_1_1sc_0_4_1Lcall_f0_r && lizzieLet60_4Lcall_f1_1es_14_1es_15_1_1sc_0_4_1Lcall_f0_d[0])}};
  
  /* buf (Ty CTf) : (lizzieLet60_4Lcall_f1_1es_14_1es_15_1_1sc_0_4_1Lcall_f0,CTf) > (lizzieLet63_1_argbuf,CTf) */
  CTf_t lizzieLet60_4Lcall_f1_1es_14_1es_15_1_1sc_0_4_1Lcall_f0_bufchan_d;
  logic lizzieLet60_4Lcall_f1_1es_14_1es_15_1_1sc_0_4_1Lcall_f0_bufchan_r;
  assign lizzieLet60_4Lcall_f1_1es_14_1es_15_1_1sc_0_4_1Lcall_f0_r = ((! lizzieLet60_4Lcall_f1_1es_14_1es_15_1_1sc_0_4_1Lcall_f0_bufchan_d[0]) || lizzieLet60_4Lcall_f1_1es_14_1es_15_1_1sc_0_4_1Lcall_f0_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet60_4Lcall_f1_1es_14_1es_15_1_1sc_0_4_1Lcall_f0_bufchan_d <= {163'd0,
                                                                            1'd0};
    else
      if (lizzieLet60_4Lcall_f1_1es_14_1es_15_1_1sc_0_4_1Lcall_f0_r)
        lizzieLet60_4Lcall_f1_1es_14_1es_15_1_1sc_0_4_1Lcall_f0_bufchan_d <= lizzieLet60_4Lcall_f1_1es_14_1es_15_1_1sc_0_4_1Lcall_f0_d;
  CTf_t lizzieLet60_4Lcall_f1_1es_14_1es_15_1_1sc_0_4_1Lcall_f0_bufchan_buf;
  assign lizzieLet60_4Lcall_f1_1es_14_1es_15_1_1sc_0_4_1Lcall_f0_bufchan_r = (! lizzieLet60_4Lcall_f1_1es_14_1es_15_1_1sc_0_4_1Lcall_f0_bufchan_buf[0]);
  assign lizzieLet63_1_argbuf_d = (lizzieLet60_4Lcall_f1_1es_14_1es_15_1_1sc_0_4_1Lcall_f0_bufchan_buf[0] ? lizzieLet60_4Lcall_f1_1es_14_1es_15_1_1sc_0_4_1Lcall_f0_bufchan_buf :
                                   lizzieLet60_4Lcall_f1_1es_14_1es_15_1_1sc_0_4_1Lcall_f0_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet60_4Lcall_f1_1es_14_1es_15_1_1sc_0_4_1Lcall_f0_bufchan_buf <= {163'd0,
                                                                              1'd0};
    else
      if ((lizzieLet63_1_argbuf_r && lizzieLet60_4Lcall_f1_1es_14_1es_15_1_1sc_0_4_1Lcall_f0_bufchan_buf[0]))
        lizzieLet60_4Lcall_f1_1es_14_1es_15_1_1sc_0_4_1Lcall_f0_bufchan_buf <= {163'd0,
                                                                                1'd0};
      else if (((! lizzieLet63_1_argbuf_r) && (! lizzieLet60_4Lcall_f1_1es_14_1es_15_1_1sc_0_4_1Lcall_f0_bufchan_buf[0])))
        lizzieLet60_4Lcall_f1_1es_14_1es_15_1_1sc_0_4_1Lcall_f0_bufchan_buf <= lizzieLet60_4Lcall_f1_1es_14_1es_15_1_1sc_0_4_1Lcall_f0_bufchan_d;
  
  /* dcon (Ty CTf,
      Dcon Lcall_f1) : [(lizzieLet60_4Lcall_f2,Pointer_QTree_Bool),
                        (es_15_destruct,Pointer_QTree_Bool),
                        (sc_0_3_destruct,Pointer_CTf),
                        (q1a8H_2_destruct,Pointer_QTree_Bool),
                        (t1a8R_2_destruct,Pointer_QTree_Bool),
                        (t1'a8W_2_destruct,Pointer_QTree_Bool)] > (lizzieLet60_4Lcall_f2_1es_15_1sc_0_3_1q1a8H_2_1t1a8R_2_1t1'a8W_2_1Lcall_f1,CTf) */
  assign \lizzieLet60_4Lcall_f2_1es_15_1sc_0_3_1q1a8H_2_1t1a8R_2_1t1'a8W_2_1Lcall_f1_d  = Lcall_f1_dc((& {lizzieLet60_4Lcall_f2_d[0],
                                                                                                          es_15_destruct_d[0],
                                                                                                          sc_0_3_destruct_d[0],
                                                                                                          q1a8H_2_destruct_d[0],
                                                                                                          t1a8R_2_destruct_d[0],
                                                                                                          \t1'a8W_2_destruct_d [0]}), lizzieLet60_4Lcall_f2_d, es_15_destruct_d, sc_0_3_destruct_d, q1a8H_2_destruct_d, t1a8R_2_destruct_d, \t1'a8W_2_destruct_d );
  assign {lizzieLet60_4Lcall_f2_r,
          es_15_destruct_r,
          sc_0_3_destruct_r,
          q1a8H_2_destruct_r,
          t1a8R_2_destruct_r,
          \t1'a8W_2_destruct_r } = {6 {(\lizzieLet60_4Lcall_f2_1es_15_1sc_0_3_1q1a8H_2_1t1a8R_2_1t1'a8W_2_1Lcall_f1_r  && \lizzieLet60_4Lcall_f2_1es_15_1sc_0_3_1q1a8H_2_1t1a8R_2_1t1'a8W_2_1Lcall_f1_d [0])}};
  
  /* buf (Ty CTf) : (lizzieLet60_4Lcall_f2_1es_15_1sc_0_3_1q1a8H_2_1t1a8R_2_1t1'a8W_2_1Lcall_f1,CTf) > (lizzieLet62_1_argbuf,CTf) */
  CTf_t \lizzieLet60_4Lcall_f2_1es_15_1sc_0_3_1q1a8H_2_1t1a8R_2_1t1'a8W_2_1Lcall_f1_bufchan_d ;
  logic \lizzieLet60_4Lcall_f2_1es_15_1sc_0_3_1q1a8H_2_1t1a8R_2_1t1'a8W_2_1Lcall_f1_bufchan_r ;
  assign \lizzieLet60_4Lcall_f2_1es_15_1sc_0_3_1q1a8H_2_1t1a8R_2_1t1'a8W_2_1Lcall_f1_r  = ((! \lizzieLet60_4Lcall_f2_1es_15_1sc_0_3_1q1a8H_2_1t1a8R_2_1t1'a8W_2_1Lcall_f1_bufchan_d [0]) || \lizzieLet60_4Lcall_f2_1es_15_1sc_0_3_1q1a8H_2_1t1a8R_2_1t1'a8W_2_1Lcall_f1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet60_4Lcall_f2_1es_15_1sc_0_3_1q1a8H_2_1t1a8R_2_1t1'a8W_2_1Lcall_f1_bufchan_d  <= {163'd0,
                                                                                                 1'd0};
    else
      if (\lizzieLet60_4Lcall_f2_1es_15_1sc_0_3_1q1a8H_2_1t1a8R_2_1t1'a8W_2_1Lcall_f1_r )
        \lizzieLet60_4Lcall_f2_1es_15_1sc_0_3_1q1a8H_2_1t1a8R_2_1t1'a8W_2_1Lcall_f1_bufchan_d  <= \lizzieLet60_4Lcall_f2_1es_15_1sc_0_3_1q1a8H_2_1t1a8R_2_1t1'a8W_2_1Lcall_f1_d ;
  CTf_t \lizzieLet60_4Lcall_f2_1es_15_1sc_0_3_1q1a8H_2_1t1a8R_2_1t1'a8W_2_1Lcall_f1_bufchan_buf ;
  assign \lizzieLet60_4Lcall_f2_1es_15_1sc_0_3_1q1a8H_2_1t1a8R_2_1t1'a8W_2_1Lcall_f1_bufchan_r  = (! \lizzieLet60_4Lcall_f2_1es_15_1sc_0_3_1q1a8H_2_1t1a8R_2_1t1'a8W_2_1Lcall_f1_bufchan_buf [0]);
  assign lizzieLet62_1_argbuf_d = (\lizzieLet60_4Lcall_f2_1es_15_1sc_0_3_1q1a8H_2_1t1a8R_2_1t1'a8W_2_1Lcall_f1_bufchan_buf [0] ? \lizzieLet60_4Lcall_f2_1es_15_1sc_0_3_1q1a8H_2_1t1a8R_2_1t1'a8W_2_1Lcall_f1_bufchan_buf  :
                                   \lizzieLet60_4Lcall_f2_1es_15_1sc_0_3_1q1a8H_2_1t1a8R_2_1t1'a8W_2_1Lcall_f1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet60_4Lcall_f2_1es_15_1sc_0_3_1q1a8H_2_1t1a8R_2_1t1'a8W_2_1Lcall_f1_bufchan_buf  <= {163'd0,
                                                                                                   1'd0};
    else
      if ((lizzieLet62_1_argbuf_r && \lizzieLet60_4Lcall_f2_1es_15_1sc_0_3_1q1a8H_2_1t1a8R_2_1t1'a8W_2_1Lcall_f1_bufchan_buf [0]))
        \lizzieLet60_4Lcall_f2_1es_15_1sc_0_3_1q1a8H_2_1t1a8R_2_1t1'a8W_2_1Lcall_f1_bufchan_buf  <= {163'd0,
                                                                                                     1'd0};
      else if (((! lizzieLet62_1_argbuf_r) && (! \lizzieLet60_4Lcall_f2_1es_15_1sc_0_3_1q1a8H_2_1t1a8R_2_1t1'a8W_2_1Lcall_f1_bufchan_buf [0])))
        \lizzieLet60_4Lcall_f2_1es_15_1sc_0_3_1q1a8H_2_1t1a8R_2_1t1'a8W_2_1Lcall_f1_bufchan_buf  <= \lizzieLet60_4Lcall_f2_1es_15_1sc_0_3_1q1a8H_2_1t1a8R_2_1t1'a8W_2_1Lcall_f1_bufchan_d ;
  
  /* dcon (Ty CTf,
      Dcon Lcall_f2) : [(lizzieLet60_4Lcall_f3,Pointer_QTree_Bool),
                        (sc_0_2_destruct,Pointer_CTf),
                        (q1a8H_1_destruct,Pointer_QTree_Bool),
                        (t1a8R_1_destruct,Pointer_QTree_Bool),
                        (t1'a8W_1_destruct,Pointer_QTree_Bool),
                        (q2a8I_1_destruct,Pointer_QTree_Bool),
                        (t2a8S_1_destruct,Pointer_QTree_Bool),
                        (t2'a8X_1_destruct,Pointer_QTree_Bool)] > (lizzieLet60_4Lcall_f3_1sc_0_2_1q1a8H_1_1t1a8R_1_1t1'a8W_1_1q2a8I_1_1t2a8S_1_1t2'a8X_1_1Lcall_f2,CTf) */
  assign \lizzieLet60_4Lcall_f3_1sc_0_2_1q1a8H_1_1t1a8R_1_1t1'a8W_1_1q2a8I_1_1t2a8S_1_1t2'a8X_1_1Lcall_f2_d  = Lcall_f2_dc((& {lizzieLet60_4Lcall_f3_d[0],
                                                                                                                               sc_0_2_destruct_d[0],
                                                                                                                               q1a8H_1_destruct_d[0],
                                                                                                                               t1a8R_1_destruct_d[0],
                                                                                                                               \t1'a8W_1_destruct_d [0],
                                                                                                                               q2a8I_1_destruct_d[0],
                                                                                                                               t2a8S_1_destruct_d[0],
                                                                                                                               \t2'a8X_1_destruct_d [0]}), lizzieLet60_4Lcall_f3_d, sc_0_2_destruct_d, q1a8H_1_destruct_d, t1a8R_1_destruct_d, \t1'a8W_1_destruct_d , q2a8I_1_destruct_d, t2a8S_1_destruct_d, \t2'a8X_1_destruct_d );
  assign {lizzieLet60_4Lcall_f3_r,
          sc_0_2_destruct_r,
          q1a8H_1_destruct_r,
          t1a8R_1_destruct_r,
          \t1'a8W_1_destruct_r ,
          q2a8I_1_destruct_r,
          t2a8S_1_destruct_r,
          \t2'a8X_1_destruct_r } = {8 {(\lizzieLet60_4Lcall_f3_1sc_0_2_1q1a8H_1_1t1a8R_1_1t1'a8W_1_1q2a8I_1_1t2a8S_1_1t2'a8X_1_1Lcall_f2_r  && \lizzieLet60_4Lcall_f3_1sc_0_2_1q1a8H_1_1t1a8R_1_1t1'a8W_1_1q2a8I_1_1t2a8S_1_1t2'a8X_1_1Lcall_f2_d [0])}};
  
  /* buf (Ty CTf) : (lizzieLet60_4Lcall_f3_1sc_0_2_1q1a8H_1_1t1a8R_1_1t1'a8W_1_1q2a8I_1_1t2a8S_1_1t2'a8X_1_1Lcall_f2,CTf) > (lizzieLet61_1_argbuf,CTf) */
  CTf_t \lizzieLet60_4Lcall_f3_1sc_0_2_1q1a8H_1_1t1a8R_1_1t1'a8W_1_1q2a8I_1_1t2a8S_1_1t2'a8X_1_1Lcall_f2_bufchan_d ;
  logic \lizzieLet60_4Lcall_f3_1sc_0_2_1q1a8H_1_1t1a8R_1_1t1'a8W_1_1q2a8I_1_1t2a8S_1_1t2'a8X_1_1Lcall_f2_bufchan_r ;
  assign \lizzieLet60_4Lcall_f3_1sc_0_2_1q1a8H_1_1t1a8R_1_1t1'a8W_1_1q2a8I_1_1t2a8S_1_1t2'a8X_1_1Lcall_f2_r  = ((! \lizzieLet60_4Lcall_f3_1sc_0_2_1q1a8H_1_1t1a8R_1_1t1'a8W_1_1q2a8I_1_1t2a8S_1_1t2'a8X_1_1Lcall_f2_bufchan_d [0]) || \lizzieLet60_4Lcall_f3_1sc_0_2_1q1a8H_1_1t1a8R_1_1t1'a8W_1_1q2a8I_1_1t2a8S_1_1t2'a8X_1_1Lcall_f2_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet60_4Lcall_f3_1sc_0_2_1q1a8H_1_1t1a8R_1_1t1'a8W_1_1q2a8I_1_1t2a8S_1_1t2'a8X_1_1Lcall_f2_bufchan_d  <= {163'd0,
                                                                                                                      1'd0};
    else
      if (\lizzieLet60_4Lcall_f3_1sc_0_2_1q1a8H_1_1t1a8R_1_1t1'a8W_1_1q2a8I_1_1t2a8S_1_1t2'a8X_1_1Lcall_f2_r )
        \lizzieLet60_4Lcall_f3_1sc_0_2_1q1a8H_1_1t1a8R_1_1t1'a8W_1_1q2a8I_1_1t2a8S_1_1t2'a8X_1_1Lcall_f2_bufchan_d  <= \lizzieLet60_4Lcall_f3_1sc_0_2_1q1a8H_1_1t1a8R_1_1t1'a8W_1_1q2a8I_1_1t2a8S_1_1t2'a8X_1_1Lcall_f2_d ;
  CTf_t \lizzieLet60_4Lcall_f3_1sc_0_2_1q1a8H_1_1t1a8R_1_1t1'a8W_1_1q2a8I_1_1t2a8S_1_1t2'a8X_1_1Lcall_f2_bufchan_buf ;
  assign \lizzieLet60_4Lcall_f3_1sc_0_2_1q1a8H_1_1t1a8R_1_1t1'a8W_1_1q2a8I_1_1t2a8S_1_1t2'a8X_1_1Lcall_f2_bufchan_r  = (! \lizzieLet60_4Lcall_f3_1sc_0_2_1q1a8H_1_1t1a8R_1_1t1'a8W_1_1q2a8I_1_1t2a8S_1_1t2'a8X_1_1Lcall_f2_bufchan_buf [0]);
  assign lizzieLet61_1_argbuf_d = (\lizzieLet60_4Lcall_f3_1sc_0_2_1q1a8H_1_1t1a8R_1_1t1'a8W_1_1q2a8I_1_1t2a8S_1_1t2'a8X_1_1Lcall_f2_bufchan_buf [0] ? \lizzieLet60_4Lcall_f3_1sc_0_2_1q1a8H_1_1t1a8R_1_1t1'a8W_1_1q2a8I_1_1t2a8S_1_1t2'a8X_1_1Lcall_f2_bufchan_buf  :
                                   \lizzieLet60_4Lcall_f3_1sc_0_2_1q1a8H_1_1t1a8R_1_1t1'a8W_1_1q2a8I_1_1t2a8S_1_1t2'a8X_1_1Lcall_f2_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet60_4Lcall_f3_1sc_0_2_1q1a8H_1_1t1a8R_1_1t1'a8W_1_1q2a8I_1_1t2a8S_1_1t2'a8X_1_1Lcall_f2_bufchan_buf  <= {163'd0,
                                                                                                                        1'd0};
    else
      if ((lizzieLet61_1_argbuf_r && \lizzieLet60_4Lcall_f3_1sc_0_2_1q1a8H_1_1t1a8R_1_1t1'a8W_1_1q2a8I_1_1t2a8S_1_1t2'a8X_1_1Lcall_f2_bufchan_buf [0]))
        \lizzieLet60_4Lcall_f3_1sc_0_2_1q1a8H_1_1t1a8R_1_1t1'a8W_1_1q2a8I_1_1t2a8S_1_1t2'a8X_1_1Lcall_f2_bufchan_buf  <= {163'd0,
                                                                                                                          1'd0};
      else if (((! lizzieLet61_1_argbuf_r) && (! \lizzieLet60_4Lcall_f3_1sc_0_2_1q1a8H_1_1t1a8R_1_1t1'a8W_1_1q2a8I_1_1t2a8S_1_1t2'a8X_1_1Lcall_f2_bufchan_buf [0])))
        \lizzieLet60_4Lcall_f3_1sc_0_2_1q1a8H_1_1t1a8R_1_1t1'a8W_1_1q2a8I_1_1t2a8S_1_1t2'a8X_1_1Lcall_f2_bufchan_buf  <= \lizzieLet60_4Lcall_f3_1sc_0_2_1q1a8H_1_1t1a8R_1_1t1'a8W_1_1q2a8I_1_1t2a8S_1_1t2'a8X_1_1Lcall_f2_bufchan_d ;
  
  /* fork (Ty Pointer_QTree_Bool) : (lizzieLet60_4Lfsbos,Pointer_QTree_Bool) > [(lizzieLet60_4Lfsbos_1_merge_merge_merge_fork_1,Pointer_QTree_Bool),
                                                                           (lizzieLet60_4Lfsbos_1_merge_merge_merge_fork_2,Pointer_QTree_Bool)] */
  logic [1:0] lizzieLet60_4Lfsbos_emitted;
  logic [1:0] lizzieLet60_4Lfsbos_done;
  assign lizzieLet60_4Lfsbos_1_merge_merge_merge_fork_1_d = {lizzieLet60_4Lfsbos_d[16:1],
                                                             (lizzieLet60_4Lfsbos_d[0] && (! lizzieLet60_4Lfsbos_emitted[0]))};
  assign lizzieLet60_4Lfsbos_1_merge_merge_merge_fork_2_d = {lizzieLet60_4Lfsbos_d[16:1],
                                                             (lizzieLet60_4Lfsbos_d[0] && (! lizzieLet60_4Lfsbos_emitted[1]))};
  assign lizzieLet60_4Lfsbos_done = (lizzieLet60_4Lfsbos_emitted | ({lizzieLet60_4Lfsbos_1_merge_merge_merge_fork_2_d[0],
                                                                     lizzieLet60_4Lfsbos_1_merge_merge_merge_fork_1_d[0]} & {lizzieLet60_4Lfsbos_1_merge_merge_merge_fork_2_r,
                                                                                                                             lizzieLet60_4Lfsbos_1_merge_merge_merge_fork_1_r}));
  assign lizzieLet60_4Lfsbos_r = (& lizzieLet60_4Lfsbos_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet60_4Lfsbos_emitted <= 2'd0;
    else
      lizzieLet60_4Lfsbos_emitted <= (lizzieLet60_4Lfsbos_r ? 2'd0 :
                                      lizzieLet60_4Lfsbos_done);
  
  /* togo (Ty Pointer_QTree_Bool) : (lizzieLet60_4Lfsbos_1_merge_merge_merge_fork_1,Pointer_QTree_Bool) > (call_f_goConst,Go) */
  assign call_f_goConst_d = lizzieLet60_4Lfsbos_1_merge_merge_merge_fork_1_d[0];
  assign lizzieLet60_4Lfsbos_1_merge_merge_merge_fork_1_r = call_f_goConst_r;
  
  /* buf (Ty Pointer_QTree_Bool) : (lizzieLet60_4Lfsbos_1_merge_merge_merge_fork_2,Pointer_QTree_Bool) > (f_resbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t lizzieLet60_4Lfsbos_1_merge_merge_merge_fork_2_bufchan_d;
  logic lizzieLet60_4Lfsbos_1_merge_merge_merge_fork_2_bufchan_r;
  assign lizzieLet60_4Lfsbos_1_merge_merge_merge_fork_2_r = ((! lizzieLet60_4Lfsbos_1_merge_merge_merge_fork_2_bufchan_d[0]) || lizzieLet60_4Lfsbos_1_merge_merge_merge_fork_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet60_4Lfsbos_1_merge_merge_merge_fork_2_bufchan_d <= {16'd0,
                                                                   1'd0};
    else
      if (lizzieLet60_4Lfsbos_1_merge_merge_merge_fork_2_r)
        lizzieLet60_4Lfsbos_1_merge_merge_merge_fork_2_bufchan_d <= lizzieLet60_4Lfsbos_1_merge_merge_merge_fork_2_d;
  Pointer_QTree_Bool_t lizzieLet60_4Lfsbos_1_merge_merge_merge_fork_2_bufchan_buf;
  assign lizzieLet60_4Lfsbos_1_merge_merge_merge_fork_2_bufchan_r = (! lizzieLet60_4Lfsbos_1_merge_merge_merge_fork_2_bufchan_buf[0]);
  assign f_resbuf_d = (lizzieLet60_4Lfsbos_1_merge_merge_merge_fork_2_bufchan_buf[0] ? lizzieLet60_4Lfsbos_1_merge_merge_merge_fork_2_bufchan_buf :
                       lizzieLet60_4Lfsbos_1_merge_merge_merge_fork_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet60_4Lfsbos_1_merge_merge_merge_fork_2_bufchan_buf <= {16'd0,
                                                                     1'd0};
    else
      if ((f_resbuf_r && lizzieLet60_4Lfsbos_1_merge_merge_merge_fork_2_bufchan_buf[0]))
        lizzieLet60_4Lfsbos_1_merge_merge_merge_fork_2_bufchan_buf <= {16'd0,
                                                                       1'd0};
      else if (((! f_resbuf_r) && (! lizzieLet60_4Lfsbos_1_merge_merge_merge_fork_2_bufchan_buf[0])))
        lizzieLet60_4Lfsbos_1_merge_merge_merge_fork_2_bufchan_buf <= lizzieLet60_4Lfsbos_1_merge_merge_merge_fork_2_bufchan_d;
  
  /* destruct (Ty CTf'''''''''''',
          Dcon Lcall_f''''''''''''0) : (lizzieLet65_1Lcall_f''''''''''''0,CTf'''''''''''') > [(es_1_1_destruct,Pointer_QTree_Bool),
                                                                                              (es_2_2_destruct,Pointer_QTree_Bool),
                                                                                              (es_3_3_destruct,Pointer_QTree_Bool),
                                                                                              (sc_0_9_destruct,Pointer_CTf'''''''''''')] */
  logic [3:0] \lizzieLet65_1Lcall_f''''''''''''0_emitted ;
  logic [3:0] \lizzieLet65_1Lcall_f''''''''''''0_done ;
  assign es_1_1_destruct_d = {\lizzieLet65_1Lcall_f''''''''''''0_d [19:4],
                              (\lizzieLet65_1Lcall_f''''''''''''0_d [0] && (! \lizzieLet65_1Lcall_f''''''''''''0_emitted [0]))};
  assign es_2_2_destruct_d = {\lizzieLet65_1Lcall_f''''''''''''0_d [35:20],
                              (\lizzieLet65_1Lcall_f''''''''''''0_d [0] && (! \lizzieLet65_1Lcall_f''''''''''''0_emitted [1]))};
  assign es_3_3_destruct_d = {\lizzieLet65_1Lcall_f''''''''''''0_d [51:36],
                              (\lizzieLet65_1Lcall_f''''''''''''0_d [0] && (! \lizzieLet65_1Lcall_f''''''''''''0_emitted [2]))};
  assign sc_0_9_destruct_d = {\lizzieLet65_1Lcall_f''''''''''''0_d [67:52],
                              (\lizzieLet65_1Lcall_f''''''''''''0_d [0] && (! \lizzieLet65_1Lcall_f''''''''''''0_emitted [3]))};
  assign \lizzieLet65_1Lcall_f''''''''''''0_done  = (\lizzieLet65_1Lcall_f''''''''''''0_emitted  | ({sc_0_9_destruct_d[0],
                                                                                                     es_3_3_destruct_d[0],
                                                                                                     es_2_2_destruct_d[0],
                                                                                                     es_1_1_destruct_d[0]} & {sc_0_9_destruct_r,
                                                                                                                              es_3_3_destruct_r,
                                                                                                                              es_2_2_destruct_r,
                                                                                                                              es_1_1_destruct_r}));
  assign \lizzieLet65_1Lcall_f''''''''''''0_r  = (& \lizzieLet65_1Lcall_f''''''''''''0_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet65_1Lcall_f''''''''''''0_emitted  <= 4'd0;
    else
      \lizzieLet65_1Lcall_f''''''''''''0_emitted  <= (\lizzieLet65_1Lcall_f''''''''''''0_r  ? 4'd0 :
                                                      \lizzieLet65_1Lcall_f''''''''''''0_done );
  
  /* destruct (Ty CTf'''''''''''',
          Dcon Lcall_f''''''''''''1) : (lizzieLet65_1Lcall_f''''''''''''1,CTf'''''''''''') > [(es_2_1_destruct,Pointer_QTree_Bool),
                                                                                              (es_3_2_destruct,Pointer_QTree_Bool),
                                                                                              (sc_0_8_destruct,Pointer_CTf''''''''''''),
                                                                                              (q1a98_3_destruct,Pointer_QTree_Bool),
                                                                                              (t1a9d_3_destruct,Pointer_QTree_Bool)] */
  logic [4:0] \lizzieLet65_1Lcall_f''''''''''''1_emitted ;
  logic [4:0] \lizzieLet65_1Lcall_f''''''''''''1_done ;
  assign es_2_1_destruct_d = {\lizzieLet65_1Lcall_f''''''''''''1_d [19:4],
                              (\lizzieLet65_1Lcall_f''''''''''''1_d [0] && (! \lizzieLet65_1Lcall_f''''''''''''1_emitted [0]))};
  assign es_3_2_destruct_d = {\lizzieLet65_1Lcall_f''''''''''''1_d [35:20],
                              (\lizzieLet65_1Lcall_f''''''''''''1_d [0] && (! \lizzieLet65_1Lcall_f''''''''''''1_emitted [1]))};
  assign sc_0_8_destruct_d = {\lizzieLet65_1Lcall_f''''''''''''1_d [51:36],
                              (\lizzieLet65_1Lcall_f''''''''''''1_d [0] && (! \lizzieLet65_1Lcall_f''''''''''''1_emitted [2]))};
  assign q1a98_3_destruct_d = {\lizzieLet65_1Lcall_f''''''''''''1_d [67:52],
                               (\lizzieLet65_1Lcall_f''''''''''''1_d [0] && (! \lizzieLet65_1Lcall_f''''''''''''1_emitted [3]))};
  assign t1a9d_3_destruct_d = {\lizzieLet65_1Lcall_f''''''''''''1_d [83:68],
                               (\lizzieLet65_1Lcall_f''''''''''''1_d [0] && (! \lizzieLet65_1Lcall_f''''''''''''1_emitted [4]))};
  assign \lizzieLet65_1Lcall_f''''''''''''1_done  = (\lizzieLet65_1Lcall_f''''''''''''1_emitted  | ({t1a9d_3_destruct_d[0],
                                                                                                     q1a98_3_destruct_d[0],
                                                                                                     sc_0_8_destruct_d[0],
                                                                                                     es_3_2_destruct_d[0],
                                                                                                     es_2_1_destruct_d[0]} & {t1a9d_3_destruct_r,
                                                                                                                              q1a98_3_destruct_r,
                                                                                                                              sc_0_8_destruct_r,
                                                                                                                              es_3_2_destruct_r,
                                                                                                                              es_2_1_destruct_r}));
  assign \lizzieLet65_1Lcall_f''''''''''''1_r  = (& \lizzieLet65_1Lcall_f''''''''''''1_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet65_1Lcall_f''''''''''''1_emitted  <= 5'd0;
    else
      \lizzieLet65_1Lcall_f''''''''''''1_emitted  <= (\lizzieLet65_1Lcall_f''''''''''''1_r  ? 5'd0 :
                                                      \lizzieLet65_1Lcall_f''''''''''''1_done );
  
  /* destruct (Ty CTf'''''''''''',
          Dcon Lcall_f''''''''''''2) : (lizzieLet65_1Lcall_f''''''''''''2,CTf'''''''''''') > [(es_3_1_destruct,Pointer_QTree_Bool),
                                                                                              (sc_0_7_destruct,Pointer_CTf''''''''''''),
                                                                                              (q1a98_2_destruct,Pointer_QTree_Bool),
                                                                                              (t1a9d_2_destruct,Pointer_QTree_Bool),
                                                                                              (q2a99_2_destruct,Pointer_QTree_Bool),
                                                                                              (t2a9e_2_destruct,Pointer_QTree_Bool)] */
  logic [5:0] \lizzieLet65_1Lcall_f''''''''''''2_emitted ;
  logic [5:0] \lizzieLet65_1Lcall_f''''''''''''2_done ;
  assign es_3_1_destruct_d = {\lizzieLet65_1Lcall_f''''''''''''2_d [19:4],
                              (\lizzieLet65_1Lcall_f''''''''''''2_d [0] && (! \lizzieLet65_1Lcall_f''''''''''''2_emitted [0]))};
  assign sc_0_7_destruct_d = {\lizzieLet65_1Lcall_f''''''''''''2_d [35:20],
                              (\lizzieLet65_1Lcall_f''''''''''''2_d [0] && (! \lizzieLet65_1Lcall_f''''''''''''2_emitted [1]))};
  assign q1a98_2_destruct_d = {\lizzieLet65_1Lcall_f''''''''''''2_d [51:36],
                               (\lizzieLet65_1Lcall_f''''''''''''2_d [0] && (! \lizzieLet65_1Lcall_f''''''''''''2_emitted [2]))};
  assign t1a9d_2_destruct_d = {\lizzieLet65_1Lcall_f''''''''''''2_d [67:52],
                               (\lizzieLet65_1Lcall_f''''''''''''2_d [0] && (! \lizzieLet65_1Lcall_f''''''''''''2_emitted [3]))};
  assign q2a99_2_destruct_d = {\lizzieLet65_1Lcall_f''''''''''''2_d [83:68],
                               (\lizzieLet65_1Lcall_f''''''''''''2_d [0] && (! \lizzieLet65_1Lcall_f''''''''''''2_emitted [4]))};
  assign t2a9e_2_destruct_d = {\lizzieLet65_1Lcall_f''''''''''''2_d [99:84],
                               (\lizzieLet65_1Lcall_f''''''''''''2_d [0] && (! \lizzieLet65_1Lcall_f''''''''''''2_emitted [5]))};
  assign \lizzieLet65_1Lcall_f''''''''''''2_done  = (\lizzieLet65_1Lcall_f''''''''''''2_emitted  | ({t2a9e_2_destruct_d[0],
                                                                                                     q2a99_2_destruct_d[0],
                                                                                                     t1a9d_2_destruct_d[0],
                                                                                                     q1a98_2_destruct_d[0],
                                                                                                     sc_0_7_destruct_d[0],
                                                                                                     es_3_1_destruct_d[0]} & {t2a9e_2_destruct_r,
                                                                                                                              q2a99_2_destruct_r,
                                                                                                                              t1a9d_2_destruct_r,
                                                                                                                              q1a98_2_destruct_r,
                                                                                                                              sc_0_7_destruct_r,
                                                                                                                              es_3_1_destruct_r}));
  assign \lizzieLet65_1Lcall_f''''''''''''2_r  = (& \lizzieLet65_1Lcall_f''''''''''''2_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet65_1Lcall_f''''''''''''2_emitted  <= 6'd0;
    else
      \lizzieLet65_1Lcall_f''''''''''''2_emitted  <= (\lizzieLet65_1Lcall_f''''''''''''2_r  ? 6'd0 :
                                                      \lizzieLet65_1Lcall_f''''''''''''2_done );
  
  /* destruct (Ty CTf'''''''''''',
          Dcon Lcall_f''''''''''''3) : (lizzieLet65_1Lcall_f''''''''''''3,CTf'''''''''''') > [(sc_0_6_destruct,Pointer_CTf''''''''''''),
                                                                                              (q1a98_1_destruct,Pointer_QTree_Bool),
                                                                                              (t1a9d_1_destruct,Pointer_QTree_Bool),
                                                                                              (q2a99_1_destruct,Pointer_QTree_Bool),
                                                                                              (t2a9e_1_destruct,Pointer_QTree_Bool),
                                                                                              (q3a9a_1_destruct,Pointer_QTree_Bool),
                                                                                              (t3a9f_1_destruct,Pointer_QTree_Bool)] */
  logic [6:0] \lizzieLet65_1Lcall_f''''''''''''3_emitted ;
  logic [6:0] \lizzieLet65_1Lcall_f''''''''''''3_done ;
  assign sc_0_6_destruct_d = {\lizzieLet65_1Lcall_f''''''''''''3_d [19:4],
                              (\lizzieLet65_1Lcall_f''''''''''''3_d [0] && (! \lizzieLet65_1Lcall_f''''''''''''3_emitted [0]))};
  assign q1a98_1_destruct_d = {\lizzieLet65_1Lcall_f''''''''''''3_d [35:20],
                               (\lizzieLet65_1Lcall_f''''''''''''3_d [0] && (! \lizzieLet65_1Lcall_f''''''''''''3_emitted [1]))};
  assign t1a9d_1_destruct_d = {\lizzieLet65_1Lcall_f''''''''''''3_d [51:36],
                               (\lizzieLet65_1Lcall_f''''''''''''3_d [0] && (! \lizzieLet65_1Lcall_f''''''''''''3_emitted [2]))};
  assign q2a99_1_destruct_d = {\lizzieLet65_1Lcall_f''''''''''''3_d [67:52],
                               (\lizzieLet65_1Lcall_f''''''''''''3_d [0] && (! \lizzieLet65_1Lcall_f''''''''''''3_emitted [3]))};
  assign t2a9e_1_destruct_d = {\lizzieLet65_1Lcall_f''''''''''''3_d [83:68],
                               (\lizzieLet65_1Lcall_f''''''''''''3_d [0] && (! \lizzieLet65_1Lcall_f''''''''''''3_emitted [4]))};
  assign q3a9a_1_destruct_d = {\lizzieLet65_1Lcall_f''''''''''''3_d [99:84],
                               (\lizzieLet65_1Lcall_f''''''''''''3_d [0] && (! \lizzieLet65_1Lcall_f''''''''''''3_emitted [5]))};
  assign t3a9f_1_destruct_d = {\lizzieLet65_1Lcall_f''''''''''''3_d [115:100],
                               (\lizzieLet65_1Lcall_f''''''''''''3_d [0] && (! \lizzieLet65_1Lcall_f''''''''''''3_emitted [6]))};
  assign \lizzieLet65_1Lcall_f''''''''''''3_done  = (\lizzieLet65_1Lcall_f''''''''''''3_emitted  | ({t3a9f_1_destruct_d[0],
                                                                                                     q3a9a_1_destruct_d[0],
                                                                                                     t2a9e_1_destruct_d[0],
                                                                                                     q2a99_1_destruct_d[0],
                                                                                                     t1a9d_1_destruct_d[0],
                                                                                                     q1a98_1_destruct_d[0],
                                                                                                     sc_0_6_destruct_d[0]} & {t3a9f_1_destruct_r,
                                                                                                                              q3a9a_1_destruct_r,
                                                                                                                              t2a9e_1_destruct_r,
                                                                                                                              q2a99_1_destruct_r,
                                                                                                                              t1a9d_1_destruct_r,
                                                                                                                              q1a98_1_destruct_r,
                                                                                                                              sc_0_6_destruct_r}));
  assign \lizzieLet65_1Lcall_f''''''''''''3_r  = (& \lizzieLet65_1Lcall_f''''''''''''3_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet65_1Lcall_f''''''''''''3_emitted  <= 7'd0;
    else
      \lizzieLet65_1Lcall_f''''''''''''3_emitted  <= (\lizzieLet65_1Lcall_f''''''''''''3_r  ? 7'd0 :
                                                      \lizzieLet65_1Lcall_f''''''''''''3_done );
  
  /* demux (Ty CTf'''''''''''',
       Ty CTf'''''''''''') : (lizzieLet65_2,CTf'''''''''''') (lizzieLet65_1,CTf'''''''''''') > [(_1,CTf''''''''''''),
                                                                                                (lizzieLet65_1Lcall_f''''''''''''3,CTf''''''''''''),
                                                                                                (lizzieLet65_1Lcall_f''''''''''''2,CTf''''''''''''),
                                                                                                (lizzieLet65_1Lcall_f''''''''''''1,CTf''''''''''''),
                                                                                                (lizzieLet65_1Lcall_f''''''''''''0,CTf'''''''''''')] */
  logic [4:0] lizzieLet65_1_onehotd;
  always_comb
    if ((lizzieLet65_2_d[0] && lizzieLet65_1_d[0]))
      unique case (lizzieLet65_2_d[3:1])
        3'd0: lizzieLet65_1_onehotd = 5'd1;
        3'd1: lizzieLet65_1_onehotd = 5'd2;
        3'd2: lizzieLet65_1_onehotd = 5'd4;
        3'd3: lizzieLet65_1_onehotd = 5'd8;
        3'd4: lizzieLet65_1_onehotd = 5'd16;
        default: lizzieLet65_1_onehotd = 5'd0;
      endcase
    else lizzieLet65_1_onehotd = 5'd0;
  assign _1_d = {lizzieLet65_1_d[115:1], lizzieLet65_1_onehotd[0]};
  assign \lizzieLet65_1Lcall_f''''''''''''3_d  = {lizzieLet65_1_d[115:1],
                                                  lizzieLet65_1_onehotd[1]};
  assign \lizzieLet65_1Lcall_f''''''''''''2_d  = {lizzieLet65_1_d[115:1],
                                                  lizzieLet65_1_onehotd[2]};
  assign \lizzieLet65_1Lcall_f''''''''''''1_d  = {lizzieLet65_1_d[115:1],
                                                  lizzieLet65_1_onehotd[3]};
  assign \lizzieLet65_1Lcall_f''''''''''''0_d  = {lizzieLet65_1_d[115:1],
                                                  lizzieLet65_1_onehotd[4]};
  assign lizzieLet65_1_r = (| (lizzieLet65_1_onehotd & {\lizzieLet65_1Lcall_f''''''''''''0_r ,
                                                        \lizzieLet65_1Lcall_f''''''''''''1_r ,
                                                        \lizzieLet65_1Lcall_f''''''''''''2_r ,
                                                        \lizzieLet65_1Lcall_f''''''''''''3_r ,
                                                        _1_r}));
  assign lizzieLet65_2_r = lizzieLet65_1_r;
  
  /* demux (Ty CTf'''''''''''',
       Ty Go) : (lizzieLet65_3,CTf'''''''''''') (go_8_goMux_data,Go) > [(_0,Go),
                                                                        (lizzieLet65_3Lcall_f''''''''''''3,Go),
                                                                        (lizzieLet65_3Lcall_f''''''''''''2,Go),
                                                                        (lizzieLet65_3Lcall_f''''''''''''1,Go),
                                                                        (lizzieLet65_3Lcall_f''''''''''''0,Go)] */
  logic [4:0] go_8_goMux_data_onehotd;
  always_comb
    if ((lizzieLet65_3_d[0] && go_8_goMux_data_d[0]))
      unique case (lizzieLet65_3_d[3:1])
        3'd0: go_8_goMux_data_onehotd = 5'd1;
        3'd1: go_8_goMux_data_onehotd = 5'd2;
        3'd2: go_8_goMux_data_onehotd = 5'd4;
        3'd3: go_8_goMux_data_onehotd = 5'd8;
        3'd4: go_8_goMux_data_onehotd = 5'd16;
        default: go_8_goMux_data_onehotd = 5'd0;
      endcase
    else go_8_goMux_data_onehotd = 5'd0;
  assign _0_d = go_8_goMux_data_onehotd[0];
  assign \lizzieLet65_3Lcall_f''''''''''''3_d  = go_8_goMux_data_onehotd[1];
  assign \lizzieLet65_3Lcall_f''''''''''''2_d  = go_8_goMux_data_onehotd[2];
  assign \lizzieLet65_3Lcall_f''''''''''''1_d  = go_8_goMux_data_onehotd[3];
  assign \lizzieLet65_3Lcall_f''''''''''''0_d  = go_8_goMux_data_onehotd[4];
  assign go_8_goMux_data_r = (| (go_8_goMux_data_onehotd & {\lizzieLet65_3Lcall_f''''''''''''0_r ,
                                                            \lizzieLet65_3Lcall_f''''''''''''1_r ,
                                                            \lizzieLet65_3Lcall_f''''''''''''2_r ,
                                                            \lizzieLet65_3Lcall_f''''''''''''3_r ,
                                                            _0_r}));
  assign lizzieLet65_3_r = go_8_goMux_data_r;
  
  /* buf (Ty Go) : (lizzieLet65_3Lcall_f''''''''''''0,Go) > (lizzieLet65_3Lcall_f''''''''''''0_1_argbuf,Go) */
  Go_t \lizzieLet65_3Lcall_f''''''''''''0_bufchan_d ;
  logic \lizzieLet65_3Lcall_f''''''''''''0_bufchan_r ;
  assign \lizzieLet65_3Lcall_f''''''''''''0_r  = ((! \lizzieLet65_3Lcall_f''''''''''''0_bufchan_d [0]) || \lizzieLet65_3Lcall_f''''''''''''0_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet65_3Lcall_f''''''''''''0_bufchan_d  <= 1'd0;
    else
      if (\lizzieLet65_3Lcall_f''''''''''''0_r )
        \lizzieLet65_3Lcall_f''''''''''''0_bufchan_d  <= \lizzieLet65_3Lcall_f''''''''''''0_d ;
  Go_t \lizzieLet65_3Lcall_f''''''''''''0_bufchan_buf ;
  assign \lizzieLet65_3Lcall_f''''''''''''0_bufchan_r  = (! \lizzieLet65_3Lcall_f''''''''''''0_bufchan_buf [0]);
  assign \lizzieLet65_3Lcall_f''''''''''''0_1_argbuf_d  = (\lizzieLet65_3Lcall_f''''''''''''0_bufchan_buf [0] ? \lizzieLet65_3Lcall_f''''''''''''0_bufchan_buf  :
                                                           \lizzieLet65_3Lcall_f''''''''''''0_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet65_3Lcall_f''''''''''''0_bufchan_buf  <= 1'd0;
    else
      if ((\lizzieLet65_3Lcall_f''''''''''''0_1_argbuf_r  && \lizzieLet65_3Lcall_f''''''''''''0_bufchan_buf [0]))
        \lizzieLet65_3Lcall_f''''''''''''0_bufchan_buf  <= 1'd0;
      else if (((! \lizzieLet65_3Lcall_f''''''''''''0_1_argbuf_r ) && (! \lizzieLet65_3Lcall_f''''''''''''0_bufchan_buf [0])))
        \lizzieLet65_3Lcall_f''''''''''''0_bufchan_buf  <= \lizzieLet65_3Lcall_f''''''''''''0_bufchan_d ;
  
  /* buf (Ty Go) : (lizzieLet65_3Lcall_f''''''''''''1,Go) > (lizzieLet65_3Lcall_f''''''''''''1_1_argbuf,Go) */
  Go_t \lizzieLet65_3Lcall_f''''''''''''1_bufchan_d ;
  logic \lizzieLet65_3Lcall_f''''''''''''1_bufchan_r ;
  assign \lizzieLet65_3Lcall_f''''''''''''1_r  = ((! \lizzieLet65_3Lcall_f''''''''''''1_bufchan_d [0]) || \lizzieLet65_3Lcall_f''''''''''''1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet65_3Lcall_f''''''''''''1_bufchan_d  <= 1'd0;
    else
      if (\lizzieLet65_3Lcall_f''''''''''''1_r )
        \lizzieLet65_3Lcall_f''''''''''''1_bufchan_d  <= \lizzieLet65_3Lcall_f''''''''''''1_d ;
  Go_t \lizzieLet65_3Lcall_f''''''''''''1_bufchan_buf ;
  assign \lizzieLet65_3Lcall_f''''''''''''1_bufchan_r  = (! \lizzieLet65_3Lcall_f''''''''''''1_bufchan_buf [0]);
  assign \lizzieLet65_3Lcall_f''''''''''''1_1_argbuf_d  = (\lizzieLet65_3Lcall_f''''''''''''1_bufchan_buf [0] ? \lizzieLet65_3Lcall_f''''''''''''1_bufchan_buf  :
                                                           \lizzieLet65_3Lcall_f''''''''''''1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet65_3Lcall_f''''''''''''1_bufchan_buf  <= 1'd0;
    else
      if ((\lizzieLet65_3Lcall_f''''''''''''1_1_argbuf_r  && \lizzieLet65_3Lcall_f''''''''''''1_bufchan_buf [0]))
        \lizzieLet65_3Lcall_f''''''''''''1_bufchan_buf  <= 1'd0;
      else if (((! \lizzieLet65_3Lcall_f''''''''''''1_1_argbuf_r ) && (! \lizzieLet65_3Lcall_f''''''''''''1_bufchan_buf [0])))
        \lizzieLet65_3Lcall_f''''''''''''1_bufchan_buf  <= \lizzieLet65_3Lcall_f''''''''''''1_bufchan_d ;
  
  /* buf (Ty Go) : (lizzieLet65_3Lcall_f''''''''''''2,Go) > (lizzieLet65_3Lcall_f''''''''''''2_1_argbuf,Go) */
  Go_t \lizzieLet65_3Lcall_f''''''''''''2_bufchan_d ;
  logic \lizzieLet65_3Lcall_f''''''''''''2_bufchan_r ;
  assign \lizzieLet65_3Lcall_f''''''''''''2_r  = ((! \lizzieLet65_3Lcall_f''''''''''''2_bufchan_d [0]) || \lizzieLet65_3Lcall_f''''''''''''2_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet65_3Lcall_f''''''''''''2_bufchan_d  <= 1'd0;
    else
      if (\lizzieLet65_3Lcall_f''''''''''''2_r )
        \lizzieLet65_3Lcall_f''''''''''''2_bufchan_d  <= \lizzieLet65_3Lcall_f''''''''''''2_d ;
  Go_t \lizzieLet65_3Lcall_f''''''''''''2_bufchan_buf ;
  assign \lizzieLet65_3Lcall_f''''''''''''2_bufchan_r  = (! \lizzieLet65_3Lcall_f''''''''''''2_bufchan_buf [0]);
  assign \lizzieLet65_3Lcall_f''''''''''''2_1_argbuf_d  = (\lizzieLet65_3Lcall_f''''''''''''2_bufchan_buf [0] ? \lizzieLet65_3Lcall_f''''''''''''2_bufchan_buf  :
                                                           \lizzieLet65_3Lcall_f''''''''''''2_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet65_3Lcall_f''''''''''''2_bufchan_buf  <= 1'd0;
    else
      if ((\lizzieLet65_3Lcall_f''''''''''''2_1_argbuf_r  && \lizzieLet65_3Lcall_f''''''''''''2_bufchan_buf [0]))
        \lizzieLet65_3Lcall_f''''''''''''2_bufchan_buf  <= 1'd0;
      else if (((! \lizzieLet65_3Lcall_f''''''''''''2_1_argbuf_r ) && (! \lizzieLet65_3Lcall_f''''''''''''2_bufchan_buf [0])))
        \lizzieLet65_3Lcall_f''''''''''''2_bufchan_buf  <= \lizzieLet65_3Lcall_f''''''''''''2_bufchan_d ;
  
  /* buf (Ty Go) : (lizzieLet65_3Lcall_f''''''''''''3,Go) > (lizzieLet65_3Lcall_f''''''''''''3_1_argbuf,Go) */
  Go_t \lizzieLet65_3Lcall_f''''''''''''3_bufchan_d ;
  logic \lizzieLet65_3Lcall_f''''''''''''3_bufchan_r ;
  assign \lizzieLet65_3Lcall_f''''''''''''3_r  = ((! \lizzieLet65_3Lcall_f''''''''''''3_bufchan_d [0]) || \lizzieLet65_3Lcall_f''''''''''''3_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet65_3Lcall_f''''''''''''3_bufchan_d  <= 1'd0;
    else
      if (\lizzieLet65_3Lcall_f''''''''''''3_r )
        \lizzieLet65_3Lcall_f''''''''''''3_bufchan_d  <= \lizzieLet65_3Lcall_f''''''''''''3_d ;
  Go_t \lizzieLet65_3Lcall_f''''''''''''3_bufchan_buf ;
  assign \lizzieLet65_3Lcall_f''''''''''''3_bufchan_r  = (! \lizzieLet65_3Lcall_f''''''''''''3_bufchan_buf [0]);
  assign \lizzieLet65_3Lcall_f''''''''''''3_1_argbuf_d  = (\lizzieLet65_3Lcall_f''''''''''''3_bufchan_buf [0] ? \lizzieLet65_3Lcall_f''''''''''''3_bufchan_buf  :
                                                           \lizzieLet65_3Lcall_f''''''''''''3_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet65_3Lcall_f''''''''''''3_bufchan_buf  <= 1'd0;
    else
      if ((\lizzieLet65_3Lcall_f''''''''''''3_1_argbuf_r  && \lizzieLet65_3Lcall_f''''''''''''3_bufchan_buf [0]))
        \lizzieLet65_3Lcall_f''''''''''''3_bufchan_buf  <= 1'd0;
      else if (((! \lizzieLet65_3Lcall_f''''''''''''3_1_argbuf_r ) && (! \lizzieLet65_3Lcall_f''''''''''''3_bufchan_buf [0])))
        \lizzieLet65_3Lcall_f''''''''''''3_bufchan_buf  <= \lizzieLet65_3Lcall_f''''''''''''3_bufchan_d ;
  
  /* demux (Ty CTf'''''''''''',
       Ty Pointer_QTree_Bool) : (lizzieLet65_4,CTf'''''''''''') (srtarg_0_1_goMux_mux,Pointer_QTree_Bool) > [(lizzieLet65_4Lf''''''''''''sbos,Pointer_QTree_Bool),
                                                                                                             (lizzieLet65_4Lcall_f''''''''''''3,Pointer_QTree_Bool),
                                                                                                             (lizzieLet65_4Lcall_f''''''''''''2,Pointer_QTree_Bool),
                                                                                                             (lizzieLet65_4Lcall_f''''''''''''1,Pointer_QTree_Bool),
                                                                                                             (lizzieLet65_4Lcall_f''''''''''''0,Pointer_QTree_Bool)] */
  logic [4:0] srtarg_0_1_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet65_4_d[0] && srtarg_0_1_goMux_mux_d[0]))
      unique case (lizzieLet65_4_d[3:1])
        3'd0: srtarg_0_1_goMux_mux_onehotd = 5'd1;
        3'd1: srtarg_0_1_goMux_mux_onehotd = 5'd2;
        3'd2: srtarg_0_1_goMux_mux_onehotd = 5'd4;
        3'd3: srtarg_0_1_goMux_mux_onehotd = 5'd8;
        3'd4: srtarg_0_1_goMux_mux_onehotd = 5'd16;
        default: srtarg_0_1_goMux_mux_onehotd = 5'd0;
      endcase
    else srtarg_0_1_goMux_mux_onehotd = 5'd0;
  assign \lizzieLet65_4Lf''''''''''''sbos_d  = {srtarg_0_1_goMux_mux_d[16:1],
                                                srtarg_0_1_goMux_mux_onehotd[0]};
  assign \lizzieLet65_4Lcall_f''''''''''''3_d  = {srtarg_0_1_goMux_mux_d[16:1],
                                                  srtarg_0_1_goMux_mux_onehotd[1]};
  assign \lizzieLet65_4Lcall_f''''''''''''2_d  = {srtarg_0_1_goMux_mux_d[16:1],
                                                  srtarg_0_1_goMux_mux_onehotd[2]};
  assign \lizzieLet65_4Lcall_f''''''''''''1_d  = {srtarg_0_1_goMux_mux_d[16:1],
                                                  srtarg_0_1_goMux_mux_onehotd[3]};
  assign \lizzieLet65_4Lcall_f''''''''''''0_d  = {srtarg_0_1_goMux_mux_d[16:1],
                                                  srtarg_0_1_goMux_mux_onehotd[4]};
  assign srtarg_0_1_goMux_mux_r = (| (srtarg_0_1_goMux_mux_onehotd & {\lizzieLet65_4Lcall_f''''''''''''0_r ,
                                                                      \lizzieLet65_4Lcall_f''''''''''''1_r ,
                                                                      \lizzieLet65_4Lcall_f''''''''''''2_r ,
                                                                      \lizzieLet65_4Lcall_f''''''''''''3_r ,
                                                                      \lizzieLet65_4Lf''''''''''''sbos_r }));
  assign lizzieLet65_4_r = srtarg_0_1_goMux_mux_r;
  
  /* dcon (Ty QTree_Bool,
      Dcon QNode_Bool) : [(lizzieLet65_4Lcall_f''''''''''''0,Pointer_QTree_Bool),
                          (es_1_1_destruct,Pointer_QTree_Bool),
                          (es_2_2_destruct,Pointer_QTree_Bool),
                          (es_3_3_destruct,Pointer_QTree_Bool)] > (lizzieLet65_4Lcall_f''''''''''''0_1es_1_1_1es_2_2_1es_3_3_1QNode_Bool,QTree_Bool) */
  assign \lizzieLet65_4Lcall_f''''''''''''0_1es_1_1_1es_2_2_1es_3_3_1QNode_Bool_d  = QNode_Bool_dc((& {\lizzieLet65_4Lcall_f''''''''''''0_d [0],
                                                                                                       es_1_1_destruct_d[0],
                                                                                                       es_2_2_destruct_d[0],
                                                                                                       es_3_3_destruct_d[0]}), \lizzieLet65_4Lcall_f''''''''''''0_d , es_1_1_destruct_d, es_2_2_destruct_d, es_3_3_destruct_d);
  assign {\lizzieLet65_4Lcall_f''''''''''''0_r ,
          es_1_1_destruct_r,
          es_2_2_destruct_r,
          es_3_3_destruct_r} = {4 {(\lizzieLet65_4Lcall_f''''''''''''0_1es_1_1_1es_2_2_1es_3_3_1QNode_Bool_r  && \lizzieLet65_4Lcall_f''''''''''''0_1es_1_1_1es_2_2_1es_3_3_1QNode_Bool_d [0])}};
  
  /* buf (Ty QTree_Bool) : (lizzieLet65_4Lcall_f''''''''''''0_1es_1_1_1es_2_2_1es_3_3_1QNode_Bool,QTree_Bool) > (lizzieLet69_1_argbuf,QTree_Bool) */
  QTree_Bool_t \lizzieLet65_4Lcall_f''''''''''''0_1es_1_1_1es_2_2_1es_3_3_1QNode_Bool_bufchan_d ;
  logic \lizzieLet65_4Lcall_f''''''''''''0_1es_1_1_1es_2_2_1es_3_3_1QNode_Bool_bufchan_r ;
  assign \lizzieLet65_4Lcall_f''''''''''''0_1es_1_1_1es_2_2_1es_3_3_1QNode_Bool_r  = ((! \lizzieLet65_4Lcall_f''''''''''''0_1es_1_1_1es_2_2_1es_3_3_1QNode_Bool_bufchan_d [0]) || \lizzieLet65_4Lcall_f''''''''''''0_1es_1_1_1es_2_2_1es_3_3_1QNode_Bool_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet65_4Lcall_f''''''''''''0_1es_1_1_1es_2_2_1es_3_3_1QNode_Bool_bufchan_d  <= {66'd0,
                                                                                            1'd0};
    else
      if (\lizzieLet65_4Lcall_f''''''''''''0_1es_1_1_1es_2_2_1es_3_3_1QNode_Bool_r )
        \lizzieLet65_4Lcall_f''''''''''''0_1es_1_1_1es_2_2_1es_3_3_1QNode_Bool_bufchan_d  <= \lizzieLet65_4Lcall_f''''''''''''0_1es_1_1_1es_2_2_1es_3_3_1QNode_Bool_d ;
  QTree_Bool_t \lizzieLet65_4Lcall_f''''''''''''0_1es_1_1_1es_2_2_1es_3_3_1QNode_Bool_bufchan_buf ;
  assign \lizzieLet65_4Lcall_f''''''''''''0_1es_1_1_1es_2_2_1es_3_3_1QNode_Bool_bufchan_r  = (! \lizzieLet65_4Lcall_f''''''''''''0_1es_1_1_1es_2_2_1es_3_3_1QNode_Bool_bufchan_buf [0]);
  assign lizzieLet69_1_argbuf_d = (\lizzieLet65_4Lcall_f''''''''''''0_1es_1_1_1es_2_2_1es_3_3_1QNode_Bool_bufchan_buf [0] ? \lizzieLet65_4Lcall_f''''''''''''0_1es_1_1_1es_2_2_1es_3_3_1QNode_Bool_bufchan_buf  :
                                   \lizzieLet65_4Lcall_f''''''''''''0_1es_1_1_1es_2_2_1es_3_3_1QNode_Bool_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet65_4Lcall_f''''''''''''0_1es_1_1_1es_2_2_1es_3_3_1QNode_Bool_bufchan_buf  <= {66'd0,
                                                                                              1'd0};
    else
      if ((lizzieLet69_1_argbuf_r && \lizzieLet65_4Lcall_f''''''''''''0_1es_1_1_1es_2_2_1es_3_3_1QNode_Bool_bufchan_buf [0]))
        \lizzieLet65_4Lcall_f''''''''''''0_1es_1_1_1es_2_2_1es_3_3_1QNode_Bool_bufchan_buf  <= {66'd0,
                                                                                                1'd0};
      else if (((! lizzieLet69_1_argbuf_r) && (! \lizzieLet65_4Lcall_f''''''''''''0_1es_1_1_1es_2_2_1es_3_3_1QNode_Bool_bufchan_buf [0])))
        \lizzieLet65_4Lcall_f''''''''''''0_1es_1_1_1es_2_2_1es_3_3_1QNode_Bool_bufchan_buf  <= \lizzieLet65_4Lcall_f''''''''''''0_1es_1_1_1es_2_2_1es_3_3_1QNode_Bool_bufchan_d ;
  
  /* dcon (Ty CTf'''''''''''',
      Dcon Lcall_f''''''''''''0) : [(lizzieLet65_4Lcall_f''''''''''''1,Pointer_QTree_Bool),
                                    (es_2_1_destruct,Pointer_QTree_Bool),
                                    (es_3_2_destruct,Pointer_QTree_Bool),
                                    (sc_0_8_destruct,Pointer_CTf'''''''''''')] > (lizzieLet65_4Lcall_f''''''''''''1_1es_2_1_1es_3_2_1sc_0_8_1Lcall_f''''''''''''0,CTf'''''''''''') */
  assign \lizzieLet65_4Lcall_f''''''''''''1_1es_2_1_1es_3_2_1sc_0_8_1Lcall_f''''''''''''0_d  = \Lcall_f''''''''''''0_dc ((& {\lizzieLet65_4Lcall_f''''''''''''1_d [0],
                                                                                                                             es_2_1_destruct_d[0],
                                                                                                                             es_3_2_destruct_d[0],
                                                                                                                             sc_0_8_destruct_d[0]}), \lizzieLet65_4Lcall_f''''''''''''1_d , es_2_1_destruct_d, es_3_2_destruct_d, sc_0_8_destruct_d);
  assign {\lizzieLet65_4Lcall_f''''''''''''1_r ,
          es_2_1_destruct_r,
          es_3_2_destruct_r,
          sc_0_8_destruct_r} = {4 {(\lizzieLet65_4Lcall_f''''''''''''1_1es_2_1_1es_3_2_1sc_0_8_1Lcall_f''''''''''''0_r  && \lizzieLet65_4Lcall_f''''''''''''1_1es_2_1_1es_3_2_1sc_0_8_1Lcall_f''''''''''''0_d [0])}};
  
  /* buf (Ty CTf'''''''''''') : (lizzieLet65_4Lcall_f''''''''''''1_1es_2_1_1es_3_2_1sc_0_8_1Lcall_f''''''''''''0,CTf'''''''''''') > (lizzieLet68_1_argbuf,CTf'''''''''''') */
  \CTf''''''''''''_t  \lizzieLet65_4Lcall_f''''''''''''1_1es_2_1_1es_3_2_1sc_0_8_1Lcall_f''''''''''''0_bufchan_d ;
  logic \lizzieLet65_4Lcall_f''''''''''''1_1es_2_1_1es_3_2_1sc_0_8_1Lcall_f''''''''''''0_bufchan_r ;
  assign \lizzieLet65_4Lcall_f''''''''''''1_1es_2_1_1es_3_2_1sc_0_8_1Lcall_f''''''''''''0_r  = ((! \lizzieLet65_4Lcall_f''''''''''''1_1es_2_1_1es_3_2_1sc_0_8_1Lcall_f''''''''''''0_bufchan_d [0]) || \lizzieLet65_4Lcall_f''''''''''''1_1es_2_1_1es_3_2_1sc_0_8_1Lcall_f''''''''''''0_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet65_4Lcall_f''''''''''''1_1es_2_1_1es_3_2_1sc_0_8_1Lcall_f''''''''''''0_bufchan_d  <= {115'd0,
                                                                                                      1'd0};
    else
      if (\lizzieLet65_4Lcall_f''''''''''''1_1es_2_1_1es_3_2_1sc_0_8_1Lcall_f''''''''''''0_r )
        \lizzieLet65_4Lcall_f''''''''''''1_1es_2_1_1es_3_2_1sc_0_8_1Lcall_f''''''''''''0_bufchan_d  <= \lizzieLet65_4Lcall_f''''''''''''1_1es_2_1_1es_3_2_1sc_0_8_1Lcall_f''''''''''''0_d ;
  \CTf''''''''''''_t  \lizzieLet65_4Lcall_f''''''''''''1_1es_2_1_1es_3_2_1sc_0_8_1Lcall_f''''''''''''0_bufchan_buf ;
  assign \lizzieLet65_4Lcall_f''''''''''''1_1es_2_1_1es_3_2_1sc_0_8_1Lcall_f''''''''''''0_bufchan_r  = (! \lizzieLet65_4Lcall_f''''''''''''1_1es_2_1_1es_3_2_1sc_0_8_1Lcall_f''''''''''''0_bufchan_buf [0]);
  assign lizzieLet68_1_argbuf_d = (\lizzieLet65_4Lcall_f''''''''''''1_1es_2_1_1es_3_2_1sc_0_8_1Lcall_f''''''''''''0_bufchan_buf [0] ? \lizzieLet65_4Lcall_f''''''''''''1_1es_2_1_1es_3_2_1sc_0_8_1Lcall_f''''''''''''0_bufchan_buf  :
                                   \lizzieLet65_4Lcall_f''''''''''''1_1es_2_1_1es_3_2_1sc_0_8_1Lcall_f''''''''''''0_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet65_4Lcall_f''''''''''''1_1es_2_1_1es_3_2_1sc_0_8_1Lcall_f''''''''''''0_bufchan_buf  <= {115'd0,
                                                                                                        1'd0};
    else
      if ((lizzieLet68_1_argbuf_r && \lizzieLet65_4Lcall_f''''''''''''1_1es_2_1_1es_3_2_1sc_0_8_1Lcall_f''''''''''''0_bufchan_buf [0]))
        \lizzieLet65_4Lcall_f''''''''''''1_1es_2_1_1es_3_2_1sc_0_8_1Lcall_f''''''''''''0_bufchan_buf  <= {115'd0,
                                                                                                          1'd0};
      else if (((! lizzieLet68_1_argbuf_r) && (! \lizzieLet65_4Lcall_f''''''''''''1_1es_2_1_1es_3_2_1sc_0_8_1Lcall_f''''''''''''0_bufchan_buf [0])))
        \lizzieLet65_4Lcall_f''''''''''''1_1es_2_1_1es_3_2_1sc_0_8_1Lcall_f''''''''''''0_bufchan_buf  <= \lizzieLet65_4Lcall_f''''''''''''1_1es_2_1_1es_3_2_1sc_0_8_1Lcall_f''''''''''''0_bufchan_d ;
  
  /* dcon (Ty CTf'''''''''''',
      Dcon Lcall_f''''''''''''1) : [(lizzieLet65_4Lcall_f''''''''''''2,Pointer_QTree_Bool),
                                    (es_3_1_destruct,Pointer_QTree_Bool),
                                    (sc_0_7_destruct,Pointer_CTf''''''''''''),
                                    (q1a98_2_destruct,Pointer_QTree_Bool),
                                    (t1a9d_2_destruct,Pointer_QTree_Bool)] > (lizzieLet65_4Lcall_f''''''''''''2_1es_3_1_1sc_0_7_1q1a98_2_1t1a9d_2_1Lcall_f''''''''''''1,CTf'''''''''''') */
  assign \lizzieLet65_4Lcall_f''''''''''''2_1es_3_1_1sc_0_7_1q1a98_2_1t1a9d_2_1Lcall_f''''''''''''1_d  = \Lcall_f''''''''''''1_dc ((& {\lizzieLet65_4Lcall_f''''''''''''2_d [0],
                                                                                                                                       es_3_1_destruct_d[0],
                                                                                                                                       sc_0_7_destruct_d[0],
                                                                                                                                       q1a98_2_destruct_d[0],
                                                                                                                                       t1a9d_2_destruct_d[0]}), \lizzieLet65_4Lcall_f''''''''''''2_d , es_3_1_destruct_d, sc_0_7_destruct_d, q1a98_2_destruct_d, t1a9d_2_destruct_d);
  assign {\lizzieLet65_4Lcall_f''''''''''''2_r ,
          es_3_1_destruct_r,
          sc_0_7_destruct_r,
          q1a98_2_destruct_r,
          t1a9d_2_destruct_r} = {5 {(\lizzieLet65_4Lcall_f''''''''''''2_1es_3_1_1sc_0_7_1q1a98_2_1t1a9d_2_1Lcall_f''''''''''''1_r  && \lizzieLet65_4Lcall_f''''''''''''2_1es_3_1_1sc_0_7_1q1a98_2_1t1a9d_2_1Lcall_f''''''''''''1_d [0])}};
  
  /* buf (Ty CTf'''''''''''') : (lizzieLet65_4Lcall_f''''''''''''2_1es_3_1_1sc_0_7_1q1a98_2_1t1a9d_2_1Lcall_f''''''''''''1,CTf'''''''''''') > (lizzieLet67_1_argbuf,CTf'''''''''''') */
  \CTf''''''''''''_t  \lizzieLet65_4Lcall_f''''''''''''2_1es_3_1_1sc_0_7_1q1a98_2_1t1a9d_2_1Lcall_f''''''''''''1_bufchan_d ;
  logic \lizzieLet65_4Lcall_f''''''''''''2_1es_3_1_1sc_0_7_1q1a98_2_1t1a9d_2_1Lcall_f''''''''''''1_bufchan_r ;
  assign \lizzieLet65_4Lcall_f''''''''''''2_1es_3_1_1sc_0_7_1q1a98_2_1t1a9d_2_1Lcall_f''''''''''''1_r  = ((! \lizzieLet65_4Lcall_f''''''''''''2_1es_3_1_1sc_0_7_1q1a98_2_1t1a9d_2_1Lcall_f''''''''''''1_bufchan_d [0]) || \lizzieLet65_4Lcall_f''''''''''''2_1es_3_1_1sc_0_7_1q1a98_2_1t1a9d_2_1Lcall_f''''''''''''1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet65_4Lcall_f''''''''''''2_1es_3_1_1sc_0_7_1q1a98_2_1t1a9d_2_1Lcall_f''''''''''''1_bufchan_d  <= {115'd0,
                                                                                                                1'd0};
    else
      if (\lizzieLet65_4Lcall_f''''''''''''2_1es_3_1_1sc_0_7_1q1a98_2_1t1a9d_2_1Lcall_f''''''''''''1_r )
        \lizzieLet65_4Lcall_f''''''''''''2_1es_3_1_1sc_0_7_1q1a98_2_1t1a9d_2_1Lcall_f''''''''''''1_bufchan_d  <= \lizzieLet65_4Lcall_f''''''''''''2_1es_3_1_1sc_0_7_1q1a98_2_1t1a9d_2_1Lcall_f''''''''''''1_d ;
  \CTf''''''''''''_t  \lizzieLet65_4Lcall_f''''''''''''2_1es_3_1_1sc_0_7_1q1a98_2_1t1a9d_2_1Lcall_f''''''''''''1_bufchan_buf ;
  assign \lizzieLet65_4Lcall_f''''''''''''2_1es_3_1_1sc_0_7_1q1a98_2_1t1a9d_2_1Lcall_f''''''''''''1_bufchan_r  = (! \lizzieLet65_4Lcall_f''''''''''''2_1es_3_1_1sc_0_7_1q1a98_2_1t1a9d_2_1Lcall_f''''''''''''1_bufchan_buf [0]);
  assign lizzieLet67_1_argbuf_d = (\lizzieLet65_4Lcall_f''''''''''''2_1es_3_1_1sc_0_7_1q1a98_2_1t1a9d_2_1Lcall_f''''''''''''1_bufchan_buf [0] ? \lizzieLet65_4Lcall_f''''''''''''2_1es_3_1_1sc_0_7_1q1a98_2_1t1a9d_2_1Lcall_f''''''''''''1_bufchan_buf  :
                                   \lizzieLet65_4Lcall_f''''''''''''2_1es_3_1_1sc_0_7_1q1a98_2_1t1a9d_2_1Lcall_f''''''''''''1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet65_4Lcall_f''''''''''''2_1es_3_1_1sc_0_7_1q1a98_2_1t1a9d_2_1Lcall_f''''''''''''1_bufchan_buf  <= {115'd0,
                                                                                                                  1'd0};
    else
      if ((lizzieLet67_1_argbuf_r && \lizzieLet65_4Lcall_f''''''''''''2_1es_3_1_1sc_0_7_1q1a98_2_1t1a9d_2_1Lcall_f''''''''''''1_bufchan_buf [0]))
        \lizzieLet65_4Lcall_f''''''''''''2_1es_3_1_1sc_0_7_1q1a98_2_1t1a9d_2_1Lcall_f''''''''''''1_bufchan_buf  <= {115'd0,
                                                                                                                    1'd0};
      else if (((! lizzieLet67_1_argbuf_r) && (! \lizzieLet65_4Lcall_f''''''''''''2_1es_3_1_1sc_0_7_1q1a98_2_1t1a9d_2_1Lcall_f''''''''''''1_bufchan_buf [0])))
        \lizzieLet65_4Lcall_f''''''''''''2_1es_3_1_1sc_0_7_1q1a98_2_1t1a9d_2_1Lcall_f''''''''''''1_bufchan_buf  <= \lizzieLet65_4Lcall_f''''''''''''2_1es_3_1_1sc_0_7_1q1a98_2_1t1a9d_2_1Lcall_f''''''''''''1_bufchan_d ;
  
  /* dcon (Ty CTf'''''''''''',
      Dcon Lcall_f''''''''''''2) : [(lizzieLet65_4Lcall_f''''''''''''3,Pointer_QTree_Bool),
                                    (sc_0_6_destruct,Pointer_CTf''''''''''''),
                                    (q1a98_1_destruct,Pointer_QTree_Bool),
                                    (t1a9d_1_destruct,Pointer_QTree_Bool),
                                    (q2a99_1_destruct,Pointer_QTree_Bool),
                                    (t2a9e_1_destruct,Pointer_QTree_Bool)] > (lizzieLet65_4Lcall_f''''''''''''3_1sc_0_6_1q1a98_1_1t1a9d_1_1q2a99_1_1t2a9e_1_1Lcall_f''''''''''''2,CTf'''''''''''') */
  assign \lizzieLet65_4Lcall_f''''''''''''3_1sc_0_6_1q1a98_1_1t1a9d_1_1q2a99_1_1t2a9e_1_1Lcall_f''''''''''''2_d  = \Lcall_f''''''''''''2_dc ((& {\lizzieLet65_4Lcall_f''''''''''''3_d [0],
                                                                                                                                                 sc_0_6_destruct_d[0],
                                                                                                                                                 q1a98_1_destruct_d[0],
                                                                                                                                                 t1a9d_1_destruct_d[0],
                                                                                                                                                 q2a99_1_destruct_d[0],
                                                                                                                                                 t2a9e_1_destruct_d[0]}), \lizzieLet65_4Lcall_f''''''''''''3_d , sc_0_6_destruct_d, q1a98_1_destruct_d, t1a9d_1_destruct_d, q2a99_1_destruct_d, t2a9e_1_destruct_d);
  assign {\lizzieLet65_4Lcall_f''''''''''''3_r ,
          sc_0_6_destruct_r,
          q1a98_1_destruct_r,
          t1a9d_1_destruct_r,
          q2a99_1_destruct_r,
          t2a9e_1_destruct_r} = {6 {(\lizzieLet65_4Lcall_f''''''''''''3_1sc_0_6_1q1a98_1_1t1a9d_1_1q2a99_1_1t2a9e_1_1Lcall_f''''''''''''2_r  && \lizzieLet65_4Lcall_f''''''''''''3_1sc_0_6_1q1a98_1_1t1a9d_1_1q2a99_1_1t2a9e_1_1Lcall_f''''''''''''2_d [0])}};
  
  /* buf (Ty CTf'''''''''''') : (lizzieLet65_4Lcall_f''''''''''''3_1sc_0_6_1q1a98_1_1t1a9d_1_1q2a99_1_1t2a9e_1_1Lcall_f''''''''''''2,CTf'''''''''''') > (lizzieLet66_1_argbuf,CTf'''''''''''') */
  \CTf''''''''''''_t  \lizzieLet65_4Lcall_f''''''''''''3_1sc_0_6_1q1a98_1_1t1a9d_1_1q2a99_1_1t2a9e_1_1Lcall_f''''''''''''2_bufchan_d ;
  logic \lizzieLet65_4Lcall_f''''''''''''3_1sc_0_6_1q1a98_1_1t1a9d_1_1q2a99_1_1t2a9e_1_1Lcall_f''''''''''''2_bufchan_r ;
  assign \lizzieLet65_4Lcall_f''''''''''''3_1sc_0_6_1q1a98_1_1t1a9d_1_1q2a99_1_1t2a9e_1_1Lcall_f''''''''''''2_r  = ((! \lizzieLet65_4Lcall_f''''''''''''3_1sc_0_6_1q1a98_1_1t1a9d_1_1q2a99_1_1t2a9e_1_1Lcall_f''''''''''''2_bufchan_d [0]) || \lizzieLet65_4Lcall_f''''''''''''3_1sc_0_6_1q1a98_1_1t1a9d_1_1q2a99_1_1t2a9e_1_1Lcall_f''''''''''''2_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet65_4Lcall_f''''''''''''3_1sc_0_6_1q1a98_1_1t1a9d_1_1q2a99_1_1t2a9e_1_1Lcall_f''''''''''''2_bufchan_d  <= {115'd0,
                                                                                                                          1'd0};
    else
      if (\lizzieLet65_4Lcall_f''''''''''''3_1sc_0_6_1q1a98_1_1t1a9d_1_1q2a99_1_1t2a9e_1_1Lcall_f''''''''''''2_r )
        \lizzieLet65_4Lcall_f''''''''''''3_1sc_0_6_1q1a98_1_1t1a9d_1_1q2a99_1_1t2a9e_1_1Lcall_f''''''''''''2_bufchan_d  <= \lizzieLet65_4Lcall_f''''''''''''3_1sc_0_6_1q1a98_1_1t1a9d_1_1q2a99_1_1t2a9e_1_1Lcall_f''''''''''''2_d ;
  \CTf''''''''''''_t  \lizzieLet65_4Lcall_f''''''''''''3_1sc_0_6_1q1a98_1_1t1a9d_1_1q2a99_1_1t2a9e_1_1Lcall_f''''''''''''2_bufchan_buf ;
  assign \lizzieLet65_4Lcall_f''''''''''''3_1sc_0_6_1q1a98_1_1t1a9d_1_1q2a99_1_1t2a9e_1_1Lcall_f''''''''''''2_bufchan_r  = (! \lizzieLet65_4Lcall_f''''''''''''3_1sc_0_6_1q1a98_1_1t1a9d_1_1q2a99_1_1t2a9e_1_1Lcall_f''''''''''''2_bufchan_buf [0]);
  assign lizzieLet66_1_argbuf_d = (\lizzieLet65_4Lcall_f''''''''''''3_1sc_0_6_1q1a98_1_1t1a9d_1_1q2a99_1_1t2a9e_1_1Lcall_f''''''''''''2_bufchan_buf [0] ? \lizzieLet65_4Lcall_f''''''''''''3_1sc_0_6_1q1a98_1_1t1a9d_1_1q2a99_1_1t2a9e_1_1Lcall_f''''''''''''2_bufchan_buf  :
                                   \lizzieLet65_4Lcall_f''''''''''''3_1sc_0_6_1q1a98_1_1t1a9d_1_1q2a99_1_1t2a9e_1_1Lcall_f''''''''''''2_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet65_4Lcall_f''''''''''''3_1sc_0_6_1q1a98_1_1t1a9d_1_1q2a99_1_1t2a9e_1_1Lcall_f''''''''''''2_bufchan_buf  <= {115'd0,
                                                                                                                            1'd0};
    else
      if ((lizzieLet66_1_argbuf_r && \lizzieLet65_4Lcall_f''''''''''''3_1sc_0_6_1q1a98_1_1t1a9d_1_1q2a99_1_1t2a9e_1_1Lcall_f''''''''''''2_bufchan_buf [0]))
        \lizzieLet65_4Lcall_f''''''''''''3_1sc_0_6_1q1a98_1_1t1a9d_1_1q2a99_1_1t2a9e_1_1Lcall_f''''''''''''2_bufchan_buf  <= {115'd0,
                                                                                                                              1'd0};
      else if (((! lizzieLet66_1_argbuf_r) && (! \lizzieLet65_4Lcall_f''''''''''''3_1sc_0_6_1q1a98_1_1t1a9d_1_1q2a99_1_1t2a9e_1_1Lcall_f''''''''''''2_bufchan_buf [0])))
        \lizzieLet65_4Lcall_f''''''''''''3_1sc_0_6_1q1a98_1_1t1a9d_1_1q2a99_1_1t2a9e_1_1Lcall_f''''''''''''2_bufchan_buf  <= \lizzieLet65_4Lcall_f''''''''''''3_1sc_0_6_1q1a98_1_1t1a9d_1_1q2a99_1_1t2a9e_1_1Lcall_f''''''''''''2_bufchan_d ;
  
  /* fork (Ty Pointer_QTree_Bool) : (lizzieLet65_4Lf''''''''''''sbos,Pointer_QTree_Bool) > [(lizzieLet65_4Lf''''''''''''sbos_1_merge_merge_fork_1,Pointer_QTree_Bool),
                                                                                       (lizzieLet65_4Lf''''''''''''sbos_1_merge_merge_fork_2,Pointer_QTree_Bool)] */
  logic [1:0] \lizzieLet65_4Lf''''''''''''sbos_emitted ;
  logic [1:0] \lizzieLet65_4Lf''''''''''''sbos_done ;
  assign \lizzieLet65_4Lf''''''''''''sbos_1_merge_merge_fork_1_d  = {\lizzieLet65_4Lf''''''''''''sbos_d [16:1],
                                                                     (\lizzieLet65_4Lf''''''''''''sbos_d [0] && (! \lizzieLet65_4Lf''''''''''''sbos_emitted [0]))};
  assign \lizzieLet65_4Lf''''''''''''sbos_1_merge_merge_fork_2_d  = {\lizzieLet65_4Lf''''''''''''sbos_d [16:1],
                                                                     (\lizzieLet65_4Lf''''''''''''sbos_d [0] && (! \lizzieLet65_4Lf''''''''''''sbos_emitted [1]))};
  assign \lizzieLet65_4Lf''''''''''''sbos_done  = (\lizzieLet65_4Lf''''''''''''sbos_emitted  | ({\lizzieLet65_4Lf''''''''''''sbos_1_merge_merge_fork_2_d [0],
                                                                                                 \lizzieLet65_4Lf''''''''''''sbos_1_merge_merge_fork_1_d [0]} & {\lizzieLet65_4Lf''''''''''''sbos_1_merge_merge_fork_2_r ,
                                                                                                                                                                 \lizzieLet65_4Lf''''''''''''sbos_1_merge_merge_fork_1_r }));
  assign \lizzieLet65_4Lf''''''''''''sbos_r  = (& \lizzieLet65_4Lf''''''''''''sbos_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet65_4Lf''''''''''''sbos_emitted  <= 2'd0;
    else
      \lizzieLet65_4Lf''''''''''''sbos_emitted  <= (\lizzieLet65_4Lf''''''''''''sbos_r  ? 2'd0 :
                                                    \lizzieLet65_4Lf''''''''''''sbos_done );
  
  /* togo (Ty Pointer_QTree_Bool) : (lizzieLet65_4Lf''''''''''''sbos_1_merge_merge_fork_1,Pointer_QTree_Bool) > (call_f''''''''''''_goConst,Go) */
  assign \call_f''''''''''''_goConst_d  = \lizzieLet65_4Lf''''''''''''sbos_1_merge_merge_fork_1_d [0];
  assign \lizzieLet65_4Lf''''''''''''sbos_1_merge_merge_fork_1_r  = \call_f''''''''''''_goConst_r ;
  
  /* mergectrl (Ty C10,Ty TupGo) : [(lvlrf2-0TupGo_1,TupGo),
                               (lvlrf2-0TupGo2,TupGo),
                               (lvlrf2-0TupGo3,TupGo),
                               (lvlrf2-0TupGo4,TupGo),
                               (lvlrf2-0TupGo5,TupGo),
                               (lvlrf2-0TupGo6,TupGo),
                               (lvlrf2-0TupGo7,TupGo),
                               (lvlrf2-0TupGo8,TupGo),
                               (lvlrf2-0TupGo9,TupGo),
                               (lvlrf2-0TupGo10,TupGo)] > (lvlrf2-0_choice,C10) (lvlrf2-0_data,TupGo) */
  logic [9:0] \lvlrf2-0TupGo_1_select_d ;
  assign \lvlrf2-0TupGo_1_select_d  = ((| \lvlrf2-0TupGo_1_select_q ) ? \lvlrf2-0TupGo_1_select_q  :
                                       (\lvlrf2-0TupGo_1_d [0] ? 10'd1 :
                                        (\lvlrf2-0TupGo2_d [0] ? 10'd2 :
                                         (\lvlrf2-0TupGo3_d [0] ? 10'd4 :
                                          (\lvlrf2-0TupGo4_d [0] ? 10'd8 :
                                           (\lvlrf2-0TupGo5_d [0] ? 10'd16 :
                                            (\lvlrf2-0TupGo6_d [0] ? 10'd32 :
                                             (\lvlrf2-0TupGo7_d [0] ? 10'd64 :
                                              (\lvlrf2-0TupGo8_d [0] ? 10'd128 :
                                               (\lvlrf2-0TupGo9_d [0] ? 10'd256 :
                                                (\lvlrf2-0TupGo10_d [0] ? 10'd512 :
                                                 10'd0)))))))))));
  logic [9:0] \lvlrf2-0TupGo_1_select_q ;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \lvlrf2-0TupGo_1_select_q  <= 10'd0;
    else
      \lvlrf2-0TupGo_1_select_q  <= (\lvlrf2-0TupGo_1_done  ? 10'd0 :
                                     \lvlrf2-0TupGo_1_select_d );
  logic [1:0] \lvlrf2-0TupGo_1_emit_q ;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \lvlrf2-0TupGo_1_emit_q  <= 2'd0;
    else
      \lvlrf2-0TupGo_1_emit_q  <= (\lvlrf2-0TupGo_1_done  ? 2'd0 :
                                   \lvlrf2-0TupGo_1_emit_d );
  logic [1:0] \lvlrf2-0TupGo_1_emit_d ;
  assign \lvlrf2-0TupGo_1_emit_d  = (\lvlrf2-0TupGo_1_emit_q  | ({\lvlrf2-0_choice_d [0],
                                                                  \lvlrf2-0_data_d [0]} & {\lvlrf2-0_choice_r ,
                                                                                           \lvlrf2-0_data_r }));
  logic \lvlrf2-0TupGo_1_done ;
  assign \lvlrf2-0TupGo_1_done  = (& \lvlrf2-0TupGo_1_emit_d );
  assign {\lvlrf2-0TupGo10_r ,
          \lvlrf2-0TupGo9_r ,
          \lvlrf2-0TupGo8_r ,
          \lvlrf2-0TupGo7_r ,
          \lvlrf2-0TupGo6_r ,
          \lvlrf2-0TupGo5_r ,
          \lvlrf2-0TupGo4_r ,
          \lvlrf2-0TupGo3_r ,
          \lvlrf2-0TupGo2_r ,
          \lvlrf2-0TupGo_1_r } = (\lvlrf2-0TupGo_1_done  ? \lvlrf2-0TupGo_1_select_d  :
                                  10'd0);
  assign \lvlrf2-0_data_d  = ((\lvlrf2-0TupGo_1_select_d [0] && (! \lvlrf2-0TupGo_1_emit_q [0])) ? \lvlrf2-0TupGo_1_d  :
                              ((\lvlrf2-0TupGo_1_select_d [1] && (! \lvlrf2-0TupGo_1_emit_q [0])) ? \lvlrf2-0TupGo2_d  :
                               ((\lvlrf2-0TupGo_1_select_d [2] && (! \lvlrf2-0TupGo_1_emit_q [0])) ? \lvlrf2-0TupGo3_d  :
                                ((\lvlrf2-0TupGo_1_select_d [3] && (! \lvlrf2-0TupGo_1_emit_q [0])) ? \lvlrf2-0TupGo4_d  :
                                 ((\lvlrf2-0TupGo_1_select_d [4] && (! \lvlrf2-0TupGo_1_emit_q [0])) ? \lvlrf2-0TupGo5_d  :
                                  ((\lvlrf2-0TupGo_1_select_d [5] && (! \lvlrf2-0TupGo_1_emit_q [0])) ? \lvlrf2-0TupGo6_d  :
                                   ((\lvlrf2-0TupGo_1_select_d [6] && (! \lvlrf2-0TupGo_1_emit_q [0])) ? \lvlrf2-0TupGo7_d  :
                                    ((\lvlrf2-0TupGo_1_select_d [7] && (! \lvlrf2-0TupGo_1_emit_q [0])) ? \lvlrf2-0TupGo8_d  :
                                     ((\lvlrf2-0TupGo_1_select_d [8] && (! \lvlrf2-0TupGo_1_emit_q [0])) ? \lvlrf2-0TupGo9_d  :
                                      ((\lvlrf2-0TupGo_1_select_d [9] && (! \lvlrf2-0TupGo_1_emit_q [0])) ? \lvlrf2-0TupGo10_d  :
                                       1'd0))))))))));
  assign \lvlrf2-0_choice_d  = ((\lvlrf2-0TupGo_1_select_d [0] && (! \lvlrf2-0TupGo_1_emit_q [1])) ? C1_10_dc(1'd1) :
                                ((\lvlrf2-0TupGo_1_select_d [1] && (! \lvlrf2-0TupGo_1_emit_q [1])) ? C2_10_dc(1'd1) :
                                 ((\lvlrf2-0TupGo_1_select_d [2] && (! \lvlrf2-0TupGo_1_emit_q [1])) ? C3_10_dc(1'd1) :
                                  ((\lvlrf2-0TupGo_1_select_d [3] && (! \lvlrf2-0TupGo_1_emit_q [1])) ? C4_10_dc(1'd1) :
                                   ((\lvlrf2-0TupGo_1_select_d [4] && (! \lvlrf2-0TupGo_1_emit_q [1])) ? C5_10_dc(1'd1) :
                                    ((\lvlrf2-0TupGo_1_select_d [5] && (! \lvlrf2-0TupGo_1_emit_q [1])) ? C6_10_dc(1'd1) :
                                     ((\lvlrf2-0TupGo_1_select_d [6] && (! \lvlrf2-0TupGo_1_emit_q [1])) ? C7_10_dc(1'd1) :
                                      ((\lvlrf2-0TupGo_1_select_d [7] && (! \lvlrf2-0TupGo_1_emit_q [1])) ? C8_10_dc(1'd1) :
                                       ((\lvlrf2-0TupGo_1_select_d [8] && (! \lvlrf2-0TupGo_1_emit_q [1])) ? C9_10_dc(1'd1) :
                                        ((\lvlrf2-0TupGo_1_select_d [9] && (! \lvlrf2-0TupGo_1_emit_q [1])) ? C10_10_dc(1'd1) :
                                         {4'd0, 1'd0}))))))))));
  
  /* dcon (Ty MyBool,
      Dcon MyTrue) : [(lvlrf2-0TupGogo_6,Go)] > (go_6_1MyTrue,MyBool) */
  assign go_6_1MyTrue_d = MyTrue_dc((& {\lvlrf2-0TupGogo_6_d [0]}), \lvlrf2-0TupGogo_6_d );
  assign {\lvlrf2-0TupGogo_6_r } = {1 {(go_6_1MyTrue_r && go_6_1MyTrue_d[0])}};
  
  /* buf (Ty Pointer_QTree_Bool) : (lvlrf2-0_1,Pointer_QTree_Bool) > (lvlrf2-0_resbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t \lvlrf2-0_1_bufchan_d ;
  logic \lvlrf2-0_1_bufchan_r ;
  assign \lvlrf2-0_1_r  = ((! \lvlrf2-0_1_bufchan_d [0]) || \lvlrf2-0_1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \lvlrf2-0_1_bufchan_d  <= {16'd0, 1'd0};
    else if (\lvlrf2-0_1_r ) \lvlrf2-0_1_bufchan_d  <= \lvlrf2-0_1_d ;
  Pointer_QTree_Bool_t \lvlrf2-0_1_bufchan_buf ;
  assign \lvlrf2-0_1_bufchan_r  = (! \lvlrf2-0_1_bufchan_buf [0]);
  assign \lvlrf2-0_resbuf_d  = (\lvlrf2-0_1_bufchan_buf [0] ? \lvlrf2-0_1_bufchan_buf  :
                                \lvlrf2-0_1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \lvlrf2-0_1_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((\lvlrf2-0_resbuf_r  && \lvlrf2-0_1_bufchan_buf [0]))
        \lvlrf2-0_1_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! \lvlrf2-0_resbuf_r ) && (! \lvlrf2-0_1_bufchan_buf [0])))
        \lvlrf2-0_1_bufchan_buf  <= \lvlrf2-0_1_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Bool) : (lvlrf2-0_10,Pointer_QTree_Bool) > (lvlrf2-0_10_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t \lvlrf2-0_10_bufchan_d ;
  logic \lvlrf2-0_10_bufchan_r ;
  assign \lvlrf2-0_10_r  = ((! \lvlrf2-0_10_bufchan_d [0]) || \lvlrf2-0_10_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \lvlrf2-0_10_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\lvlrf2-0_10_r ) \lvlrf2-0_10_bufchan_d  <= \lvlrf2-0_10_d ;
  Pointer_QTree_Bool_t \lvlrf2-0_10_bufchan_buf ;
  assign \lvlrf2-0_10_bufchan_r  = (! \lvlrf2-0_10_bufchan_buf [0]);
  assign \lvlrf2-0_10_argbuf_d  = (\lvlrf2-0_10_bufchan_buf [0] ? \lvlrf2-0_10_bufchan_buf  :
                                   \lvlrf2-0_10_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \lvlrf2-0_10_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((\lvlrf2-0_10_argbuf_r  && \lvlrf2-0_10_bufchan_buf [0]))
        \lvlrf2-0_10_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! \lvlrf2-0_10_argbuf_r ) && (! \lvlrf2-0_10_bufchan_buf [0])))
        \lvlrf2-0_10_bufchan_buf  <= \lvlrf2-0_10_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Bool) : (lvlrf2-0_10_argbuf,Pointer_QTree_Bool) > (lizzieLet27_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t \lvlrf2-0_10_argbuf_bufchan_d ;
  logic \lvlrf2-0_10_argbuf_bufchan_r ;
  assign \lvlrf2-0_10_argbuf_r  = ((! \lvlrf2-0_10_argbuf_bufchan_d [0]) || \lvlrf2-0_10_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lvlrf2-0_10_argbuf_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\lvlrf2-0_10_argbuf_r )
        \lvlrf2-0_10_argbuf_bufchan_d  <= \lvlrf2-0_10_argbuf_d ;
  Pointer_QTree_Bool_t \lvlrf2-0_10_argbuf_bufchan_buf ;
  assign \lvlrf2-0_10_argbuf_bufchan_r  = (! \lvlrf2-0_10_argbuf_bufchan_buf [0]);
  assign lizzieLet27_1_argbuf_d = (\lvlrf2-0_10_argbuf_bufchan_buf [0] ? \lvlrf2-0_10_argbuf_bufchan_buf  :
                                   \lvlrf2-0_10_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lvlrf2-0_10_argbuf_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((lizzieLet27_1_argbuf_r && \lvlrf2-0_10_argbuf_bufchan_buf [0]))
        \lvlrf2-0_10_argbuf_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! lizzieLet27_1_argbuf_r) && (! \lvlrf2-0_10_argbuf_bufchan_buf [0])))
        \lvlrf2-0_10_argbuf_bufchan_buf  <= \lvlrf2-0_10_argbuf_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Bool) : (lvlrf2-0_2,Pointer_QTree_Bool) > (lvlrf2-0_2_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t \lvlrf2-0_2_bufchan_d ;
  logic \lvlrf2-0_2_bufchan_r ;
  assign \lvlrf2-0_2_r  = ((! \lvlrf2-0_2_bufchan_d [0]) || \lvlrf2-0_2_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \lvlrf2-0_2_bufchan_d  <= {16'd0, 1'd0};
    else if (\lvlrf2-0_2_r ) \lvlrf2-0_2_bufchan_d  <= \lvlrf2-0_2_d ;
  Pointer_QTree_Bool_t \lvlrf2-0_2_bufchan_buf ;
  assign \lvlrf2-0_2_bufchan_r  = (! \lvlrf2-0_2_bufchan_buf [0]);
  assign \lvlrf2-0_2_argbuf_d  = (\lvlrf2-0_2_bufchan_buf [0] ? \lvlrf2-0_2_bufchan_buf  :
                                  \lvlrf2-0_2_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \lvlrf2-0_2_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((\lvlrf2-0_2_argbuf_r  && \lvlrf2-0_2_bufchan_buf [0]))
        \lvlrf2-0_2_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! \lvlrf2-0_2_argbuf_r ) && (! \lvlrf2-0_2_bufchan_buf [0])))
        \lvlrf2-0_2_bufchan_buf  <= \lvlrf2-0_2_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Bool) : (lvlrf2-0_2_argbuf,Pointer_QTree_Bool) > (lizzieLet5_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t \lvlrf2-0_2_argbuf_bufchan_d ;
  logic \lvlrf2-0_2_argbuf_bufchan_r ;
  assign \lvlrf2-0_2_argbuf_r  = ((! \lvlrf2-0_2_argbuf_bufchan_d [0]) || \lvlrf2-0_2_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lvlrf2-0_2_argbuf_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\lvlrf2-0_2_argbuf_r )
        \lvlrf2-0_2_argbuf_bufchan_d  <= \lvlrf2-0_2_argbuf_d ;
  Pointer_QTree_Bool_t \lvlrf2-0_2_argbuf_bufchan_buf ;
  assign \lvlrf2-0_2_argbuf_bufchan_r  = (! \lvlrf2-0_2_argbuf_bufchan_buf [0]);
  assign lizzieLet5_1_argbuf_d = (\lvlrf2-0_2_argbuf_bufchan_buf [0] ? \lvlrf2-0_2_argbuf_bufchan_buf  :
                                  \lvlrf2-0_2_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lvlrf2-0_2_argbuf_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((lizzieLet5_1_argbuf_r && \lvlrf2-0_2_argbuf_bufchan_buf [0]))
        \lvlrf2-0_2_argbuf_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! lizzieLet5_1_argbuf_r) && (! \lvlrf2-0_2_argbuf_bufchan_buf [0])))
        \lvlrf2-0_2_argbuf_bufchan_buf  <= \lvlrf2-0_2_argbuf_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Bool) : (lvlrf2-0_3,Pointer_QTree_Bool) > (lvlrf2-0_3_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t \lvlrf2-0_3_bufchan_d ;
  logic \lvlrf2-0_3_bufchan_r ;
  assign \lvlrf2-0_3_r  = ((! \lvlrf2-0_3_bufchan_d [0]) || \lvlrf2-0_3_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \lvlrf2-0_3_bufchan_d  <= {16'd0, 1'd0};
    else if (\lvlrf2-0_3_r ) \lvlrf2-0_3_bufchan_d  <= \lvlrf2-0_3_d ;
  Pointer_QTree_Bool_t \lvlrf2-0_3_bufchan_buf ;
  assign \lvlrf2-0_3_bufchan_r  = (! \lvlrf2-0_3_bufchan_buf [0]);
  assign \lvlrf2-0_3_argbuf_d  = (\lvlrf2-0_3_bufchan_buf [0] ? \lvlrf2-0_3_bufchan_buf  :
                                  \lvlrf2-0_3_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \lvlrf2-0_3_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((\lvlrf2-0_3_argbuf_r  && \lvlrf2-0_3_bufchan_buf [0]))
        \lvlrf2-0_3_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! \lvlrf2-0_3_argbuf_r ) && (! \lvlrf2-0_3_bufchan_buf [0])))
        \lvlrf2-0_3_bufchan_buf  <= \lvlrf2-0_3_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Bool) : (lvlrf2-0_3_argbuf,Pointer_QTree_Bool) > (lizzieLet48_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t \lvlrf2-0_3_argbuf_bufchan_d ;
  logic \lvlrf2-0_3_argbuf_bufchan_r ;
  assign \lvlrf2-0_3_argbuf_r  = ((! \lvlrf2-0_3_argbuf_bufchan_d [0]) || \lvlrf2-0_3_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lvlrf2-0_3_argbuf_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\lvlrf2-0_3_argbuf_r )
        \lvlrf2-0_3_argbuf_bufchan_d  <= \lvlrf2-0_3_argbuf_d ;
  Pointer_QTree_Bool_t \lvlrf2-0_3_argbuf_bufchan_buf ;
  assign \lvlrf2-0_3_argbuf_bufchan_r  = (! \lvlrf2-0_3_argbuf_bufchan_buf [0]);
  assign lizzieLet48_1_argbuf_d = (\lvlrf2-0_3_argbuf_bufchan_buf [0] ? \lvlrf2-0_3_argbuf_bufchan_buf  :
                                   \lvlrf2-0_3_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lvlrf2-0_3_argbuf_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((lizzieLet48_1_argbuf_r && \lvlrf2-0_3_argbuf_bufchan_buf [0]))
        \lvlrf2-0_3_argbuf_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! lizzieLet48_1_argbuf_r) && (! \lvlrf2-0_3_argbuf_bufchan_buf [0])))
        \lvlrf2-0_3_argbuf_bufchan_buf  <= \lvlrf2-0_3_argbuf_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Bool) : (lvlrf2-0_4,Pointer_QTree_Bool) > (lvlrf2-0_4_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t \lvlrf2-0_4_bufchan_d ;
  logic \lvlrf2-0_4_bufchan_r ;
  assign \lvlrf2-0_4_r  = ((! \lvlrf2-0_4_bufchan_d [0]) || \lvlrf2-0_4_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \lvlrf2-0_4_bufchan_d  <= {16'd0, 1'd0};
    else if (\lvlrf2-0_4_r ) \lvlrf2-0_4_bufchan_d  <= \lvlrf2-0_4_d ;
  Pointer_QTree_Bool_t \lvlrf2-0_4_bufchan_buf ;
  assign \lvlrf2-0_4_bufchan_r  = (! \lvlrf2-0_4_bufchan_buf [0]);
  assign \lvlrf2-0_4_argbuf_d  = (\lvlrf2-0_4_bufchan_buf [0] ? \lvlrf2-0_4_bufchan_buf  :
                                  \lvlrf2-0_4_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \lvlrf2-0_4_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((\lvlrf2-0_4_argbuf_r  && \lvlrf2-0_4_bufchan_buf [0]))
        \lvlrf2-0_4_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! \lvlrf2-0_4_argbuf_r ) && (! \lvlrf2-0_4_bufchan_buf [0])))
        \lvlrf2-0_4_bufchan_buf  <= \lvlrf2-0_4_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Bool) : (lvlrf2-0_4_argbuf,Pointer_QTree_Bool) > (lizzieLet49_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t \lvlrf2-0_4_argbuf_bufchan_d ;
  logic \lvlrf2-0_4_argbuf_bufchan_r ;
  assign \lvlrf2-0_4_argbuf_r  = ((! \lvlrf2-0_4_argbuf_bufchan_d [0]) || \lvlrf2-0_4_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lvlrf2-0_4_argbuf_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\lvlrf2-0_4_argbuf_r )
        \lvlrf2-0_4_argbuf_bufchan_d  <= \lvlrf2-0_4_argbuf_d ;
  Pointer_QTree_Bool_t \lvlrf2-0_4_argbuf_bufchan_buf ;
  assign \lvlrf2-0_4_argbuf_bufchan_r  = (! \lvlrf2-0_4_argbuf_bufchan_buf [0]);
  assign lizzieLet49_1_argbuf_d = (\lvlrf2-0_4_argbuf_bufchan_buf [0] ? \lvlrf2-0_4_argbuf_bufchan_buf  :
                                   \lvlrf2-0_4_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lvlrf2-0_4_argbuf_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((lizzieLet49_1_argbuf_r && \lvlrf2-0_4_argbuf_bufchan_buf [0]))
        \lvlrf2-0_4_argbuf_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! lizzieLet49_1_argbuf_r) && (! \lvlrf2-0_4_argbuf_bufchan_buf [0])))
        \lvlrf2-0_4_argbuf_bufchan_buf  <= \lvlrf2-0_4_argbuf_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Bool) : (lvlrf2-0_5,Pointer_QTree_Bool) > (lvlrf2-0_5_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t \lvlrf2-0_5_bufchan_d ;
  logic \lvlrf2-0_5_bufchan_r ;
  assign \lvlrf2-0_5_r  = ((! \lvlrf2-0_5_bufchan_d [0]) || \lvlrf2-0_5_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \lvlrf2-0_5_bufchan_d  <= {16'd0, 1'd0};
    else if (\lvlrf2-0_5_r ) \lvlrf2-0_5_bufchan_d  <= \lvlrf2-0_5_d ;
  Pointer_QTree_Bool_t \lvlrf2-0_5_bufchan_buf ;
  assign \lvlrf2-0_5_bufchan_r  = (! \lvlrf2-0_5_bufchan_buf [0]);
  assign \lvlrf2-0_5_argbuf_d  = (\lvlrf2-0_5_bufchan_buf [0] ? \lvlrf2-0_5_bufchan_buf  :
                                  \lvlrf2-0_5_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \lvlrf2-0_5_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((\lvlrf2-0_5_argbuf_r  && \lvlrf2-0_5_bufchan_buf [0]))
        \lvlrf2-0_5_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! \lvlrf2-0_5_argbuf_r ) && (! \lvlrf2-0_5_bufchan_buf [0])))
        \lvlrf2-0_5_bufchan_buf  <= \lvlrf2-0_5_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Bool) : (lvlrf2-0_5_argbuf,Pointer_QTree_Bool) > (lizzieLet16_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t \lvlrf2-0_5_argbuf_bufchan_d ;
  logic \lvlrf2-0_5_argbuf_bufchan_r ;
  assign \lvlrf2-0_5_argbuf_r  = ((! \lvlrf2-0_5_argbuf_bufchan_d [0]) || \lvlrf2-0_5_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lvlrf2-0_5_argbuf_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\lvlrf2-0_5_argbuf_r )
        \lvlrf2-0_5_argbuf_bufchan_d  <= \lvlrf2-0_5_argbuf_d ;
  Pointer_QTree_Bool_t \lvlrf2-0_5_argbuf_bufchan_buf ;
  assign \lvlrf2-0_5_argbuf_bufchan_r  = (! \lvlrf2-0_5_argbuf_bufchan_buf [0]);
  assign lizzieLet16_1_argbuf_d = (\lvlrf2-0_5_argbuf_bufchan_buf [0] ? \lvlrf2-0_5_argbuf_bufchan_buf  :
                                   \lvlrf2-0_5_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lvlrf2-0_5_argbuf_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((lizzieLet16_1_argbuf_r && \lvlrf2-0_5_argbuf_bufchan_buf [0]))
        \lvlrf2-0_5_argbuf_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! lizzieLet16_1_argbuf_r) && (! \lvlrf2-0_5_argbuf_bufchan_buf [0])))
        \lvlrf2-0_5_argbuf_bufchan_buf  <= \lvlrf2-0_5_argbuf_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Bool) : (lvlrf2-0_6,Pointer_QTree_Bool) > (lvlrf2-0_6_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t \lvlrf2-0_6_bufchan_d ;
  logic \lvlrf2-0_6_bufchan_r ;
  assign \lvlrf2-0_6_r  = ((! \lvlrf2-0_6_bufchan_d [0]) || \lvlrf2-0_6_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \lvlrf2-0_6_bufchan_d  <= {16'd0, 1'd0};
    else if (\lvlrf2-0_6_r ) \lvlrf2-0_6_bufchan_d  <= \lvlrf2-0_6_d ;
  Pointer_QTree_Bool_t \lvlrf2-0_6_bufchan_buf ;
  assign \lvlrf2-0_6_bufchan_r  = (! \lvlrf2-0_6_bufchan_buf [0]);
  assign \lvlrf2-0_6_argbuf_d  = (\lvlrf2-0_6_bufchan_buf [0] ? \lvlrf2-0_6_bufchan_buf  :
                                  \lvlrf2-0_6_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \lvlrf2-0_6_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((\lvlrf2-0_6_argbuf_r  && \lvlrf2-0_6_bufchan_buf [0]))
        \lvlrf2-0_6_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! \lvlrf2-0_6_argbuf_r ) && (! \lvlrf2-0_6_bufchan_buf [0])))
        \lvlrf2-0_6_bufchan_buf  <= \lvlrf2-0_6_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Bool) : (lvlrf2-0_6_argbuf,Pointer_QTree_Bool) > (lizzieLet17_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t \lvlrf2-0_6_argbuf_bufchan_d ;
  logic \lvlrf2-0_6_argbuf_bufchan_r ;
  assign \lvlrf2-0_6_argbuf_r  = ((! \lvlrf2-0_6_argbuf_bufchan_d [0]) || \lvlrf2-0_6_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lvlrf2-0_6_argbuf_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\lvlrf2-0_6_argbuf_r )
        \lvlrf2-0_6_argbuf_bufchan_d  <= \lvlrf2-0_6_argbuf_d ;
  Pointer_QTree_Bool_t \lvlrf2-0_6_argbuf_bufchan_buf ;
  assign \lvlrf2-0_6_argbuf_bufchan_r  = (! \lvlrf2-0_6_argbuf_bufchan_buf [0]);
  assign lizzieLet17_1_argbuf_d = (\lvlrf2-0_6_argbuf_bufchan_buf [0] ? \lvlrf2-0_6_argbuf_bufchan_buf  :
                                   \lvlrf2-0_6_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lvlrf2-0_6_argbuf_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((lizzieLet17_1_argbuf_r && \lvlrf2-0_6_argbuf_bufchan_buf [0]))
        \lvlrf2-0_6_argbuf_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! lizzieLet17_1_argbuf_r) && (! \lvlrf2-0_6_argbuf_bufchan_buf [0])))
        \lvlrf2-0_6_argbuf_bufchan_buf  <= \lvlrf2-0_6_argbuf_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Bool) : (lvlrf2-0_7,Pointer_QTree_Bool) > (lvlrf2-0_7_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t \lvlrf2-0_7_bufchan_d ;
  logic \lvlrf2-0_7_bufchan_r ;
  assign \lvlrf2-0_7_r  = ((! \lvlrf2-0_7_bufchan_d [0]) || \lvlrf2-0_7_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \lvlrf2-0_7_bufchan_d  <= {16'd0, 1'd0};
    else if (\lvlrf2-0_7_r ) \lvlrf2-0_7_bufchan_d  <= \lvlrf2-0_7_d ;
  Pointer_QTree_Bool_t \lvlrf2-0_7_bufchan_buf ;
  assign \lvlrf2-0_7_bufchan_r  = (! \lvlrf2-0_7_bufchan_buf [0]);
  assign \lvlrf2-0_7_argbuf_d  = (\lvlrf2-0_7_bufchan_buf [0] ? \lvlrf2-0_7_bufchan_buf  :
                                  \lvlrf2-0_7_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \lvlrf2-0_7_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((\lvlrf2-0_7_argbuf_r  && \lvlrf2-0_7_bufchan_buf [0]))
        \lvlrf2-0_7_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! \lvlrf2-0_7_argbuf_r ) && (! \lvlrf2-0_7_bufchan_buf [0])))
        \lvlrf2-0_7_bufchan_buf  <= \lvlrf2-0_7_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Bool) : (lvlrf2-0_7_argbuf,Pointer_QTree_Bool) > (lizzieLet21_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t \lvlrf2-0_7_argbuf_bufchan_d ;
  logic \lvlrf2-0_7_argbuf_bufchan_r ;
  assign \lvlrf2-0_7_argbuf_r  = ((! \lvlrf2-0_7_argbuf_bufchan_d [0]) || \lvlrf2-0_7_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lvlrf2-0_7_argbuf_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\lvlrf2-0_7_argbuf_r )
        \lvlrf2-0_7_argbuf_bufchan_d  <= \lvlrf2-0_7_argbuf_d ;
  Pointer_QTree_Bool_t \lvlrf2-0_7_argbuf_bufchan_buf ;
  assign \lvlrf2-0_7_argbuf_bufchan_r  = (! \lvlrf2-0_7_argbuf_bufchan_buf [0]);
  assign lizzieLet21_1_argbuf_d = (\lvlrf2-0_7_argbuf_bufchan_buf [0] ? \lvlrf2-0_7_argbuf_bufchan_buf  :
                                   \lvlrf2-0_7_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lvlrf2-0_7_argbuf_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((lizzieLet21_1_argbuf_r && \lvlrf2-0_7_argbuf_bufchan_buf [0]))
        \lvlrf2-0_7_argbuf_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! lizzieLet21_1_argbuf_r) && (! \lvlrf2-0_7_argbuf_bufchan_buf [0])))
        \lvlrf2-0_7_argbuf_bufchan_buf  <= \lvlrf2-0_7_argbuf_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Bool) : (lvlrf2-0_8,Pointer_QTree_Bool) > (lvlrf2-0_8_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t \lvlrf2-0_8_bufchan_d ;
  logic \lvlrf2-0_8_bufchan_r ;
  assign \lvlrf2-0_8_r  = ((! \lvlrf2-0_8_bufchan_d [0]) || \lvlrf2-0_8_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \lvlrf2-0_8_bufchan_d  <= {16'd0, 1'd0};
    else if (\lvlrf2-0_8_r ) \lvlrf2-0_8_bufchan_d  <= \lvlrf2-0_8_d ;
  Pointer_QTree_Bool_t \lvlrf2-0_8_bufchan_buf ;
  assign \lvlrf2-0_8_bufchan_r  = (! \lvlrf2-0_8_bufchan_buf [0]);
  assign \lvlrf2-0_8_argbuf_d  = (\lvlrf2-0_8_bufchan_buf [0] ? \lvlrf2-0_8_bufchan_buf  :
                                  \lvlrf2-0_8_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \lvlrf2-0_8_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((\lvlrf2-0_8_argbuf_r  && \lvlrf2-0_8_bufchan_buf [0]))
        \lvlrf2-0_8_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! \lvlrf2-0_8_argbuf_r ) && (! \lvlrf2-0_8_bufchan_buf [0])))
        \lvlrf2-0_8_bufchan_buf  <= \lvlrf2-0_8_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Bool) : (lvlrf2-0_8_argbuf,Pointer_QTree_Bool) > (lizzieLet22_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t \lvlrf2-0_8_argbuf_bufchan_d ;
  logic \lvlrf2-0_8_argbuf_bufchan_r ;
  assign \lvlrf2-0_8_argbuf_r  = ((! \lvlrf2-0_8_argbuf_bufchan_d [0]) || \lvlrf2-0_8_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lvlrf2-0_8_argbuf_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\lvlrf2-0_8_argbuf_r )
        \lvlrf2-0_8_argbuf_bufchan_d  <= \lvlrf2-0_8_argbuf_d ;
  Pointer_QTree_Bool_t \lvlrf2-0_8_argbuf_bufchan_buf ;
  assign \lvlrf2-0_8_argbuf_bufchan_r  = (! \lvlrf2-0_8_argbuf_bufchan_buf [0]);
  assign lizzieLet22_1_argbuf_d = (\lvlrf2-0_8_argbuf_bufchan_buf [0] ? \lvlrf2-0_8_argbuf_bufchan_buf  :
                                   \lvlrf2-0_8_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lvlrf2-0_8_argbuf_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((lizzieLet22_1_argbuf_r && \lvlrf2-0_8_argbuf_bufchan_buf [0]))
        \lvlrf2-0_8_argbuf_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! lizzieLet22_1_argbuf_r) && (! \lvlrf2-0_8_argbuf_bufchan_buf [0])))
        \lvlrf2-0_8_argbuf_bufchan_buf  <= \lvlrf2-0_8_argbuf_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Bool) : (lvlrf2-0_9,Pointer_QTree_Bool) > (lvlrf2-0_9_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t \lvlrf2-0_9_bufchan_d ;
  logic \lvlrf2-0_9_bufchan_r ;
  assign \lvlrf2-0_9_r  = ((! \lvlrf2-0_9_bufchan_d [0]) || \lvlrf2-0_9_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \lvlrf2-0_9_bufchan_d  <= {16'd0, 1'd0};
    else if (\lvlrf2-0_9_r ) \lvlrf2-0_9_bufchan_d  <= \lvlrf2-0_9_d ;
  Pointer_QTree_Bool_t \lvlrf2-0_9_bufchan_buf ;
  assign \lvlrf2-0_9_bufchan_r  = (! \lvlrf2-0_9_bufchan_buf [0]);
  assign \lvlrf2-0_9_argbuf_d  = (\lvlrf2-0_9_bufchan_buf [0] ? \lvlrf2-0_9_bufchan_buf  :
                                  \lvlrf2-0_9_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \lvlrf2-0_9_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((\lvlrf2-0_9_argbuf_r  && \lvlrf2-0_9_bufchan_buf [0]))
        \lvlrf2-0_9_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! \lvlrf2-0_9_argbuf_r ) && (! \lvlrf2-0_9_bufchan_buf [0])))
        \lvlrf2-0_9_bufchan_buf  <= \lvlrf2-0_9_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Bool) : (lvlrf2-0_9_argbuf,Pointer_QTree_Bool) > (lizzieLet26_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t \lvlrf2-0_9_argbuf_bufchan_d ;
  logic \lvlrf2-0_9_argbuf_bufchan_r ;
  assign \lvlrf2-0_9_argbuf_r  = ((! \lvlrf2-0_9_argbuf_bufchan_d [0]) || \lvlrf2-0_9_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lvlrf2-0_9_argbuf_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\lvlrf2-0_9_argbuf_r )
        \lvlrf2-0_9_argbuf_bufchan_d  <= \lvlrf2-0_9_argbuf_d ;
  Pointer_QTree_Bool_t \lvlrf2-0_9_argbuf_bufchan_buf ;
  assign \lvlrf2-0_9_argbuf_bufchan_r  = (! \lvlrf2-0_9_argbuf_bufchan_buf [0]);
  assign lizzieLet26_1_argbuf_d = (\lvlrf2-0_9_argbuf_bufchan_buf [0] ? \lvlrf2-0_9_argbuf_bufchan_buf  :
                                   \lvlrf2-0_9_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lvlrf2-0_9_argbuf_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((lizzieLet26_1_argbuf_r && \lvlrf2-0_9_argbuf_bufchan_buf [0]))
        \lvlrf2-0_9_argbuf_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! lizzieLet26_1_argbuf_r) && (! \lvlrf2-0_9_argbuf_bufchan_buf [0])))
        \lvlrf2-0_9_argbuf_bufchan_buf  <= \lvlrf2-0_9_argbuf_bufchan_d ;
  
  /* demux (Ty C10,
       Ty Pointer_QTree_Bool) : (lvlrf2-0_choice,C10) (writeQTree_BoollizzieLet59_1_argbuf_rwb,Pointer_QTree_Bool) > [(lvlrf2-0_1,Pointer_QTree_Bool),
                                                                                                                      (lvlrf2-0_2,Pointer_QTree_Bool),
                                                                                                                      (lvlrf2-0_3,Pointer_QTree_Bool),
                                                                                                                      (lvlrf2-0_4,Pointer_QTree_Bool),
                                                                                                                      (lvlrf2-0_5,Pointer_QTree_Bool),
                                                                                                                      (lvlrf2-0_6,Pointer_QTree_Bool),
                                                                                                                      (lvlrf2-0_7,Pointer_QTree_Bool),
                                                                                                                      (lvlrf2-0_8,Pointer_QTree_Bool),
                                                                                                                      (lvlrf2-0_9,Pointer_QTree_Bool),
                                                                                                                      (lvlrf2-0_10,Pointer_QTree_Bool)] */
  logic [9:0] writeQTree_BoollizzieLet59_1_argbuf_rwb_onehotd;
  always_comb
    if ((\lvlrf2-0_choice_d [0] && writeQTree_BoollizzieLet59_1_argbuf_rwb_d[0]))
      unique case (\lvlrf2-0_choice_d [4:1])
        4'd0: writeQTree_BoollizzieLet59_1_argbuf_rwb_onehotd = 10'd1;
        4'd1: writeQTree_BoollizzieLet59_1_argbuf_rwb_onehotd = 10'd2;
        4'd2: writeQTree_BoollizzieLet59_1_argbuf_rwb_onehotd = 10'd4;
        4'd3: writeQTree_BoollizzieLet59_1_argbuf_rwb_onehotd = 10'd8;
        4'd4: writeQTree_BoollizzieLet59_1_argbuf_rwb_onehotd = 10'd16;
        4'd5: writeQTree_BoollizzieLet59_1_argbuf_rwb_onehotd = 10'd32;
        4'd6: writeQTree_BoollizzieLet59_1_argbuf_rwb_onehotd = 10'd64;
        4'd7: writeQTree_BoollizzieLet59_1_argbuf_rwb_onehotd = 10'd128;
        4'd8: writeQTree_BoollizzieLet59_1_argbuf_rwb_onehotd = 10'd256;
        4'd9: writeQTree_BoollizzieLet59_1_argbuf_rwb_onehotd = 10'd512;
        default: writeQTree_BoollizzieLet59_1_argbuf_rwb_onehotd = 10'd0;
      endcase
    else writeQTree_BoollizzieLet59_1_argbuf_rwb_onehotd = 10'd0;
  assign \lvlrf2-0_1_d  = {writeQTree_BoollizzieLet59_1_argbuf_rwb_d[16:1],
                           writeQTree_BoollizzieLet59_1_argbuf_rwb_onehotd[0]};
  assign \lvlrf2-0_2_d  = {writeQTree_BoollizzieLet59_1_argbuf_rwb_d[16:1],
                           writeQTree_BoollizzieLet59_1_argbuf_rwb_onehotd[1]};
  assign \lvlrf2-0_3_d  = {writeQTree_BoollizzieLet59_1_argbuf_rwb_d[16:1],
                           writeQTree_BoollizzieLet59_1_argbuf_rwb_onehotd[2]};
  assign \lvlrf2-0_4_d  = {writeQTree_BoollizzieLet59_1_argbuf_rwb_d[16:1],
                           writeQTree_BoollizzieLet59_1_argbuf_rwb_onehotd[3]};
  assign \lvlrf2-0_5_d  = {writeQTree_BoollizzieLet59_1_argbuf_rwb_d[16:1],
                           writeQTree_BoollizzieLet59_1_argbuf_rwb_onehotd[4]};
  assign \lvlrf2-0_6_d  = {writeQTree_BoollizzieLet59_1_argbuf_rwb_d[16:1],
                           writeQTree_BoollizzieLet59_1_argbuf_rwb_onehotd[5]};
  assign \lvlrf2-0_7_d  = {writeQTree_BoollizzieLet59_1_argbuf_rwb_d[16:1],
                           writeQTree_BoollizzieLet59_1_argbuf_rwb_onehotd[6]};
  assign \lvlrf2-0_8_d  = {writeQTree_BoollizzieLet59_1_argbuf_rwb_d[16:1],
                           writeQTree_BoollizzieLet59_1_argbuf_rwb_onehotd[7]};
  assign \lvlrf2-0_9_d  = {writeQTree_BoollizzieLet59_1_argbuf_rwb_d[16:1],
                           writeQTree_BoollizzieLet59_1_argbuf_rwb_onehotd[8]};
  assign \lvlrf2-0_10_d  = {writeQTree_BoollizzieLet59_1_argbuf_rwb_d[16:1],
                            writeQTree_BoollizzieLet59_1_argbuf_rwb_onehotd[9]};
  assign writeQTree_BoollizzieLet59_1_argbuf_rwb_r = (| (writeQTree_BoollizzieLet59_1_argbuf_rwb_onehotd & {\lvlrf2-0_10_r ,
                                                                                                            \lvlrf2-0_9_r ,
                                                                                                            \lvlrf2-0_8_r ,
                                                                                                            \lvlrf2-0_7_r ,
                                                                                                            \lvlrf2-0_6_r ,
                                                                                                            \lvlrf2-0_5_r ,
                                                                                                            \lvlrf2-0_4_r ,
                                                                                                            \lvlrf2-0_3_r ,
                                                                                                            \lvlrf2-0_2_r ,
                                                                                                            \lvlrf2-0_1_r }));
  assign \lvlrf2-0_choice_r  = writeQTree_BoollizzieLet59_1_argbuf_rwb_r;
  
  /* destruct (Ty TupGo,
          Dcon TupGo) : (lvlrf2-0_data,TupGo) > [(lvlrf2-0TupGogo_6,Go)] */
  assign \lvlrf2-0TupGogo_6_d  = \lvlrf2-0_data_d [0];
  assign \lvlrf2-0_data_r  = \lvlrf2-0TupGogo_6_r ;
  
  /* buf (Ty Pointer_QTree_Bool) : (lvlrf2-0_resbuf,Pointer_QTree_Bool) > (lizzieLet4_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t \lvlrf2-0_resbuf_bufchan_d ;
  logic \lvlrf2-0_resbuf_bufchan_r ;
  assign \lvlrf2-0_resbuf_r  = ((! \lvlrf2-0_resbuf_bufchan_d [0]) || \lvlrf2-0_resbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \lvlrf2-0_resbuf_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\lvlrf2-0_resbuf_r )
        \lvlrf2-0_resbuf_bufchan_d  <= \lvlrf2-0_resbuf_d ;
  Pointer_QTree_Bool_t \lvlrf2-0_resbuf_bufchan_buf ;
  assign \lvlrf2-0_resbuf_bufchan_r  = (! \lvlrf2-0_resbuf_bufchan_buf [0]);
  assign lizzieLet4_1_argbuf_d = (\lvlrf2-0_resbuf_bufchan_buf [0] ? \lvlrf2-0_resbuf_bufchan_buf  :
                                  \lvlrf2-0_resbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lvlrf2-0_resbuf_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((lizzieLet4_1_argbuf_r && \lvlrf2-0_resbuf_bufchan_buf [0]))
        \lvlrf2-0_resbuf_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! lizzieLet4_1_argbuf_r) && (! \lvlrf2-0_resbuf_bufchan_buf [0])))
        \lvlrf2-0_resbuf_bufchan_buf  <= \lvlrf2-0_resbuf_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Bool) : (m1a84_1,Pointer_QTree_Bool) > (m1a84_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t m1a84_1_bufchan_d;
  logic m1a84_1_bufchan_r;
  assign m1a84_1_r = ((! m1a84_1_bufchan_d[0]) || m1a84_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m1a84_1_bufchan_d <= {16'd0, 1'd0};
    else if (m1a84_1_r) m1a84_1_bufchan_d <= m1a84_1_d;
  Pointer_QTree_Bool_t m1a84_1_bufchan_buf;
  assign m1a84_1_bufchan_r = (! m1a84_1_bufchan_buf[0]);
  assign m1a84_1_argbuf_d = (m1a84_1_bufchan_buf[0] ? m1a84_1_bufchan_buf :
                             m1a84_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m1a84_1_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((m1a84_1_argbuf_r && m1a84_1_bufchan_buf[0]))
        m1a84_1_bufchan_buf <= {16'd0, 1'd0};
      else if (((! m1a84_1_argbuf_r) && (! m1a84_1_bufchan_buf[0])))
        m1a84_1_bufchan_buf <= m1a84_1_bufchan_d;
  
  /* fork (Ty Pointer_QTree_Bool) : (m1a84_goMux_mux,Pointer_QTree_Bool) > [(m1a84_1,Pointer_QTree_Bool),
                                                                       (m1a84_2,Pointer_QTree_Bool)] */
  logic [1:0] m1a84_goMux_mux_emitted;
  logic [1:0] m1a84_goMux_mux_done;
  assign m1a84_1_d = {m1a84_goMux_mux_d[16:1],
                      (m1a84_goMux_mux_d[0] && (! m1a84_goMux_mux_emitted[0]))};
  assign m1a84_2_d = {m1a84_goMux_mux_d[16:1],
                      (m1a84_goMux_mux_d[0] && (! m1a84_goMux_mux_emitted[1]))};
  assign m1a84_goMux_mux_done = (m1a84_goMux_mux_emitted | ({m1a84_2_d[0],
                                                             m1a84_1_d[0]} & {m1a84_2_r,
                                                                              m1a84_1_r}));
  assign m1a84_goMux_mux_r = (& m1a84_goMux_mux_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m1a84_goMux_mux_emitted <= 2'd0;
    else
      m1a84_goMux_mux_emitted <= (m1a84_goMux_mux_r ? 2'd0 :
                                  m1a84_goMux_mux_done);
  
  /* buf (Ty Pointer_QTree_Bool) : (m2a85_1,Pointer_QTree_Bool) > (m2a85_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t m2a85_1_bufchan_d;
  logic m2a85_1_bufchan_r;
  assign m2a85_1_r = ((! m2a85_1_bufchan_d[0]) || m2a85_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m2a85_1_bufchan_d <= {16'd0, 1'd0};
    else if (m2a85_1_r) m2a85_1_bufchan_d <= m2a85_1_d;
  Pointer_QTree_Bool_t m2a85_1_bufchan_buf;
  assign m2a85_1_bufchan_r = (! m2a85_1_bufchan_buf[0]);
  assign m2a85_1_argbuf_d = (m2a85_1_bufchan_buf[0] ? m2a85_1_bufchan_buf :
                             m2a85_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m2a85_1_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((m2a85_1_argbuf_r && m2a85_1_bufchan_buf[0]))
        m2a85_1_bufchan_buf <= {16'd0, 1'd0};
      else if (((! m2a85_1_argbuf_r) && (! m2a85_1_bufchan_buf[0])))
        m2a85_1_bufchan_buf <= m2a85_1_bufchan_d;
  
  /* fork (Ty Pointer_QTree_Bool) : (m2a85_goMux_mux,Pointer_QTree_Bool) > [(m2a85_1,Pointer_QTree_Bool),
                                                                       (m2a85_2,Pointer_QTree_Bool)] */
  logic [1:0] m2a85_goMux_mux_emitted;
  logic [1:0] m2a85_goMux_mux_done;
  assign m2a85_1_d = {m2a85_goMux_mux_d[16:1],
                      (m2a85_goMux_mux_d[0] && (! m2a85_goMux_mux_emitted[0]))};
  assign m2a85_2_d = {m2a85_goMux_mux_d[16:1],
                      (m2a85_goMux_mux_d[0] && (! m2a85_goMux_mux_emitted[1]))};
  assign m2a85_goMux_mux_done = (m2a85_goMux_mux_emitted | ({m2a85_2_d[0],
                                                             m2a85_1_d[0]} & {m2a85_2_r,
                                                                              m2a85_1_r}));
  assign m2a85_goMux_mux_r = (& m2a85_goMux_mux_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m2a85_goMux_mux_emitted <= 2'd0;
    else
      m2a85_goMux_mux_emitted <= (m2a85_goMux_mux_r ? 2'd0 :
                                  m2a85_goMux_mux_done);
  
  /* buf (Ty Pointer_QTree_Bool) : (m3a86_1,Pointer_QTree_Bool) > (m3a86_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t m3a86_1_bufchan_d;
  logic m3a86_1_bufchan_r;
  assign m3a86_1_r = ((! m3a86_1_bufchan_d[0]) || m3a86_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m3a86_1_bufchan_d <= {16'd0, 1'd0};
    else if (m3a86_1_r) m3a86_1_bufchan_d <= m3a86_1_d;
  Pointer_QTree_Bool_t m3a86_1_bufchan_buf;
  assign m3a86_1_bufchan_r = (! m3a86_1_bufchan_buf[0]);
  assign m3a86_1_argbuf_d = (m3a86_1_bufchan_buf[0] ? m3a86_1_bufchan_buf :
                             m3a86_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m3a86_1_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((m3a86_1_argbuf_r && m3a86_1_bufchan_buf[0]))
        m3a86_1_bufchan_buf <= {16'd0, 1'd0};
      else if (((! m3a86_1_argbuf_r) && (! m3a86_1_bufchan_buf[0])))
        m3a86_1_bufchan_buf <= m3a86_1_bufchan_d;
  
  /* fork (Ty Pointer_QTree_Bool) : (m3a86_goMux_mux,Pointer_QTree_Bool) > [(m3a86_1,Pointer_QTree_Bool),
                                                                       (m3a86_2,Pointer_QTree_Bool)] */
  logic [1:0] m3a86_goMux_mux_emitted;
  logic [1:0] m3a86_goMux_mux_done;
  assign m3a86_1_d = {m3a86_goMux_mux_d[16:1],
                      (m3a86_goMux_mux_d[0] && (! m3a86_goMux_mux_emitted[0]))};
  assign m3a86_2_d = {m3a86_goMux_mux_d[16:1],
                      (m3a86_goMux_mux_d[0] && (! m3a86_goMux_mux_emitted[1]))};
  assign m3a86_goMux_mux_done = (m3a86_goMux_mux_emitted | ({m3a86_2_d[0],
                                                             m3a86_1_d[0]} & {m3a86_2_r,
                                                                              m3a86_1_r}));
  assign m3a86_goMux_mux_r = (& m3a86_goMux_mux_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m3a86_goMux_mux_emitted <= 2'd0;
    else
      m3a86_goMux_mux_emitted <= (m3a86_goMux_mux_r ? 2'd0 :
                                  m3a86_goMux_mux_done);
  
  /* buf (Ty Pointer_QTree_Bool) : (q1a8H_3_destruct,Pointer_QTree_Bool) > (q1a8H_3_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t q1a8H_3_destruct_bufchan_d;
  logic q1a8H_3_destruct_bufchan_r;
  assign q1a8H_3_destruct_r = ((! q1a8H_3_destruct_bufchan_d[0]) || q1a8H_3_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q1a8H_3_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q1a8H_3_destruct_r)
        q1a8H_3_destruct_bufchan_d <= q1a8H_3_destruct_d;
  Pointer_QTree_Bool_t q1a8H_3_destruct_bufchan_buf;
  assign q1a8H_3_destruct_bufchan_r = (! q1a8H_3_destruct_bufchan_buf[0]);
  assign q1a8H_3_1_argbuf_d = (q1a8H_3_destruct_bufchan_buf[0] ? q1a8H_3_destruct_bufchan_buf :
                               q1a8H_3_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q1a8H_3_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q1a8H_3_1_argbuf_r && q1a8H_3_destruct_bufchan_buf[0]))
        q1a8H_3_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q1a8H_3_1_argbuf_r) && (! q1a8H_3_destruct_bufchan_buf[0])))
        q1a8H_3_destruct_bufchan_buf <= q1a8H_3_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (q1a98_3_destruct,Pointer_QTree_Bool) > (q1a98_3_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t q1a98_3_destruct_bufchan_d;
  logic q1a98_3_destruct_bufchan_r;
  assign q1a98_3_destruct_r = ((! q1a98_3_destruct_bufchan_d[0]) || q1a98_3_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q1a98_3_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q1a98_3_destruct_r)
        q1a98_3_destruct_bufchan_d <= q1a98_3_destruct_d;
  Pointer_QTree_Bool_t q1a98_3_destruct_bufchan_buf;
  assign q1a98_3_destruct_bufchan_r = (! q1a98_3_destruct_bufchan_buf[0]);
  assign q1a98_3_1_argbuf_d = (q1a98_3_destruct_bufchan_buf[0] ? q1a98_3_destruct_bufchan_buf :
                               q1a98_3_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q1a98_3_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q1a98_3_1_argbuf_r && q1a98_3_destruct_bufchan_buf[0]))
        q1a98_3_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q1a98_3_1_argbuf_r) && (! q1a98_3_destruct_bufchan_buf[0])))
        q1a98_3_destruct_bufchan_buf <= q1a98_3_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (q2a8I_2_destruct,Pointer_QTree_Bool) > (q2a8I_2_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t q2a8I_2_destruct_bufchan_d;
  logic q2a8I_2_destruct_bufchan_r;
  assign q2a8I_2_destruct_r = ((! q2a8I_2_destruct_bufchan_d[0]) || q2a8I_2_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q2a8I_2_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q2a8I_2_destruct_r)
        q2a8I_2_destruct_bufchan_d <= q2a8I_2_destruct_d;
  Pointer_QTree_Bool_t q2a8I_2_destruct_bufchan_buf;
  assign q2a8I_2_destruct_bufchan_r = (! q2a8I_2_destruct_bufchan_buf[0]);
  assign q2a8I_2_1_argbuf_d = (q2a8I_2_destruct_bufchan_buf[0] ? q2a8I_2_destruct_bufchan_buf :
                               q2a8I_2_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q2a8I_2_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q2a8I_2_1_argbuf_r && q2a8I_2_destruct_bufchan_buf[0]))
        q2a8I_2_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q2a8I_2_1_argbuf_r) && (! q2a8I_2_destruct_bufchan_buf[0])))
        q2a8I_2_destruct_bufchan_buf <= q2a8I_2_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (q2a99_2_destruct,Pointer_QTree_Bool) > (q2a99_2_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t q2a99_2_destruct_bufchan_d;
  logic q2a99_2_destruct_bufchan_r;
  assign q2a99_2_destruct_r = ((! q2a99_2_destruct_bufchan_d[0]) || q2a99_2_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q2a99_2_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q2a99_2_destruct_r)
        q2a99_2_destruct_bufchan_d <= q2a99_2_destruct_d;
  Pointer_QTree_Bool_t q2a99_2_destruct_bufchan_buf;
  assign q2a99_2_destruct_bufchan_r = (! q2a99_2_destruct_bufchan_buf[0]);
  assign q2a99_2_1_argbuf_d = (q2a99_2_destruct_bufchan_buf[0] ? q2a99_2_destruct_bufchan_buf :
                               q2a99_2_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q2a99_2_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q2a99_2_1_argbuf_r && q2a99_2_destruct_bufchan_buf[0]))
        q2a99_2_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q2a99_2_1_argbuf_r) && (! q2a99_2_destruct_bufchan_buf[0])))
        q2a99_2_destruct_bufchan_buf <= q2a99_2_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (q3a8J_1_destruct,Pointer_QTree_Bool) > (q3a8J_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t q3a8J_1_destruct_bufchan_d;
  logic q3a8J_1_destruct_bufchan_r;
  assign q3a8J_1_destruct_r = ((! q3a8J_1_destruct_bufchan_d[0]) || q3a8J_1_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q3a8J_1_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q3a8J_1_destruct_r)
        q3a8J_1_destruct_bufchan_d <= q3a8J_1_destruct_d;
  Pointer_QTree_Bool_t q3a8J_1_destruct_bufchan_buf;
  assign q3a8J_1_destruct_bufchan_r = (! q3a8J_1_destruct_bufchan_buf[0]);
  assign q3a8J_1_1_argbuf_d = (q3a8J_1_destruct_bufchan_buf[0] ? q3a8J_1_destruct_bufchan_buf :
                               q3a8J_1_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q3a8J_1_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q3a8J_1_1_argbuf_r && q3a8J_1_destruct_bufchan_buf[0]))
        q3a8J_1_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q3a8J_1_1_argbuf_r) && (! q3a8J_1_destruct_bufchan_buf[0])))
        q3a8J_1_destruct_bufchan_buf <= q3a8J_1_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (q3a9a_1_destruct,Pointer_QTree_Bool) > (q3a9a_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t q3a9a_1_destruct_bufchan_d;
  logic q3a9a_1_destruct_bufchan_r;
  assign q3a9a_1_destruct_r = ((! q3a9a_1_destruct_bufchan_d[0]) || q3a9a_1_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q3a9a_1_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q3a9a_1_destruct_r)
        q3a9a_1_destruct_bufchan_d <= q3a9a_1_destruct_d;
  Pointer_QTree_Bool_t q3a9a_1_destruct_bufchan_buf;
  assign q3a9a_1_destruct_bufchan_r = (! q3a9a_1_destruct_bufchan_buf[0]);
  assign q3a9a_1_1_argbuf_d = (q3a9a_1_destruct_bufchan_buf[0] ? q3a9a_1_destruct_bufchan_buf :
                               q3a9a_1_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q3a9a_1_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q3a9a_1_1_argbuf_r && q3a9a_1_destruct_bufchan_buf[0]))
        q3a9a_1_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q3a9a_1_1_argbuf_r) && (! q3a9a_1_destruct_bufchan_buf[0])))
        q3a9a_1_destruct_bufchan_buf <= q3a9a_1_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (q4a90_1,Pointer_QTree_Bool) > (q4a90_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t q4a90_1_bufchan_d;
  logic q4a90_1_bufchan_r;
  assign q4a90_1_r = ((! q4a90_1_bufchan_d[0]) || q4a90_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q4a90_1_bufchan_d <= {16'd0, 1'd0};
    else if (q4a90_1_r) q4a90_1_bufchan_d <= q4a90_1_d;
  Pointer_QTree_Bool_t q4a90_1_bufchan_buf;
  assign q4a90_1_bufchan_r = (! q4a90_1_bufchan_buf[0]);
  assign q4a90_1_argbuf_d = (q4a90_1_bufchan_buf[0] ? q4a90_1_bufchan_buf :
                             q4a90_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q4a90_1_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q4a90_1_argbuf_r && q4a90_1_bufchan_buf[0]))
        q4a90_1_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q4a90_1_argbuf_r) && (! q4a90_1_bufchan_buf[0])))
        q4a90_1_bufchan_buf <= q4a90_1_bufchan_d;
  
  /* fork (Ty Pointer_QTree_Bool) : (q4a90_goMux_mux,Pointer_QTree_Bool) > [(q4a90_1,Pointer_QTree_Bool),
                                                                       (q4a90_2,Pointer_QTree_Bool)] */
  logic [1:0] q4a90_goMux_mux_emitted;
  logic [1:0] q4a90_goMux_mux_done;
  assign q4a90_1_d = {q4a90_goMux_mux_d[16:1],
                      (q4a90_goMux_mux_d[0] && (! q4a90_goMux_mux_emitted[0]))};
  assign q4a90_2_d = {q4a90_goMux_mux_d[16:1],
                      (q4a90_goMux_mux_d[0] && (! q4a90_goMux_mux_emitted[1]))};
  assign q4a90_goMux_mux_done = (q4a90_goMux_mux_emitted | ({q4a90_2_d[0],
                                                             q4a90_1_d[0]} & {q4a90_2_r,
                                                                              q4a90_1_r}));
  assign q4a90_goMux_mux_r = (& q4a90_goMux_mux_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q4a90_goMux_mux_emitted <= 2'd0;
    else
      q4a90_goMux_mux_emitted <= (q4a90_goMux_mux_r ? 2'd0 :
                                  q4a90_goMux_mux_done);
  
  /* buf (Ty CTf'''''''''''') : (readPointer_CTf''''''''''''scfarg_0_1_1_argbuf,CTf'''''''''''') > (readPointer_CTf''''''''''''scfarg_0_1_1_argbuf_rwb,CTf'''''''''''') */
  \CTf''''''''''''_t  \readPointer_CTf''''''''''''scfarg_0_1_1_argbuf_bufchan_d ;
  logic \readPointer_CTf''''''''''''scfarg_0_1_1_argbuf_bufchan_r ;
  assign \readPointer_CTf''''''''''''scfarg_0_1_1_argbuf_r  = ((! \readPointer_CTf''''''''''''scfarg_0_1_1_argbuf_bufchan_d [0]) || \readPointer_CTf''''''''''''scfarg_0_1_1_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \readPointer_CTf''''''''''''scfarg_0_1_1_argbuf_bufchan_d  <= {115'd0,
                                                                     1'd0};
    else
      if (\readPointer_CTf''''''''''''scfarg_0_1_1_argbuf_r )
        \readPointer_CTf''''''''''''scfarg_0_1_1_argbuf_bufchan_d  <= \readPointer_CTf''''''''''''scfarg_0_1_1_argbuf_d ;
  \CTf''''''''''''_t  \readPointer_CTf''''''''''''scfarg_0_1_1_argbuf_bufchan_buf ;
  assign \readPointer_CTf''''''''''''scfarg_0_1_1_argbuf_bufchan_r  = (! \readPointer_CTf''''''''''''scfarg_0_1_1_argbuf_bufchan_buf [0]);
  assign \readPointer_CTf''''''''''''scfarg_0_1_1_argbuf_rwb_d  = (\readPointer_CTf''''''''''''scfarg_0_1_1_argbuf_bufchan_buf [0] ? \readPointer_CTf''''''''''''scfarg_0_1_1_argbuf_bufchan_buf  :
                                                                   \readPointer_CTf''''''''''''scfarg_0_1_1_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \readPointer_CTf''''''''''''scfarg_0_1_1_argbuf_bufchan_buf  <= {115'd0,
                                                                       1'd0};
    else
      if ((\readPointer_CTf''''''''''''scfarg_0_1_1_argbuf_rwb_r  && \readPointer_CTf''''''''''''scfarg_0_1_1_argbuf_bufchan_buf [0]))
        \readPointer_CTf''''''''''''scfarg_0_1_1_argbuf_bufchan_buf  <= {115'd0,
                                                                         1'd0};
      else if (((! \readPointer_CTf''''''''''''scfarg_0_1_1_argbuf_rwb_r ) && (! \readPointer_CTf''''''''''''scfarg_0_1_1_argbuf_bufchan_buf [0])))
        \readPointer_CTf''''''''''''scfarg_0_1_1_argbuf_bufchan_buf  <= \readPointer_CTf''''''''''''scfarg_0_1_1_argbuf_bufchan_d ;
  
  /* fork (Ty CTf'''''''''''') : (readPointer_CTf''''''''''''scfarg_0_1_1_argbuf_rwb,CTf'''''''''''') > [(lizzieLet65_1,CTf''''''''''''),
                                                                                                    (lizzieLet65_2,CTf''''''''''''),
                                                                                                    (lizzieLet65_3,CTf''''''''''''),
                                                                                                    (lizzieLet65_4,CTf'''''''''''')] */
  logic [3:0] \readPointer_CTf''''''''''''scfarg_0_1_1_argbuf_rwb_emitted ;
  logic [3:0] \readPointer_CTf''''''''''''scfarg_0_1_1_argbuf_rwb_done ;
  assign lizzieLet65_1_d = {\readPointer_CTf''''''''''''scfarg_0_1_1_argbuf_rwb_d [115:1],
                            (\readPointer_CTf''''''''''''scfarg_0_1_1_argbuf_rwb_d [0] && (! \readPointer_CTf''''''''''''scfarg_0_1_1_argbuf_rwb_emitted [0]))};
  assign lizzieLet65_2_d = {\readPointer_CTf''''''''''''scfarg_0_1_1_argbuf_rwb_d [115:1],
                            (\readPointer_CTf''''''''''''scfarg_0_1_1_argbuf_rwb_d [0] && (! \readPointer_CTf''''''''''''scfarg_0_1_1_argbuf_rwb_emitted [1]))};
  assign lizzieLet65_3_d = {\readPointer_CTf''''''''''''scfarg_0_1_1_argbuf_rwb_d [115:1],
                            (\readPointer_CTf''''''''''''scfarg_0_1_1_argbuf_rwb_d [0] && (! \readPointer_CTf''''''''''''scfarg_0_1_1_argbuf_rwb_emitted [2]))};
  assign lizzieLet65_4_d = {\readPointer_CTf''''''''''''scfarg_0_1_1_argbuf_rwb_d [115:1],
                            (\readPointer_CTf''''''''''''scfarg_0_1_1_argbuf_rwb_d [0] && (! \readPointer_CTf''''''''''''scfarg_0_1_1_argbuf_rwb_emitted [3]))};
  assign \readPointer_CTf''''''''''''scfarg_0_1_1_argbuf_rwb_done  = (\readPointer_CTf''''''''''''scfarg_0_1_1_argbuf_rwb_emitted  | ({lizzieLet65_4_d[0],
                                                                                                                                       lizzieLet65_3_d[0],
                                                                                                                                       lizzieLet65_2_d[0],
                                                                                                                                       lizzieLet65_1_d[0]} & {lizzieLet65_4_r,
                                                                                                                                                              lizzieLet65_3_r,
                                                                                                                                                              lizzieLet65_2_r,
                                                                                                                                                              lizzieLet65_1_r}));
  assign \readPointer_CTf''''''''''''scfarg_0_1_1_argbuf_rwb_r  = (& \readPointer_CTf''''''''''''scfarg_0_1_1_argbuf_rwb_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \readPointer_CTf''''''''''''scfarg_0_1_1_argbuf_rwb_emitted  <= 4'd0;
    else
      \readPointer_CTf''''''''''''scfarg_0_1_1_argbuf_rwb_emitted  <= (\readPointer_CTf''''''''''''scfarg_0_1_1_argbuf_rwb_r  ? 4'd0 :
                                                                       \readPointer_CTf''''''''''''scfarg_0_1_1_argbuf_rwb_done );
  
  /* buf (Ty CTf) : (readPointer_CTfscfarg_0_1_argbuf,CTf) > (readPointer_CTfscfarg_0_1_argbuf_rwb,CTf) */
  CTf_t readPointer_CTfscfarg_0_1_argbuf_bufchan_d;
  logic readPointer_CTfscfarg_0_1_argbuf_bufchan_r;
  assign readPointer_CTfscfarg_0_1_argbuf_r = ((! readPointer_CTfscfarg_0_1_argbuf_bufchan_d[0]) || readPointer_CTfscfarg_0_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_CTfscfarg_0_1_argbuf_bufchan_d <= {163'd0, 1'd0};
    else
      if (readPointer_CTfscfarg_0_1_argbuf_r)
        readPointer_CTfscfarg_0_1_argbuf_bufchan_d <= readPointer_CTfscfarg_0_1_argbuf_d;
  CTf_t readPointer_CTfscfarg_0_1_argbuf_bufchan_buf;
  assign readPointer_CTfscfarg_0_1_argbuf_bufchan_r = (! readPointer_CTfscfarg_0_1_argbuf_bufchan_buf[0]);
  assign readPointer_CTfscfarg_0_1_argbuf_rwb_d = (readPointer_CTfscfarg_0_1_argbuf_bufchan_buf[0] ? readPointer_CTfscfarg_0_1_argbuf_bufchan_buf :
                                                   readPointer_CTfscfarg_0_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_CTfscfarg_0_1_argbuf_bufchan_buf <= {163'd0, 1'd0};
    else
      if ((readPointer_CTfscfarg_0_1_argbuf_rwb_r && readPointer_CTfscfarg_0_1_argbuf_bufchan_buf[0]))
        readPointer_CTfscfarg_0_1_argbuf_bufchan_buf <= {163'd0, 1'd0};
      else if (((! readPointer_CTfscfarg_0_1_argbuf_rwb_r) && (! readPointer_CTfscfarg_0_1_argbuf_bufchan_buf[0])))
        readPointer_CTfscfarg_0_1_argbuf_bufchan_buf <= readPointer_CTfscfarg_0_1_argbuf_bufchan_d;
  
  /* fork (Ty CTf) : (readPointer_CTfscfarg_0_1_argbuf_rwb,CTf) > [(lizzieLet60_1,CTf),
                                                              (lizzieLet60_2,CTf),
                                                              (lizzieLet60_3,CTf),
                                                              (lizzieLet60_4,CTf)] */
  logic [3:0] readPointer_CTfscfarg_0_1_argbuf_rwb_emitted;
  logic [3:0] readPointer_CTfscfarg_0_1_argbuf_rwb_done;
  assign lizzieLet60_1_d = {readPointer_CTfscfarg_0_1_argbuf_rwb_d[163:1],
                            (readPointer_CTfscfarg_0_1_argbuf_rwb_d[0] && (! readPointer_CTfscfarg_0_1_argbuf_rwb_emitted[0]))};
  assign lizzieLet60_2_d = {readPointer_CTfscfarg_0_1_argbuf_rwb_d[163:1],
                            (readPointer_CTfscfarg_0_1_argbuf_rwb_d[0] && (! readPointer_CTfscfarg_0_1_argbuf_rwb_emitted[1]))};
  assign lizzieLet60_3_d = {readPointer_CTfscfarg_0_1_argbuf_rwb_d[163:1],
                            (readPointer_CTfscfarg_0_1_argbuf_rwb_d[0] && (! readPointer_CTfscfarg_0_1_argbuf_rwb_emitted[2]))};
  assign lizzieLet60_4_d = {readPointer_CTfscfarg_0_1_argbuf_rwb_d[163:1],
                            (readPointer_CTfscfarg_0_1_argbuf_rwb_d[0] && (! readPointer_CTfscfarg_0_1_argbuf_rwb_emitted[3]))};
  assign readPointer_CTfscfarg_0_1_argbuf_rwb_done = (readPointer_CTfscfarg_0_1_argbuf_rwb_emitted | ({lizzieLet60_4_d[0],
                                                                                                       lizzieLet60_3_d[0],
                                                                                                       lizzieLet60_2_d[0],
                                                                                                       lizzieLet60_1_d[0]} & {lizzieLet60_4_r,
                                                                                                                              lizzieLet60_3_r,
                                                                                                                              lizzieLet60_2_r,
                                                                                                                              lizzieLet60_1_r}));
  assign readPointer_CTfscfarg_0_1_argbuf_rwb_r = (& readPointer_CTfscfarg_0_1_argbuf_rwb_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_CTfscfarg_0_1_argbuf_rwb_emitted <= 4'd0;
    else
      readPointer_CTfscfarg_0_1_argbuf_rwb_emitted <= (readPointer_CTfscfarg_0_1_argbuf_rwb_r ? 4'd0 :
                                                       readPointer_CTfscfarg_0_1_argbuf_rwb_done);
  
  /* buf (Ty QTree_Bool) : (readPointer_QTree_Boolm1a84_1_argbuf,QTree_Bool) > (readPointer_QTree_Boolm1a84_1_argbuf_rwb,QTree_Bool) */
  QTree_Bool_t readPointer_QTree_Boolm1a84_1_argbuf_bufchan_d;
  logic readPointer_QTree_Boolm1a84_1_argbuf_bufchan_r;
  assign readPointer_QTree_Boolm1a84_1_argbuf_r = ((! readPointer_QTree_Boolm1a84_1_argbuf_bufchan_d[0]) || readPointer_QTree_Boolm1a84_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Boolm1a84_1_argbuf_bufchan_d <= {66'd0, 1'd0};
    else
      if (readPointer_QTree_Boolm1a84_1_argbuf_r)
        readPointer_QTree_Boolm1a84_1_argbuf_bufchan_d <= readPointer_QTree_Boolm1a84_1_argbuf_d;
  QTree_Bool_t readPointer_QTree_Boolm1a84_1_argbuf_bufchan_buf;
  assign readPointer_QTree_Boolm1a84_1_argbuf_bufchan_r = (! readPointer_QTree_Boolm1a84_1_argbuf_bufchan_buf[0]);
  assign readPointer_QTree_Boolm1a84_1_argbuf_rwb_d = (readPointer_QTree_Boolm1a84_1_argbuf_bufchan_buf[0] ? readPointer_QTree_Boolm1a84_1_argbuf_bufchan_buf :
                                                       readPointer_QTree_Boolm1a84_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Boolm1a84_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((readPointer_QTree_Boolm1a84_1_argbuf_rwb_r && readPointer_QTree_Boolm1a84_1_argbuf_bufchan_buf[0]))
        readPointer_QTree_Boolm1a84_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
      else if (((! readPointer_QTree_Boolm1a84_1_argbuf_rwb_r) && (! readPointer_QTree_Boolm1a84_1_argbuf_bufchan_buf[0])))
        readPointer_QTree_Boolm1a84_1_argbuf_bufchan_buf <= readPointer_QTree_Boolm1a84_1_argbuf_bufchan_d;
  
  /* fork (Ty QTree_Bool) : (readPointer_QTree_Boolm1a84_1_argbuf_rwb,QTree_Bool) > [(lizzieLet0_1,QTree_Bool),
                                                                                (lizzieLet0_2,QTree_Bool),
                                                                                (lizzieLet0_3,QTree_Bool),
                                                                                (lizzieLet0_4,QTree_Bool),
                                                                                (lizzieLet0_5,QTree_Bool),
                                                                                (lizzieLet0_6,QTree_Bool),
                                                                                (lizzieLet0_7,QTree_Bool),
                                                                                (lizzieLet0_8,QTree_Bool),
                                                                                (lizzieLet0_9,QTree_Bool)] */
  logic [8:0] readPointer_QTree_Boolm1a84_1_argbuf_rwb_emitted;
  logic [8:0] readPointer_QTree_Boolm1a84_1_argbuf_rwb_done;
  assign lizzieLet0_1_d = {readPointer_QTree_Boolm1a84_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_Boolm1a84_1_argbuf_rwb_d[0] && (! readPointer_QTree_Boolm1a84_1_argbuf_rwb_emitted[0]))};
  assign lizzieLet0_2_d = {readPointer_QTree_Boolm1a84_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_Boolm1a84_1_argbuf_rwb_d[0] && (! readPointer_QTree_Boolm1a84_1_argbuf_rwb_emitted[1]))};
  assign lizzieLet0_3_d = {readPointer_QTree_Boolm1a84_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_Boolm1a84_1_argbuf_rwb_d[0] && (! readPointer_QTree_Boolm1a84_1_argbuf_rwb_emitted[2]))};
  assign lizzieLet0_4_d = {readPointer_QTree_Boolm1a84_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_Boolm1a84_1_argbuf_rwb_d[0] && (! readPointer_QTree_Boolm1a84_1_argbuf_rwb_emitted[3]))};
  assign lizzieLet0_5_d = {readPointer_QTree_Boolm1a84_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_Boolm1a84_1_argbuf_rwb_d[0] && (! readPointer_QTree_Boolm1a84_1_argbuf_rwb_emitted[4]))};
  assign lizzieLet0_6_d = {readPointer_QTree_Boolm1a84_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_Boolm1a84_1_argbuf_rwb_d[0] && (! readPointer_QTree_Boolm1a84_1_argbuf_rwb_emitted[5]))};
  assign lizzieLet0_7_d = {readPointer_QTree_Boolm1a84_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_Boolm1a84_1_argbuf_rwb_d[0] && (! readPointer_QTree_Boolm1a84_1_argbuf_rwb_emitted[6]))};
  assign lizzieLet0_8_d = {readPointer_QTree_Boolm1a84_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_Boolm1a84_1_argbuf_rwb_d[0] && (! readPointer_QTree_Boolm1a84_1_argbuf_rwb_emitted[7]))};
  assign lizzieLet0_9_d = {readPointer_QTree_Boolm1a84_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_Boolm1a84_1_argbuf_rwb_d[0] && (! readPointer_QTree_Boolm1a84_1_argbuf_rwb_emitted[8]))};
  assign readPointer_QTree_Boolm1a84_1_argbuf_rwb_done = (readPointer_QTree_Boolm1a84_1_argbuf_rwb_emitted | ({lizzieLet0_9_d[0],
                                                                                                               lizzieLet0_8_d[0],
                                                                                                               lizzieLet0_7_d[0],
                                                                                                               lizzieLet0_6_d[0],
                                                                                                               lizzieLet0_5_d[0],
                                                                                                               lizzieLet0_4_d[0],
                                                                                                               lizzieLet0_3_d[0],
                                                                                                               lizzieLet0_2_d[0],
                                                                                                               lizzieLet0_1_d[0]} & {lizzieLet0_9_r,
                                                                                                                                     lizzieLet0_8_r,
                                                                                                                                     lizzieLet0_7_r,
                                                                                                                                     lizzieLet0_6_r,
                                                                                                                                     lizzieLet0_5_r,
                                                                                                                                     lizzieLet0_4_r,
                                                                                                                                     lizzieLet0_3_r,
                                                                                                                                     lizzieLet0_2_r,
                                                                                                                                     lizzieLet0_1_r}));
  assign readPointer_QTree_Boolm1a84_1_argbuf_rwb_r = (& readPointer_QTree_Boolm1a84_1_argbuf_rwb_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Boolm1a84_1_argbuf_rwb_emitted <= 9'd0;
    else
      readPointer_QTree_Boolm1a84_1_argbuf_rwb_emitted <= (readPointer_QTree_Boolm1a84_1_argbuf_rwb_r ? 9'd0 :
                                                           readPointer_QTree_Boolm1a84_1_argbuf_rwb_done);
  
  /* buf (Ty QTree_Bool) : (readPointer_QTree_Boolm2a85_1_argbuf,QTree_Bool) > (readPointer_QTree_Boolm2a85_1_argbuf_rwb,QTree_Bool) */
  QTree_Bool_t readPointer_QTree_Boolm2a85_1_argbuf_bufchan_d;
  logic readPointer_QTree_Boolm2a85_1_argbuf_bufchan_r;
  assign readPointer_QTree_Boolm2a85_1_argbuf_r = ((! readPointer_QTree_Boolm2a85_1_argbuf_bufchan_d[0]) || readPointer_QTree_Boolm2a85_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Boolm2a85_1_argbuf_bufchan_d <= {66'd0, 1'd0};
    else
      if (readPointer_QTree_Boolm2a85_1_argbuf_r)
        readPointer_QTree_Boolm2a85_1_argbuf_bufchan_d <= readPointer_QTree_Boolm2a85_1_argbuf_d;
  QTree_Bool_t readPointer_QTree_Boolm2a85_1_argbuf_bufchan_buf;
  assign readPointer_QTree_Boolm2a85_1_argbuf_bufchan_r = (! readPointer_QTree_Boolm2a85_1_argbuf_bufchan_buf[0]);
  assign readPointer_QTree_Boolm2a85_1_argbuf_rwb_d = (readPointer_QTree_Boolm2a85_1_argbuf_bufchan_buf[0] ? readPointer_QTree_Boolm2a85_1_argbuf_bufchan_buf :
                                                       readPointer_QTree_Boolm2a85_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Boolm2a85_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((readPointer_QTree_Boolm2a85_1_argbuf_rwb_r && readPointer_QTree_Boolm2a85_1_argbuf_bufchan_buf[0]))
        readPointer_QTree_Boolm2a85_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
      else if (((! readPointer_QTree_Boolm2a85_1_argbuf_rwb_r) && (! readPointer_QTree_Boolm2a85_1_argbuf_bufchan_buf[0])))
        readPointer_QTree_Boolm2a85_1_argbuf_bufchan_buf <= readPointer_QTree_Boolm2a85_1_argbuf_bufchan_d;
  
  /* buf (Ty QTree_Bool) : (readPointer_QTree_Boolm3a86_1_argbuf,QTree_Bool) > (readPointer_QTree_Boolm3a86_1_argbuf_rwb,QTree_Bool) */
  QTree_Bool_t readPointer_QTree_Boolm3a86_1_argbuf_bufchan_d;
  logic readPointer_QTree_Boolm3a86_1_argbuf_bufchan_r;
  assign readPointer_QTree_Boolm3a86_1_argbuf_r = ((! readPointer_QTree_Boolm3a86_1_argbuf_bufchan_d[0]) || readPointer_QTree_Boolm3a86_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Boolm3a86_1_argbuf_bufchan_d <= {66'd0, 1'd0};
    else
      if (readPointer_QTree_Boolm3a86_1_argbuf_r)
        readPointer_QTree_Boolm3a86_1_argbuf_bufchan_d <= readPointer_QTree_Boolm3a86_1_argbuf_d;
  QTree_Bool_t readPointer_QTree_Boolm3a86_1_argbuf_bufchan_buf;
  assign readPointer_QTree_Boolm3a86_1_argbuf_bufchan_r = (! readPointer_QTree_Boolm3a86_1_argbuf_bufchan_buf[0]);
  assign readPointer_QTree_Boolm3a86_1_argbuf_rwb_d = (readPointer_QTree_Boolm3a86_1_argbuf_bufchan_buf[0] ? readPointer_QTree_Boolm3a86_1_argbuf_bufchan_buf :
                                                       readPointer_QTree_Boolm3a86_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Boolm3a86_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((readPointer_QTree_Boolm3a86_1_argbuf_rwb_r && readPointer_QTree_Boolm3a86_1_argbuf_bufchan_buf[0]))
        readPointer_QTree_Boolm3a86_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
      else if (((! readPointer_QTree_Boolm3a86_1_argbuf_rwb_r) && (! readPointer_QTree_Boolm3a86_1_argbuf_bufchan_buf[0])))
        readPointer_QTree_Boolm3a86_1_argbuf_bufchan_buf <= readPointer_QTree_Boolm3a86_1_argbuf_bufchan_d;
  
  /* buf (Ty QTree_Bool) : (readPointer_QTree_Boolq4a90_1_argbuf,QTree_Bool) > (readPointer_QTree_Boolq4a90_1_argbuf_rwb,QTree_Bool) */
  QTree_Bool_t readPointer_QTree_Boolq4a90_1_argbuf_bufchan_d;
  logic readPointer_QTree_Boolq4a90_1_argbuf_bufchan_r;
  assign readPointer_QTree_Boolq4a90_1_argbuf_r = ((! readPointer_QTree_Boolq4a90_1_argbuf_bufchan_d[0]) || readPointer_QTree_Boolq4a90_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Boolq4a90_1_argbuf_bufchan_d <= {66'd0, 1'd0};
    else
      if (readPointer_QTree_Boolq4a90_1_argbuf_r)
        readPointer_QTree_Boolq4a90_1_argbuf_bufchan_d <= readPointer_QTree_Boolq4a90_1_argbuf_d;
  QTree_Bool_t readPointer_QTree_Boolq4a90_1_argbuf_bufchan_buf;
  assign readPointer_QTree_Boolq4a90_1_argbuf_bufchan_r = (! readPointer_QTree_Boolq4a90_1_argbuf_bufchan_buf[0]);
  assign readPointer_QTree_Boolq4a90_1_argbuf_rwb_d = (readPointer_QTree_Boolq4a90_1_argbuf_bufchan_buf[0] ? readPointer_QTree_Boolq4a90_1_argbuf_bufchan_buf :
                                                       readPointer_QTree_Boolq4a90_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Boolq4a90_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((readPointer_QTree_Boolq4a90_1_argbuf_rwb_r && readPointer_QTree_Boolq4a90_1_argbuf_bufchan_buf[0]))
        readPointer_QTree_Boolq4a90_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
      else if (((! readPointer_QTree_Boolq4a90_1_argbuf_rwb_r) && (! readPointer_QTree_Boolq4a90_1_argbuf_bufchan_buf[0])))
        readPointer_QTree_Boolq4a90_1_argbuf_bufchan_buf <= readPointer_QTree_Boolq4a90_1_argbuf_bufchan_d;
  
  /* fork (Ty QTree_Bool) : (readPointer_QTree_Boolq4a90_1_argbuf_rwb,QTree_Bool) > [(lizzieLet45_1,QTree_Bool),
                                                                                (lizzieLet45_2,QTree_Bool),
                                                                                (lizzieLet45_3,QTree_Bool),
                                                                                (lizzieLet45_4,QTree_Bool),
                                                                                (lizzieLet45_5,QTree_Bool),
                                                                                (lizzieLet45_6,QTree_Bool),
                                                                                (lizzieLet45_7,QTree_Bool)] */
  logic [6:0] readPointer_QTree_Boolq4a90_1_argbuf_rwb_emitted;
  logic [6:0] readPointer_QTree_Boolq4a90_1_argbuf_rwb_done;
  assign lizzieLet45_1_d = {readPointer_QTree_Boolq4a90_1_argbuf_rwb_d[66:1],
                            (readPointer_QTree_Boolq4a90_1_argbuf_rwb_d[0] && (! readPointer_QTree_Boolq4a90_1_argbuf_rwb_emitted[0]))};
  assign lizzieLet45_2_d = {readPointer_QTree_Boolq4a90_1_argbuf_rwb_d[66:1],
                            (readPointer_QTree_Boolq4a90_1_argbuf_rwb_d[0] && (! readPointer_QTree_Boolq4a90_1_argbuf_rwb_emitted[1]))};
  assign lizzieLet45_3_d = {readPointer_QTree_Boolq4a90_1_argbuf_rwb_d[66:1],
                            (readPointer_QTree_Boolq4a90_1_argbuf_rwb_d[0] && (! readPointer_QTree_Boolq4a90_1_argbuf_rwb_emitted[2]))};
  assign lizzieLet45_4_d = {readPointer_QTree_Boolq4a90_1_argbuf_rwb_d[66:1],
                            (readPointer_QTree_Boolq4a90_1_argbuf_rwb_d[0] && (! readPointer_QTree_Boolq4a90_1_argbuf_rwb_emitted[3]))};
  assign lizzieLet45_5_d = {readPointer_QTree_Boolq4a90_1_argbuf_rwb_d[66:1],
                            (readPointer_QTree_Boolq4a90_1_argbuf_rwb_d[0] && (! readPointer_QTree_Boolq4a90_1_argbuf_rwb_emitted[4]))};
  assign lizzieLet45_6_d = {readPointer_QTree_Boolq4a90_1_argbuf_rwb_d[66:1],
                            (readPointer_QTree_Boolq4a90_1_argbuf_rwb_d[0] && (! readPointer_QTree_Boolq4a90_1_argbuf_rwb_emitted[5]))};
  assign lizzieLet45_7_d = {readPointer_QTree_Boolq4a90_1_argbuf_rwb_d[66:1],
                            (readPointer_QTree_Boolq4a90_1_argbuf_rwb_d[0] && (! readPointer_QTree_Boolq4a90_1_argbuf_rwb_emitted[6]))};
  assign readPointer_QTree_Boolq4a90_1_argbuf_rwb_done = (readPointer_QTree_Boolq4a90_1_argbuf_rwb_emitted | ({lizzieLet45_7_d[0],
                                                                                                               lizzieLet45_6_d[0],
                                                                                                               lizzieLet45_5_d[0],
                                                                                                               lizzieLet45_4_d[0],
                                                                                                               lizzieLet45_3_d[0],
                                                                                                               lizzieLet45_2_d[0],
                                                                                                               lizzieLet45_1_d[0]} & {lizzieLet45_7_r,
                                                                                                                                      lizzieLet45_6_r,
                                                                                                                                      lizzieLet45_5_r,
                                                                                                                                      lizzieLet45_4_r,
                                                                                                                                      lizzieLet45_3_r,
                                                                                                                                      lizzieLet45_2_r,
                                                                                                                                      lizzieLet45_1_r}));
  assign readPointer_QTree_Boolq4a90_1_argbuf_rwb_r = (& readPointer_QTree_Boolq4a90_1_argbuf_rwb_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Boolq4a90_1_argbuf_rwb_emitted <= 7'd0;
    else
      readPointer_QTree_Boolq4a90_1_argbuf_rwb_emitted <= (readPointer_QTree_Boolq4a90_1_argbuf_rwb_r ? 7'd0 :
                                                           readPointer_QTree_Boolq4a90_1_argbuf_rwb_done);
  
  /* buf (Ty QTree_Bool) : (readPointer_QTree_Boolt4a91_1_argbuf,QTree_Bool) > (readPointer_QTree_Boolt4a91_1_argbuf_rwb,QTree_Bool) */
  QTree_Bool_t readPointer_QTree_Boolt4a91_1_argbuf_bufchan_d;
  logic readPointer_QTree_Boolt4a91_1_argbuf_bufchan_r;
  assign readPointer_QTree_Boolt4a91_1_argbuf_r = ((! readPointer_QTree_Boolt4a91_1_argbuf_bufchan_d[0]) || readPointer_QTree_Boolt4a91_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Boolt4a91_1_argbuf_bufchan_d <= {66'd0, 1'd0};
    else
      if (readPointer_QTree_Boolt4a91_1_argbuf_r)
        readPointer_QTree_Boolt4a91_1_argbuf_bufchan_d <= readPointer_QTree_Boolt4a91_1_argbuf_d;
  QTree_Bool_t readPointer_QTree_Boolt4a91_1_argbuf_bufchan_buf;
  assign readPointer_QTree_Boolt4a91_1_argbuf_bufchan_r = (! readPointer_QTree_Boolt4a91_1_argbuf_bufchan_buf[0]);
  assign readPointer_QTree_Boolt4a91_1_argbuf_rwb_d = (readPointer_QTree_Boolt4a91_1_argbuf_bufchan_buf[0] ? readPointer_QTree_Boolt4a91_1_argbuf_bufchan_buf :
                                                       readPointer_QTree_Boolt4a91_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Boolt4a91_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((readPointer_QTree_Boolt4a91_1_argbuf_rwb_r && readPointer_QTree_Boolt4a91_1_argbuf_bufchan_buf[0]))
        readPointer_QTree_Boolt4a91_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
      else if (((! readPointer_QTree_Boolt4a91_1_argbuf_rwb_r) && (! readPointer_QTree_Boolt4a91_1_argbuf_bufchan_buf[0])))
        readPointer_QTree_Boolt4a91_1_argbuf_bufchan_buf <= readPointer_QTree_Boolt4a91_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CTf) : (sc_0_5_destruct,Pointer_CTf) > (sc_0_5_1_argbuf,Pointer_CTf) */
  Pointer_CTf_t sc_0_5_destruct_bufchan_d;
  logic sc_0_5_destruct_bufchan_r;
  assign sc_0_5_destruct_r = ((! sc_0_5_destruct_bufchan_d[0]) || sc_0_5_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) sc_0_5_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (sc_0_5_destruct_r)
        sc_0_5_destruct_bufchan_d <= sc_0_5_destruct_d;
  Pointer_CTf_t sc_0_5_destruct_bufchan_buf;
  assign sc_0_5_destruct_bufchan_r = (! sc_0_5_destruct_bufchan_buf[0]);
  assign sc_0_5_1_argbuf_d = (sc_0_5_destruct_bufchan_buf[0] ? sc_0_5_destruct_bufchan_buf :
                              sc_0_5_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) sc_0_5_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((sc_0_5_1_argbuf_r && sc_0_5_destruct_bufchan_buf[0]))
        sc_0_5_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! sc_0_5_1_argbuf_r) && (! sc_0_5_destruct_bufchan_buf[0])))
        sc_0_5_destruct_bufchan_buf <= sc_0_5_destruct_bufchan_d;
  
  /* buf (Ty Pointer_CTf'''''''''''') : (sc_0_9_destruct,Pointer_CTf'''''''''''') > (sc_0_9_1_argbuf,Pointer_CTf'''''''''''') */
  \Pointer_CTf''''''''''''_t  sc_0_9_destruct_bufchan_d;
  logic sc_0_9_destruct_bufchan_r;
  assign sc_0_9_destruct_r = ((! sc_0_9_destruct_bufchan_d[0]) || sc_0_9_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) sc_0_9_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (sc_0_9_destruct_r)
        sc_0_9_destruct_bufchan_d <= sc_0_9_destruct_d;
  \Pointer_CTf''''''''''''_t  sc_0_9_destruct_bufchan_buf;
  assign sc_0_9_destruct_bufchan_r = (! sc_0_9_destruct_bufchan_buf[0]);
  assign sc_0_9_1_argbuf_d = (sc_0_9_destruct_bufchan_buf[0] ? sc_0_9_destruct_bufchan_buf :
                              sc_0_9_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) sc_0_9_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((sc_0_9_1_argbuf_r && sc_0_9_destruct_bufchan_buf[0]))
        sc_0_9_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! sc_0_9_1_argbuf_r) && (! sc_0_9_destruct_bufchan_buf[0])))
        sc_0_9_destruct_bufchan_buf <= sc_0_9_destruct_bufchan_d;
  
  /* buf (Ty Pointer_CTf'''''''''''') : (scfarg_0_1_goMux_mux,Pointer_CTf'''''''''''') > (scfarg_0_1_1_argbuf,Pointer_CTf'''''''''''') */
  \Pointer_CTf''''''''''''_t  scfarg_0_1_goMux_mux_bufchan_d;
  logic scfarg_0_1_goMux_mux_bufchan_r;
  assign scfarg_0_1_goMux_mux_r = ((! scfarg_0_1_goMux_mux_bufchan_d[0]) || scfarg_0_1_goMux_mux_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      scfarg_0_1_goMux_mux_bufchan_d <= {16'd0, 1'd0};
    else
      if (scfarg_0_1_goMux_mux_r)
        scfarg_0_1_goMux_mux_bufchan_d <= scfarg_0_1_goMux_mux_d;
  \Pointer_CTf''''''''''''_t  scfarg_0_1_goMux_mux_bufchan_buf;
  assign scfarg_0_1_goMux_mux_bufchan_r = (! scfarg_0_1_goMux_mux_bufchan_buf[0]);
  assign scfarg_0_1_1_argbuf_d = (scfarg_0_1_goMux_mux_bufchan_buf[0] ? scfarg_0_1_goMux_mux_bufchan_buf :
                                  scfarg_0_1_goMux_mux_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      scfarg_0_1_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((scfarg_0_1_1_argbuf_r && scfarg_0_1_goMux_mux_bufchan_buf[0]))
        scfarg_0_1_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
      else if (((! scfarg_0_1_1_argbuf_r) && (! scfarg_0_1_goMux_mux_bufchan_buf[0])))
        scfarg_0_1_goMux_mux_bufchan_buf <= scfarg_0_1_goMux_mux_bufchan_d;
  
  /* buf (Ty Pointer_CTf) : (scfarg_0_goMux_mux,Pointer_CTf) > (scfarg_0_1_argbuf,Pointer_CTf) */
  Pointer_CTf_t scfarg_0_goMux_mux_bufchan_d;
  logic scfarg_0_goMux_mux_bufchan_r;
  assign scfarg_0_goMux_mux_r = ((! scfarg_0_goMux_mux_bufchan_d[0]) || scfarg_0_goMux_mux_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) scfarg_0_goMux_mux_bufchan_d <= {16'd0, 1'd0};
    else
      if (scfarg_0_goMux_mux_r)
        scfarg_0_goMux_mux_bufchan_d <= scfarg_0_goMux_mux_d;
  Pointer_CTf_t scfarg_0_goMux_mux_bufchan_buf;
  assign scfarg_0_goMux_mux_bufchan_r = (! scfarg_0_goMux_mux_bufchan_buf[0]);
  assign scfarg_0_1_argbuf_d = (scfarg_0_goMux_mux_bufchan_buf[0] ? scfarg_0_goMux_mux_bufchan_buf :
                                scfarg_0_goMux_mux_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      scfarg_0_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((scfarg_0_1_argbuf_r && scfarg_0_goMux_mux_bufchan_buf[0]))
        scfarg_0_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
      else if (((! scfarg_0_1_argbuf_r) && (! scfarg_0_goMux_mux_bufchan_buf[0])))
        scfarg_0_goMux_mux_bufchan_buf <= scfarg_0_goMux_mux_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (t1'a8W_3_destruct,Pointer_QTree_Bool) > (t1'a8W_3_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t \t1'a8W_3_destruct_bufchan_d ;
  logic \t1'a8W_3_destruct_bufchan_r ;
  assign \t1'a8W_3_destruct_r  = ((! \t1'a8W_3_destruct_bufchan_d [0]) || \t1'a8W_3_destruct_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \t1'a8W_3_destruct_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\t1'a8W_3_destruct_r )
        \t1'a8W_3_destruct_bufchan_d  <= \t1'a8W_3_destruct_d ;
  Pointer_QTree_Bool_t \t1'a8W_3_destruct_bufchan_buf ;
  assign \t1'a8W_3_destruct_bufchan_r  = (! \t1'a8W_3_destruct_bufchan_buf [0]);
  assign \t1'a8W_3_1_argbuf_d  = (\t1'a8W_3_destruct_bufchan_buf [0] ? \t1'a8W_3_destruct_bufchan_buf  :
                                  \t1'a8W_3_destruct_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \t1'a8W_3_destruct_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((\t1'a8W_3_1_argbuf_r  && \t1'a8W_3_destruct_bufchan_buf [0]))
        \t1'a8W_3_destruct_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! \t1'a8W_3_1_argbuf_r ) && (! \t1'a8W_3_destruct_bufchan_buf [0])))
        \t1'a8W_3_destruct_bufchan_buf  <= \t1'a8W_3_destruct_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Bool) : (t1a8M_destruct,Pointer_QTree_Bool) > (t1a8M_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t t1a8M_destruct_bufchan_d;
  logic t1a8M_destruct_bufchan_r;
  assign t1a8M_destruct_r = ((! t1a8M_destruct_bufchan_d[0]) || t1a8M_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t1a8M_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (t1a8M_destruct_r) t1a8M_destruct_bufchan_d <= t1a8M_destruct_d;
  Pointer_QTree_Bool_t t1a8M_destruct_bufchan_buf;
  assign t1a8M_destruct_bufchan_r = (! t1a8M_destruct_bufchan_buf[0]);
  assign t1a8M_1_argbuf_d = (t1a8M_destruct_bufchan_buf[0] ? t1a8M_destruct_bufchan_buf :
                             t1a8M_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t1a8M_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((t1a8M_1_argbuf_r && t1a8M_destruct_bufchan_buf[0]))
        t1a8M_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! t1a8M_1_argbuf_r) && (! t1a8M_destruct_bufchan_buf[0])))
        t1a8M_destruct_bufchan_buf <= t1a8M_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (t1a8R_3_destruct,Pointer_QTree_Bool) > (t1a8R_3_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t t1a8R_3_destruct_bufchan_d;
  logic t1a8R_3_destruct_bufchan_r;
  assign t1a8R_3_destruct_r = ((! t1a8R_3_destruct_bufchan_d[0]) || t1a8R_3_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t1a8R_3_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (t1a8R_3_destruct_r)
        t1a8R_3_destruct_bufchan_d <= t1a8R_3_destruct_d;
  Pointer_QTree_Bool_t t1a8R_3_destruct_bufchan_buf;
  assign t1a8R_3_destruct_bufchan_r = (! t1a8R_3_destruct_bufchan_buf[0]);
  assign t1a8R_3_1_argbuf_d = (t1a8R_3_destruct_bufchan_buf[0] ? t1a8R_3_destruct_bufchan_buf :
                               t1a8R_3_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t1a8R_3_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((t1a8R_3_1_argbuf_r && t1a8R_3_destruct_bufchan_buf[0]))
        t1a8R_3_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! t1a8R_3_1_argbuf_r) && (! t1a8R_3_destruct_bufchan_buf[0])))
        t1a8R_3_destruct_bufchan_buf <= t1a8R_3_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (t1a8i_destruct,Pointer_QTree_Bool) > (t1a8i_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t t1a8i_destruct_bufchan_d;
  logic t1a8i_destruct_bufchan_r;
  assign t1a8i_destruct_r = ((! t1a8i_destruct_bufchan_d[0]) || t1a8i_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t1a8i_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (t1a8i_destruct_r) t1a8i_destruct_bufchan_d <= t1a8i_destruct_d;
  Pointer_QTree_Bool_t t1a8i_destruct_bufchan_buf;
  assign t1a8i_destruct_bufchan_r = (! t1a8i_destruct_bufchan_buf[0]);
  assign t1a8i_1_argbuf_d = (t1a8i_destruct_bufchan_buf[0] ? t1a8i_destruct_bufchan_buf :
                             t1a8i_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t1a8i_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((t1a8i_1_argbuf_r && t1a8i_destruct_bufchan_buf[0]))
        t1a8i_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! t1a8i_1_argbuf_r) && (! t1a8i_destruct_bufchan_buf[0])))
        t1a8i_destruct_bufchan_buf <= t1a8i_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (t1a9d_3_destruct,Pointer_QTree_Bool) > (t1a9d_3_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t t1a9d_3_destruct_bufchan_d;
  logic t1a9d_3_destruct_bufchan_r;
  assign t1a9d_3_destruct_r = ((! t1a9d_3_destruct_bufchan_d[0]) || t1a9d_3_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t1a9d_3_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (t1a9d_3_destruct_r)
        t1a9d_3_destruct_bufchan_d <= t1a9d_3_destruct_d;
  Pointer_QTree_Bool_t t1a9d_3_destruct_bufchan_buf;
  assign t1a9d_3_destruct_bufchan_r = (! t1a9d_3_destruct_bufchan_buf[0]);
  assign t1a9d_3_1_argbuf_d = (t1a9d_3_destruct_bufchan_buf[0] ? t1a9d_3_destruct_bufchan_buf :
                               t1a9d_3_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t1a9d_3_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((t1a9d_3_1_argbuf_r && t1a9d_3_destruct_bufchan_buf[0]))
        t1a9d_3_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! t1a9d_3_1_argbuf_r) && (! t1a9d_3_destruct_bufchan_buf[0])))
        t1a9d_3_destruct_bufchan_buf <= t1a9d_3_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (t2'a8X_2_destruct,Pointer_QTree_Bool) > (t2'a8X_2_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t \t2'a8X_2_destruct_bufchan_d ;
  logic \t2'a8X_2_destruct_bufchan_r ;
  assign \t2'a8X_2_destruct_r  = ((! \t2'a8X_2_destruct_bufchan_d [0]) || \t2'a8X_2_destruct_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \t2'a8X_2_destruct_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\t2'a8X_2_destruct_r )
        \t2'a8X_2_destruct_bufchan_d  <= \t2'a8X_2_destruct_d ;
  Pointer_QTree_Bool_t \t2'a8X_2_destruct_bufchan_buf ;
  assign \t2'a8X_2_destruct_bufchan_r  = (! \t2'a8X_2_destruct_bufchan_buf [0]);
  assign \t2'a8X_2_1_argbuf_d  = (\t2'a8X_2_destruct_bufchan_buf [0] ? \t2'a8X_2_destruct_bufchan_buf  :
                                  \t2'a8X_2_destruct_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \t2'a8X_2_destruct_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((\t2'a8X_2_1_argbuf_r  && \t2'a8X_2_destruct_bufchan_buf [0]))
        \t2'a8X_2_destruct_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! \t2'a8X_2_1_argbuf_r ) && (! \t2'a8X_2_destruct_bufchan_buf [0])))
        \t2'a8X_2_destruct_bufchan_buf  <= \t2'a8X_2_destruct_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Bool) : (t2a8N_destruct,Pointer_QTree_Bool) > (t2a8N_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t t2a8N_destruct_bufchan_d;
  logic t2a8N_destruct_bufchan_r;
  assign t2a8N_destruct_r = ((! t2a8N_destruct_bufchan_d[0]) || t2a8N_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t2a8N_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (t2a8N_destruct_r) t2a8N_destruct_bufchan_d <= t2a8N_destruct_d;
  Pointer_QTree_Bool_t t2a8N_destruct_bufchan_buf;
  assign t2a8N_destruct_bufchan_r = (! t2a8N_destruct_bufchan_buf[0]);
  assign t2a8N_1_argbuf_d = (t2a8N_destruct_bufchan_buf[0] ? t2a8N_destruct_bufchan_buf :
                             t2a8N_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t2a8N_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((t2a8N_1_argbuf_r && t2a8N_destruct_bufchan_buf[0]))
        t2a8N_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! t2a8N_1_argbuf_r) && (! t2a8N_destruct_bufchan_buf[0])))
        t2a8N_destruct_bufchan_buf <= t2a8N_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (t2a8S_2_destruct,Pointer_QTree_Bool) > (t2a8S_2_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t t2a8S_2_destruct_bufchan_d;
  logic t2a8S_2_destruct_bufchan_r;
  assign t2a8S_2_destruct_r = ((! t2a8S_2_destruct_bufchan_d[0]) || t2a8S_2_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t2a8S_2_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (t2a8S_2_destruct_r)
        t2a8S_2_destruct_bufchan_d <= t2a8S_2_destruct_d;
  Pointer_QTree_Bool_t t2a8S_2_destruct_bufchan_buf;
  assign t2a8S_2_destruct_bufchan_r = (! t2a8S_2_destruct_bufchan_buf[0]);
  assign t2a8S_2_1_argbuf_d = (t2a8S_2_destruct_bufchan_buf[0] ? t2a8S_2_destruct_bufchan_buf :
                               t2a8S_2_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t2a8S_2_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((t2a8S_2_1_argbuf_r && t2a8S_2_destruct_bufchan_buf[0]))
        t2a8S_2_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! t2a8S_2_1_argbuf_r) && (! t2a8S_2_destruct_bufchan_buf[0])))
        t2a8S_2_destruct_bufchan_buf <= t2a8S_2_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (t2a8j_destruct,Pointer_QTree_Bool) > (t2a8j_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t t2a8j_destruct_bufchan_d;
  logic t2a8j_destruct_bufchan_r;
  assign t2a8j_destruct_r = ((! t2a8j_destruct_bufchan_d[0]) || t2a8j_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t2a8j_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (t2a8j_destruct_r) t2a8j_destruct_bufchan_d <= t2a8j_destruct_d;
  Pointer_QTree_Bool_t t2a8j_destruct_bufchan_buf;
  assign t2a8j_destruct_bufchan_r = (! t2a8j_destruct_bufchan_buf[0]);
  assign t2a8j_1_argbuf_d = (t2a8j_destruct_bufchan_buf[0] ? t2a8j_destruct_bufchan_buf :
                             t2a8j_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t2a8j_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((t2a8j_1_argbuf_r && t2a8j_destruct_bufchan_buf[0]))
        t2a8j_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! t2a8j_1_argbuf_r) && (! t2a8j_destruct_bufchan_buf[0])))
        t2a8j_destruct_bufchan_buf <= t2a8j_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (t2a9e_2_destruct,Pointer_QTree_Bool) > (t2a9e_2_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t t2a9e_2_destruct_bufchan_d;
  logic t2a9e_2_destruct_bufchan_r;
  assign t2a9e_2_destruct_r = ((! t2a9e_2_destruct_bufchan_d[0]) || t2a9e_2_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t2a9e_2_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (t2a9e_2_destruct_r)
        t2a9e_2_destruct_bufchan_d <= t2a9e_2_destruct_d;
  Pointer_QTree_Bool_t t2a9e_2_destruct_bufchan_buf;
  assign t2a9e_2_destruct_bufchan_r = (! t2a9e_2_destruct_bufchan_buf[0]);
  assign t2a9e_2_1_argbuf_d = (t2a9e_2_destruct_bufchan_buf[0] ? t2a9e_2_destruct_bufchan_buf :
                               t2a9e_2_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t2a9e_2_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((t2a9e_2_1_argbuf_r && t2a9e_2_destruct_bufchan_buf[0]))
        t2a9e_2_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! t2a9e_2_1_argbuf_r) && (! t2a9e_2_destruct_bufchan_buf[0])))
        t2a9e_2_destruct_bufchan_buf <= t2a9e_2_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (t3'a8Y_1_destruct,Pointer_QTree_Bool) > (t3'a8Y_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t \t3'a8Y_1_destruct_bufchan_d ;
  logic \t3'a8Y_1_destruct_bufchan_r ;
  assign \t3'a8Y_1_destruct_r  = ((! \t3'a8Y_1_destruct_bufchan_d [0]) || \t3'a8Y_1_destruct_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \t3'a8Y_1_destruct_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\t3'a8Y_1_destruct_r )
        \t3'a8Y_1_destruct_bufchan_d  <= \t3'a8Y_1_destruct_d ;
  Pointer_QTree_Bool_t \t3'a8Y_1_destruct_bufchan_buf ;
  assign \t3'a8Y_1_destruct_bufchan_r  = (! \t3'a8Y_1_destruct_bufchan_buf [0]);
  assign \t3'a8Y_1_1_argbuf_d  = (\t3'a8Y_1_destruct_bufchan_buf [0] ? \t3'a8Y_1_destruct_bufchan_buf  :
                                  \t3'a8Y_1_destruct_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \t3'a8Y_1_destruct_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((\t3'a8Y_1_1_argbuf_r  && \t3'a8Y_1_destruct_bufchan_buf [0]))
        \t3'a8Y_1_destruct_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! \t3'a8Y_1_1_argbuf_r ) && (! \t3'a8Y_1_destruct_bufchan_buf [0])))
        \t3'a8Y_1_destruct_bufchan_buf  <= \t3'a8Y_1_destruct_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Bool) : (t3a8O_destruct,Pointer_QTree_Bool) > (t3a8O_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t t3a8O_destruct_bufchan_d;
  logic t3a8O_destruct_bufchan_r;
  assign t3a8O_destruct_r = ((! t3a8O_destruct_bufchan_d[0]) || t3a8O_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t3a8O_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (t3a8O_destruct_r) t3a8O_destruct_bufchan_d <= t3a8O_destruct_d;
  Pointer_QTree_Bool_t t3a8O_destruct_bufchan_buf;
  assign t3a8O_destruct_bufchan_r = (! t3a8O_destruct_bufchan_buf[0]);
  assign t3a8O_1_argbuf_d = (t3a8O_destruct_bufchan_buf[0] ? t3a8O_destruct_bufchan_buf :
                             t3a8O_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t3a8O_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((t3a8O_1_argbuf_r && t3a8O_destruct_bufchan_buf[0]))
        t3a8O_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! t3a8O_1_argbuf_r) && (! t3a8O_destruct_bufchan_buf[0])))
        t3a8O_destruct_bufchan_buf <= t3a8O_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (t3a8T_1_destruct,Pointer_QTree_Bool) > (t3a8T_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t t3a8T_1_destruct_bufchan_d;
  logic t3a8T_1_destruct_bufchan_r;
  assign t3a8T_1_destruct_r = ((! t3a8T_1_destruct_bufchan_d[0]) || t3a8T_1_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t3a8T_1_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (t3a8T_1_destruct_r)
        t3a8T_1_destruct_bufchan_d <= t3a8T_1_destruct_d;
  Pointer_QTree_Bool_t t3a8T_1_destruct_bufchan_buf;
  assign t3a8T_1_destruct_bufchan_r = (! t3a8T_1_destruct_bufchan_buf[0]);
  assign t3a8T_1_1_argbuf_d = (t3a8T_1_destruct_bufchan_buf[0] ? t3a8T_1_destruct_bufchan_buf :
                               t3a8T_1_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t3a8T_1_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((t3a8T_1_1_argbuf_r && t3a8T_1_destruct_bufchan_buf[0]))
        t3a8T_1_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! t3a8T_1_1_argbuf_r) && (! t3a8T_1_destruct_bufchan_buf[0])))
        t3a8T_1_destruct_bufchan_buf <= t3a8T_1_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (t3a8k_destruct,Pointer_QTree_Bool) > (t3a8k_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t t3a8k_destruct_bufchan_d;
  logic t3a8k_destruct_bufchan_r;
  assign t3a8k_destruct_r = ((! t3a8k_destruct_bufchan_d[0]) || t3a8k_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t3a8k_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (t3a8k_destruct_r) t3a8k_destruct_bufchan_d <= t3a8k_destruct_d;
  Pointer_QTree_Bool_t t3a8k_destruct_bufchan_buf;
  assign t3a8k_destruct_bufchan_r = (! t3a8k_destruct_bufchan_buf[0]);
  assign t3a8k_1_argbuf_d = (t3a8k_destruct_bufchan_buf[0] ? t3a8k_destruct_bufchan_buf :
                             t3a8k_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t3a8k_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((t3a8k_1_argbuf_r && t3a8k_destruct_bufchan_buf[0]))
        t3a8k_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! t3a8k_1_argbuf_r) && (! t3a8k_destruct_bufchan_buf[0])))
        t3a8k_destruct_bufchan_buf <= t3a8k_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (t3a9f_1_destruct,Pointer_QTree_Bool) > (t3a9f_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t t3a9f_1_destruct_bufchan_d;
  logic t3a9f_1_destruct_bufchan_r;
  assign t3a9f_1_destruct_r = ((! t3a9f_1_destruct_bufchan_d[0]) || t3a9f_1_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t3a9f_1_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (t3a9f_1_destruct_r)
        t3a9f_1_destruct_bufchan_d <= t3a9f_1_destruct_d;
  Pointer_QTree_Bool_t t3a9f_1_destruct_bufchan_buf;
  assign t3a9f_1_destruct_bufchan_r = (! t3a9f_1_destruct_bufchan_buf[0]);
  assign t3a9f_1_1_argbuf_d = (t3a9f_1_destruct_bufchan_buf[0] ? t3a9f_1_destruct_bufchan_buf :
                               t3a9f_1_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t3a9f_1_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((t3a9f_1_1_argbuf_r && t3a9f_1_destruct_bufchan_buf[0]))
        t3a9f_1_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! t3a9f_1_1_argbuf_r) && (! t3a9f_1_destruct_bufchan_buf[0])))
        t3a9f_1_destruct_bufchan_buf <= t3a9f_1_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (t4'a8Z_destruct,Pointer_QTree_Bool) > (t4'a8Z_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t \t4'a8Z_destruct_bufchan_d ;
  logic \t4'a8Z_destruct_bufchan_r ;
  assign \t4'a8Z_destruct_r  = ((! \t4'a8Z_destruct_bufchan_d [0]) || \t4'a8Z_destruct_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \t4'a8Z_destruct_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\t4'a8Z_destruct_r )
        \t4'a8Z_destruct_bufchan_d  <= \t4'a8Z_destruct_d ;
  Pointer_QTree_Bool_t \t4'a8Z_destruct_bufchan_buf ;
  assign \t4'a8Z_destruct_bufchan_r  = (! \t4'a8Z_destruct_bufchan_buf [0]);
  assign \t4'a8Z_1_argbuf_d  = (\t4'a8Z_destruct_bufchan_buf [0] ? \t4'a8Z_destruct_bufchan_buf  :
                                \t4'a8Z_destruct_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \t4'a8Z_destruct_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((\t4'a8Z_1_argbuf_r  && \t4'a8Z_destruct_bufchan_buf [0]))
        \t4'a8Z_destruct_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! \t4'a8Z_1_argbuf_r ) && (! \t4'a8Z_destruct_bufchan_buf [0])))
        \t4'a8Z_destruct_bufchan_buf  <= \t4'a8Z_destruct_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Bool) : (t4a8P_destruct,Pointer_QTree_Bool) > (t4a8P_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t t4a8P_destruct_bufchan_d;
  logic t4a8P_destruct_bufchan_r;
  assign t4a8P_destruct_r = ((! t4a8P_destruct_bufchan_d[0]) || t4a8P_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t4a8P_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (t4a8P_destruct_r) t4a8P_destruct_bufchan_d <= t4a8P_destruct_d;
  Pointer_QTree_Bool_t t4a8P_destruct_bufchan_buf;
  assign t4a8P_destruct_bufchan_r = (! t4a8P_destruct_bufchan_buf[0]);
  assign t4a8P_1_argbuf_d = (t4a8P_destruct_bufchan_buf[0] ? t4a8P_destruct_bufchan_buf :
                             t4a8P_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t4a8P_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((t4a8P_1_argbuf_r && t4a8P_destruct_bufchan_buf[0]))
        t4a8P_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! t4a8P_1_argbuf_r) && (! t4a8P_destruct_bufchan_buf[0])))
        t4a8P_destruct_bufchan_buf <= t4a8P_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (t4a8l_destruct,Pointer_QTree_Bool) > (t4a8l_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t t4a8l_destruct_bufchan_d;
  logic t4a8l_destruct_bufchan_r;
  assign t4a8l_destruct_r = ((! t4a8l_destruct_bufchan_d[0]) || t4a8l_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t4a8l_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (t4a8l_destruct_r) t4a8l_destruct_bufchan_d <= t4a8l_destruct_d;
  Pointer_QTree_Bool_t t4a8l_destruct_bufchan_buf;
  assign t4a8l_destruct_bufchan_r = (! t4a8l_destruct_bufchan_buf[0]);
  assign t4a8l_1_argbuf_d = (t4a8l_destruct_bufchan_buf[0] ? t4a8l_destruct_bufchan_buf :
                             t4a8l_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t4a8l_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((t4a8l_1_argbuf_r && t4a8l_destruct_bufchan_buf[0]))
        t4a8l_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! t4a8l_1_argbuf_r) && (! t4a8l_destruct_bufchan_buf[0])))
        t4a8l_destruct_bufchan_buf <= t4a8l_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (t4a91_1,Pointer_QTree_Bool) > (t4a91_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t t4a91_1_bufchan_d;
  logic t4a91_1_bufchan_r;
  assign t4a91_1_r = ((! t4a91_1_bufchan_d[0]) || t4a91_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t4a91_1_bufchan_d <= {16'd0, 1'd0};
    else if (t4a91_1_r) t4a91_1_bufchan_d <= t4a91_1_d;
  Pointer_QTree_Bool_t t4a91_1_bufchan_buf;
  assign t4a91_1_bufchan_r = (! t4a91_1_bufchan_buf[0]);
  assign t4a91_1_argbuf_d = (t4a91_1_bufchan_buf[0] ? t4a91_1_bufchan_buf :
                             t4a91_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t4a91_1_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((t4a91_1_argbuf_r && t4a91_1_bufchan_buf[0]))
        t4a91_1_bufchan_buf <= {16'd0, 1'd0};
      else if (((! t4a91_1_argbuf_r) && (! t4a91_1_bufchan_buf[0])))
        t4a91_1_bufchan_buf <= t4a91_1_bufchan_d;
  
  /* fork (Ty Pointer_QTree_Bool) : (t4a91_goMux_mux,Pointer_QTree_Bool) > [(t4a91_1,Pointer_QTree_Bool),
                                                                       (t4a91_2,Pointer_QTree_Bool)] */
  logic [1:0] t4a91_goMux_mux_emitted;
  logic [1:0] t4a91_goMux_mux_done;
  assign t4a91_1_d = {t4a91_goMux_mux_d[16:1],
                      (t4a91_goMux_mux_d[0] && (! t4a91_goMux_mux_emitted[0]))};
  assign t4a91_2_d = {t4a91_goMux_mux_d[16:1],
                      (t4a91_goMux_mux_d[0] && (! t4a91_goMux_mux_emitted[1]))};
  assign t4a91_goMux_mux_done = (t4a91_goMux_mux_emitted | ({t4a91_2_d[0],
                                                             t4a91_1_d[0]} & {t4a91_2_r,
                                                                              t4a91_1_r}));
  assign t4a91_goMux_mux_r = (& t4a91_goMux_mux_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t4a91_goMux_mux_emitted <= 2'd0;
    else
      t4a91_goMux_mux_emitted <= (t4a91_goMux_mux_r ? 2'd0 :
                                  t4a91_goMux_mux_done);
  
  /* buf (Ty Pointer_QTree_Bool) : (t5a9g_destruct,Pointer_QTree_Bool) > (t5a9g_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t t5a9g_destruct_bufchan_d;
  logic t5a9g_destruct_bufchan_r;
  assign t5a9g_destruct_r = ((! t5a9g_destruct_bufchan_d[0]) || t5a9g_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t5a9g_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (t5a9g_destruct_r) t5a9g_destruct_bufchan_d <= t5a9g_destruct_d;
  Pointer_QTree_Bool_t t5a9g_destruct_bufchan_buf;
  assign t5a9g_destruct_bufchan_r = (! t5a9g_destruct_bufchan_buf[0]);
  assign t5a9g_1_argbuf_d = (t5a9g_destruct_bufchan_buf[0] ? t5a9g_destruct_bufchan_buf :
                             t5a9g_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t5a9g_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((t5a9g_1_argbuf_r && t5a9g_destruct_bufchan_buf[0]))
        t5a9g_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! t5a9g_1_argbuf_r) && (! t5a9g_destruct_bufchan_buf[0])))
        t5a9g_destruct_bufchan_buf <= t5a9g_destruct_bufchan_d;
  
  /* buf (Ty Pointer_CTf'''''''''''') : (writeCTf''''''''''''lizzieLet54_1_argbuf,Pointer_CTf'''''''''''') > (writeCTf''''''''''''lizzieLet54_1_argbuf_rwb,Pointer_CTf'''''''''''') */
  \Pointer_CTf''''''''''''_t  \writeCTf''''''''''''lizzieLet54_1_argbuf_bufchan_d ;
  logic \writeCTf''''''''''''lizzieLet54_1_argbuf_bufchan_r ;
  assign \writeCTf''''''''''''lizzieLet54_1_argbuf_r  = ((! \writeCTf''''''''''''lizzieLet54_1_argbuf_bufchan_d [0]) || \writeCTf''''''''''''lizzieLet54_1_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf''''''''''''lizzieLet54_1_argbuf_bufchan_d  <= {16'd0,
                                                               1'd0};
    else
      if (\writeCTf''''''''''''lizzieLet54_1_argbuf_r )
        \writeCTf''''''''''''lizzieLet54_1_argbuf_bufchan_d  <= \writeCTf''''''''''''lizzieLet54_1_argbuf_d ;
  \Pointer_CTf''''''''''''_t  \writeCTf''''''''''''lizzieLet54_1_argbuf_bufchan_buf ;
  assign \writeCTf''''''''''''lizzieLet54_1_argbuf_bufchan_r  = (! \writeCTf''''''''''''lizzieLet54_1_argbuf_bufchan_buf [0]);
  assign \writeCTf''''''''''''lizzieLet54_1_argbuf_rwb_d  = (\writeCTf''''''''''''lizzieLet54_1_argbuf_bufchan_buf [0] ? \writeCTf''''''''''''lizzieLet54_1_argbuf_bufchan_buf  :
                                                             \writeCTf''''''''''''lizzieLet54_1_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf''''''''''''lizzieLet54_1_argbuf_bufchan_buf  <= {16'd0,
                                                                 1'd0};
    else
      if ((\writeCTf''''''''''''lizzieLet54_1_argbuf_rwb_r  && \writeCTf''''''''''''lizzieLet54_1_argbuf_bufchan_buf [0]))
        \writeCTf''''''''''''lizzieLet54_1_argbuf_bufchan_buf  <= {16'd0,
                                                                   1'd0};
      else if (((! \writeCTf''''''''''''lizzieLet54_1_argbuf_rwb_r ) && (! \writeCTf''''''''''''lizzieLet54_1_argbuf_bufchan_buf [0])))
        \writeCTf''''''''''''lizzieLet54_1_argbuf_bufchan_buf  <= \writeCTf''''''''''''lizzieLet54_1_argbuf_bufchan_d ;
  
  /* buf (Ty Pointer_CTf'''''''''''') : (writeCTf''''''''''''lizzieLet54_1_argbuf_rwb,Pointer_CTf'''''''''''') > (sca3_1_1_argbuf,Pointer_CTf'''''''''''') */
  \Pointer_CTf''''''''''''_t  \writeCTf''''''''''''lizzieLet54_1_argbuf_rwb_bufchan_d ;
  logic \writeCTf''''''''''''lizzieLet54_1_argbuf_rwb_bufchan_r ;
  assign \writeCTf''''''''''''lizzieLet54_1_argbuf_rwb_r  = ((! \writeCTf''''''''''''lizzieLet54_1_argbuf_rwb_bufchan_d [0]) || \writeCTf''''''''''''lizzieLet54_1_argbuf_rwb_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf''''''''''''lizzieLet54_1_argbuf_rwb_bufchan_d  <= {16'd0,
                                                                   1'd0};
    else
      if (\writeCTf''''''''''''lizzieLet54_1_argbuf_rwb_r )
        \writeCTf''''''''''''lizzieLet54_1_argbuf_rwb_bufchan_d  <= \writeCTf''''''''''''lizzieLet54_1_argbuf_rwb_d ;
  \Pointer_CTf''''''''''''_t  \writeCTf''''''''''''lizzieLet54_1_argbuf_rwb_bufchan_buf ;
  assign \writeCTf''''''''''''lizzieLet54_1_argbuf_rwb_bufchan_r  = (! \writeCTf''''''''''''lizzieLet54_1_argbuf_rwb_bufchan_buf [0]);
  assign sca3_1_1_argbuf_d = (\writeCTf''''''''''''lizzieLet54_1_argbuf_rwb_bufchan_buf [0] ? \writeCTf''''''''''''lizzieLet54_1_argbuf_rwb_bufchan_buf  :
                              \writeCTf''''''''''''lizzieLet54_1_argbuf_rwb_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf''''''''''''lizzieLet54_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                     1'd0};
    else
      if ((sca3_1_1_argbuf_r && \writeCTf''''''''''''lizzieLet54_1_argbuf_rwb_bufchan_buf [0]))
        \writeCTf''''''''''''lizzieLet54_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                       1'd0};
      else if (((! sca3_1_1_argbuf_r) && (! \writeCTf''''''''''''lizzieLet54_1_argbuf_rwb_bufchan_buf [0])))
        \writeCTf''''''''''''lizzieLet54_1_argbuf_rwb_bufchan_buf  <= \writeCTf''''''''''''lizzieLet54_1_argbuf_rwb_bufchan_d ;
  
  /* buf (Ty Pointer_CTf'''''''''''') : (writeCTf''''''''''''lizzieLet58_1_argbuf,Pointer_CTf'''''''''''') > (writeCTf''''''''''''lizzieLet58_1_argbuf_rwb,Pointer_CTf'''''''''''') */
  \Pointer_CTf''''''''''''_t  \writeCTf''''''''''''lizzieLet58_1_argbuf_bufchan_d ;
  logic \writeCTf''''''''''''lizzieLet58_1_argbuf_bufchan_r ;
  assign \writeCTf''''''''''''lizzieLet58_1_argbuf_r  = ((! \writeCTf''''''''''''lizzieLet58_1_argbuf_bufchan_d [0]) || \writeCTf''''''''''''lizzieLet58_1_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf''''''''''''lizzieLet58_1_argbuf_bufchan_d  <= {16'd0,
                                                               1'd0};
    else
      if (\writeCTf''''''''''''lizzieLet58_1_argbuf_r )
        \writeCTf''''''''''''lizzieLet58_1_argbuf_bufchan_d  <= \writeCTf''''''''''''lizzieLet58_1_argbuf_d ;
  \Pointer_CTf''''''''''''_t  \writeCTf''''''''''''lizzieLet58_1_argbuf_bufchan_buf ;
  assign \writeCTf''''''''''''lizzieLet58_1_argbuf_bufchan_r  = (! \writeCTf''''''''''''lizzieLet58_1_argbuf_bufchan_buf [0]);
  assign \writeCTf''''''''''''lizzieLet58_1_argbuf_rwb_d  = (\writeCTf''''''''''''lizzieLet58_1_argbuf_bufchan_buf [0] ? \writeCTf''''''''''''lizzieLet58_1_argbuf_bufchan_buf  :
                                                             \writeCTf''''''''''''lizzieLet58_1_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf''''''''''''lizzieLet58_1_argbuf_bufchan_buf  <= {16'd0,
                                                                 1'd0};
    else
      if ((\writeCTf''''''''''''lizzieLet58_1_argbuf_rwb_r  && \writeCTf''''''''''''lizzieLet58_1_argbuf_bufchan_buf [0]))
        \writeCTf''''''''''''lizzieLet58_1_argbuf_bufchan_buf  <= {16'd0,
                                                                   1'd0};
      else if (((! \writeCTf''''''''''''lizzieLet58_1_argbuf_rwb_r ) && (! \writeCTf''''''''''''lizzieLet58_1_argbuf_bufchan_buf [0])))
        \writeCTf''''''''''''lizzieLet58_1_argbuf_bufchan_buf  <= \writeCTf''''''''''''lizzieLet58_1_argbuf_bufchan_d ;
  
  /* buf (Ty Pointer_CTf'''''''''''') : (writeCTf''''''''''''lizzieLet58_1_argbuf_rwb,Pointer_CTf'''''''''''') > (lizzieLet7_1_1_argbuf,Pointer_CTf'''''''''''') */
  \Pointer_CTf''''''''''''_t  \writeCTf''''''''''''lizzieLet58_1_argbuf_rwb_bufchan_d ;
  logic \writeCTf''''''''''''lizzieLet58_1_argbuf_rwb_bufchan_r ;
  assign \writeCTf''''''''''''lizzieLet58_1_argbuf_rwb_r  = ((! \writeCTf''''''''''''lizzieLet58_1_argbuf_rwb_bufchan_d [0]) || \writeCTf''''''''''''lizzieLet58_1_argbuf_rwb_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf''''''''''''lizzieLet58_1_argbuf_rwb_bufchan_d  <= {16'd0,
                                                                   1'd0};
    else
      if (\writeCTf''''''''''''lizzieLet58_1_argbuf_rwb_r )
        \writeCTf''''''''''''lizzieLet58_1_argbuf_rwb_bufchan_d  <= \writeCTf''''''''''''lizzieLet58_1_argbuf_rwb_d ;
  \Pointer_CTf''''''''''''_t  \writeCTf''''''''''''lizzieLet58_1_argbuf_rwb_bufchan_buf ;
  assign \writeCTf''''''''''''lizzieLet58_1_argbuf_rwb_bufchan_r  = (! \writeCTf''''''''''''lizzieLet58_1_argbuf_rwb_bufchan_buf [0]);
  assign lizzieLet7_1_1_argbuf_d = (\writeCTf''''''''''''lizzieLet58_1_argbuf_rwb_bufchan_buf [0] ? \writeCTf''''''''''''lizzieLet58_1_argbuf_rwb_bufchan_buf  :
                                    \writeCTf''''''''''''lizzieLet58_1_argbuf_rwb_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf''''''''''''lizzieLet58_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                     1'd0};
    else
      if ((lizzieLet7_1_1_argbuf_r && \writeCTf''''''''''''lizzieLet58_1_argbuf_rwb_bufchan_buf [0]))
        \writeCTf''''''''''''lizzieLet58_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                       1'd0};
      else if (((! lizzieLet7_1_1_argbuf_r) && (! \writeCTf''''''''''''lizzieLet58_1_argbuf_rwb_bufchan_buf [0])))
        \writeCTf''''''''''''lizzieLet58_1_argbuf_rwb_bufchan_buf  <= \writeCTf''''''''''''lizzieLet58_1_argbuf_rwb_bufchan_d ;
  
  /* buf (Ty Pointer_CTf'''''''''''') : (writeCTf''''''''''''lizzieLet66_1_argbuf,Pointer_CTf'''''''''''') > (writeCTf''''''''''''lizzieLet66_1_argbuf_rwb,Pointer_CTf'''''''''''') */
  \Pointer_CTf''''''''''''_t  \writeCTf''''''''''''lizzieLet66_1_argbuf_bufchan_d ;
  logic \writeCTf''''''''''''lizzieLet66_1_argbuf_bufchan_r ;
  assign \writeCTf''''''''''''lizzieLet66_1_argbuf_r  = ((! \writeCTf''''''''''''lizzieLet66_1_argbuf_bufchan_d [0]) || \writeCTf''''''''''''lizzieLet66_1_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf''''''''''''lizzieLet66_1_argbuf_bufchan_d  <= {16'd0,
                                                               1'd0};
    else
      if (\writeCTf''''''''''''lizzieLet66_1_argbuf_r )
        \writeCTf''''''''''''lizzieLet66_1_argbuf_bufchan_d  <= \writeCTf''''''''''''lizzieLet66_1_argbuf_d ;
  \Pointer_CTf''''''''''''_t  \writeCTf''''''''''''lizzieLet66_1_argbuf_bufchan_buf ;
  assign \writeCTf''''''''''''lizzieLet66_1_argbuf_bufchan_r  = (! \writeCTf''''''''''''lizzieLet66_1_argbuf_bufchan_buf [0]);
  assign \writeCTf''''''''''''lizzieLet66_1_argbuf_rwb_d  = (\writeCTf''''''''''''lizzieLet66_1_argbuf_bufchan_buf [0] ? \writeCTf''''''''''''lizzieLet66_1_argbuf_bufchan_buf  :
                                                             \writeCTf''''''''''''lizzieLet66_1_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf''''''''''''lizzieLet66_1_argbuf_bufchan_buf  <= {16'd0,
                                                                 1'd0};
    else
      if ((\writeCTf''''''''''''lizzieLet66_1_argbuf_rwb_r  && \writeCTf''''''''''''lizzieLet66_1_argbuf_bufchan_buf [0]))
        \writeCTf''''''''''''lizzieLet66_1_argbuf_bufchan_buf  <= {16'd0,
                                                                   1'd0};
      else if (((! \writeCTf''''''''''''lizzieLet66_1_argbuf_rwb_r ) && (! \writeCTf''''''''''''lizzieLet66_1_argbuf_bufchan_buf [0])))
        \writeCTf''''''''''''lizzieLet66_1_argbuf_bufchan_buf  <= \writeCTf''''''''''''lizzieLet66_1_argbuf_bufchan_d ;
  
  /* buf (Ty Pointer_CTf'''''''''''') : (writeCTf''''''''''''lizzieLet66_1_argbuf_rwb,Pointer_CTf'''''''''''') > (sca2_1_1_argbuf,Pointer_CTf'''''''''''') */
  \Pointer_CTf''''''''''''_t  \writeCTf''''''''''''lizzieLet66_1_argbuf_rwb_bufchan_d ;
  logic \writeCTf''''''''''''lizzieLet66_1_argbuf_rwb_bufchan_r ;
  assign \writeCTf''''''''''''lizzieLet66_1_argbuf_rwb_r  = ((! \writeCTf''''''''''''lizzieLet66_1_argbuf_rwb_bufchan_d [0]) || \writeCTf''''''''''''lizzieLet66_1_argbuf_rwb_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf''''''''''''lizzieLet66_1_argbuf_rwb_bufchan_d  <= {16'd0,
                                                                   1'd0};
    else
      if (\writeCTf''''''''''''lizzieLet66_1_argbuf_rwb_r )
        \writeCTf''''''''''''lizzieLet66_1_argbuf_rwb_bufchan_d  <= \writeCTf''''''''''''lizzieLet66_1_argbuf_rwb_d ;
  \Pointer_CTf''''''''''''_t  \writeCTf''''''''''''lizzieLet66_1_argbuf_rwb_bufchan_buf ;
  assign \writeCTf''''''''''''lizzieLet66_1_argbuf_rwb_bufchan_r  = (! \writeCTf''''''''''''lizzieLet66_1_argbuf_rwb_bufchan_buf [0]);
  assign sca2_1_1_argbuf_d = (\writeCTf''''''''''''lizzieLet66_1_argbuf_rwb_bufchan_buf [0] ? \writeCTf''''''''''''lizzieLet66_1_argbuf_rwb_bufchan_buf  :
                              \writeCTf''''''''''''lizzieLet66_1_argbuf_rwb_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf''''''''''''lizzieLet66_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                     1'd0};
    else
      if ((sca2_1_1_argbuf_r && \writeCTf''''''''''''lizzieLet66_1_argbuf_rwb_bufchan_buf [0]))
        \writeCTf''''''''''''lizzieLet66_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                       1'd0};
      else if (((! sca2_1_1_argbuf_r) && (! \writeCTf''''''''''''lizzieLet66_1_argbuf_rwb_bufchan_buf [0])))
        \writeCTf''''''''''''lizzieLet66_1_argbuf_rwb_bufchan_buf  <= \writeCTf''''''''''''lizzieLet66_1_argbuf_rwb_bufchan_d ;
  
  /* buf (Ty Pointer_CTf'''''''''''') : (writeCTf''''''''''''lizzieLet67_1_argbuf,Pointer_CTf'''''''''''') > (writeCTf''''''''''''lizzieLet67_1_argbuf_rwb,Pointer_CTf'''''''''''') */
  \Pointer_CTf''''''''''''_t  \writeCTf''''''''''''lizzieLet67_1_argbuf_bufchan_d ;
  logic \writeCTf''''''''''''lizzieLet67_1_argbuf_bufchan_r ;
  assign \writeCTf''''''''''''lizzieLet67_1_argbuf_r  = ((! \writeCTf''''''''''''lizzieLet67_1_argbuf_bufchan_d [0]) || \writeCTf''''''''''''lizzieLet67_1_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf''''''''''''lizzieLet67_1_argbuf_bufchan_d  <= {16'd0,
                                                               1'd0};
    else
      if (\writeCTf''''''''''''lizzieLet67_1_argbuf_r )
        \writeCTf''''''''''''lizzieLet67_1_argbuf_bufchan_d  <= \writeCTf''''''''''''lizzieLet67_1_argbuf_d ;
  \Pointer_CTf''''''''''''_t  \writeCTf''''''''''''lizzieLet67_1_argbuf_bufchan_buf ;
  assign \writeCTf''''''''''''lizzieLet67_1_argbuf_bufchan_r  = (! \writeCTf''''''''''''lizzieLet67_1_argbuf_bufchan_buf [0]);
  assign \writeCTf''''''''''''lizzieLet67_1_argbuf_rwb_d  = (\writeCTf''''''''''''lizzieLet67_1_argbuf_bufchan_buf [0] ? \writeCTf''''''''''''lizzieLet67_1_argbuf_bufchan_buf  :
                                                             \writeCTf''''''''''''lizzieLet67_1_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf''''''''''''lizzieLet67_1_argbuf_bufchan_buf  <= {16'd0,
                                                                 1'd0};
    else
      if ((\writeCTf''''''''''''lizzieLet67_1_argbuf_rwb_r  && \writeCTf''''''''''''lizzieLet67_1_argbuf_bufchan_buf [0]))
        \writeCTf''''''''''''lizzieLet67_1_argbuf_bufchan_buf  <= {16'd0,
                                                                   1'd0};
      else if (((! \writeCTf''''''''''''lizzieLet67_1_argbuf_rwb_r ) && (! \writeCTf''''''''''''lizzieLet67_1_argbuf_bufchan_buf [0])))
        \writeCTf''''''''''''lizzieLet67_1_argbuf_bufchan_buf  <= \writeCTf''''''''''''lizzieLet67_1_argbuf_bufchan_d ;
  
  /* buf (Ty Pointer_CTf'''''''''''') : (writeCTf''''''''''''lizzieLet67_1_argbuf_rwb,Pointer_CTf'''''''''''') > (sca1_1_1_argbuf,Pointer_CTf'''''''''''') */
  \Pointer_CTf''''''''''''_t  \writeCTf''''''''''''lizzieLet67_1_argbuf_rwb_bufchan_d ;
  logic \writeCTf''''''''''''lizzieLet67_1_argbuf_rwb_bufchan_r ;
  assign \writeCTf''''''''''''lizzieLet67_1_argbuf_rwb_r  = ((! \writeCTf''''''''''''lizzieLet67_1_argbuf_rwb_bufchan_d [0]) || \writeCTf''''''''''''lizzieLet67_1_argbuf_rwb_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf''''''''''''lizzieLet67_1_argbuf_rwb_bufchan_d  <= {16'd0,
                                                                   1'd0};
    else
      if (\writeCTf''''''''''''lizzieLet67_1_argbuf_rwb_r )
        \writeCTf''''''''''''lizzieLet67_1_argbuf_rwb_bufchan_d  <= \writeCTf''''''''''''lizzieLet67_1_argbuf_rwb_d ;
  \Pointer_CTf''''''''''''_t  \writeCTf''''''''''''lizzieLet67_1_argbuf_rwb_bufchan_buf ;
  assign \writeCTf''''''''''''lizzieLet67_1_argbuf_rwb_bufchan_r  = (! \writeCTf''''''''''''lizzieLet67_1_argbuf_rwb_bufchan_buf [0]);
  assign sca1_1_1_argbuf_d = (\writeCTf''''''''''''lizzieLet67_1_argbuf_rwb_bufchan_buf [0] ? \writeCTf''''''''''''lizzieLet67_1_argbuf_rwb_bufchan_buf  :
                              \writeCTf''''''''''''lizzieLet67_1_argbuf_rwb_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf''''''''''''lizzieLet67_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                     1'd0};
    else
      if ((sca1_1_1_argbuf_r && \writeCTf''''''''''''lizzieLet67_1_argbuf_rwb_bufchan_buf [0]))
        \writeCTf''''''''''''lizzieLet67_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                       1'd0};
      else if (((! sca1_1_1_argbuf_r) && (! \writeCTf''''''''''''lizzieLet67_1_argbuf_rwb_bufchan_buf [0])))
        \writeCTf''''''''''''lizzieLet67_1_argbuf_rwb_bufchan_buf  <= \writeCTf''''''''''''lizzieLet67_1_argbuf_rwb_bufchan_d ;
  
  /* buf (Ty Pointer_CTf'''''''''''') : (writeCTf''''''''''''lizzieLet68_1_argbuf,Pointer_CTf'''''''''''') > (writeCTf''''''''''''lizzieLet68_1_argbuf_rwb,Pointer_CTf'''''''''''') */
  \Pointer_CTf''''''''''''_t  \writeCTf''''''''''''lizzieLet68_1_argbuf_bufchan_d ;
  logic \writeCTf''''''''''''lizzieLet68_1_argbuf_bufchan_r ;
  assign \writeCTf''''''''''''lizzieLet68_1_argbuf_r  = ((! \writeCTf''''''''''''lizzieLet68_1_argbuf_bufchan_d [0]) || \writeCTf''''''''''''lizzieLet68_1_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf''''''''''''lizzieLet68_1_argbuf_bufchan_d  <= {16'd0,
                                                               1'd0};
    else
      if (\writeCTf''''''''''''lizzieLet68_1_argbuf_r )
        \writeCTf''''''''''''lizzieLet68_1_argbuf_bufchan_d  <= \writeCTf''''''''''''lizzieLet68_1_argbuf_d ;
  \Pointer_CTf''''''''''''_t  \writeCTf''''''''''''lizzieLet68_1_argbuf_bufchan_buf ;
  assign \writeCTf''''''''''''lizzieLet68_1_argbuf_bufchan_r  = (! \writeCTf''''''''''''lizzieLet68_1_argbuf_bufchan_buf [0]);
  assign \writeCTf''''''''''''lizzieLet68_1_argbuf_rwb_d  = (\writeCTf''''''''''''lizzieLet68_1_argbuf_bufchan_buf [0] ? \writeCTf''''''''''''lizzieLet68_1_argbuf_bufchan_buf  :
                                                             \writeCTf''''''''''''lizzieLet68_1_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf''''''''''''lizzieLet68_1_argbuf_bufchan_buf  <= {16'd0,
                                                                 1'd0};
    else
      if ((\writeCTf''''''''''''lizzieLet68_1_argbuf_rwb_r  && \writeCTf''''''''''''lizzieLet68_1_argbuf_bufchan_buf [0]))
        \writeCTf''''''''''''lizzieLet68_1_argbuf_bufchan_buf  <= {16'd0,
                                                                   1'd0};
      else if (((! \writeCTf''''''''''''lizzieLet68_1_argbuf_rwb_r ) && (! \writeCTf''''''''''''lizzieLet68_1_argbuf_bufchan_buf [0])))
        \writeCTf''''''''''''lizzieLet68_1_argbuf_bufchan_buf  <= \writeCTf''''''''''''lizzieLet68_1_argbuf_bufchan_d ;
  
  /* buf (Ty Pointer_CTf'''''''''''') : (writeCTf''''''''''''lizzieLet68_1_argbuf_rwb,Pointer_CTf'''''''''''') > (sca0_1_1_argbuf,Pointer_CTf'''''''''''') */
  \Pointer_CTf''''''''''''_t  \writeCTf''''''''''''lizzieLet68_1_argbuf_rwb_bufchan_d ;
  logic \writeCTf''''''''''''lizzieLet68_1_argbuf_rwb_bufchan_r ;
  assign \writeCTf''''''''''''lizzieLet68_1_argbuf_rwb_r  = ((! \writeCTf''''''''''''lizzieLet68_1_argbuf_rwb_bufchan_d [0]) || \writeCTf''''''''''''lizzieLet68_1_argbuf_rwb_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf''''''''''''lizzieLet68_1_argbuf_rwb_bufchan_d  <= {16'd0,
                                                                   1'd0};
    else
      if (\writeCTf''''''''''''lizzieLet68_1_argbuf_rwb_r )
        \writeCTf''''''''''''lizzieLet68_1_argbuf_rwb_bufchan_d  <= \writeCTf''''''''''''lizzieLet68_1_argbuf_rwb_d ;
  \Pointer_CTf''''''''''''_t  \writeCTf''''''''''''lizzieLet68_1_argbuf_rwb_bufchan_buf ;
  assign \writeCTf''''''''''''lizzieLet68_1_argbuf_rwb_bufchan_r  = (! \writeCTf''''''''''''lizzieLet68_1_argbuf_rwb_bufchan_buf [0]);
  assign sca0_1_1_argbuf_d = (\writeCTf''''''''''''lizzieLet68_1_argbuf_rwb_bufchan_buf [0] ? \writeCTf''''''''''''lizzieLet68_1_argbuf_rwb_bufchan_buf  :
                              \writeCTf''''''''''''lizzieLet68_1_argbuf_rwb_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf''''''''''''lizzieLet68_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                     1'd0};
    else
      if ((sca0_1_1_argbuf_r && \writeCTf''''''''''''lizzieLet68_1_argbuf_rwb_bufchan_buf [0]))
        \writeCTf''''''''''''lizzieLet68_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                       1'd0};
      else if (((! sca0_1_1_argbuf_r) && (! \writeCTf''''''''''''lizzieLet68_1_argbuf_rwb_bufchan_buf [0])))
        \writeCTf''''''''''''lizzieLet68_1_argbuf_rwb_bufchan_buf  <= \writeCTf''''''''''''lizzieLet68_1_argbuf_rwb_bufchan_d ;
  
  /* buf (Ty Pointer_CTf) : (writeCTflizzieLet41_1_argbuf,Pointer_CTf) > (writeCTflizzieLet41_1_argbuf_rwb,Pointer_CTf) */
  Pointer_CTf_t writeCTflizzieLet41_1_argbuf_bufchan_d;
  logic writeCTflizzieLet41_1_argbuf_bufchan_r;
  assign writeCTflizzieLet41_1_argbuf_r = ((! writeCTflizzieLet41_1_argbuf_bufchan_d[0]) || writeCTflizzieLet41_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTflizzieLet41_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCTflizzieLet41_1_argbuf_r)
        writeCTflizzieLet41_1_argbuf_bufchan_d <= writeCTflizzieLet41_1_argbuf_d;
  Pointer_CTf_t writeCTflizzieLet41_1_argbuf_bufchan_buf;
  assign writeCTflizzieLet41_1_argbuf_bufchan_r = (! writeCTflizzieLet41_1_argbuf_bufchan_buf[0]);
  assign writeCTflizzieLet41_1_argbuf_rwb_d = (writeCTflizzieLet41_1_argbuf_bufchan_buf[0] ? writeCTflizzieLet41_1_argbuf_bufchan_buf :
                                               writeCTflizzieLet41_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTflizzieLet41_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeCTflizzieLet41_1_argbuf_rwb_r && writeCTflizzieLet41_1_argbuf_bufchan_buf[0]))
        writeCTflizzieLet41_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeCTflizzieLet41_1_argbuf_rwb_r) && (! writeCTflizzieLet41_1_argbuf_bufchan_buf[0])))
        writeCTflizzieLet41_1_argbuf_bufchan_buf <= writeCTflizzieLet41_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CTf) : (writeCTflizzieLet41_1_argbuf_rwb,Pointer_CTf) > (sca3_1_argbuf,Pointer_CTf) */
  Pointer_CTf_t writeCTflizzieLet41_1_argbuf_rwb_bufchan_d;
  logic writeCTflizzieLet41_1_argbuf_rwb_bufchan_r;
  assign writeCTflizzieLet41_1_argbuf_rwb_r = ((! writeCTflizzieLet41_1_argbuf_rwb_bufchan_d[0]) || writeCTflizzieLet41_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTflizzieLet41_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCTflizzieLet41_1_argbuf_rwb_r)
        writeCTflizzieLet41_1_argbuf_rwb_bufchan_d <= writeCTflizzieLet41_1_argbuf_rwb_d;
  Pointer_CTf_t writeCTflizzieLet41_1_argbuf_rwb_bufchan_buf;
  assign writeCTflizzieLet41_1_argbuf_rwb_bufchan_r = (! writeCTflizzieLet41_1_argbuf_rwb_bufchan_buf[0]);
  assign sca3_1_argbuf_d = (writeCTflizzieLet41_1_argbuf_rwb_bufchan_buf[0] ? writeCTflizzieLet41_1_argbuf_rwb_bufchan_buf :
                            writeCTflizzieLet41_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTflizzieLet41_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((sca3_1_argbuf_r && writeCTflizzieLet41_1_argbuf_rwb_bufchan_buf[0]))
        writeCTflizzieLet41_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
      else if (((! sca3_1_argbuf_r) && (! writeCTflizzieLet41_1_argbuf_rwb_bufchan_buf[0])))
        writeCTflizzieLet41_1_argbuf_rwb_bufchan_buf <= writeCTflizzieLet41_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CTf) : (writeCTflizzieLet57_1_argbuf,Pointer_CTf) > (writeCTflizzieLet57_1_argbuf_rwb,Pointer_CTf) */
  Pointer_CTf_t writeCTflizzieLet57_1_argbuf_bufchan_d;
  logic writeCTflizzieLet57_1_argbuf_bufchan_r;
  assign writeCTflizzieLet57_1_argbuf_r = ((! writeCTflizzieLet57_1_argbuf_bufchan_d[0]) || writeCTflizzieLet57_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTflizzieLet57_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCTflizzieLet57_1_argbuf_r)
        writeCTflizzieLet57_1_argbuf_bufchan_d <= writeCTflizzieLet57_1_argbuf_d;
  Pointer_CTf_t writeCTflizzieLet57_1_argbuf_bufchan_buf;
  assign writeCTflizzieLet57_1_argbuf_bufchan_r = (! writeCTflizzieLet57_1_argbuf_bufchan_buf[0]);
  assign writeCTflizzieLet57_1_argbuf_rwb_d = (writeCTflizzieLet57_1_argbuf_bufchan_buf[0] ? writeCTflizzieLet57_1_argbuf_bufchan_buf :
                                               writeCTflizzieLet57_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTflizzieLet57_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeCTflizzieLet57_1_argbuf_rwb_r && writeCTflizzieLet57_1_argbuf_bufchan_buf[0]))
        writeCTflizzieLet57_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeCTflizzieLet57_1_argbuf_rwb_r) && (! writeCTflizzieLet57_1_argbuf_bufchan_buf[0])))
        writeCTflizzieLet57_1_argbuf_bufchan_buf <= writeCTflizzieLet57_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CTf) : (writeCTflizzieLet57_1_argbuf_rwb,Pointer_CTf) > (lizzieLet33_1_argbuf,Pointer_CTf) */
  Pointer_CTf_t writeCTflizzieLet57_1_argbuf_rwb_bufchan_d;
  logic writeCTflizzieLet57_1_argbuf_rwb_bufchan_r;
  assign writeCTflizzieLet57_1_argbuf_rwb_r = ((! writeCTflizzieLet57_1_argbuf_rwb_bufchan_d[0]) || writeCTflizzieLet57_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTflizzieLet57_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCTflizzieLet57_1_argbuf_rwb_r)
        writeCTflizzieLet57_1_argbuf_rwb_bufchan_d <= writeCTflizzieLet57_1_argbuf_rwb_d;
  Pointer_CTf_t writeCTflizzieLet57_1_argbuf_rwb_bufchan_buf;
  assign writeCTflizzieLet57_1_argbuf_rwb_bufchan_r = (! writeCTflizzieLet57_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet33_1_argbuf_d = (writeCTflizzieLet57_1_argbuf_rwb_bufchan_buf[0] ? writeCTflizzieLet57_1_argbuf_rwb_bufchan_buf :
                                   writeCTflizzieLet57_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTflizzieLet57_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet33_1_argbuf_r && writeCTflizzieLet57_1_argbuf_rwb_bufchan_buf[0]))
        writeCTflizzieLet57_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet33_1_argbuf_r) && (! writeCTflizzieLet57_1_argbuf_rwb_bufchan_buf[0])))
        writeCTflizzieLet57_1_argbuf_rwb_bufchan_buf <= writeCTflizzieLet57_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CTf) : (writeCTflizzieLet61_1_argbuf,Pointer_CTf) > (writeCTflizzieLet61_1_argbuf_rwb,Pointer_CTf) */
  Pointer_CTf_t writeCTflizzieLet61_1_argbuf_bufchan_d;
  logic writeCTflizzieLet61_1_argbuf_bufchan_r;
  assign writeCTflizzieLet61_1_argbuf_r = ((! writeCTflizzieLet61_1_argbuf_bufchan_d[0]) || writeCTflizzieLet61_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTflizzieLet61_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCTflizzieLet61_1_argbuf_r)
        writeCTflizzieLet61_1_argbuf_bufchan_d <= writeCTflizzieLet61_1_argbuf_d;
  Pointer_CTf_t writeCTflizzieLet61_1_argbuf_bufchan_buf;
  assign writeCTflizzieLet61_1_argbuf_bufchan_r = (! writeCTflizzieLet61_1_argbuf_bufchan_buf[0]);
  assign writeCTflizzieLet61_1_argbuf_rwb_d = (writeCTflizzieLet61_1_argbuf_bufchan_buf[0] ? writeCTflizzieLet61_1_argbuf_bufchan_buf :
                                               writeCTflizzieLet61_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTflizzieLet61_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeCTflizzieLet61_1_argbuf_rwb_r && writeCTflizzieLet61_1_argbuf_bufchan_buf[0]))
        writeCTflizzieLet61_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeCTflizzieLet61_1_argbuf_rwb_r) && (! writeCTflizzieLet61_1_argbuf_bufchan_buf[0])))
        writeCTflizzieLet61_1_argbuf_bufchan_buf <= writeCTflizzieLet61_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CTf) : (writeCTflizzieLet61_1_argbuf_rwb,Pointer_CTf) > (sca2_1_argbuf,Pointer_CTf) */
  Pointer_CTf_t writeCTflizzieLet61_1_argbuf_rwb_bufchan_d;
  logic writeCTflizzieLet61_1_argbuf_rwb_bufchan_r;
  assign writeCTflizzieLet61_1_argbuf_rwb_r = ((! writeCTflizzieLet61_1_argbuf_rwb_bufchan_d[0]) || writeCTflizzieLet61_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTflizzieLet61_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCTflizzieLet61_1_argbuf_rwb_r)
        writeCTflizzieLet61_1_argbuf_rwb_bufchan_d <= writeCTflizzieLet61_1_argbuf_rwb_d;
  Pointer_CTf_t writeCTflizzieLet61_1_argbuf_rwb_bufchan_buf;
  assign writeCTflizzieLet61_1_argbuf_rwb_bufchan_r = (! writeCTflizzieLet61_1_argbuf_rwb_bufchan_buf[0]);
  assign sca2_1_argbuf_d = (writeCTflizzieLet61_1_argbuf_rwb_bufchan_buf[0] ? writeCTflizzieLet61_1_argbuf_rwb_bufchan_buf :
                            writeCTflizzieLet61_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTflizzieLet61_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((sca2_1_argbuf_r && writeCTflizzieLet61_1_argbuf_rwb_bufchan_buf[0]))
        writeCTflizzieLet61_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
      else if (((! sca2_1_argbuf_r) && (! writeCTflizzieLet61_1_argbuf_rwb_bufchan_buf[0])))
        writeCTflizzieLet61_1_argbuf_rwb_bufchan_buf <= writeCTflizzieLet61_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CTf) : (writeCTflizzieLet62_1_argbuf,Pointer_CTf) > (writeCTflizzieLet62_1_argbuf_rwb,Pointer_CTf) */
  Pointer_CTf_t writeCTflizzieLet62_1_argbuf_bufchan_d;
  logic writeCTflizzieLet62_1_argbuf_bufchan_r;
  assign writeCTflizzieLet62_1_argbuf_r = ((! writeCTflizzieLet62_1_argbuf_bufchan_d[0]) || writeCTflizzieLet62_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTflizzieLet62_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCTflizzieLet62_1_argbuf_r)
        writeCTflizzieLet62_1_argbuf_bufchan_d <= writeCTflizzieLet62_1_argbuf_d;
  Pointer_CTf_t writeCTflizzieLet62_1_argbuf_bufchan_buf;
  assign writeCTflizzieLet62_1_argbuf_bufchan_r = (! writeCTflizzieLet62_1_argbuf_bufchan_buf[0]);
  assign writeCTflizzieLet62_1_argbuf_rwb_d = (writeCTflizzieLet62_1_argbuf_bufchan_buf[0] ? writeCTflizzieLet62_1_argbuf_bufchan_buf :
                                               writeCTflizzieLet62_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTflizzieLet62_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeCTflizzieLet62_1_argbuf_rwb_r && writeCTflizzieLet62_1_argbuf_bufchan_buf[0]))
        writeCTflizzieLet62_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeCTflizzieLet62_1_argbuf_rwb_r) && (! writeCTflizzieLet62_1_argbuf_bufchan_buf[0])))
        writeCTflizzieLet62_1_argbuf_bufchan_buf <= writeCTflizzieLet62_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CTf) : (writeCTflizzieLet62_1_argbuf_rwb,Pointer_CTf) > (sca1_1_argbuf,Pointer_CTf) */
  Pointer_CTf_t writeCTflizzieLet62_1_argbuf_rwb_bufchan_d;
  logic writeCTflizzieLet62_1_argbuf_rwb_bufchan_r;
  assign writeCTflizzieLet62_1_argbuf_rwb_r = ((! writeCTflizzieLet62_1_argbuf_rwb_bufchan_d[0]) || writeCTflizzieLet62_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTflizzieLet62_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCTflizzieLet62_1_argbuf_rwb_r)
        writeCTflizzieLet62_1_argbuf_rwb_bufchan_d <= writeCTflizzieLet62_1_argbuf_rwb_d;
  Pointer_CTf_t writeCTflizzieLet62_1_argbuf_rwb_bufchan_buf;
  assign writeCTflizzieLet62_1_argbuf_rwb_bufchan_r = (! writeCTflizzieLet62_1_argbuf_rwb_bufchan_buf[0]);
  assign sca1_1_argbuf_d = (writeCTflizzieLet62_1_argbuf_rwb_bufchan_buf[0] ? writeCTflizzieLet62_1_argbuf_rwb_bufchan_buf :
                            writeCTflizzieLet62_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTflizzieLet62_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((sca1_1_argbuf_r && writeCTflizzieLet62_1_argbuf_rwb_bufchan_buf[0]))
        writeCTflizzieLet62_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
      else if (((! sca1_1_argbuf_r) && (! writeCTflizzieLet62_1_argbuf_rwb_bufchan_buf[0])))
        writeCTflizzieLet62_1_argbuf_rwb_bufchan_buf <= writeCTflizzieLet62_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CTf) : (writeCTflizzieLet63_1_argbuf,Pointer_CTf) > (writeCTflizzieLet63_1_argbuf_rwb,Pointer_CTf) */
  Pointer_CTf_t writeCTflizzieLet63_1_argbuf_bufchan_d;
  logic writeCTflizzieLet63_1_argbuf_bufchan_r;
  assign writeCTflizzieLet63_1_argbuf_r = ((! writeCTflizzieLet63_1_argbuf_bufchan_d[0]) || writeCTflizzieLet63_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTflizzieLet63_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCTflizzieLet63_1_argbuf_r)
        writeCTflizzieLet63_1_argbuf_bufchan_d <= writeCTflizzieLet63_1_argbuf_d;
  Pointer_CTf_t writeCTflizzieLet63_1_argbuf_bufchan_buf;
  assign writeCTflizzieLet63_1_argbuf_bufchan_r = (! writeCTflizzieLet63_1_argbuf_bufchan_buf[0]);
  assign writeCTflizzieLet63_1_argbuf_rwb_d = (writeCTflizzieLet63_1_argbuf_bufchan_buf[0] ? writeCTflizzieLet63_1_argbuf_bufchan_buf :
                                               writeCTflizzieLet63_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTflizzieLet63_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeCTflizzieLet63_1_argbuf_rwb_r && writeCTflizzieLet63_1_argbuf_bufchan_buf[0]))
        writeCTflizzieLet63_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeCTflizzieLet63_1_argbuf_rwb_r) && (! writeCTflizzieLet63_1_argbuf_bufchan_buf[0])))
        writeCTflizzieLet63_1_argbuf_bufchan_buf <= writeCTflizzieLet63_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CTf) : (writeCTflizzieLet63_1_argbuf_rwb,Pointer_CTf) > (sca0_1_argbuf,Pointer_CTf) */
  Pointer_CTf_t writeCTflizzieLet63_1_argbuf_rwb_bufchan_d;
  logic writeCTflizzieLet63_1_argbuf_rwb_bufchan_r;
  assign writeCTflizzieLet63_1_argbuf_rwb_r = ((! writeCTflizzieLet63_1_argbuf_rwb_bufchan_d[0]) || writeCTflizzieLet63_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTflizzieLet63_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCTflizzieLet63_1_argbuf_rwb_r)
        writeCTflizzieLet63_1_argbuf_rwb_bufchan_d <= writeCTflizzieLet63_1_argbuf_rwb_d;
  Pointer_CTf_t writeCTflizzieLet63_1_argbuf_rwb_bufchan_buf;
  assign writeCTflizzieLet63_1_argbuf_rwb_bufchan_r = (! writeCTflizzieLet63_1_argbuf_rwb_bufchan_buf[0]);
  assign sca0_1_argbuf_d = (writeCTflizzieLet63_1_argbuf_rwb_bufchan_buf[0] ? writeCTflizzieLet63_1_argbuf_rwb_bufchan_buf :
                            writeCTflizzieLet63_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTflizzieLet63_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((sca0_1_argbuf_r && writeCTflizzieLet63_1_argbuf_rwb_bufchan_buf[0]))
        writeCTflizzieLet63_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
      else if (((! sca0_1_argbuf_r) && (! writeCTflizzieLet63_1_argbuf_rwb_bufchan_buf[0])))
        writeCTflizzieLet63_1_argbuf_rwb_bufchan_buf <= writeCTflizzieLet63_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet10_1_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet10_1_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet10_1_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet10_1_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet10_1_1_argbuf_r = ((! writeQTree_BoollizzieLet10_1_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet10_1_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet10_1_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet10_1_1_argbuf_r)
        writeQTree_BoollizzieLet10_1_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet10_1_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet10_1_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet10_1_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet10_1_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet10_1_1_argbuf_rwb_d = (writeQTree_BoollizzieLet10_1_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet10_1_1_argbuf_bufchan_buf :
                                                        writeQTree_BoollizzieLet10_1_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet10_1_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet10_1_1_argbuf_rwb_r && writeQTree_BoollizzieLet10_1_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet10_1_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet10_1_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet10_1_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet10_1_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet10_1_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet10_1_1_argbuf_rwb,Pointer_QTree_Bool) > (lizzieLet12_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet10_1_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet10_1_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet10_1_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet10_1_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet10_1_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet10_1_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                              1'd0};
    else
      if (writeQTree_BoollizzieLet10_1_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet10_1_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet10_1_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet10_1_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet10_1_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet10_1_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet12_1_argbuf_d = (writeQTree_BoollizzieLet10_1_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet10_1_1_argbuf_rwb_bufchan_buf :
                                   writeQTree_BoollizzieLet10_1_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet10_1_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
    else
      if ((lizzieLet12_1_argbuf_r && writeQTree_BoollizzieLet10_1_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet10_1_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                  1'd0};
      else if (((! lizzieLet12_1_argbuf_r) && (! writeQTree_BoollizzieLet10_1_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet10_1_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet10_1_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet11_1_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet11_1_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet11_1_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet11_1_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet11_1_1_argbuf_r = ((! writeQTree_BoollizzieLet11_1_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet11_1_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet11_1_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet11_1_1_argbuf_r)
        writeQTree_BoollizzieLet11_1_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet11_1_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet11_1_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet11_1_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet11_1_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet11_1_1_argbuf_rwb_d = (writeQTree_BoollizzieLet11_1_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet11_1_1_argbuf_bufchan_buf :
                                                        writeQTree_BoollizzieLet11_1_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet11_1_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet11_1_1_argbuf_rwb_r && writeQTree_BoollizzieLet11_1_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet11_1_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet11_1_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet11_1_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet11_1_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet11_1_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet11_1_1_argbuf_rwb,Pointer_QTree_Bool) > (lizzieLet13_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet11_1_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet11_1_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet11_1_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet11_1_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet11_1_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet11_1_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                              1'd0};
    else
      if (writeQTree_BoollizzieLet11_1_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet11_1_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet11_1_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet11_1_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet11_1_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet11_1_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet13_1_argbuf_d = (writeQTree_BoollizzieLet11_1_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet11_1_1_argbuf_rwb_bufchan_buf :
                                   writeQTree_BoollizzieLet11_1_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet11_1_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
    else
      if ((lizzieLet13_1_argbuf_r && writeQTree_BoollizzieLet11_1_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet11_1_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                  1'd0};
      else if (((! lizzieLet13_1_argbuf_r) && (! writeQTree_BoollizzieLet11_1_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet11_1_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet11_1_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet12_1_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet12_1_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet12_1_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet12_1_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet12_1_1_argbuf_r = ((! writeQTree_BoollizzieLet12_1_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet12_1_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet12_1_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet12_1_1_argbuf_r)
        writeQTree_BoollizzieLet12_1_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet12_1_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet12_1_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet12_1_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet12_1_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet12_1_1_argbuf_rwb_d = (writeQTree_BoollizzieLet12_1_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet12_1_1_argbuf_bufchan_buf :
                                                        writeQTree_BoollizzieLet12_1_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet12_1_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet12_1_1_argbuf_rwb_r && writeQTree_BoollizzieLet12_1_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet12_1_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet12_1_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet12_1_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet12_1_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet12_1_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet12_1_1_argbuf_rwb,Pointer_QTree_Bool) > (lizzieLet14_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet12_1_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet12_1_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet12_1_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet12_1_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet12_1_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet12_1_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                              1'd0};
    else
      if (writeQTree_BoollizzieLet12_1_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet12_1_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet12_1_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet12_1_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet12_1_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet12_1_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet14_1_argbuf_d = (writeQTree_BoollizzieLet12_1_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet12_1_1_argbuf_rwb_bufchan_buf :
                                   writeQTree_BoollizzieLet12_1_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet12_1_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
    else
      if ((lizzieLet14_1_argbuf_r && writeQTree_BoollizzieLet12_1_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet12_1_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                  1'd0};
      else if (((! lizzieLet14_1_argbuf_r) && (! writeQTree_BoollizzieLet12_1_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet12_1_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet12_1_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet15_1_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet15_1_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet15_1_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet15_1_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet15_1_1_argbuf_r = ((! writeQTree_BoollizzieLet15_1_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet15_1_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet15_1_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet15_1_1_argbuf_r)
        writeQTree_BoollizzieLet15_1_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet15_1_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet15_1_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet15_1_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet15_1_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet15_1_1_argbuf_rwb_d = (writeQTree_BoollizzieLet15_1_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet15_1_1_argbuf_bufchan_buf :
                                                        writeQTree_BoollizzieLet15_1_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet15_1_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet15_1_1_argbuf_rwb_r && writeQTree_BoollizzieLet15_1_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet15_1_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet15_1_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet15_1_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet15_1_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet15_1_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet15_1_1_argbuf_rwb,Pointer_QTree_Bool) > (lizzieLet15_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet15_1_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet15_1_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet15_1_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet15_1_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet15_1_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet15_1_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                              1'd0};
    else
      if (writeQTree_BoollizzieLet15_1_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet15_1_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet15_1_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet15_1_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet15_1_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet15_1_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet15_1_argbuf_d = (writeQTree_BoollizzieLet15_1_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet15_1_1_argbuf_rwb_bufchan_buf :
                                   writeQTree_BoollizzieLet15_1_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet15_1_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
    else
      if ((lizzieLet15_1_argbuf_r && writeQTree_BoollizzieLet15_1_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet15_1_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                  1'd0};
      else if (((! lizzieLet15_1_argbuf_r) && (! writeQTree_BoollizzieLet15_1_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet15_1_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet15_1_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet18_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet18_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet18_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet18_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet18_1_argbuf_r = ((! writeQTree_BoollizzieLet18_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet18_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet18_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet18_1_argbuf_r)
        writeQTree_BoollizzieLet18_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet18_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet18_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet18_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet18_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet18_1_argbuf_rwb_d = (writeQTree_BoollizzieLet18_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet18_1_argbuf_bufchan_buf :
                                                      writeQTree_BoollizzieLet18_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet18_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet18_1_argbuf_rwb_r && writeQTree_BoollizzieLet18_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet18_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet18_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet18_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet18_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet18_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet18_1_argbuf_rwb,Pointer_QTree_Bool) > (lizzieLet16_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet18_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet18_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet18_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet18_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet18_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet18_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet18_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet18_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet18_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet18_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet18_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet18_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet16_1_1_argbuf_d = (writeQTree_BoollizzieLet18_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet18_1_argbuf_rwb_bufchan_buf :
                                     writeQTree_BoollizzieLet18_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet18_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                              1'd0};
    else
      if ((lizzieLet16_1_1_argbuf_r && writeQTree_BoollizzieLet18_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet18_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
      else if (((! lizzieLet16_1_1_argbuf_r) && (! writeQTree_BoollizzieLet18_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet18_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet18_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet19_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet19_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet19_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet19_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet19_1_argbuf_r = ((! writeQTree_BoollizzieLet19_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet19_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet19_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet19_1_argbuf_r)
        writeQTree_BoollizzieLet19_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet19_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet19_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet19_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet19_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet19_1_argbuf_rwb_d = (writeQTree_BoollizzieLet19_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet19_1_argbuf_bufchan_buf :
                                                      writeQTree_BoollizzieLet19_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet19_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet19_1_argbuf_rwb_r && writeQTree_BoollizzieLet19_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet19_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet19_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet19_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet19_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet19_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet19_1_argbuf_rwb,Pointer_QTree_Bool) > (lizzieLet17_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet19_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet19_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet19_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet19_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet19_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet19_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet19_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet19_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet19_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet19_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet19_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet19_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet17_1_1_argbuf_d = (writeQTree_BoollizzieLet19_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet19_1_argbuf_rwb_bufchan_buf :
                                     writeQTree_BoollizzieLet19_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet19_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                              1'd0};
    else
      if ((lizzieLet17_1_1_argbuf_r && writeQTree_BoollizzieLet19_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet19_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
      else if (((! lizzieLet17_1_1_argbuf_r) && (! writeQTree_BoollizzieLet19_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet19_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet19_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet23_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet23_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet23_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet23_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet23_1_argbuf_r = ((! writeQTree_BoollizzieLet23_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet23_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet23_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet23_1_argbuf_r)
        writeQTree_BoollizzieLet23_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet23_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet23_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet23_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet23_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet23_1_argbuf_rwb_d = (writeQTree_BoollizzieLet23_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet23_1_argbuf_bufchan_buf :
                                                      writeQTree_BoollizzieLet23_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet23_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet23_1_argbuf_rwb_r && writeQTree_BoollizzieLet23_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet23_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet23_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet23_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet23_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet23_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet23_1_argbuf_rwb,Pointer_QTree_Bool) > (lizzieLet18_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet23_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet23_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet23_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet23_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet23_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet23_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet23_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet23_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet23_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet23_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet23_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet23_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet18_1_1_argbuf_d = (writeQTree_BoollizzieLet23_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet23_1_argbuf_rwb_bufchan_buf :
                                     writeQTree_BoollizzieLet23_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet23_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                              1'd0};
    else
      if ((lizzieLet18_1_1_argbuf_r && writeQTree_BoollizzieLet23_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet23_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
      else if (((! lizzieLet18_1_1_argbuf_r) && (! writeQTree_BoollizzieLet23_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet23_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet23_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet24_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet24_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet24_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet24_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet24_1_argbuf_r = ((! writeQTree_BoollizzieLet24_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet24_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet24_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet24_1_argbuf_r)
        writeQTree_BoollizzieLet24_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet24_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet24_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet24_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet24_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet24_1_argbuf_rwb_d = (writeQTree_BoollizzieLet24_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet24_1_argbuf_bufchan_buf :
                                                      writeQTree_BoollizzieLet24_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet24_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet24_1_argbuf_rwb_r && writeQTree_BoollizzieLet24_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet24_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet24_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet24_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet24_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet24_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet24_1_argbuf_rwb,Pointer_QTree_Bool) > (lizzieLet19_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet24_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet24_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet24_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet24_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet24_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet24_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet24_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet24_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet24_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet24_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet24_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet24_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet19_1_1_argbuf_d = (writeQTree_BoollizzieLet24_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet24_1_argbuf_rwb_bufchan_buf :
                                     writeQTree_BoollizzieLet24_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet24_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                              1'd0};
    else
      if ((lizzieLet19_1_1_argbuf_r && writeQTree_BoollizzieLet24_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet24_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
      else if (((! lizzieLet19_1_1_argbuf_r) && (! writeQTree_BoollizzieLet24_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet24_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet24_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet28_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet28_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet28_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet28_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet28_1_argbuf_r = ((! writeQTree_BoollizzieLet28_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet28_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet28_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet28_1_argbuf_r)
        writeQTree_BoollizzieLet28_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet28_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet28_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet28_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet28_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet28_1_argbuf_rwb_d = (writeQTree_BoollizzieLet28_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet28_1_argbuf_bufchan_buf :
                                                      writeQTree_BoollizzieLet28_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet28_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet28_1_argbuf_rwb_r && writeQTree_BoollizzieLet28_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet28_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet28_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet28_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet28_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet28_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet28_1_argbuf_rwb,Pointer_QTree_Bool) > (lizzieLet20_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet28_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet28_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet28_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet28_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet28_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet28_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet28_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet28_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet28_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet28_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet28_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet28_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet20_1_argbuf_d = (writeQTree_BoollizzieLet28_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet28_1_argbuf_rwb_bufchan_buf :
                                   writeQTree_BoollizzieLet28_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet28_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                              1'd0};
    else
      if ((lizzieLet20_1_argbuf_r && writeQTree_BoollizzieLet28_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet28_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
      else if (((! lizzieLet20_1_argbuf_r) && (! writeQTree_BoollizzieLet28_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet28_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet28_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet29_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet29_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet29_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet29_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet29_1_argbuf_r = ((! writeQTree_BoollizzieLet29_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet29_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet29_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet29_1_argbuf_r)
        writeQTree_BoollizzieLet29_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet29_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet29_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet29_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet29_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet29_1_argbuf_rwb_d = (writeQTree_BoollizzieLet29_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet29_1_argbuf_bufchan_buf :
                                                      writeQTree_BoollizzieLet29_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet29_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet29_1_argbuf_rwb_r && writeQTree_BoollizzieLet29_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet29_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet29_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet29_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet29_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet29_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet29_1_argbuf_rwb,Pointer_QTree_Bool) > (lizzieLet21_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet29_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet29_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet29_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet29_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet29_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet29_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet29_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet29_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet29_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet29_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet29_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet29_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet21_1_1_argbuf_d = (writeQTree_BoollizzieLet29_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet29_1_argbuf_rwb_bufchan_buf :
                                     writeQTree_BoollizzieLet29_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet29_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                              1'd0};
    else
      if ((lizzieLet21_1_1_argbuf_r && writeQTree_BoollizzieLet29_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet29_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
      else if (((! lizzieLet21_1_1_argbuf_r) && (! writeQTree_BoollizzieLet29_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet29_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet29_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet30_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet30_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet30_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet30_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet30_1_argbuf_r = ((! writeQTree_BoollizzieLet30_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet30_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet30_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet30_1_argbuf_r)
        writeQTree_BoollizzieLet30_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet30_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet30_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet30_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet30_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet30_1_argbuf_rwb_d = (writeQTree_BoollizzieLet30_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet30_1_argbuf_bufchan_buf :
                                                      writeQTree_BoollizzieLet30_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet30_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet30_1_argbuf_rwb_r && writeQTree_BoollizzieLet30_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet30_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet30_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet30_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet30_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet30_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet30_1_argbuf_rwb,Pointer_QTree_Bool) > (lizzieLet22_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet30_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet30_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet30_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet30_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet30_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet30_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet30_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet30_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet30_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet30_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet30_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet30_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet22_1_1_argbuf_d = (writeQTree_BoollizzieLet30_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet30_1_argbuf_rwb_bufchan_buf :
                                     writeQTree_BoollizzieLet30_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet30_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                              1'd0};
    else
      if ((lizzieLet22_1_1_argbuf_r && writeQTree_BoollizzieLet30_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet30_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
      else if (((! lizzieLet22_1_1_argbuf_r) && (! writeQTree_BoollizzieLet30_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet30_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet30_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet31_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet31_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet31_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet31_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet31_1_argbuf_r = ((! writeQTree_BoollizzieLet31_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet31_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet31_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet31_1_argbuf_r)
        writeQTree_BoollizzieLet31_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet31_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet31_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet31_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet31_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet31_1_argbuf_rwb_d = (writeQTree_BoollizzieLet31_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet31_1_argbuf_bufchan_buf :
                                                      writeQTree_BoollizzieLet31_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet31_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet31_1_argbuf_rwb_r && writeQTree_BoollizzieLet31_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet31_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet31_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet31_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet31_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet31_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet31_1_argbuf_rwb,Pointer_QTree_Bool) > (lizzieLet23_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet31_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet31_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet31_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet31_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet31_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet31_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet31_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet31_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet31_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet31_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet31_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet31_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet23_1_1_argbuf_d = (writeQTree_BoollizzieLet31_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet31_1_argbuf_rwb_bufchan_buf :
                                     writeQTree_BoollizzieLet31_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet31_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                              1'd0};
    else
      if ((lizzieLet23_1_1_argbuf_r && writeQTree_BoollizzieLet31_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet31_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
      else if (((! lizzieLet23_1_1_argbuf_r) && (! writeQTree_BoollizzieLet31_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet31_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet31_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet34_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet34_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet34_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet34_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet34_1_argbuf_r = ((! writeQTree_BoollizzieLet34_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet34_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet34_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet34_1_argbuf_r)
        writeQTree_BoollizzieLet34_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet34_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet34_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet34_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet34_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet34_1_argbuf_rwb_d = (writeQTree_BoollizzieLet34_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet34_1_argbuf_bufchan_buf :
                                                      writeQTree_BoollizzieLet34_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet34_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet34_1_argbuf_rwb_r && writeQTree_BoollizzieLet34_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet34_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet34_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet34_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet34_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet34_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet34_1_argbuf_rwb,Pointer_QTree_Bool) > (lizzieLet24_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet34_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet34_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet34_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet34_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet34_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet34_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet34_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet34_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet34_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet34_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet34_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet34_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet24_1_1_argbuf_d = (writeQTree_BoollizzieLet34_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet34_1_argbuf_rwb_bufchan_buf :
                                     writeQTree_BoollizzieLet34_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet34_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                              1'd0};
    else
      if ((lizzieLet24_1_1_argbuf_r && writeQTree_BoollizzieLet34_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet34_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
      else if (((! lizzieLet24_1_1_argbuf_r) && (! writeQTree_BoollizzieLet34_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet34_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet34_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet35_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet35_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet35_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet35_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet35_1_argbuf_r = ((! writeQTree_BoollizzieLet35_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet35_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet35_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet35_1_argbuf_r)
        writeQTree_BoollizzieLet35_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet35_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet35_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet35_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet35_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet35_1_argbuf_rwb_d = (writeQTree_BoollizzieLet35_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet35_1_argbuf_bufchan_buf :
                                                      writeQTree_BoollizzieLet35_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet35_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet35_1_argbuf_rwb_r && writeQTree_BoollizzieLet35_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet35_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet35_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet35_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet35_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet35_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet35_1_argbuf_rwb,Pointer_QTree_Bool) > (lizzieLet25_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet35_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet35_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet35_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet35_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet35_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet35_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet35_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet35_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet35_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet35_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet35_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet35_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet25_1_argbuf_d = (writeQTree_BoollizzieLet35_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet35_1_argbuf_rwb_bufchan_buf :
                                   writeQTree_BoollizzieLet35_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet35_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                              1'd0};
    else
      if ((lizzieLet25_1_argbuf_r && writeQTree_BoollizzieLet35_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet35_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
      else if (((! lizzieLet25_1_argbuf_r) && (! writeQTree_BoollizzieLet35_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet35_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet35_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet36_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet36_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet36_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet36_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet36_1_argbuf_r = ((! writeQTree_BoollizzieLet36_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet36_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet36_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet36_1_argbuf_r)
        writeQTree_BoollizzieLet36_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet36_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet36_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet36_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet36_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet36_1_argbuf_rwb_d = (writeQTree_BoollizzieLet36_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet36_1_argbuf_bufchan_buf :
                                                      writeQTree_BoollizzieLet36_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet36_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet36_1_argbuf_rwb_r && writeQTree_BoollizzieLet36_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet36_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet36_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet36_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet36_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet36_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet36_1_argbuf_rwb,Pointer_QTree_Bool) > (lizzieLet26_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet36_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet36_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet36_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet36_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet36_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet36_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet36_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet36_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet36_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet36_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet36_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet36_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet26_1_1_argbuf_d = (writeQTree_BoollizzieLet36_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet36_1_argbuf_rwb_bufchan_buf :
                                     writeQTree_BoollizzieLet36_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet36_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                              1'd0};
    else
      if ((lizzieLet26_1_1_argbuf_r && writeQTree_BoollizzieLet36_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet36_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
      else if (((! lizzieLet26_1_1_argbuf_r) && (! writeQTree_BoollizzieLet36_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet36_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet36_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet37_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet37_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet37_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet37_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet37_1_argbuf_r = ((! writeQTree_BoollizzieLet37_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet37_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet37_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet37_1_argbuf_r)
        writeQTree_BoollizzieLet37_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet37_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet37_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet37_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet37_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet37_1_argbuf_rwb_d = (writeQTree_BoollizzieLet37_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet37_1_argbuf_bufchan_buf :
                                                      writeQTree_BoollizzieLet37_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet37_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet37_1_argbuf_rwb_r && writeQTree_BoollizzieLet37_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet37_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet37_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet37_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet37_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet37_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet37_1_argbuf_rwb,Pointer_QTree_Bool) > (lizzieLet27_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet37_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet37_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet37_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet37_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet37_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet37_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet37_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet37_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet37_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet37_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet37_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet37_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet27_1_1_argbuf_d = (writeQTree_BoollizzieLet37_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet37_1_argbuf_rwb_bufchan_buf :
                                     writeQTree_BoollizzieLet37_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet37_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                              1'd0};
    else
      if ((lizzieLet27_1_1_argbuf_r && writeQTree_BoollizzieLet37_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet37_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
      else if (((! lizzieLet27_1_1_argbuf_r) && (! writeQTree_BoollizzieLet37_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet37_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet37_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet39_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet39_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet39_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet39_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet39_1_argbuf_r = ((! writeQTree_BoollizzieLet39_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet39_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet39_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet39_1_argbuf_r)
        writeQTree_BoollizzieLet39_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet39_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet39_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet39_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet39_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet39_1_argbuf_rwb_d = (writeQTree_BoollizzieLet39_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet39_1_argbuf_bufchan_buf :
                                                      writeQTree_BoollizzieLet39_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet39_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet39_1_argbuf_rwb_r && writeQTree_BoollizzieLet39_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet39_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet39_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet39_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet39_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet39_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet39_1_argbuf_rwb,Pointer_QTree_Bool) > (lizzieLet28_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet39_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet39_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet39_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet39_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet39_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet39_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet39_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet39_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet39_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet39_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet39_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet39_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet28_1_1_argbuf_d = (writeQTree_BoollizzieLet39_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet39_1_argbuf_rwb_bufchan_buf :
                                     writeQTree_BoollizzieLet39_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet39_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                              1'd0};
    else
      if ((lizzieLet28_1_1_argbuf_r && writeQTree_BoollizzieLet39_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet39_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
      else if (((! lizzieLet28_1_1_argbuf_r) && (! writeQTree_BoollizzieLet39_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet39_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet39_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet3_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet3_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet3_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet3_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet3_1_argbuf_r = ((! writeQTree_BoollizzieLet3_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet3_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet3_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet3_1_argbuf_r)
        writeQTree_BoollizzieLet3_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet3_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet3_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet3_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet3_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet3_1_argbuf_rwb_d = (writeQTree_BoollizzieLet3_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet3_1_argbuf_bufchan_buf :
                                                     writeQTree_BoollizzieLet3_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet3_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet3_1_argbuf_rwb_r && writeQTree_BoollizzieLet3_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet3_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet3_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet3_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet3_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet3_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet3_1_argbuf_rwb,Pointer_QTree_Bool) > (lizzieLet8_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet3_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet3_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet3_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet3_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet3_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet3_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet3_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet3_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet3_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet3_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet3_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet3_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet8_1_argbuf_d = (writeQTree_BoollizzieLet3_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet3_1_argbuf_rwb_bufchan_buf :
                                  writeQTree_BoollizzieLet3_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet3_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((lizzieLet8_1_argbuf_r && writeQTree_BoollizzieLet3_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet3_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! lizzieLet8_1_argbuf_r) && (! writeQTree_BoollizzieLet3_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet3_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet3_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet40_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet40_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet40_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet40_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet40_1_argbuf_r = ((! writeQTree_BoollizzieLet40_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet40_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet40_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet40_1_argbuf_r)
        writeQTree_BoollizzieLet40_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet40_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet40_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet40_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet40_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet40_1_argbuf_rwb_d = (writeQTree_BoollizzieLet40_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet40_1_argbuf_bufchan_buf :
                                                      writeQTree_BoollizzieLet40_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet40_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet40_1_argbuf_rwb_r && writeQTree_BoollizzieLet40_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet40_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet40_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet40_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet40_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet40_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet40_1_argbuf_rwb,Pointer_QTree_Bool) > (lizzieLet29_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet40_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet40_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet40_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet40_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet40_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet40_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet40_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet40_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet40_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet40_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet40_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet40_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet29_1_1_argbuf_d = (writeQTree_BoollizzieLet40_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet40_1_argbuf_rwb_bufchan_buf :
                                     writeQTree_BoollizzieLet40_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet40_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                              1'd0};
    else
      if ((lizzieLet29_1_1_argbuf_r && writeQTree_BoollizzieLet40_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet40_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
      else if (((! lizzieLet29_1_1_argbuf_r) && (! writeQTree_BoollizzieLet40_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet40_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet40_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet42_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet42_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet42_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet42_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet42_1_argbuf_r = ((! writeQTree_BoollizzieLet42_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet42_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet42_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet42_1_argbuf_r)
        writeQTree_BoollizzieLet42_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet42_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet42_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet42_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet42_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet42_1_argbuf_rwb_d = (writeQTree_BoollizzieLet42_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet42_1_argbuf_bufchan_buf :
                                                      writeQTree_BoollizzieLet42_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet42_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet42_1_argbuf_rwb_r && writeQTree_BoollizzieLet42_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet42_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet42_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet42_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet42_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet42_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet42_1_argbuf_rwb,Pointer_QTree_Bool) > (lizzieLet30_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet42_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet42_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet42_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet42_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet42_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet42_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet42_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet42_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet42_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet42_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet42_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet42_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet30_1_1_argbuf_d = (writeQTree_BoollizzieLet42_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet42_1_argbuf_rwb_bufchan_buf :
                                     writeQTree_BoollizzieLet42_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet42_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                              1'd0};
    else
      if ((lizzieLet30_1_1_argbuf_r && writeQTree_BoollizzieLet42_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet42_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
      else if (((! lizzieLet30_1_1_argbuf_r) && (! writeQTree_BoollizzieLet42_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet42_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet42_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet43_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet43_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet43_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet43_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet43_1_argbuf_r = ((! writeQTree_BoollizzieLet43_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet43_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet43_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet43_1_argbuf_r)
        writeQTree_BoollizzieLet43_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet43_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet43_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet43_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet43_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet43_1_argbuf_rwb_d = (writeQTree_BoollizzieLet43_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet43_1_argbuf_bufchan_buf :
                                                      writeQTree_BoollizzieLet43_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet43_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet43_1_argbuf_rwb_r && writeQTree_BoollizzieLet43_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet43_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet43_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet43_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet43_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet43_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet43_1_argbuf_rwb,Pointer_QTree_Bool) > (lizzieLet31_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet43_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet43_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet43_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet43_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet43_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet43_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet43_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet43_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet43_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet43_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet43_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet43_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet31_1_1_argbuf_d = (writeQTree_BoollizzieLet43_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet43_1_argbuf_rwb_bufchan_buf :
                                     writeQTree_BoollizzieLet43_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet43_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                              1'd0};
    else
      if ((lizzieLet31_1_1_argbuf_r && writeQTree_BoollizzieLet43_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet43_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
      else if (((! lizzieLet31_1_1_argbuf_r) && (! writeQTree_BoollizzieLet43_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet43_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet43_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet44_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet44_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet44_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet44_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet44_1_argbuf_r = ((! writeQTree_BoollizzieLet44_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet44_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet44_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet44_1_argbuf_r)
        writeQTree_BoollizzieLet44_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet44_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet44_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet44_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet44_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet44_1_argbuf_rwb_d = (writeQTree_BoollizzieLet44_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet44_1_argbuf_bufchan_buf :
                                                      writeQTree_BoollizzieLet44_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet44_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet44_1_argbuf_rwb_r && writeQTree_BoollizzieLet44_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet44_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet44_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet44_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet44_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet44_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet44_1_argbuf_rwb,Pointer_QTree_Bool) > (lizzieLet32_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet44_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet44_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet44_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet44_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet44_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet44_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet44_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet44_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet44_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet44_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet44_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet44_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet32_1_argbuf_d = (writeQTree_BoollizzieLet44_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet44_1_argbuf_rwb_bufchan_buf :
                                   writeQTree_BoollizzieLet44_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet44_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                              1'd0};
    else
      if ((lizzieLet32_1_argbuf_r && writeQTree_BoollizzieLet44_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet44_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
      else if (((! lizzieLet32_1_argbuf_r) && (! writeQTree_BoollizzieLet44_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet44_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet44_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet47_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet47_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet47_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet47_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet47_1_argbuf_r = ((! writeQTree_BoollizzieLet47_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet47_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet47_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet47_1_argbuf_r)
        writeQTree_BoollizzieLet47_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet47_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet47_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet47_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet47_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet47_1_argbuf_rwb_d = (writeQTree_BoollizzieLet47_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet47_1_argbuf_bufchan_buf :
                                                      writeQTree_BoollizzieLet47_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet47_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet47_1_argbuf_rwb_r && writeQTree_BoollizzieLet47_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet47_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet47_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet47_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet47_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet47_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet47_1_argbuf_rwb,Pointer_QTree_Bool) > (lizzieLet1_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet47_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet47_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet47_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet47_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet47_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet47_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet47_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet47_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet47_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet47_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet47_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet47_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet1_1_1_argbuf_d = (writeQTree_BoollizzieLet47_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet47_1_argbuf_rwb_bufchan_buf :
                                    writeQTree_BoollizzieLet47_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet47_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                              1'd0};
    else
      if ((lizzieLet1_1_1_argbuf_r && writeQTree_BoollizzieLet47_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet47_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
      else if (((! lizzieLet1_1_1_argbuf_r) && (! writeQTree_BoollizzieLet47_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet47_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet47_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet50_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet50_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet50_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet50_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet50_1_argbuf_r = ((! writeQTree_BoollizzieLet50_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet50_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet50_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet50_1_argbuf_r)
        writeQTree_BoollizzieLet50_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet50_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet50_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet50_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet50_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet50_1_argbuf_rwb_d = (writeQTree_BoollizzieLet50_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet50_1_argbuf_bufchan_buf :
                                                      writeQTree_BoollizzieLet50_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet50_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet50_1_argbuf_rwb_r && writeQTree_BoollizzieLet50_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet50_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet50_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet50_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet50_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet50_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet50_1_argbuf_rwb,Pointer_QTree_Bool) > (lizzieLet2_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet50_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet50_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet50_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet50_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet50_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet50_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet50_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet50_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet50_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet50_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet50_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet50_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet2_1_1_argbuf_d = (writeQTree_BoollizzieLet50_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet50_1_argbuf_rwb_bufchan_buf :
                                    writeQTree_BoollizzieLet50_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet50_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                              1'd0};
    else
      if ((lizzieLet2_1_1_argbuf_r && writeQTree_BoollizzieLet50_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet50_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
      else if (((! lizzieLet2_1_1_argbuf_r) && (! writeQTree_BoollizzieLet50_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet50_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet50_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet51_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet51_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet51_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet51_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet51_1_argbuf_r = ((! writeQTree_BoollizzieLet51_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet51_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet51_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet51_1_argbuf_r)
        writeQTree_BoollizzieLet51_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet51_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet51_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet51_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet51_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet51_1_argbuf_rwb_d = (writeQTree_BoollizzieLet51_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet51_1_argbuf_bufchan_buf :
                                                      writeQTree_BoollizzieLet51_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet51_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet51_1_argbuf_rwb_r && writeQTree_BoollizzieLet51_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet51_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet51_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet51_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet51_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet51_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet51_1_argbuf_rwb,Pointer_QTree_Bool) > (lizzieLet3_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet51_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet51_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet51_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet51_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet51_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet51_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet51_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet51_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet51_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet51_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet51_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet51_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet3_1_1_argbuf_d = (writeQTree_BoollizzieLet51_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet51_1_argbuf_rwb_bufchan_buf :
                                    writeQTree_BoollizzieLet51_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet51_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                              1'd0};
    else
      if ((lizzieLet3_1_1_argbuf_r && writeQTree_BoollizzieLet51_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet51_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
      else if (((! lizzieLet3_1_1_argbuf_r) && (! writeQTree_BoollizzieLet51_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet51_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet51_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet53_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet53_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet53_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet53_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet53_1_argbuf_r = ((! writeQTree_BoollizzieLet53_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet53_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet53_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet53_1_argbuf_r)
        writeQTree_BoollizzieLet53_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet53_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet53_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet53_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet53_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet53_1_argbuf_rwb_d = (writeQTree_BoollizzieLet53_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet53_1_argbuf_bufchan_buf :
                                                      writeQTree_BoollizzieLet53_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet53_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet53_1_argbuf_rwb_r && writeQTree_BoollizzieLet53_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet53_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet53_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet53_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet53_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet53_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet53_1_argbuf_rwb,Pointer_QTree_Bool) > (lizzieLet4_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet53_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet53_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet53_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet53_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet53_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet53_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet53_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet53_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet53_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet53_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet53_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet53_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet4_1_1_argbuf_d = (writeQTree_BoollizzieLet53_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet53_1_argbuf_rwb_bufchan_buf :
                                    writeQTree_BoollizzieLet53_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet53_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                              1'd0};
    else
      if ((lizzieLet4_1_1_argbuf_r && writeQTree_BoollizzieLet53_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet53_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
      else if (((! lizzieLet4_1_1_argbuf_r) && (! writeQTree_BoollizzieLet53_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet53_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet53_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet55_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet55_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet55_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet55_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet55_1_argbuf_r = ((! writeQTree_BoollizzieLet55_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet55_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet55_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet55_1_argbuf_r)
        writeQTree_BoollizzieLet55_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet55_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet55_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet55_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet55_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet55_1_argbuf_rwb_d = (writeQTree_BoollizzieLet55_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet55_1_argbuf_bufchan_buf :
                                                      writeQTree_BoollizzieLet55_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet55_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet55_1_argbuf_rwb_r && writeQTree_BoollizzieLet55_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet55_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet55_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet55_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet55_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet55_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet55_1_argbuf_rwb,Pointer_QTree_Bool) > (lizzieLet5_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet55_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet55_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet55_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet55_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet55_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet55_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet55_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet55_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet55_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet55_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet55_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet55_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet5_1_1_argbuf_d = (writeQTree_BoollizzieLet55_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet55_1_argbuf_rwb_bufchan_buf :
                                    writeQTree_BoollizzieLet55_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet55_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                              1'd0};
    else
      if ((lizzieLet5_1_1_argbuf_r && writeQTree_BoollizzieLet55_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet55_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
      else if (((! lizzieLet5_1_1_argbuf_r) && (! writeQTree_BoollizzieLet55_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet55_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet55_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet56_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet56_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet56_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet56_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet56_1_argbuf_r = ((! writeQTree_BoollizzieLet56_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet56_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet56_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet56_1_argbuf_r)
        writeQTree_BoollizzieLet56_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet56_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet56_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet56_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet56_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet56_1_argbuf_rwb_d = (writeQTree_BoollizzieLet56_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet56_1_argbuf_bufchan_buf :
                                                      writeQTree_BoollizzieLet56_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet56_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet56_1_argbuf_rwb_r && writeQTree_BoollizzieLet56_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet56_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet56_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet56_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet56_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet56_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet56_1_argbuf_rwb,Pointer_QTree_Bool) > (lizzieLet6_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet56_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet56_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet56_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet56_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet56_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet56_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet56_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet56_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet56_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet56_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet56_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet56_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet6_1_1_argbuf_d = (writeQTree_BoollizzieLet56_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet56_1_argbuf_rwb_bufchan_buf :
                                    writeQTree_BoollizzieLet56_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet56_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                              1'd0};
    else
      if ((lizzieLet6_1_1_argbuf_r && writeQTree_BoollizzieLet56_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet56_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
      else if (((! lizzieLet6_1_1_argbuf_r) && (! writeQTree_BoollizzieLet56_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet56_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet56_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet59_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet59_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet59_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet59_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet59_1_argbuf_r = ((! writeQTree_BoollizzieLet59_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet59_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet59_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet59_1_argbuf_r)
        writeQTree_BoollizzieLet59_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet59_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet59_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet59_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet59_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet59_1_argbuf_rwb_d = (writeQTree_BoollizzieLet59_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet59_1_argbuf_bufchan_buf :
                                                      writeQTree_BoollizzieLet59_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet59_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet59_1_argbuf_rwb_r && writeQTree_BoollizzieLet59_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet59_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet59_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet59_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet59_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet59_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet64_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet64_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet64_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet64_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet64_1_argbuf_r = ((! writeQTree_BoollizzieLet64_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet64_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet64_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet64_1_argbuf_r)
        writeQTree_BoollizzieLet64_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet64_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet64_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet64_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet64_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet64_1_argbuf_rwb_d = (writeQTree_BoollizzieLet64_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet64_1_argbuf_bufchan_buf :
                                                      writeQTree_BoollizzieLet64_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet64_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet64_1_argbuf_rwb_r && writeQTree_BoollizzieLet64_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet64_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet64_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet64_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet64_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet64_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet64_1_argbuf_rwb,Pointer_QTree_Bool) > (contRet_0_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet64_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet64_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet64_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet64_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet64_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet64_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet64_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet64_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet64_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet64_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet64_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet64_1_argbuf_rwb_bufchan_buf[0]);
  assign contRet_0_1_argbuf_d = (writeQTree_BoollizzieLet64_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet64_1_argbuf_rwb_bufchan_buf :
                                 writeQTree_BoollizzieLet64_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet64_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                              1'd0};
    else
      if ((contRet_0_1_argbuf_r && writeQTree_BoollizzieLet64_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet64_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
      else if (((! contRet_0_1_argbuf_r) && (! writeQTree_BoollizzieLet64_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet64_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet64_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet69_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet69_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet69_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet69_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet69_1_argbuf_r = ((! writeQTree_BoollizzieLet69_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet69_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet69_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet69_1_argbuf_r)
        writeQTree_BoollizzieLet69_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet69_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet69_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet69_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet69_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet69_1_argbuf_rwb_d = (writeQTree_BoollizzieLet69_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet69_1_argbuf_bufchan_buf :
                                                      writeQTree_BoollizzieLet69_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet69_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet69_1_argbuf_rwb_r && writeQTree_BoollizzieLet69_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet69_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet69_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet69_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet69_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet69_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet69_1_argbuf_rwb,Pointer_QTree_Bool) > (contRet_0_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet69_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet69_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet69_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet69_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet69_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet69_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet69_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet69_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet69_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet69_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet69_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet69_1_argbuf_rwb_bufchan_buf[0]);
  assign contRet_0_1_1_argbuf_d = (writeQTree_BoollizzieLet69_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet69_1_argbuf_rwb_bufchan_buf :
                                   writeQTree_BoollizzieLet69_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet69_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                              1'd0};
    else
      if ((contRet_0_1_1_argbuf_r && writeQTree_BoollizzieLet69_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet69_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
      else if (((! contRet_0_1_1_argbuf_r) && (! writeQTree_BoollizzieLet69_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet69_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet69_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet6_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet6_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet6_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet6_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet6_1_argbuf_r = ((! writeQTree_BoollizzieLet6_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet6_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet6_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet6_1_argbuf_r)
        writeQTree_BoollizzieLet6_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet6_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet6_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet6_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet6_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet6_1_argbuf_rwb_d = (writeQTree_BoollizzieLet6_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet6_1_argbuf_bufchan_buf :
                                                     writeQTree_BoollizzieLet6_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet6_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet6_1_argbuf_rwb_r && writeQTree_BoollizzieLet6_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet6_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet6_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet6_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet6_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet6_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet6_1_argbuf_rwb,Pointer_QTree_Bool) > (lizzieLet9_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet6_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet6_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet6_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet6_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet6_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet6_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet6_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet6_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet6_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet6_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet6_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet6_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet9_1_argbuf_d = (writeQTree_BoollizzieLet6_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet6_1_argbuf_rwb_bufchan_buf :
                                  writeQTree_BoollizzieLet6_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet6_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((lizzieLet9_1_argbuf_r && writeQTree_BoollizzieLet6_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet6_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! lizzieLet9_1_argbuf_r) && (! writeQTree_BoollizzieLet6_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet6_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet6_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet7_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet7_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet7_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet7_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet7_1_argbuf_r = ((! writeQTree_BoollizzieLet7_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet7_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet7_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet7_1_argbuf_r)
        writeQTree_BoollizzieLet7_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet7_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet7_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet7_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet7_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet7_1_argbuf_rwb_d = (writeQTree_BoollizzieLet7_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet7_1_argbuf_bufchan_buf :
                                                     writeQTree_BoollizzieLet7_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet7_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet7_1_argbuf_rwb_r && writeQTree_BoollizzieLet7_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet7_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet7_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet7_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet7_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet7_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet7_1_argbuf_rwb,Pointer_QTree_Bool) > (lizzieLet10_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet7_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet7_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet7_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet7_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet7_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet7_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet7_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet7_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet7_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet7_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet7_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet7_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet10_1_argbuf_d = (writeQTree_BoollizzieLet7_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet7_1_argbuf_rwb_bufchan_buf :
                                   writeQTree_BoollizzieLet7_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet7_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((lizzieLet10_1_argbuf_r && writeQTree_BoollizzieLet7_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet7_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! lizzieLet10_1_argbuf_r) && (! writeQTree_BoollizzieLet7_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet7_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet7_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet9_1_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet9_1_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet9_1_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet9_1_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet9_1_1_argbuf_r = ((! writeQTree_BoollizzieLet9_1_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet9_1_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet9_1_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet9_1_1_argbuf_r)
        writeQTree_BoollizzieLet9_1_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet9_1_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet9_1_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet9_1_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet9_1_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet9_1_1_argbuf_rwb_d = (writeQTree_BoollizzieLet9_1_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet9_1_1_argbuf_bufchan_buf :
                                                       writeQTree_BoollizzieLet9_1_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet9_1_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet9_1_1_argbuf_rwb_r && writeQTree_BoollizzieLet9_1_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet9_1_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet9_1_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet9_1_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet9_1_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet9_1_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet9_1_1_argbuf_rwb,Pointer_QTree_Bool) > (lizzieLet11_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet9_1_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet9_1_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet9_1_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet9_1_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet9_1_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet9_1_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                             1'd0};
    else
      if (writeQTree_BoollizzieLet9_1_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet9_1_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet9_1_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet9_1_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet9_1_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet9_1_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet11_1_argbuf_d = (writeQTree_BoollizzieLet9_1_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet9_1_1_argbuf_rwb_bufchan_buf :
                                   writeQTree_BoollizzieLet9_1_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet9_1_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
    else
      if ((lizzieLet11_1_argbuf_r && writeQTree_BoollizzieLet9_1_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet9_1_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                 1'd0};
      else if (((! lizzieLet11_1_argbuf_r) && (! writeQTree_BoollizzieLet9_1_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet9_1_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet9_1_1_argbuf_rwb_bufchan_d;
endmodule