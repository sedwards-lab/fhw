`timescale 1ns/1ns
import mMaskAdd_package::*;

module mMaskAdd(
  input logic clk,
  input logic reset,
  input Go_t \\QTree_Int_src_d ,
  output logic \\QTree_Int_src_r ,
  input QTree_Int_t dummy_write_QTree_Int_d,
  output logic dummy_write_QTree_Int_r,
  input Go_t \\MaskQTree_src_d ,
  output logic \\MaskQTree_src_r ,
  input MaskQTree_t dummy_write_MaskQTree_d,
  output logic dummy_write_MaskQTree_r,
  input Go_t sourceGo_d,
  output logic sourceGo_r,
  input Pointer_MaskQTree_t m1a92_0_d,
  output logic m1a92_0_r,
  input Pointer_QTree_Int_t m2a93_1_d,
  output logic m2a93_1_r,
  input Pointer_QTree_Int_t m3a94_2_d,
  output logic m3a94_2_r,
  output \Word16#_t  forkHP1_QTree_Int_snk_dout,
  input logic forkHP1_QTree_Int_snk_rout,
  output Pointer_QTree_Int_t dummy_write_QTree_Int_sink_dout,
  input logic dummy_write_QTree_Int_sink_rout,
  output \Word16#_t  forkHP1_MaskQTree_snk_dout,
  input logic forkHP1_MaskQTree_snk_rout,
  output Pointer_MaskQTree_t dummy_write_MaskQTree_sink_dout,
  input logic dummy_write_MaskQTree_sink_rout,
  output Int_t \es_6_1I#_dout ,
  input logic \es_6_1I#_rout 
  );
  /* --define=INPUTS=((__05CQTree_Int_src, 0, 1, Go), (dummy_write_QTree_Int, 66, 73786976294838206464, QTree_Int), (__05CMaskQTree_src, 0, 1, Go), (dummy_write_MaskQTree, 66, 73786976294838206464, MaskQTree), (sourceGo, 0, 1, Go), (m1a92_0, 16, 65536, Pointer_MaskQTree), (m2a93_1, 16, 65536, Pointer_QTree_Int), (m3a94_2, 16, 65536, Pointer_QTree_Int)) */
  /* --define=TAPS=() */
  /* --define=OUTPUTS=((forkHP1_QTree_Int_snk, 16, 65536, Word16__023), (dummy_write_QTree_Int_sink, 16, 65536, Pointer_QTree_Int), (forkHP1_MaskQTree_snk, 16, 65536, Word16__023), (dummy_write_MaskQTree_sink, 16, 65536, Pointer_MaskQTree), (es_6_1I__023, 32, 4294967296, Int)) */
  /* TYPE_START
CT__024wmAdd_Int 16 3 (0,[0]) (1,[16p,0,16p,16p,16p,16p,16p,16p]) (2,[16p,16p,0,16p,16p,16p,16p]) (3,[16p,16p,16p,0,16p,16p]) (4,[16p,16p,16p,16p])
QTree_Int 16 2 (0,[0]) (1,[32]) (2,[16p,16p,16p,16p]) (3,[0])
CT__024wnnz_Int 16 3 (0,[0]) (1,[16p,16p,16p,16p]) (2,[32,16p,16p,16p]) (3,[32,32,16p,16p]) (4,[32,32,32,16p])
CTmain_mask_Int 16 3 (0,[0]) (1,[16p,16p,16p,16p,16p,16p,16p]) (2,[16p,16p,16p,16p,16p,16p]) (3,[16p,16p,16p,16p,16p]) (4,[16p,16p,16p,16p])
MaskQTree 16 2 (0,[0]) (1,[0]) (2,[16p,16p,16p,16p])
TupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int 16 0 (0,[0,0,16p,16p])
TupGo___Pointer_QTree_Int 16 0 (0,[0,16p])
TupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT__024wmAdd_Int 16 0 (0,[0,0,16p,16p,16p])
TupGo___Pointer_QTree_Int___Pointer_CT__024wnnz_Int 16 0 (0,[0,16p,16p])
TupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Int 16 0 (0,[0,16p,16p,16p])
TupGo___Pointer_QTree_Int___Pointer_MaskQTree 16 0 (0,[0,16p,16p])
TYPE_END */
  /*  */
  /*  */
  Go_t go_1_d;
  logic go_1_r;
  Go_t go_2_d;
  logic go_2_r;
  Go_t go_3_d;
  logic go_3_r;
  Go_t go_4_d;
  logic go_4_r;
  Go_t go__5_d;
  logic go__5_r;
  Go_t go__6_d;
  logic go__6_r;
  Go_t go__7_d;
  logic go__7_r;
  Go_t go__8_d;
  logic go__8_r;
  Go_t go__9_d;
  logic go__9_r;
  Go_t go__10_d;
  logic go__10_r;
  \Word16#_t  initHP_CT$wmAdd_Int_d;
  logic initHP_CT$wmAdd_Int_r;
  \Word16#_t  incrHP_CT$wmAdd_Int_d;
  logic incrHP_CT$wmAdd_Int_r;
  Go_t incrHP_mergeCT$wmAdd_Int_d;
  logic incrHP_mergeCT$wmAdd_Int_r;
  Go_t incrHP_CT$wmAdd_Int1_d;
  logic incrHP_CT$wmAdd_Int1_r;
  Go_t incrHP_CT$wmAdd_Int2_d;
  logic incrHP_CT$wmAdd_Int2_r;
  \Word16#_t  addHP_CT$wmAdd_Int_d;
  logic addHP_CT$wmAdd_Int_r;
  \Word16#_t  mergeHP_CT$wmAdd_Int_d;
  logic mergeHP_CT$wmAdd_Int_r;
  Go_t incrHP_mergeCT$wmAdd_Int_buf_d;
  logic incrHP_mergeCT$wmAdd_Int_buf_r;
  \Word16#_t  mergeHP_CT$wmAdd_Int_buf_d;
  logic mergeHP_CT$wmAdd_Int_buf_r;
  \Word16#_t  forkHP1_CT$wmAdd_Int_d;
  logic forkHP1_CT$wmAdd_Int_r;
  \Word16#_t  forkHP1_CT$wmAdd_In2_d;
  logic forkHP1_CT$wmAdd_In2_r;
  \Word16#_t  forkHP1_CT$wmAdd_In3_d;
  logic forkHP1_CT$wmAdd_In3_r;
  C2_t memMergeChoice_CT$wmAdd_Int_d;
  logic memMergeChoice_CT$wmAdd_Int_r;
  MemIn_CT$wmAdd_Int_t memMergeIn_CT$wmAdd_Int_d;
  logic memMergeIn_CT$wmAdd_Int_r;
  MemOut_CT$wmAdd_Int_t memOut_CT$wmAdd_Int_d;
  logic memOut_CT$wmAdd_Int_r;
  MemOut_CT$wmAdd_Int_t memReadOut_CT$wmAdd_Int_d;
  logic memReadOut_CT$wmAdd_Int_r;
  MemOut_CT$wmAdd_Int_t memWriteOut_CT$wmAdd_Int_d;
  logic memWriteOut_CT$wmAdd_Int_r;
  MemIn_CT$wmAdd_Int_t memMergeIn_CT$wmAdd_Int_dbuf_d;
  logic memMergeIn_CT$wmAdd_Int_dbuf_r;
  MemIn_CT$wmAdd_Int_t memMergeIn_CT$wmAdd_Int_rbuf_d;
  logic memMergeIn_CT$wmAdd_Int_rbuf_r;
  MemOut_CT$wmAdd_Int_t memOut_CT$wmAdd_Int_dbuf_d;
  logic memOut_CT$wmAdd_Int_dbuf_r;
  MemOut_CT$wmAdd_Int_t memOut_CT$wmAdd_Int_rbuf_d;
  logic memOut_CT$wmAdd_Int_rbuf_r;
  \Word16#_t  destructReadIn_CT$wmAdd_Int_d;
  logic destructReadIn_CT$wmAdd_Int_r;
  MemIn_CT$wmAdd_Int_t dconReadIn_CT$wmAdd_Int_d;
  logic dconReadIn_CT$wmAdd_Int_r;
  CT$wmAdd_Int_t readPointer_CT$wmAdd_Intscfarg_0_1_argbuf_d;
  logic readPointer_CT$wmAdd_Intscfarg_0_1_argbuf_r;
  C5_t writeMerge_choice_CT$wmAdd_Int_d;
  logic writeMerge_choice_CT$wmAdd_Int_r;
  CT$wmAdd_Int_t writeMerge_data_CT$wmAdd_Int_d;
  logic writeMerge_data_CT$wmAdd_Int_r;
  Pointer_CT$wmAdd_Int_t writeCT$wmAdd_IntlizzieLet0_1_argbuf_d;
  logic writeCT$wmAdd_IntlizzieLet0_1_argbuf_r;
  Pointer_CT$wmAdd_Int_t writeCT$wmAdd_IntlizzieLet23_1_argbuf_d;
  logic writeCT$wmAdd_IntlizzieLet23_1_argbuf_r;
  Pointer_CT$wmAdd_Int_t writeCT$wmAdd_IntlizzieLet24_1_argbuf_d;
  logic writeCT$wmAdd_IntlizzieLet24_1_argbuf_r;
  Pointer_CT$wmAdd_Int_t writeCT$wmAdd_IntlizzieLet25_1_argbuf_d;
  logic writeCT$wmAdd_IntlizzieLet25_1_argbuf_r;
  Pointer_CT$wmAdd_Int_t writeCT$wmAdd_IntlizzieLet9_1_1_argbuf_d;
  logic writeCT$wmAdd_IntlizzieLet9_1_1_argbuf_r;
  MemIn_CT$wmAdd_Int_t dconWriteIn_CT$wmAdd_Int_d;
  logic dconWriteIn_CT$wmAdd_Int_r;
  Pointer_CT$wmAdd_Int_t dconPtr_CT$wmAdd_Int_d;
  logic dconPtr_CT$wmAdd_Int_r;
  Pointer_CT$wmAdd_Int_t _78_d;
  logic _78_r;
  assign _78_r = 1'd1;
  Pointer_CT$wmAdd_Int_t demuxWriteResult_CT$wmAdd_Int_d;
  logic demuxWriteResult_CT$wmAdd_Int_r;
  \Word16#_t  initHP_QTree_Int_d;
  logic initHP_QTree_Int_r;
  \Word16#_t  incrHP_QTree_Int_d;
  logic incrHP_QTree_Int_r;
  Go_t incrHP_mergeQTree_Int_d;
  logic incrHP_mergeQTree_Int_r;
  Go_t incrHP_QTree_Int1_d;
  logic incrHP_QTree_Int1_r;
  Go_t incrHP_QTree_Int2_d;
  logic incrHP_QTree_Int2_r;
  \Word16#_t  addHP_QTree_Int_d;
  logic addHP_QTree_Int_r;
  \Word16#_t  mergeHP_QTree_Int_d;
  logic mergeHP_QTree_Int_r;
  Go_t incrHP_mergeQTree_Int_buf_d;
  logic incrHP_mergeQTree_Int_buf_r;
  \Word16#_t  mergeHP_QTree_Int_buf_d;
  logic mergeHP_QTree_Int_buf_r;
  Go_t go_1_dummy_write_QTree_Int_d;
  logic go_1_dummy_write_QTree_Int_r;
  Go_t go_2_dummy_write_QTree_Int_d;
  logic go_2_dummy_write_QTree_Int_r;
  \Word16#_t  forkHP1_QTree_Int_d;
  logic forkHP1_QTree_Int_r;
  \Word16#_t  forkHP1_QTree_Int_snk_d;
  logic forkHP1_QTree_Int_snk_r;
  \Word16#_t  forkHP1_QTree_In3_d;
  logic forkHP1_QTree_In3_r;
  \Word16#_t  forkHP1_QTree_In4_d;
  logic forkHP1_QTree_In4_r;
  C2_t memMergeChoice_QTree_Int_d;
  logic memMergeChoice_QTree_Int_r;
  MemIn_QTree_Int_t memMergeIn_QTree_Int_d;
  logic memMergeIn_QTree_Int_r;
  MemOut_QTree_Int_t memOut_QTree_Int_d;
  logic memOut_QTree_Int_r;
  MemOut_QTree_Int_t memReadOut_QTree_Int_d;
  logic memReadOut_QTree_Int_r;
  MemOut_QTree_Int_t memWriteOut_QTree_Int_d;
  logic memWriteOut_QTree_Int_r;
  MemIn_QTree_Int_t memMergeIn_QTree_Int_dbuf_d;
  logic memMergeIn_QTree_Int_dbuf_r;
  MemIn_QTree_Int_t memMergeIn_QTree_Int_rbuf_d;
  logic memMergeIn_QTree_Int_rbuf_r;
  MemOut_QTree_Int_t memOut_QTree_Int_dbuf_d;
  logic memOut_QTree_Int_dbuf_r;
  MemOut_QTree_Int_t memOut_QTree_Int_rbuf_d;
  logic memOut_QTree_Int_rbuf_r;
  C4_t readMerge_choice_QTree_Int_d;
  logic readMerge_choice_QTree_Int_r;
  Pointer_QTree_Int_t readMerge_data_QTree_Int_d;
  logic readMerge_data_QTree_Int_r;
  QTree_Int_t readPointer_QTree_Intma8q_1_argbuf_d;
  logic readPointer_QTree_Intma8q_1_argbuf_r;
  QTree_Int_t readPointer_QTree_Intw1sif_1_1_argbuf_d;
  logic readPointer_QTree_Intw1sif_1_1_argbuf_r;
  QTree_Int_t readPointer_QTree_Intw2sig_1_1_argbuf_d;
  logic readPointer_QTree_Intw2sig_1_1_argbuf_r;
  QTree_Int_t readPointer_QTree_Intwsij_1_1_argbuf_d;
  logic readPointer_QTree_Intwsij_1_1_argbuf_r;
  \Word16#_t  destructReadIn_QTree_Int_d;
  logic destructReadIn_QTree_Int_r;
  MemIn_QTree_Int_t dconReadIn_QTree_Int_d;
  logic dconReadIn_QTree_Int_r;
  QTree_Int_t destructReadOut_QTree_Int_d;
  logic destructReadOut_QTree_Int_r;
  C13_t writeMerge_choice_QTree_Int_d;
  logic writeMerge_choice_QTree_Int_r;
  QTree_Int_t writeMerge_data_QTree_Int_d;
  logic writeMerge_data_QTree_Int_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet10_1_1_argbuf_d;
  logic writeQTree_IntlizzieLet10_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet11_1_1_argbuf_d;
  logic writeQTree_IntlizzieLet11_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet15_1_argbuf_d;
  logic writeQTree_IntlizzieLet15_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet17_1_argbuf_d;
  logic writeQTree_IntlizzieLet17_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet18_1_argbuf_d;
  logic writeQTree_IntlizzieLet18_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet20_1_argbuf_d;
  logic writeQTree_IntlizzieLet20_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet26_1_argbuf_d;
  logic writeQTree_IntlizzieLet26_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet35_1_argbuf_d;
  logic writeQTree_IntlizzieLet35_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet4_1_argbuf_d;
  logic writeQTree_IntlizzieLet4_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet5_1_argbuf_d;
  logic writeQTree_IntlizzieLet5_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet6_1_argbuf_d;
  logic writeQTree_IntlizzieLet6_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet8_1_1_argbuf_d;
  logic writeQTree_IntlizzieLet8_1_1_argbuf_r;
  Pointer_QTree_Int_t dummy_write_QTree_Int_sink_d;
  logic dummy_write_QTree_Int_sink_r;
  MemIn_QTree_Int_t dconWriteIn_QTree_Int_d;
  logic dconWriteIn_QTree_Int_r;
  Pointer_QTree_Int_t dconPtr_QTree_Int_d;
  logic dconPtr_QTree_Int_r;
  Pointer_QTree_Int_t _77_d;
  logic _77_r;
  assign _77_r = 1'd1;
  Pointer_QTree_Int_t demuxWriteResult_QTree_Int_d;
  logic demuxWriteResult_QTree_Int_r;
  \Word16#_t  initHP_CT$wnnz_Int_d;
  logic initHP_CT$wnnz_Int_r;
  \Word16#_t  incrHP_CT$wnnz_Int_d;
  logic incrHP_CT$wnnz_Int_r;
  Go_t incrHP_mergeCT$wnnz_Int_d;
  logic incrHP_mergeCT$wnnz_Int_r;
  Go_t incrHP_CT$wnnz_Int1_d;
  logic incrHP_CT$wnnz_Int1_r;
  Go_t incrHP_CT$wnnz_Int2_d;
  logic incrHP_CT$wnnz_Int2_r;
  \Word16#_t  addHP_CT$wnnz_Int_d;
  logic addHP_CT$wnnz_Int_r;
  \Word16#_t  mergeHP_CT$wnnz_Int_d;
  logic mergeHP_CT$wnnz_Int_r;
  Go_t incrHP_mergeCT$wnnz_Int_buf_d;
  logic incrHP_mergeCT$wnnz_Int_buf_r;
  \Word16#_t  mergeHP_CT$wnnz_Int_buf_d;
  logic mergeHP_CT$wnnz_Int_buf_r;
  \Word16#_t  forkHP1_CT$wnnz_Int_d;
  logic forkHP1_CT$wnnz_Int_r;
  \Word16#_t  forkHP1_CT$wnnz_In2_d;
  logic forkHP1_CT$wnnz_In2_r;
  \Word16#_t  forkHP1_CT$wnnz_In3_d;
  logic forkHP1_CT$wnnz_In3_r;
  C2_t memMergeChoice_CT$wnnz_Int_d;
  logic memMergeChoice_CT$wnnz_Int_r;
  MemIn_CT$wnnz_Int_t memMergeIn_CT$wnnz_Int_d;
  logic memMergeIn_CT$wnnz_Int_r;
  MemOut_CT$wnnz_Int_t memOut_CT$wnnz_Int_d;
  logic memOut_CT$wnnz_Int_r;
  MemOut_CT$wnnz_Int_t memReadOut_CT$wnnz_Int_d;
  logic memReadOut_CT$wnnz_Int_r;
  MemOut_CT$wnnz_Int_t memWriteOut_CT$wnnz_Int_d;
  logic memWriteOut_CT$wnnz_Int_r;
  MemIn_CT$wnnz_Int_t memMergeIn_CT$wnnz_Int_dbuf_d;
  logic memMergeIn_CT$wnnz_Int_dbuf_r;
  MemIn_CT$wnnz_Int_t memMergeIn_CT$wnnz_Int_rbuf_d;
  logic memMergeIn_CT$wnnz_Int_rbuf_r;
  MemOut_CT$wnnz_Int_t memOut_CT$wnnz_Int_dbuf_d;
  logic memOut_CT$wnnz_Int_dbuf_r;
  MemOut_CT$wnnz_Int_t memOut_CT$wnnz_Int_rbuf_d;
  logic memOut_CT$wnnz_Int_rbuf_r;
  \Word16#_t  destructReadIn_CT$wnnz_Int_d;
  logic destructReadIn_CT$wnnz_Int_r;
  MemIn_CT$wnnz_Int_t dconReadIn_CT$wnnz_Int_d;
  logic dconReadIn_CT$wnnz_Int_r;
  CT$wnnz_Int_t readPointer_CT$wnnz_Intscfarg_0_1_1_argbuf_d;
  logic readPointer_CT$wnnz_Intscfarg_0_1_1_argbuf_r;
  C5_t writeMerge_choice_CT$wnnz_Int_d;
  logic writeMerge_choice_CT$wnnz_Int_r;
  CT$wnnz_Int_t writeMerge_data_CT$wnnz_Int_d;
  logic writeMerge_data_CT$wnnz_Int_r;
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet13_1_1_argbuf_d;
  logic writeCT$wnnz_IntlizzieLet13_1_1_argbuf_r;
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet1_1_argbuf_d;
  logic writeCT$wnnz_IntlizzieLet1_1_argbuf_r;
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet28_1_argbuf_d;
  logic writeCT$wnnz_IntlizzieLet28_1_argbuf_r;
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet29_1_argbuf_d;
  logic writeCT$wnnz_IntlizzieLet29_1_argbuf_r;
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet30_1_argbuf_d;
  logic writeCT$wnnz_IntlizzieLet30_1_argbuf_r;
  MemIn_CT$wnnz_Int_t dconWriteIn_CT$wnnz_Int_d;
  logic dconWriteIn_CT$wnnz_Int_r;
  Pointer_CT$wnnz_Int_t dconPtr_CT$wnnz_Int_d;
  logic dconPtr_CT$wnnz_Int_r;
  Pointer_CT$wnnz_Int_t _76_d;
  logic _76_r;
  assign _76_r = 1'd1;
  Pointer_CT$wnnz_Int_t demuxWriteResult_CT$wnnz_Int_d;
  logic demuxWriteResult_CT$wnnz_Int_r;
  \Word16#_t  initHP_CTmain_mask_Int_d;
  logic initHP_CTmain_mask_Int_r;
  \Word16#_t  incrHP_CTmain_mask_Int_d;
  logic incrHP_CTmain_mask_Int_r;
  Go_t incrHP_mergeCTmain_mask_Int_d;
  logic incrHP_mergeCTmain_mask_Int_r;
  Go_t incrHP_CTmain_mask_Int1_d;
  logic incrHP_CTmain_mask_Int1_r;
  Go_t incrHP_CTmain_mask_Int2_d;
  logic incrHP_CTmain_mask_Int2_r;
  \Word16#_t  addHP_CTmain_mask_Int_d;
  logic addHP_CTmain_mask_Int_r;
  \Word16#_t  mergeHP_CTmain_mask_Int_d;
  logic mergeHP_CTmain_mask_Int_r;
  Go_t incrHP_mergeCTmain_mask_Int_buf_d;
  logic incrHP_mergeCTmain_mask_Int_buf_r;
  \Word16#_t  mergeHP_CTmain_mask_Int_buf_d;
  logic mergeHP_CTmain_mask_Int_buf_r;
  \Word16#_t  forkHP1_CTmain_mask_Int_d;
  logic forkHP1_CTmain_mask_Int_r;
  \Word16#_t  forkHP1_CTmain_mask_In2_d;
  logic forkHP1_CTmain_mask_In2_r;
  \Word16#_t  forkHP1_CTmain_mask_In3_d;
  logic forkHP1_CTmain_mask_In3_r;
  C2_t memMergeChoice_CTmain_mask_Int_d;
  logic memMergeChoice_CTmain_mask_Int_r;
  MemIn_CTmain_mask_Int_t memMergeIn_CTmain_mask_Int_d;
  logic memMergeIn_CTmain_mask_Int_r;
  MemOut_CTmain_mask_Int_t memOut_CTmain_mask_Int_d;
  logic memOut_CTmain_mask_Int_r;
  MemOut_CTmain_mask_Int_t memReadOut_CTmain_mask_Int_d;
  logic memReadOut_CTmain_mask_Int_r;
  MemOut_CTmain_mask_Int_t memWriteOut_CTmain_mask_Int_d;
  logic memWriteOut_CTmain_mask_Int_r;
  MemIn_CTmain_mask_Int_t memMergeIn_CTmain_mask_Int_dbuf_d;
  logic memMergeIn_CTmain_mask_Int_dbuf_r;
  MemIn_CTmain_mask_Int_t memMergeIn_CTmain_mask_Int_rbuf_d;
  logic memMergeIn_CTmain_mask_Int_rbuf_r;
  MemOut_CTmain_mask_Int_t memOut_CTmain_mask_Int_dbuf_d;
  logic memOut_CTmain_mask_Int_dbuf_r;
  MemOut_CTmain_mask_Int_t memOut_CTmain_mask_Int_rbuf_d;
  logic memOut_CTmain_mask_Int_rbuf_r;
  \Word16#_t  destructReadIn_CTmain_mask_Int_d;
  logic destructReadIn_CTmain_mask_Int_r;
  MemIn_CTmain_mask_Int_t dconReadIn_CTmain_mask_Int_d;
  logic dconReadIn_CTmain_mask_Int_r;
  CTmain_mask_Int_t readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf_d;
  logic readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf_r;
  C5_t writeMerge_choice_CTmain_mask_Int_d;
  logic writeMerge_choice_CTmain_mask_Int_r;
  CTmain_mask_Int_t writeMerge_data_CTmain_mask_Int_d;
  logic writeMerge_data_CTmain_mask_Int_r;
  Pointer_CTmain_mask_Int_t writeCTmain_mask_IntlizzieLet19_1_argbuf_d;
  logic writeCTmain_mask_IntlizzieLet19_1_argbuf_r;
  Pointer_CTmain_mask_Int_t writeCTmain_mask_IntlizzieLet21_1_argbuf_d;
  logic writeCTmain_mask_IntlizzieLet21_1_argbuf_r;
  Pointer_CTmain_mask_Int_t writeCTmain_mask_IntlizzieLet32_1_argbuf_d;
  logic writeCTmain_mask_IntlizzieLet32_1_argbuf_r;
  Pointer_CTmain_mask_Int_t writeCTmain_mask_IntlizzieLet33_1_argbuf_d;
  logic writeCTmain_mask_IntlizzieLet33_1_argbuf_r;
  Pointer_CTmain_mask_Int_t writeCTmain_mask_IntlizzieLet34_1_argbuf_d;
  logic writeCTmain_mask_IntlizzieLet34_1_argbuf_r;
  MemIn_CTmain_mask_Int_t dconWriteIn_CTmain_mask_Int_d;
  logic dconWriteIn_CTmain_mask_Int_r;
  Pointer_CTmain_mask_Int_t dconPtr_CTmain_mask_Int_d;
  logic dconPtr_CTmain_mask_Int_r;
  Pointer_CTmain_mask_Int_t _75_d;
  logic _75_r;
  assign _75_r = 1'd1;
  Pointer_CTmain_mask_Int_t demuxWriteResult_CTmain_mask_Int_d;
  logic demuxWriteResult_CTmain_mask_Int_r;
  \Word16#_t  initHP_MaskQTree_d;
  logic initHP_MaskQTree_r;
  \Word16#_t  incrHP_MaskQTree_d;
  logic incrHP_MaskQTree_r;
  Go_t incrHP_mergeMaskQTree_d;
  logic incrHP_mergeMaskQTree_r;
  Go_t incrHP_MaskQTree1_d;
  logic incrHP_MaskQTree1_r;
  Go_t incrHP_MaskQTree2_d;
  logic incrHP_MaskQTree2_r;
  \Word16#_t  addHP_MaskQTree_d;
  logic addHP_MaskQTree_r;
  \Word16#_t  mergeHP_MaskQTree_d;
  logic mergeHP_MaskQTree_r;
  Go_t incrHP_mergeMaskQTree_buf_d;
  logic incrHP_mergeMaskQTree_buf_r;
  \Word16#_t  mergeHP_MaskQTree_buf_d;
  logic mergeHP_MaskQTree_buf_r;
  Go_t go_1_dummy_write_MaskQTree_d;
  logic go_1_dummy_write_MaskQTree_r;
  Go_t go_2_dummy_write_MaskQTree_d;
  logic go_2_dummy_write_MaskQTree_r;
  \Word16#_t  forkHP1_MaskQTree_d;
  logic forkHP1_MaskQTree_r;
  \Word16#_t  forkHP1_MaskQTree_snk_d;
  logic forkHP1_MaskQTree_snk_r;
  \Word16#_t  forkHP1_MaskQTre3_d;
  logic forkHP1_MaskQTre3_r;
  \Word16#_t  forkHP1_MaskQTre4_d;
  logic forkHP1_MaskQTre4_r;
  C2_t memMergeChoice_MaskQTree_d;
  logic memMergeChoice_MaskQTree_r;
  MemIn_MaskQTree_t memMergeIn_MaskQTree_d;
  logic memMergeIn_MaskQTree_r;
  MemOut_MaskQTree_t memOut_MaskQTree_d;
  logic memOut_MaskQTree_r;
  MemOut_MaskQTree_t memReadOut_MaskQTree_d;
  logic memReadOut_MaskQTree_r;
  MemOut_MaskQTree_t memWriteOut_MaskQTree_d;
  logic memWriteOut_MaskQTree_r;
  MemIn_MaskQTree_t memMergeIn_MaskQTree_dbuf_d;
  logic memMergeIn_MaskQTree_dbuf_r;
  MemIn_MaskQTree_t memMergeIn_MaskQTree_rbuf_d;
  logic memMergeIn_MaskQTree_rbuf_r;
  MemOut_MaskQTree_t memOut_MaskQTree_dbuf_d;
  logic memOut_MaskQTree_dbuf_r;
  MemOut_MaskQTree_t memOut_MaskQTree_rbuf_d;
  logic memOut_MaskQTree_rbuf_r;
  \Word16#_t  destructReadIn_MaskQTree_d;
  logic destructReadIn_MaskQTree_r;
  MemIn_MaskQTree_t dconReadIn_MaskQTree_d;
  logic dconReadIn_MaskQTree_r;
  MaskQTree_t readPointer_MaskQTreemska8r_1_argbuf_d;
  logic readPointer_MaskQTreemska8r_1_argbuf_r;
  MemIn_MaskQTree_t dconWriteIn_MaskQTree_d;
  logic dconWriteIn_MaskQTree_r;
  Pointer_MaskQTree_t dconPtr_MaskQTree_d;
  logic dconPtr_MaskQTree_r;
  Pointer_MaskQTree_t _74_d;
  logic _74_r;
  assign _74_r = 1'd1;
  Pointer_MaskQTree_t dummy_write_MaskQTree_sink_d;
  logic dummy_write_MaskQTree_sink_r;
  Go_t \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgo_4_d ;
  logic \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgo_4_r ;
  MyDTInt_Int_Int_t \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intwsie_d ;
  logic \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intwsie_r ;
  Pointer_QTree_Int_t \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw1sif_d ;
  logic \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw1sif_r ;
  Pointer_QTree_Int_t \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw2sig_d ;
  logic \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw2sig_r ;
  Go_t go_4_1_d;
  logic go_4_1_r;
  Go_t go_4_2_d;
  logic go_4_2_r;
  Pointer_QTree_Int_t w1sif_1_argbuf_d;
  logic w1sif_1_argbuf_r;
  Pointer_QTree_Int_t w2sig_1_argbuf_d;
  logic w2sig_1_argbuf_r;
  MyDTInt_Int_Int_t wsie_1_argbuf_d;
  logic wsie_1_argbuf_r;
  Pointer_QTree_Int_t es_1_1_argbuf_d;
  logic es_1_1_argbuf_r;
  Go_t \$wnnz_IntTupGo___Pointer_QTree_Intgo_5_d ;
  logic \$wnnz_IntTupGo___Pointer_QTree_Intgo_5_r ;
  Pointer_QTree_Int_t \$wnnz_IntTupGo___Pointer_QTree_Intwsij_d ;
  logic \$wnnz_IntTupGo___Pointer_QTree_Intwsij_r ;
  Go_t go_5_1_d;
  logic go_5_1_r;
  Go_t go_5_2_d;
  logic go_5_2_r;
  Pointer_QTree_Int_t wsij_1_argbuf_d;
  logic wsij_1_argbuf_r;
  Int_t \es_6_1I#_d ;
  logic \es_6_1I#_r ;
  MyDTInt_Int_Int_t applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_d;
  logic applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_r;
  Int_t applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg2_d;
  logic applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg2_r;
  Int_t applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg1_d;
  logic applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg1_r;
  MyDTInt_Int_Int_t arg0_1_d;
  logic arg0_1_r;
  MyDTInt_Int_Int_t arg0_2_d;
  logic arg0_2_r;
  MyDTInt_Int_Int_t arg0_3_d;
  logic arg0_3_r;
  QTree_Int_t es_0_2_1QVal_Int_d;
  logic es_0_2_1QVal_Int_r;
  Int_t \arg0_1Dcon_$fNumInt_$c+_d ;
  logic \arg0_1Dcon_$fNumInt_$c+_r ;
  Int_t \arg0_2Dcon_$fNumInt_$c+_d ;
  logic \arg0_2Dcon_$fNumInt_$c+_r ;
  Int_t \arg0_2Dcon_$fNumInt_$c+_1_d ;
  logic \arg0_2Dcon_$fNumInt_$c+_1_r ;
  Int_t \arg0_2Dcon_$fNumInt_$c+_2_d ;
  logic \arg0_2Dcon_$fNumInt_$c+_2_r ;
  Int_t \arg0_2Dcon_$fNumInt_$c+_3_d ;
  logic \arg0_2Dcon_$fNumInt_$c+_3_r ;
  Int_t \arg0_2Dcon_$fNumInt_$c+_4_d ;
  logic \arg0_2Dcon_$fNumInt_$c+_4_r ;
  \Int#_t  xa1lV_destruct_d;
  logic xa1lV_destruct_r;
  Int_t \arg0_2Dcon_$fNumInt_$c+_1I#_d ;
  logic \arg0_2Dcon_$fNumInt_$c+_1I#_r ;
  Int_t \arg0_2Dcon_$fNumInt_$c+_3I#_d ;
  logic \arg0_2Dcon_$fNumInt_$c+_3I#_r ;
  Int_t \arg0_2Dcon_$fNumInt_$c+_3I#_1_d ;
  logic \arg0_2Dcon_$fNumInt_$c+_3I#_1_r ;
  Int_t \arg0_2Dcon_$fNumInt_$c+_3I#_2_d ;
  logic \arg0_2Dcon_$fNumInt_$c+_3I#_2_r ;
  Int_t \arg0_2Dcon_$fNumInt_$c+_3I#_3_d ;
  logic \arg0_2Dcon_$fNumInt_$c+_3I#_3_r ;
  Int_t \arg0_2Dcon_$fNumInt_$c+_3I#_4_d ;
  logic \arg0_2Dcon_$fNumInt_$c+_3I#_4_r ;
  \Int#_t  ya1lW_destruct_d;
  logic ya1lW_destruct_r;
  Int_t \arg0_2Dcon_$fNumInt_$c+_3I#_1I#_d ;
  logic \arg0_2Dcon_$fNumInt_$c+_3I#_1I#_r ;
  \Int#_t  \arg0_2Dcon_$fNumInt_$c+_3I#_3I#_d ;
  logic \arg0_2Dcon_$fNumInt_$c+_3I#_3I#_r ;
  \Int#_t  \arg0_2Dcon_$fNumInt_$c+_3I#_3I#_1ya1lW_1_Add32_d ;
  logic \arg0_2Dcon_$fNumInt_$c+_3I#_3I#_1ya1lW_1_Add32_r ;
  Int_t \es_0_1_1I#_d ;
  logic \es_0_1_1I#_r ;
  Int_t \es_0_1_1I#_mux_d ;
  logic \es_0_1_1I#_mux_r ;
  Int_t \es_0_1_1I#_mux_mux_d ;
  logic \es_0_1_1I#_mux_mux_r ;
  Int_t \es_0_1_1I#_mux_mux_mux_d ;
  logic \es_0_1_1I#_mux_mux_mux_r ;
  Go_t call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Intgo_6_d;
  logic call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Intgo_6_r;
  MyDTInt_Int_Int_t call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Intwsie_1_d;
  logic call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Intwsie_1_r;
  Pointer_QTree_Int_t call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Intw1sif_1_d;
  logic call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Intw1sif_1_r;
  Pointer_QTree_Int_t call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Intw2sig_1_d;
  logic call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Intw2sig_1_r;
  Pointer_CT$wmAdd_Int_t call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Intsc_0_d;
  logic call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Intsc_0_r;
  Go_t call_$wmAdd_Int_initBufi_d;
  logic call_$wmAdd_Int_initBufi_r;
  C5_t go_6_goMux_choice_d;
  logic go_6_goMux_choice_r;
  Go_t go_6_goMux_data_d;
  logic go_6_goMux_data_r;
  Go_t call_$wmAdd_Int_unlockFork1_d;
  logic call_$wmAdd_Int_unlockFork1_r;
  Go_t call_$wmAdd_Int_unlockFork2_d;
  logic call_$wmAdd_Int_unlockFork2_r;
  Go_t call_$wmAdd_Int_unlockFork3_d;
  logic call_$wmAdd_Int_unlockFork3_r;
  Go_t call_$wmAdd_Int_unlockFork4_d;
  logic call_$wmAdd_Int_unlockFork4_r;
  Go_t call_$wmAdd_Int_unlockFork5_d;
  logic call_$wmAdd_Int_unlockFork5_r;
  Go_t call_$wmAdd_Int_initBuf_d;
  logic call_$wmAdd_Int_initBuf_r;
  Go_t call_$wmAdd_Int_goMux1_d;
  logic call_$wmAdd_Int_goMux1_r;
  MyDTInt_Int_Int_t call_$wmAdd_Int_goMux2_d;
  logic call_$wmAdd_Int_goMux2_r;
  Pointer_QTree_Int_t call_$wmAdd_Int_goMux3_d;
  logic call_$wmAdd_Int_goMux3_r;
  Pointer_QTree_Int_t call_$wmAdd_Int_goMux4_d;
  logic call_$wmAdd_Int_goMux4_r;
  Pointer_CT$wmAdd_Int_t call_$wmAdd_Int_goMux5_d;
  logic call_$wmAdd_Int_goMux5_r;
  Go_t call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intgo_7_d;
  logic call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intgo_7_r;
  Pointer_QTree_Int_t call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intwsij_1_d;
  logic call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intwsij_1_r;
  Pointer_CT$wnnz_Int_t call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intsc_0_1_d;
  logic call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intsc_0_1_r;
  Go_t call_$wnnz_Int_initBufi_d;
  logic call_$wnnz_Int_initBufi_r;
  C5_t go_7_goMux_choice_d;
  logic go_7_goMux_choice_r;
  Go_t go_7_goMux_data_d;
  logic go_7_goMux_data_r;
  Go_t call_$wnnz_Int_unlockFork1_d;
  logic call_$wnnz_Int_unlockFork1_r;
  Go_t call_$wnnz_Int_unlockFork2_d;
  logic call_$wnnz_Int_unlockFork2_r;
  Go_t call_$wnnz_Int_unlockFork3_d;
  logic call_$wnnz_Int_unlockFork3_r;
  Go_t call_$wnnz_Int_initBuf_d;
  logic call_$wnnz_Int_initBuf_r;
  Go_t call_$wnnz_Int_goMux1_d;
  logic call_$wnnz_Int_goMux1_r;
  Pointer_QTree_Int_t call_$wnnz_Int_goMux2_d;
  logic call_$wnnz_Int_goMux2_r;
  Pointer_CT$wnnz_Int_t call_$wnnz_Int_goMux3_d;
  logic call_$wnnz_Int_goMux3_r;
  Go_t call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Intgo_8_d;
  logic call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Intgo_8_r;
  Pointer_QTree_Int_t call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Intma8q_d;
  logic call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Intma8q_r;
  Pointer_MaskQTree_t call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Intmska8r_d;
  logic call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Intmska8r_r;
  Pointer_CTmain_mask_Int_t call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Intsc_0_2_d;
  logic call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Intsc_0_2_r;
  Go_t call_main_mask_Int_initBufi_d;
  logic call_main_mask_Int_initBufi_r;
  C5_t go_8_goMux_choice_d;
  logic go_8_goMux_choice_r;
  Go_t go_8_goMux_data_d;
  logic go_8_goMux_data_r;
  Go_t call_main_mask_Int_unlockFork1_d;
  logic call_main_mask_Int_unlockFork1_r;
  Go_t call_main_mask_Int_unlockFork2_d;
  logic call_main_mask_Int_unlockFork2_r;
  Go_t call_main_mask_Int_unlockFork3_d;
  logic call_main_mask_Int_unlockFork3_r;
  Go_t call_main_mask_Int_unlockFork4_d;
  logic call_main_mask_Int_unlockFork4_r;
  Go_t call_main_mask_Int_initBuf_d;
  logic call_main_mask_Int_initBuf_r;
  Go_t call_main_mask_Int_goMux1_d;
  logic call_main_mask_Int_goMux1_r;
  Pointer_QTree_Int_t call_main_mask_Int_goMux2_d;
  logic call_main_mask_Int_goMux2_r;
  Pointer_MaskQTree_t call_main_mask_Int_goMux3_d;
  logic call_main_mask_Int_goMux3_r;
  Pointer_CTmain_mask_Int_t call_main_mask_Int_goMux4_d;
  logic call_main_mask_Int_goMux4_r;
  Int_t applyfnInt_Int_Int_5_resbuf_d;
  logic applyfnInt_Int_Int_5_resbuf_r;
  QTree_Int_t lizzieLet4_1_argbuf_d;
  logic lizzieLet4_1_argbuf_r;
  \Int#_t  contRet_0_1_1_argbuf_d;
  logic contRet_0_1_1_argbuf_r;
  \Int#_t  es_4_3_1lizzieLet27_4Lcall_$wnnz_Int0_1_Add32_d;
  logic es_4_3_1lizzieLet27_4Lcall_$wnnz_Int0_1_Add32_r;
  MyDTInt_Int_Int_t \go_1Dcon_$fNumInt_$c+_d ;
  logic \go_1Dcon_$fNumInt_$c+_r ;
  C10_t go_10_goMux_choice_1_d;
  logic go_10_goMux_choice_1_r;
  C10_t go_10_goMux_choice_2_d;
  logic go_10_goMux_choice_2_r;
  Pointer_QTree_Int_t srtarg_0_goMux_mux_d;
  logic srtarg_0_goMux_mux_r;
  Pointer_CT$wmAdd_Int_t scfarg_0_goMux_mux_d;
  logic scfarg_0_goMux_mux_r;
  C4_t go_11_goMux_choice_1_d;
  logic go_11_goMux_choice_1_r;
  C4_t go_11_goMux_choice_2_d;
  logic go_11_goMux_choice_2_r;
  \Int#_t  srtarg_0_1_goMux_mux_d;
  logic srtarg_0_1_goMux_mux_r;
  Pointer_CT$wnnz_Int_t scfarg_0_1_goMux_mux_d;
  logic scfarg_0_1_goMux_mux_r;
  C6_t go_12_goMux_choice_1_d;
  logic go_12_goMux_choice_1_r;
  C6_t go_12_goMux_choice_2_d;
  logic go_12_goMux_choice_2_r;
  Pointer_QTree_Int_t srtarg_0_2_goMux_mux_d;
  logic srtarg_0_2_goMux_mux_r;
  Pointer_CTmain_mask_Int_t scfarg_0_2_goMux_mux_d;
  logic scfarg_0_2_goMux_mux_r;
  MyDTInt_Int_Int_t es_3_1_argbuf_d;
  logic es_3_1_argbuf_r;
  Go_t go_2_argbuf_d;
  logic go_2_argbuf_r;
  TupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_t \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1_d ;
  logic \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1_r ;
  Go_t go_3_argbuf_d;
  logic go_3_argbuf_r;
  TupGo___Pointer_QTree_Int___Pointer_MaskQTree_t main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree_1_d;
  logic main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree_1_r;
  Go_t go_4_argbuf_d;
  logic go_4_argbuf_r;
  CT$wmAdd_Int_t go_4_1L$wmAdd_Intsbos_d;
  logic go_4_1L$wmAdd_Intsbos_r;
  CT$wmAdd_Int_t lizzieLet0_1_argbuf_d;
  logic lizzieLet0_1_argbuf_r;
  Go_t go_4_2_argbuf_d;
  logic go_4_2_argbuf_r;
  TupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Int_t call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Int_1_d;
  logic call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Int_1_r;
  TupGo___Pointer_QTree_Int_t \$wnnz_IntTupGo___Pointer_QTree_Int_1_d ;
  logic \$wnnz_IntTupGo___Pointer_QTree_Int_1_r ;
  CT$wnnz_Int_t go_5_1L$wnnz_Intsbos_d;
  logic go_5_1L$wnnz_Intsbos_r;
  CT$wnnz_Int_t lizzieLet1_1_argbuf_d;
  logic lizzieLet1_1_argbuf_r;
  Go_t go_5_2_argbuf_d;
  logic go_5_2_argbuf_r;
  TupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_t call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_d;
  logic call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_r;
  C5_t go_6_goMux_choice_1_d;
  logic go_6_goMux_choice_1_r;
  C5_t go_6_goMux_choice_2_d;
  logic go_6_goMux_choice_2_r;
  C5_t go_6_goMux_choice_3_d;
  logic go_6_goMux_choice_3_r;
  C5_t go_6_goMux_choice_4_d;
  logic go_6_goMux_choice_4_r;
  MyDTInt_Int_Int_t wsie_1_goMux_mux_d;
  logic wsie_1_goMux_mux_r;
  Pointer_QTree_Int_t w1sif_1_goMux_mux_d;
  logic w1sif_1_goMux_mux_r;
  Pointer_QTree_Int_t w2sig_1_goMux_mux_d;
  logic w2sig_1_goMux_mux_r;
  Pointer_CT$wmAdd_Int_t sc_0_goMux_mux_d;
  logic sc_0_goMux_mux_r;
  C5_t go_7_goMux_choice_1_d;
  logic go_7_goMux_choice_1_r;
  C5_t go_7_goMux_choice_2_d;
  logic go_7_goMux_choice_2_r;
  Pointer_QTree_Int_t wsij_1_goMux_mux_d;
  logic wsij_1_goMux_mux_r;
  Pointer_CT$wnnz_Int_t sc_0_1_goMux_mux_d;
  logic sc_0_1_goMux_mux_r;
  C5_t go_8_goMux_choice_1_d;
  logic go_8_goMux_choice_1_r;
  C5_t go_8_goMux_choice_2_d;
  logic go_8_goMux_choice_2_r;
  C5_t go_8_goMux_choice_3_d;
  logic go_8_goMux_choice_3_r;
  Pointer_QTree_Int_t ma8q_goMux_mux_d;
  logic ma8q_goMux_mux_r;
  Pointer_MaskQTree_t mska8r_goMux_mux_d;
  logic mska8r_goMux_mux_r;
  Pointer_CTmain_mask_Int_t sc_0_2_goMux_mux_d;
  logic sc_0_2_goMux_mux_r;
  CTmain_mask_Int_t go_9_1Lmain_mask_Intsbos_d;
  logic go_9_1Lmain_mask_Intsbos_r;
  CTmain_mask_Int_t lizzieLet21_1_argbuf_d;
  logic lizzieLet21_1_argbuf_r;
  Go_t go_9_2_argbuf_d;
  logic go_9_2_argbuf_r;
  TupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Int_t call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Int_1_d;
  logic call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Int_1_r;
  Pointer_QTree_Int_t q1a8C_destruct_d;
  logic q1a8C_destruct_r;
  Pointer_QTree_Int_t q2a8D_destruct_d;
  logic q2a8D_destruct_r;
  Pointer_QTree_Int_t q3a8E_destruct_d;
  logic q3a8E_destruct_r;
  Pointer_QTree_Int_t q4a8F_destruct_d;
  logic q4a8F_destruct_r;
  QTree_Int_t _73_d;
  logic _73_r;
  assign _73_r = 1'd1;
  QTree_Int_t _72_d;
  logic _72_r;
  assign _72_r = 1'd1;
  QTree_Int_t lizzieLet12_1_1QNode_Int_d;
  logic lizzieLet12_1_1QNode_Int_r;
  QTree_Int_t _71_d;
  logic _71_r;
  assign _71_r = 1'd1;
  Go_t lizzieLet12_1_3QNone_Int_d;
  logic lizzieLet12_1_3QNone_Int_r;
  Go_t lizzieLet12_1_3QVal_Int_d;
  logic lizzieLet12_1_3QVal_Int_r;
  Go_t lizzieLet12_1_3QNode_Int_d;
  logic lizzieLet12_1_3QNode_Int_r;
  Go_t lizzieLet12_1_3QError_Int_d;
  logic lizzieLet12_1_3QError_Int_r;
  Go_t lizzieLet12_1_3QError_Int_1_d;
  logic lizzieLet12_1_3QError_Int_1_r;
  Go_t lizzieLet12_1_3QError_Int_2_d;
  logic lizzieLet12_1_3QError_Int_2_r;
  Go_t lizzieLet12_1_3QError_Int_1_argbuf_d;
  logic lizzieLet12_1_3QError_Int_1_argbuf_r;
  \Int#_t  lizzieLet12_1_3QError_Int_1_argbuf_0_d;
  logic lizzieLet12_1_3QError_Int_1_argbuf_0_r;
  \Int#_t  lizzieLet5_2_1_argbuf_d;
  logic lizzieLet5_2_1_argbuf_r;
  Go_t lizzieLet12_1_3QError_Int_2_argbuf_d;
  logic lizzieLet12_1_3QError_Int_2_argbuf_r;
  Go_t lizzieLet12_1_3QNode_Int_1_argbuf_d;
  logic lizzieLet12_1_3QNode_Int_1_argbuf_r;
  Go_t lizzieLet12_1_3QNone_Int_1_d;
  logic lizzieLet12_1_3QNone_Int_1_r;
  Go_t lizzieLet12_1_3QNone_Int_2_d;
  logic lizzieLet12_1_3QNone_Int_2_r;
  Go_t lizzieLet12_1_3QNone_Int_1_argbuf_d;
  logic lizzieLet12_1_3QNone_Int_1_argbuf_r;
  \Int#_t  lizzieLet12_1_3QNone_Int_1_argbuf_0_d;
  logic lizzieLet12_1_3QNone_Int_1_argbuf_0_r;
  \Int#_t  lizzieLet5_1_1_argbuf_d;
  logic lizzieLet5_1_1_argbuf_r;
  Go_t lizzieLet12_1_3QNone_Int_2_argbuf_d;
  logic lizzieLet12_1_3QNone_Int_2_argbuf_r;
  C4_t go_11_goMux_choice_d;
  logic go_11_goMux_choice_r;
  Go_t go_11_goMux_data_d;
  logic go_11_goMux_data_r;
  Go_t lizzieLet12_1_3QVal_Int_1_d;
  logic lizzieLet12_1_3QVal_Int_1_r;
  Go_t lizzieLet12_1_3QVal_Int_2_d;
  logic lizzieLet12_1_3QVal_Int_2_r;
  Go_t lizzieLet12_1_3QVal_Int_1_argbuf_d;
  logic lizzieLet12_1_3QVal_Int_1_argbuf_r;
  \Int#_t  lizzieLet12_1_3QVal_Int_1_argbuf_1_d;
  logic lizzieLet12_1_3QVal_Int_1_argbuf_1_r;
  \Int#_t  lizzieLet6_1_1_argbuf_d;
  logic lizzieLet6_1_1_argbuf_r;
  Go_t lizzieLet12_1_3QVal_Int_2_argbuf_d;
  logic lizzieLet12_1_3QVal_Int_2_argbuf_r;
  Pointer_CT$wnnz_Int_t lizzieLet12_1_4QNone_Int_d;
  logic lizzieLet12_1_4QNone_Int_r;
  Pointer_CT$wnnz_Int_t lizzieLet12_1_4QVal_Int_d;
  logic lizzieLet12_1_4QVal_Int_r;
  Pointer_CT$wnnz_Int_t lizzieLet12_1_4QNode_Int_d;
  logic lizzieLet12_1_4QNode_Int_r;
  Pointer_CT$wnnz_Int_t lizzieLet12_1_4QError_Int_d;
  logic lizzieLet12_1_4QError_Int_r;
  Pointer_CT$wnnz_Int_t lizzieLet12_1_4QError_Int_1_argbuf_d;
  logic lizzieLet12_1_4QError_Int_1_argbuf_r;
  CT$wnnz_Int_t lizzieLet12_1_4QNode_Int_1q4a8F_1q3a8E_1q2a8D_1Lcall_$wnnz_Int3_d;
  logic lizzieLet12_1_4QNode_Int_1q4a8F_1q3a8E_1q2a8D_1Lcall_$wnnz_Int3_r;
  CT$wnnz_Int_t lizzieLet13_1_1_argbuf_d;
  logic lizzieLet13_1_1_argbuf_r;
  Pointer_CT$wnnz_Int_t lizzieLet12_1_4QNone_Int_1_argbuf_d;
  logic lizzieLet12_1_4QNone_Int_1_argbuf_r;
  Pointer_CT$wnnz_Int_t lizzieLet12_1_4QVal_Int_1_argbuf_d;
  logic lizzieLet12_1_4QVal_Int_1_argbuf_r;
  Pointer_MaskQTree_t q1a8s_destruct_d;
  logic q1a8s_destruct_r;
  Pointer_MaskQTree_t q2a8t_destruct_d;
  logic q2a8t_destruct_r;
  Pointer_MaskQTree_t q3a8u_destruct_d;
  logic q3a8u_destruct_r;
  Pointer_MaskQTree_t q4a8v_destruct_d;
  logic q4a8v_destruct_r;
  MaskQTree_t _70_d;
  logic _70_r;
  assign _70_r = 1'd1;
  MaskQTree_t _69_d;
  logic _69_r;
  assign _69_r = 1'd1;
  MaskQTree_t lizzieLet14_1_1MQNode_d;
  logic lizzieLet14_1_1MQNode_r;
  Go_t lizzieLet14_1_3MQNone_d;
  logic lizzieLet14_1_3MQNone_r;
  Go_t lizzieLet14_1_3MQVal_d;
  logic lizzieLet14_1_3MQVal_r;
  Go_t lizzieLet14_1_3MQNode_d;
  logic lizzieLet14_1_3MQNode_r;
  Go_t lizzieLet14_1_3MQNone_1_d;
  logic lizzieLet14_1_3MQNone_1_r;
  Go_t lizzieLet14_1_3MQNone_2_d;
  logic lizzieLet14_1_3MQNone_2_r;
  QTree_Int_t lizzieLet14_1_3MQNone_1QNone_Int_d;
  logic lizzieLet14_1_3MQNone_1QNone_Int_r;
  QTree_Int_t lizzieLet15_1_argbuf_d;
  logic lizzieLet15_1_argbuf_r;
  Go_t lizzieLet14_1_3MQNone_2_argbuf_d;
  logic lizzieLet14_1_3MQNone_2_argbuf_r;
  C6_t go_12_goMux_choice_d;
  logic go_12_goMux_choice_r;
  Go_t go_12_goMux_data_d;
  logic go_12_goMux_data_r;
  Go_t lizzieLet14_1_3MQVal_1_argbuf_d;
  logic lizzieLet14_1_3MQVal_1_argbuf_r;
  QTree_Int_t _68_d;
  logic _68_r;
  assign _68_r = 1'd1;
  QTree_Int_t _67_d;
  logic _67_r;
  assign _67_r = 1'd1;
  QTree_Int_t lizzieLet14_1_4MQNode_d;
  logic lizzieLet14_1_4MQNode_r;
  QTree_Int_t lizzieLet14_1_4MQNode_1_d;
  logic lizzieLet14_1_4MQNode_1_r;
  QTree_Int_t lizzieLet14_1_4MQNode_2_d;
  logic lizzieLet14_1_4MQNode_2_r;
  QTree_Int_t lizzieLet14_1_4MQNode_3_d;
  logic lizzieLet14_1_4MQNode_3_r;
  QTree_Int_t lizzieLet14_1_4MQNode_4_d;
  logic lizzieLet14_1_4MQNode_4_r;
  QTree_Int_t lizzieLet14_1_4MQNode_5_d;
  logic lizzieLet14_1_4MQNode_5_r;
  QTree_Int_t lizzieLet14_1_4MQNode_6_d;
  logic lizzieLet14_1_4MQNode_6_r;
  QTree_Int_t lizzieLet14_1_4MQNode_7_d;
  logic lizzieLet14_1_4MQNode_7_r;
  QTree_Int_t lizzieLet14_1_4MQNode_8_d;
  logic lizzieLet14_1_4MQNode_8_r;
  Pointer_QTree_Int_t t1a8x_destruct_d;
  logic t1a8x_destruct_r;
  Pointer_QTree_Int_t t2a8y_destruct_d;
  logic t2a8y_destruct_r;
  Pointer_QTree_Int_t t3a8z_destruct_d;
  logic t3a8z_destruct_r;
  Pointer_QTree_Int_t t4a8A_destruct_d;
  logic t4a8A_destruct_r;
  QTree_Int_t _66_d;
  logic _66_r;
  assign _66_r = 1'd1;
  QTree_Int_t _65_d;
  logic _65_r;
  assign _65_r = 1'd1;
  QTree_Int_t lizzieLet14_1_4MQNode_1QNode_Int_d;
  logic lizzieLet14_1_4MQNode_1QNode_Int_r;
  QTree_Int_t _64_d;
  logic _64_r;
  assign _64_r = 1'd1;
  Go_t lizzieLet14_1_4MQNode_3QNone_Int_d;
  logic lizzieLet14_1_4MQNode_3QNone_Int_r;
  Go_t lizzieLet14_1_4MQNode_3QVal_Int_d;
  logic lizzieLet14_1_4MQNode_3QVal_Int_r;
  Go_t lizzieLet14_1_4MQNode_3QNode_Int_d;
  logic lizzieLet14_1_4MQNode_3QNode_Int_r;
  Go_t lizzieLet14_1_4MQNode_3QError_Int_d;
  logic lizzieLet14_1_4MQNode_3QError_Int_r;
  Go_t lizzieLet14_1_4MQNode_3QError_Int_1_d;
  logic lizzieLet14_1_4MQNode_3QError_Int_1_r;
  Go_t lizzieLet14_1_4MQNode_3QError_Int_2_d;
  logic lizzieLet14_1_4MQNode_3QError_Int_2_r;
  QTree_Int_t lizzieLet14_1_4MQNode_3QError_Int_1QError_Int_d;
  logic lizzieLet14_1_4MQNode_3QError_Int_1QError_Int_r;
  QTree_Int_t lizzieLet20_1_argbuf_d;
  logic lizzieLet20_1_argbuf_r;
  Go_t lizzieLet14_1_4MQNode_3QError_Int_2_argbuf_d;
  logic lizzieLet14_1_4MQNode_3QError_Int_2_argbuf_r;
  Go_t lizzieLet14_1_4MQNode_3QNode_Int_1_argbuf_d;
  logic lizzieLet14_1_4MQNode_3QNode_Int_1_argbuf_r;
  Go_t lizzieLet14_1_4MQNode_3QNone_Int_1_d;
  logic lizzieLet14_1_4MQNode_3QNone_Int_1_r;
  Go_t lizzieLet14_1_4MQNode_3QNone_Int_2_d;
  logic lizzieLet14_1_4MQNode_3QNone_Int_2_r;
  QTree_Int_t lizzieLet14_1_4MQNode_3QNone_Int_1QNone_Int_d;
  logic lizzieLet14_1_4MQNode_3QNone_Int_1QNone_Int_r;
  QTree_Int_t lizzieLet17_1_argbuf_d;
  logic lizzieLet17_1_argbuf_r;
  Go_t lizzieLet14_1_4MQNode_3QNone_Int_2_argbuf_d;
  logic lizzieLet14_1_4MQNode_3QNone_Int_2_argbuf_r;
  Go_t lizzieLet14_1_4MQNode_3QVal_Int_1_d;
  logic lizzieLet14_1_4MQNode_3QVal_Int_1_r;
  Go_t lizzieLet14_1_4MQNode_3QVal_Int_2_d;
  logic lizzieLet14_1_4MQNode_3QVal_Int_2_r;
  QTree_Int_t lizzieLet14_1_4MQNode_3QVal_Int_1QError_Int_d;
  logic lizzieLet14_1_4MQNode_3QVal_Int_1QError_Int_r;
  QTree_Int_t lizzieLet18_1_argbuf_d;
  logic lizzieLet18_1_argbuf_r;
  Go_t lizzieLet14_1_4MQNode_3QVal_Int_2_argbuf_d;
  logic lizzieLet14_1_4MQNode_3QVal_Int_2_argbuf_r;
  Pointer_CTmain_mask_Int_t lizzieLet14_1_4MQNode_4QNone_Int_d;
  logic lizzieLet14_1_4MQNode_4QNone_Int_r;
  Pointer_CTmain_mask_Int_t lizzieLet14_1_4MQNode_4QVal_Int_d;
  logic lizzieLet14_1_4MQNode_4QVal_Int_r;
  Pointer_CTmain_mask_Int_t lizzieLet14_1_4MQNode_4QNode_Int_d;
  logic lizzieLet14_1_4MQNode_4QNode_Int_r;
  Pointer_CTmain_mask_Int_t lizzieLet14_1_4MQNode_4QError_Int_d;
  logic lizzieLet14_1_4MQNode_4QError_Int_r;
  Pointer_CTmain_mask_Int_t lizzieLet14_1_4MQNode_4QError_Int_1_argbuf_d;
  logic lizzieLet14_1_4MQNode_4QError_Int_1_argbuf_r;
  CTmain_mask_Int_t lizzieLet14_1_4MQNode_4QNode_Int_1t1a8x_1lizzieLet14_1_4MQNode_5QNode_Int_1t2a8y_1lizzieLet14_1_4MQNode_6QNode_Int_1t3a8z_1lizzieLet14_1_4MQNode_7QNode_Int_1Lcall_main_mask_Int3_d;
  logic lizzieLet14_1_4MQNode_4QNode_Int_1t1a8x_1lizzieLet14_1_4MQNode_5QNode_Int_1t2a8y_1lizzieLet14_1_4MQNode_6QNode_Int_1t3a8z_1lizzieLet14_1_4MQNode_7QNode_Int_1Lcall_main_mask_Int3_r;
  CTmain_mask_Int_t lizzieLet19_1_argbuf_d;
  logic lizzieLet19_1_argbuf_r;
  Pointer_CTmain_mask_Int_t lizzieLet14_1_4MQNode_4QNone_Int_1_argbuf_d;
  logic lizzieLet14_1_4MQNode_4QNone_Int_1_argbuf_r;
  Pointer_CTmain_mask_Int_t lizzieLet14_1_4MQNode_4QVal_Int_1_argbuf_d;
  logic lizzieLet14_1_4MQNode_4QVal_Int_1_argbuf_r;
  Pointer_MaskQTree_t _63_d;
  logic _63_r;
  assign _63_r = 1'd1;
  Pointer_MaskQTree_t _62_d;
  logic _62_r;
  assign _62_r = 1'd1;
  Pointer_MaskQTree_t lizzieLet14_1_4MQNode_5QNode_Int_d;
  logic lizzieLet14_1_4MQNode_5QNode_Int_r;
  Pointer_MaskQTree_t _61_d;
  logic _61_r;
  assign _61_r = 1'd1;
  Pointer_MaskQTree_t _60_d;
  logic _60_r;
  assign _60_r = 1'd1;
  Pointer_MaskQTree_t _59_d;
  logic _59_r;
  assign _59_r = 1'd1;
  Pointer_MaskQTree_t lizzieLet14_1_4MQNode_6QNode_Int_d;
  logic lizzieLet14_1_4MQNode_6QNode_Int_r;
  Pointer_MaskQTree_t _58_d;
  logic _58_r;
  assign _58_r = 1'd1;
  Pointer_MaskQTree_t _57_d;
  logic _57_r;
  assign _57_r = 1'd1;
  Pointer_MaskQTree_t _56_d;
  logic _56_r;
  assign _56_r = 1'd1;
  Pointer_MaskQTree_t lizzieLet14_1_4MQNode_7QNode_Int_d;
  logic lizzieLet14_1_4MQNode_7QNode_Int_r;
  Pointer_MaskQTree_t _55_d;
  logic _55_r;
  assign _55_r = 1'd1;
  Pointer_MaskQTree_t _54_d;
  logic _54_r;
  assign _54_r = 1'd1;
  Pointer_MaskQTree_t _53_d;
  logic _53_r;
  assign _53_r = 1'd1;
  Pointer_MaskQTree_t lizzieLet14_1_4MQNode_8QNode_Int_d;
  logic lizzieLet14_1_4MQNode_8QNode_Int_r;
  Pointer_MaskQTree_t _52_d;
  logic _52_r;
  assign _52_r = 1'd1;
  Pointer_MaskQTree_t lizzieLet14_1_4MQNode_8QNode_Int_1_argbuf_d;
  logic lizzieLet14_1_4MQNode_8QNode_Int_1_argbuf_r;
  Pointer_QTree_Int_t _51_d;
  logic _51_r;
  assign _51_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet14_1_5MQVal_d;
  logic lizzieLet14_1_5MQVal_r;
  Pointer_QTree_Int_t _50_d;
  logic _50_r;
  assign _50_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet14_1_5MQVal_1_argbuf_d;
  logic lizzieLet14_1_5MQVal_1_argbuf_r;
  Pointer_CTmain_mask_Int_t lizzieLet14_1_6MQNone_d;
  logic lizzieLet14_1_6MQNone_r;
  Pointer_CTmain_mask_Int_t lizzieLet14_1_6MQVal_d;
  logic lizzieLet14_1_6MQVal_r;
  Pointer_CTmain_mask_Int_t lizzieLet14_1_6MQNode_d;
  logic lizzieLet14_1_6MQNode_r;
  Pointer_CTmain_mask_Int_t lizzieLet14_1_6MQNone_1_argbuf_d;
  logic lizzieLet14_1_6MQNone_1_argbuf_r;
  Pointer_CTmain_mask_Int_t lizzieLet14_1_6MQVal_1_argbuf_d;
  logic lizzieLet14_1_6MQVal_1_argbuf_r;
  Pointer_QTree_Int_t es_2_destruct_d;
  logic es_2_destruct_r;
  Pointer_QTree_Int_t es_3_2_destruct_d;
  logic es_3_2_destruct_r;
  Pointer_QTree_Int_t es_4_2_destruct_d;
  logic es_4_2_destruct_r;
  Pointer_CT$wmAdd_Int_t sc_0_6_destruct_d;
  logic sc_0_6_destruct_r;
  Pointer_QTree_Int_t es_3_1_destruct_d;
  logic es_3_1_destruct_r;
  Pointer_QTree_Int_t es_4_1_destruct_d;
  logic es_4_1_destruct_r;
  Pointer_CT$wmAdd_Int_t sc_0_5_destruct_d;
  logic sc_0_5_destruct_r;
  MyDTInt_Int_Int_t wsie_4_destruct_d;
  logic wsie_4_destruct_r;
  Pointer_QTree_Int_t q1a8h_3_destruct_d;
  logic q1a8h_3_destruct_r;
  Pointer_QTree_Int_t t1a8m_3_destruct_d;
  logic t1a8m_3_destruct_r;
  Pointer_QTree_Int_t es_4_destruct_d;
  logic es_4_destruct_r;
  Pointer_CT$wmAdd_Int_t sc_0_4_destruct_d;
  logic sc_0_4_destruct_r;
  MyDTInt_Int_Int_t wsie_3_destruct_d;
  logic wsie_3_destruct_r;
  Pointer_QTree_Int_t q1a8h_2_destruct_d;
  logic q1a8h_2_destruct_r;
  Pointer_QTree_Int_t t1a8m_2_destruct_d;
  logic t1a8m_2_destruct_r;
  Pointer_QTree_Int_t q2a8i_2_destruct_d;
  logic q2a8i_2_destruct_r;
  Pointer_QTree_Int_t t2a8n_2_destruct_d;
  logic t2a8n_2_destruct_r;
  Pointer_CT$wmAdd_Int_t sc_0_3_destruct_d;
  logic sc_0_3_destruct_r;
  MyDTInt_Int_Int_t wsie_2_destruct_d;
  logic wsie_2_destruct_r;
  Pointer_QTree_Int_t q1a8h_1_destruct_d;
  logic q1a8h_1_destruct_r;
  Pointer_QTree_Int_t t1a8m_1_destruct_d;
  logic t1a8m_1_destruct_r;
  Pointer_QTree_Int_t q2a8i_1_destruct_d;
  logic q2a8i_1_destruct_r;
  Pointer_QTree_Int_t t2a8n_1_destruct_d;
  logic t2a8n_1_destruct_r;
  Pointer_QTree_Int_t q3a8j_1_destruct_d;
  logic q3a8j_1_destruct_r;
  Pointer_QTree_Int_t t3a8o_1_destruct_d;
  logic t3a8o_1_destruct_r;
  CT$wmAdd_Int_t _49_d;
  logic _49_r;
  assign _49_r = 1'd1;
  CT$wmAdd_Int_t lizzieLet22_1Lcall_$wmAdd_Int3_d;
  logic lizzieLet22_1Lcall_$wmAdd_Int3_r;
  CT$wmAdd_Int_t lizzieLet22_1Lcall_$wmAdd_Int2_d;
  logic lizzieLet22_1Lcall_$wmAdd_Int2_r;
  CT$wmAdd_Int_t lizzieLet22_1Lcall_$wmAdd_Int1_d;
  logic lizzieLet22_1Lcall_$wmAdd_Int1_r;
  CT$wmAdd_Int_t lizzieLet22_1Lcall_$wmAdd_Int0_d;
  logic lizzieLet22_1Lcall_$wmAdd_Int0_r;
  Go_t _48_d;
  logic _48_r;
  assign _48_r = 1'd1;
  Go_t lizzieLet22_3Lcall_$wmAdd_Int3_d;
  logic lizzieLet22_3Lcall_$wmAdd_Int3_r;
  Go_t lizzieLet22_3Lcall_$wmAdd_Int2_d;
  logic lizzieLet22_3Lcall_$wmAdd_Int2_r;
  Go_t lizzieLet22_3Lcall_$wmAdd_Int1_d;
  logic lizzieLet22_3Lcall_$wmAdd_Int1_r;
  Go_t lizzieLet22_3Lcall_$wmAdd_Int0_d;
  logic lizzieLet22_3Lcall_$wmAdd_Int0_r;
  Go_t lizzieLet22_3Lcall_$wmAdd_Int0_1_argbuf_d;
  logic lizzieLet22_3Lcall_$wmAdd_Int0_1_argbuf_r;
  Go_t lizzieLet22_3Lcall_$wmAdd_Int1_1_argbuf_d;
  logic lizzieLet22_3Lcall_$wmAdd_Int1_1_argbuf_r;
  Go_t lizzieLet22_3Lcall_$wmAdd_Int2_1_argbuf_d;
  logic lizzieLet22_3Lcall_$wmAdd_Int2_1_argbuf_r;
  Go_t lizzieLet22_3Lcall_$wmAdd_Int3_1_argbuf_d;
  logic lizzieLet22_3Lcall_$wmAdd_Int3_1_argbuf_r;
  Pointer_QTree_Int_t lizzieLet22_4L$wmAdd_Intsbos_d;
  logic lizzieLet22_4L$wmAdd_Intsbos_r;
  Pointer_QTree_Int_t lizzieLet22_4Lcall_$wmAdd_Int3_d;
  logic lizzieLet22_4Lcall_$wmAdd_Int3_r;
  Pointer_QTree_Int_t lizzieLet22_4Lcall_$wmAdd_Int2_d;
  logic lizzieLet22_4Lcall_$wmAdd_Int2_r;
  Pointer_QTree_Int_t lizzieLet22_4Lcall_$wmAdd_Int1_d;
  logic lizzieLet22_4Lcall_$wmAdd_Int1_r;
  Pointer_QTree_Int_t lizzieLet22_4Lcall_$wmAdd_Int0_d;
  logic lizzieLet22_4Lcall_$wmAdd_Int0_r;
  Pointer_QTree_Int_t lizzieLet22_4L$wmAdd_Intsbos_1_merge_merge_fork_1_d;
  logic lizzieLet22_4L$wmAdd_Intsbos_1_merge_merge_fork_1_r;
  Pointer_QTree_Int_t lizzieLet22_4L$wmAdd_Intsbos_1_merge_merge_fork_2_d;
  logic lizzieLet22_4L$wmAdd_Intsbos_1_merge_merge_fork_2_r;
  Go_t call_$wmAdd_Int_goConst_d;
  logic call_$wmAdd_Int_goConst_r;
  Pointer_QTree_Int_t \$wmAdd_Int_resbuf_d ;
  logic \$wmAdd_Int_resbuf_r ;
  QTree_Int_t lizzieLet22_4Lcall_$wmAdd_Int0_1es_2_1es_3_2_1es_4_2_1QNode_Int_d;
  logic lizzieLet22_4Lcall_$wmAdd_Int0_1es_2_1es_3_2_1es_4_2_1QNode_Int_r;
  QTree_Int_t lizzieLet26_1_argbuf_d;
  logic lizzieLet26_1_argbuf_r;
  CT$wmAdd_Int_t lizzieLet22_4Lcall_$wmAdd_Int1_1es_3_1_1es_4_1_1sc_0_5_1Lcall_$wmAdd_Int0_d;
  logic lizzieLet22_4Lcall_$wmAdd_Int1_1es_3_1_1es_4_1_1sc_0_5_1Lcall_$wmAdd_Int0_r;
  CT$wmAdd_Int_t lizzieLet25_1_argbuf_d;
  logic lizzieLet25_1_argbuf_r;
  CT$wmAdd_Int_t lizzieLet22_4Lcall_$wmAdd_Int2_1es_4_1sc_0_4_1wsie_3_1q1a8h_2_1t1a8m_2_1Lcall_$wmAdd_Int1_d;
  logic lizzieLet22_4Lcall_$wmAdd_Int2_1es_4_1sc_0_4_1wsie_3_1q1a8h_2_1t1a8m_2_1Lcall_$wmAdd_Int1_r;
  CT$wmAdd_Int_t lizzieLet24_1_argbuf_d;
  logic lizzieLet24_1_argbuf_r;
  CT$wmAdd_Int_t lizzieLet22_4Lcall_$wmAdd_Int3_1sc_0_3_1wsie_2_1q1a8h_1_1t1a8m_1_1q2a8i_1_1t2a8n_1_1Lcall_$wmAdd_Int2_d;
  logic lizzieLet22_4Lcall_$wmAdd_Int3_1sc_0_3_1wsie_2_1q1a8h_1_1t1a8m_1_1q2a8i_1_1t2a8n_1_1Lcall_$wmAdd_Int2_r;
  CT$wmAdd_Int_t lizzieLet23_1_argbuf_d;
  logic lizzieLet23_1_argbuf_r;
  \Int#_t  wwsim_4_destruct_d;
  logic wwsim_4_destruct_r;
  \Int#_t  ww1XiS_2_destruct_d;
  logic ww1XiS_2_destruct_r;
  \Int#_t  ww2XiV_1_destruct_d;
  logic ww2XiV_1_destruct_r;
  Pointer_CT$wnnz_Int_t sc_0_10_destruct_d;
  logic sc_0_10_destruct_r;
  \Int#_t  wwsim_3_destruct_d;
  logic wwsim_3_destruct_r;
  \Int#_t  ww1XiS_1_destruct_d;
  logic ww1XiS_1_destruct_r;
  Pointer_CT$wnnz_Int_t sc_0_9_destruct_d;
  logic sc_0_9_destruct_r;
  Pointer_QTree_Int_t q4a8F_3_destruct_d;
  logic q4a8F_3_destruct_r;
  \Int#_t  wwsim_2_destruct_d;
  logic wwsim_2_destruct_r;
  Pointer_CT$wnnz_Int_t sc_0_8_destruct_d;
  logic sc_0_8_destruct_r;
  Pointer_QTree_Int_t q4a8F_2_destruct_d;
  logic q4a8F_2_destruct_r;
  Pointer_QTree_Int_t q3a8E_2_destruct_d;
  logic q3a8E_2_destruct_r;
  Pointer_CT$wnnz_Int_t sc_0_7_destruct_d;
  logic sc_0_7_destruct_r;
  Pointer_QTree_Int_t q4a8F_1_destruct_d;
  logic q4a8F_1_destruct_r;
  Pointer_QTree_Int_t q3a8E_1_destruct_d;
  logic q3a8E_1_destruct_r;
  Pointer_QTree_Int_t q2a8D_1_destruct_d;
  logic q2a8D_1_destruct_r;
  CT$wnnz_Int_t _47_d;
  logic _47_r;
  assign _47_r = 1'd1;
  CT$wnnz_Int_t lizzieLet27_1Lcall_$wnnz_Int3_d;
  logic lizzieLet27_1Lcall_$wnnz_Int3_r;
  CT$wnnz_Int_t lizzieLet27_1Lcall_$wnnz_Int2_d;
  logic lizzieLet27_1Lcall_$wnnz_Int2_r;
  CT$wnnz_Int_t lizzieLet27_1Lcall_$wnnz_Int1_d;
  logic lizzieLet27_1Lcall_$wnnz_Int1_r;
  CT$wnnz_Int_t lizzieLet27_1Lcall_$wnnz_Int0_d;
  logic lizzieLet27_1Lcall_$wnnz_Int0_r;
  Go_t _46_d;
  logic _46_r;
  assign _46_r = 1'd1;
  Go_t lizzieLet27_3Lcall_$wnnz_Int3_d;
  logic lizzieLet27_3Lcall_$wnnz_Int3_r;
  Go_t lizzieLet27_3Lcall_$wnnz_Int2_d;
  logic lizzieLet27_3Lcall_$wnnz_Int2_r;
  Go_t lizzieLet27_3Lcall_$wnnz_Int1_d;
  logic lizzieLet27_3Lcall_$wnnz_Int1_r;
  Go_t lizzieLet27_3Lcall_$wnnz_Int0_d;
  logic lizzieLet27_3Lcall_$wnnz_Int0_r;
  Go_t lizzieLet27_3Lcall_$wnnz_Int0_1_argbuf_d;
  logic lizzieLet27_3Lcall_$wnnz_Int0_1_argbuf_r;
  Go_t lizzieLet27_3Lcall_$wnnz_Int1_1_argbuf_d;
  logic lizzieLet27_3Lcall_$wnnz_Int1_1_argbuf_r;
  Go_t lizzieLet27_3Lcall_$wnnz_Int2_1_argbuf_d;
  logic lizzieLet27_3Lcall_$wnnz_Int2_1_argbuf_r;
  Go_t lizzieLet27_3Lcall_$wnnz_Int3_1_argbuf_d;
  logic lizzieLet27_3Lcall_$wnnz_Int3_1_argbuf_r;
  \Int#_t  lizzieLet27_4L$wnnz_Intsbos_d;
  logic lizzieLet27_4L$wnnz_Intsbos_r;
  \Int#_t  lizzieLet27_4Lcall_$wnnz_Int3_d;
  logic lizzieLet27_4Lcall_$wnnz_Int3_r;
  \Int#_t  lizzieLet27_4Lcall_$wnnz_Int2_d;
  logic lizzieLet27_4Lcall_$wnnz_Int2_r;
  \Int#_t  lizzieLet27_4Lcall_$wnnz_Int1_d;
  logic lizzieLet27_4Lcall_$wnnz_Int1_r;
  \Int#_t  lizzieLet27_4Lcall_$wnnz_Int0_d;
  logic lizzieLet27_4Lcall_$wnnz_Int0_r;
  \Int#_t  lizzieLet27_4L$wnnz_Intsbos_1_merge_merge_fork_1_d;
  logic lizzieLet27_4L$wnnz_Intsbos_1_merge_merge_fork_1_r;
  \Int#_t  lizzieLet27_4L$wnnz_Intsbos_1_merge_merge_fork_2_d;
  logic lizzieLet27_4L$wnnz_Intsbos_1_merge_merge_fork_2_r;
  Go_t call_$wnnz_Int_goConst_d;
  logic call_$wnnz_Int_goConst_r;
  \Int#_t  \$wnnz_Int_resbuf_d ;
  logic \$wnnz_Int_resbuf_r ;
  CT$wnnz_Int_t lizzieLet27_4Lcall_$wnnz_Int3_1sc_0_7_1q4a8F_1_1q3a8E_1_1Lcall_$wnnz_Int2_d;
  logic lizzieLet27_4Lcall_$wnnz_Int3_1sc_0_7_1q4a8F_1_1q3a8E_1_1Lcall_$wnnz_Int2_r;
  CT$wnnz_Int_t lizzieLet28_1_argbuf_d;
  logic lizzieLet28_1_argbuf_r;
  Pointer_QTree_Int_t q1a8h_destruct_d;
  logic q1a8h_destruct_r;
  Pointer_QTree_Int_t q2a8i_destruct_d;
  logic q2a8i_destruct_r;
  Pointer_QTree_Int_t q3a8j_destruct_d;
  logic q3a8j_destruct_r;
  Pointer_QTree_Int_t q4a8k_destruct_d;
  logic q4a8k_destruct_r;
  Int_t v1a8b_destruct_d;
  logic v1a8b_destruct_r;
  QTree_Int_t _45_d;
  logic _45_r;
  assign _45_r = 1'd1;
  QTree_Int_t lizzieLet2_1QVal_Int_d;
  logic lizzieLet2_1QVal_Int_r;
  QTree_Int_t lizzieLet2_1QNode_Int_d;
  logic lizzieLet2_1QNode_Int_r;
  QTree_Int_t _44_d;
  logic _44_r;
  assign _44_r = 1'd1;
  Go_t lizzieLet2_3QNone_Int_d;
  logic lizzieLet2_3QNone_Int_r;
  Go_t lizzieLet2_3QVal_Int_d;
  logic lizzieLet2_3QVal_Int_r;
  Go_t lizzieLet2_3QNode_Int_d;
  logic lizzieLet2_3QNode_Int_r;
  Go_t lizzieLet2_3QError_Int_d;
  logic lizzieLet2_3QError_Int_r;
  Go_t lizzieLet2_3QError_Int_1_d;
  logic lizzieLet2_3QError_Int_1_r;
  Go_t lizzieLet2_3QError_Int_2_d;
  logic lizzieLet2_3QError_Int_2_r;
  QTree_Int_t lizzieLet2_3QError_Int_1QError_Int_d;
  logic lizzieLet2_3QError_Int_1QError_Int_r;
  QTree_Int_t lizzieLet11_1_1_argbuf_d;
  logic lizzieLet11_1_1_argbuf_r;
  Go_t lizzieLet2_3QError_Int_2_argbuf_d;
  logic lizzieLet2_3QError_Int_2_argbuf_r;
  Go_t lizzieLet2_3QNone_Int_1_argbuf_d;
  logic lizzieLet2_3QNone_Int_1_argbuf_r;
  C10_t go_10_goMux_choice_d;
  logic go_10_goMux_choice_r;
  Go_t go_10_goMux_data_d;
  logic go_10_goMux_data_r;
  QTree_Int_t _43_d;
  logic _43_r;
  assign _43_r = 1'd1;
  QTree_Int_t lizzieLet2_4QVal_Int_d;
  logic lizzieLet2_4QVal_Int_r;
  QTree_Int_t lizzieLet2_4QNode_Int_d;
  logic lizzieLet2_4QNode_Int_r;
  QTree_Int_t _42_d;
  logic _42_r;
  assign _42_r = 1'd1;
  QTree_Int_t lizzieLet2_4QNode_Int_1_d;
  logic lizzieLet2_4QNode_Int_1_r;
  QTree_Int_t lizzieLet2_4QNode_Int_2_d;
  logic lizzieLet2_4QNode_Int_2_r;
  QTree_Int_t lizzieLet2_4QNode_Int_3_d;
  logic lizzieLet2_4QNode_Int_3_r;
  QTree_Int_t lizzieLet2_4QNode_Int_4_d;
  logic lizzieLet2_4QNode_Int_4_r;
  QTree_Int_t lizzieLet2_4QNode_Int_5_d;
  logic lizzieLet2_4QNode_Int_5_r;
  QTree_Int_t lizzieLet2_4QNode_Int_6_d;
  logic lizzieLet2_4QNode_Int_6_r;
  QTree_Int_t lizzieLet2_4QNode_Int_7_d;
  logic lizzieLet2_4QNode_Int_7_r;
  QTree_Int_t lizzieLet2_4QNode_Int_8_d;
  logic lizzieLet2_4QNode_Int_8_r;
  QTree_Int_t lizzieLet2_4QNode_Int_9_d;
  logic lizzieLet2_4QNode_Int_9_r;
  QTree_Int_t lizzieLet2_4QNode_Int_10_d;
  logic lizzieLet2_4QNode_Int_10_r;
  Pointer_QTree_Int_t _41_d;
  logic _41_r;
  assign _41_r = 1'd1;
  Pointer_QTree_Int_t _40_d;
  logic _40_r;
  assign _40_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet2_4QNode_Int_10QNode_Int_d;
  logic lizzieLet2_4QNode_Int_10QNode_Int_r;
  Pointer_QTree_Int_t _39_d;
  logic _39_r;
  assign _39_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet2_4QNode_Int_10QNode_Int_1_argbuf_d;
  logic lizzieLet2_4QNode_Int_10QNode_Int_1_argbuf_r;
  Pointer_QTree_Int_t t1a8m_destruct_d;
  logic t1a8m_destruct_r;
  Pointer_QTree_Int_t t2a8n_destruct_d;
  logic t2a8n_destruct_r;
  Pointer_QTree_Int_t t3a8o_destruct_d;
  logic t3a8o_destruct_r;
  Pointer_QTree_Int_t t4a8p_destruct_d;
  logic t4a8p_destruct_r;
  QTree_Int_t _38_d;
  logic _38_r;
  assign _38_r = 1'd1;
  QTree_Int_t _37_d;
  logic _37_r;
  assign _37_r = 1'd1;
  QTree_Int_t lizzieLet2_4QNode_Int_1QNode_Int_d;
  logic lizzieLet2_4QNode_Int_1QNode_Int_r;
  QTree_Int_t _36_d;
  logic _36_r;
  assign _36_r = 1'd1;
  Go_t lizzieLet2_4QNode_Int_3QNone_Int_d;
  logic lizzieLet2_4QNode_Int_3QNone_Int_r;
  Go_t lizzieLet2_4QNode_Int_3QVal_Int_d;
  logic lizzieLet2_4QNode_Int_3QVal_Int_r;
  Go_t lizzieLet2_4QNode_Int_3QNode_Int_d;
  logic lizzieLet2_4QNode_Int_3QNode_Int_r;
  Go_t lizzieLet2_4QNode_Int_3QError_Int_d;
  logic lizzieLet2_4QNode_Int_3QError_Int_r;
  Go_t lizzieLet2_4QNode_Int_3QError_Int_1_d;
  logic lizzieLet2_4QNode_Int_3QError_Int_1_r;
  Go_t lizzieLet2_4QNode_Int_3QError_Int_2_d;
  logic lizzieLet2_4QNode_Int_3QError_Int_2_r;
  QTree_Int_t lizzieLet2_4QNode_Int_3QError_Int_1QError_Int_d;
  logic lizzieLet2_4QNode_Int_3QError_Int_1QError_Int_r;
  QTree_Int_t lizzieLet10_1_1_argbuf_d;
  logic lizzieLet10_1_1_argbuf_r;
  Go_t lizzieLet2_4QNode_Int_3QError_Int_2_argbuf_d;
  logic lizzieLet2_4QNode_Int_3QError_Int_2_argbuf_r;
  Go_t lizzieLet2_4QNode_Int_3QNode_Int_1_argbuf_d;
  logic lizzieLet2_4QNode_Int_3QNode_Int_1_argbuf_r;
  Go_t lizzieLet2_4QNode_Int_3QNone_Int_1_argbuf_d;
  logic lizzieLet2_4QNode_Int_3QNone_Int_1_argbuf_r;
  Go_t lizzieLet2_4QNode_Int_3QVal_Int_1_d;
  logic lizzieLet2_4QNode_Int_3QVal_Int_1_r;
  Go_t lizzieLet2_4QNode_Int_3QVal_Int_2_d;
  logic lizzieLet2_4QNode_Int_3QVal_Int_2_r;
  QTree_Int_t lizzieLet2_4QNode_Int_3QVal_Int_1QError_Int_d;
  logic lizzieLet2_4QNode_Int_3QVal_Int_1QError_Int_r;
  QTree_Int_t lizzieLet8_1_1_argbuf_d;
  logic lizzieLet8_1_1_argbuf_r;
  Go_t lizzieLet2_4QNode_Int_3QVal_Int_2_argbuf_d;
  logic lizzieLet2_4QNode_Int_3QVal_Int_2_argbuf_r;
  Pointer_CT$wmAdd_Int_t lizzieLet2_4QNode_Int_4QNone_Int_d;
  logic lizzieLet2_4QNode_Int_4QNone_Int_r;
  Pointer_CT$wmAdd_Int_t lizzieLet2_4QNode_Int_4QVal_Int_d;
  logic lizzieLet2_4QNode_Int_4QVal_Int_r;
  Pointer_CT$wmAdd_Int_t lizzieLet2_4QNode_Int_4QNode_Int_d;
  logic lizzieLet2_4QNode_Int_4QNode_Int_r;
  Pointer_CT$wmAdd_Int_t lizzieLet2_4QNode_Int_4QError_Int_d;
  logic lizzieLet2_4QNode_Int_4QError_Int_r;
  Pointer_CT$wmAdd_Int_t lizzieLet2_4QNode_Int_4QError_Int_1_argbuf_d;
  logic lizzieLet2_4QNode_Int_4QError_Int_1_argbuf_r;
  CT$wmAdd_Int_t lizzieLet2_4QNode_Int_4QNode_Int_1lizzieLet2_4QNode_Int_6QNode_Int_1lizzieLet2_4QNode_Int_7QNode_Int_1t1a8m_1lizzieLet2_4QNode_Int_8QNode_Int_1t2a8n_1lizzieLet2_4QNode_Int_9QNode_Int_1t3a8o_1Lcall_$wmAdd_Int3_d;
  logic lizzieLet2_4QNode_Int_4QNode_Int_1lizzieLet2_4QNode_Int_6QNode_Int_1lizzieLet2_4QNode_Int_7QNode_Int_1t1a8m_1lizzieLet2_4QNode_Int_8QNode_Int_1t2a8n_1lizzieLet2_4QNode_Int_9QNode_Int_1t3a8o_1Lcall_$wmAdd_Int3_r;
  CT$wmAdd_Int_t lizzieLet9_1_1_argbuf_d;
  logic lizzieLet9_1_1_argbuf_r;
  Pointer_CT$wmAdd_Int_t lizzieLet2_4QNode_Int_4QNone_Int_1_argbuf_d;
  logic lizzieLet2_4QNode_Int_4QNone_Int_1_argbuf_r;
  Pointer_CT$wmAdd_Int_t lizzieLet2_4QNode_Int_4QVal_Int_1_argbuf_d;
  logic lizzieLet2_4QNode_Int_4QVal_Int_1_argbuf_r;
  Pointer_QTree_Int_t lizzieLet2_4QNode_Int_5QNone_Int_d;
  logic lizzieLet2_4QNode_Int_5QNone_Int_r;
  Pointer_QTree_Int_t _35_d;
  logic _35_r;
  assign _35_r = 1'd1;
  Pointer_QTree_Int_t _34_d;
  logic _34_r;
  assign _34_r = 1'd1;
  Pointer_QTree_Int_t _33_d;
  logic _33_r;
  assign _33_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet2_4QNode_Int_5QNone_Int_1_argbuf_d;
  logic lizzieLet2_4QNode_Int_5QNone_Int_1_argbuf_r;
  MyDTInt_Int_Int_t _32_d;
  logic _32_r;
  assign _32_r = 1'd1;
  MyDTInt_Int_Int_t _31_d;
  logic _31_r;
  assign _31_r = 1'd1;
  MyDTInt_Int_Int_t lizzieLet2_4QNode_Int_6QNode_Int_d;
  logic lizzieLet2_4QNode_Int_6QNode_Int_r;
  MyDTInt_Int_Int_t _30_d;
  logic _30_r;
  assign _30_r = 1'd1;
  MyDTInt_Int_Int_t lizzieLet2_4QNode_Int_6QNode_Int_1_d;
  logic lizzieLet2_4QNode_Int_6QNode_Int_1_r;
  MyDTInt_Int_Int_t lizzieLet2_4QNode_Int_6QNode_Int_2_d;
  logic lizzieLet2_4QNode_Int_6QNode_Int_2_r;
  MyDTInt_Int_Int_t lizzieLet2_4QNode_Int_6QNode_Int_2_argbuf_d;
  logic lizzieLet2_4QNode_Int_6QNode_Int_2_argbuf_r;
  Pointer_QTree_Int_t _29_d;
  logic _29_r;
  assign _29_r = 1'd1;
  Pointer_QTree_Int_t _28_d;
  logic _28_r;
  assign _28_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet2_4QNode_Int_7QNode_Int_d;
  logic lizzieLet2_4QNode_Int_7QNode_Int_r;
  Pointer_QTree_Int_t _27_d;
  logic _27_r;
  assign _27_r = 1'd1;
  Pointer_QTree_Int_t _26_d;
  logic _26_r;
  assign _26_r = 1'd1;
  Pointer_QTree_Int_t _25_d;
  logic _25_r;
  assign _25_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet2_4QNode_Int_8QNode_Int_d;
  logic lizzieLet2_4QNode_Int_8QNode_Int_r;
  Pointer_QTree_Int_t _24_d;
  logic _24_r;
  assign _24_r = 1'd1;
  Pointer_QTree_Int_t _23_d;
  logic _23_r;
  assign _23_r = 1'd1;
  Pointer_QTree_Int_t _22_d;
  logic _22_r;
  assign _22_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet2_4QNode_Int_9QNode_Int_d;
  logic lizzieLet2_4QNode_Int_9QNode_Int_r;
  Pointer_QTree_Int_t _21_d;
  logic _21_r;
  assign _21_r = 1'd1;
  QTree_Int_t lizzieLet2_4QVal_Int_1_d;
  logic lizzieLet2_4QVal_Int_1_r;
  QTree_Int_t lizzieLet2_4QVal_Int_2_d;
  logic lizzieLet2_4QVal_Int_2_r;
  QTree_Int_t lizzieLet2_4QVal_Int_3_d;
  logic lizzieLet2_4QVal_Int_3_r;
  QTree_Int_t lizzieLet2_4QVal_Int_4_d;
  logic lizzieLet2_4QVal_Int_4_r;
  QTree_Int_t lizzieLet2_4QVal_Int_5_d;
  logic lizzieLet2_4QVal_Int_5_r;
  QTree_Int_t lizzieLet2_4QVal_Int_6_d;
  logic lizzieLet2_4QVal_Int_6_r;
  QTree_Int_t lizzieLet2_4QVal_Int_7_d;
  logic lizzieLet2_4QVal_Int_7_r;
  Int_t va8c_destruct_d;
  logic va8c_destruct_r;
  QTree_Int_t _20_d;
  logic _20_r;
  assign _20_r = 1'd1;
  QTree_Int_t lizzieLet2_4QVal_Int_1QVal_Int_d;
  logic lizzieLet2_4QVal_Int_1QVal_Int_r;
  QTree_Int_t _19_d;
  logic _19_r;
  assign _19_r = 1'd1;
  QTree_Int_t _18_d;
  logic _18_r;
  assign _18_r = 1'd1;
  Go_t lizzieLet2_4QVal_Int_3QNone_Int_d;
  logic lizzieLet2_4QVal_Int_3QNone_Int_r;
  Go_t lizzieLet2_4QVal_Int_3QVal_Int_d;
  logic lizzieLet2_4QVal_Int_3QVal_Int_r;
  Go_t lizzieLet2_4QVal_Int_3QNode_Int_d;
  logic lizzieLet2_4QVal_Int_3QNode_Int_r;
  Go_t lizzieLet2_4QVal_Int_3QError_Int_d;
  logic lizzieLet2_4QVal_Int_3QError_Int_r;
  Go_t lizzieLet2_4QVal_Int_3QError_Int_1_d;
  logic lizzieLet2_4QVal_Int_3QError_Int_1_r;
  Go_t lizzieLet2_4QVal_Int_3QError_Int_2_d;
  logic lizzieLet2_4QVal_Int_3QError_Int_2_r;
  QTree_Int_t lizzieLet2_4QVal_Int_3QError_Int_1QError_Int_d;
  logic lizzieLet2_4QVal_Int_3QError_Int_1QError_Int_r;
  QTree_Int_t lizzieLet6_1_argbuf_d;
  logic lizzieLet6_1_argbuf_r;
  Go_t lizzieLet2_4QVal_Int_3QError_Int_2_argbuf_d;
  logic lizzieLet2_4QVal_Int_3QError_Int_2_argbuf_r;
  Go_t lizzieLet2_4QVal_Int_3QNode_Int_1_d;
  logic lizzieLet2_4QVal_Int_3QNode_Int_1_r;
  Go_t lizzieLet2_4QVal_Int_3QNode_Int_2_d;
  logic lizzieLet2_4QVal_Int_3QNode_Int_2_r;
  QTree_Int_t lizzieLet2_4QVal_Int_3QNode_Int_1QError_Int_d;
  logic lizzieLet2_4QVal_Int_3QNode_Int_1QError_Int_r;
  QTree_Int_t lizzieLet5_1_argbuf_d;
  logic lizzieLet5_1_argbuf_r;
  Go_t lizzieLet2_4QVal_Int_3QNode_Int_2_argbuf_d;
  logic lizzieLet2_4QVal_Int_3QNode_Int_2_argbuf_r;
  Go_t lizzieLet2_4QVal_Int_3QNone_Int_1_argbuf_d;
  logic lizzieLet2_4QVal_Int_3QNone_Int_1_argbuf_r;
  Go_t lizzieLet2_4QVal_Int_3QVal_Int_1_argbuf_d;
  logic lizzieLet2_4QVal_Int_3QVal_Int_1_argbuf_r;
  Pointer_CT$wmAdd_Int_t lizzieLet2_4QVal_Int_4QNone_Int_d;
  logic lizzieLet2_4QVal_Int_4QNone_Int_r;
  Pointer_CT$wmAdd_Int_t lizzieLet2_4QVal_Int_4QVal_Int_d;
  logic lizzieLet2_4QVal_Int_4QVal_Int_r;
  Pointer_CT$wmAdd_Int_t lizzieLet2_4QVal_Int_4QNode_Int_d;
  logic lizzieLet2_4QVal_Int_4QNode_Int_r;
  Pointer_CT$wmAdd_Int_t lizzieLet2_4QVal_Int_4QError_Int_d;
  logic lizzieLet2_4QVal_Int_4QError_Int_r;
  Pointer_CT$wmAdd_Int_t lizzieLet2_4QVal_Int_4QError_Int_1_argbuf_d;
  logic lizzieLet2_4QVal_Int_4QError_Int_1_argbuf_r;
  Pointer_CT$wmAdd_Int_t lizzieLet2_4QVal_Int_4QNode_Int_1_argbuf_d;
  logic lizzieLet2_4QVal_Int_4QNode_Int_1_argbuf_r;
  Pointer_CT$wmAdd_Int_t lizzieLet2_4QVal_Int_4QNone_Int_1_argbuf_d;
  logic lizzieLet2_4QVal_Int_4QNone_Int_1_argbuf_r;
  Pointer_CT$wmAdd_Int_t lizzieLet2_4QVal_Int_4QVal_Int_1_argbuf_d;
  logic lizzieLet2_4QVal_Int_4QVal_Int_1_argbuf_r;
  Pointer_QTree_Int_t lizzieLet2_4QVal_Int_5QNone_Int_d;
  logic lizzieLet2_4QVal_Int_5QNone_Int_r;
  Pointer_QTree_Int_t _17_d;
  logic _17_r;
  assign _17_r = 1'd1;
  Pointer_QTree_Int_t _16_d;
  logic _16_r;
  assign _16_r = 1'd1;
  Pointer_QTree_Int_t _15_d;
  logic _15_r;
  assign _15_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet2_4QVal_Int_5QNone_Int_1_argbuf_d;
  logic lizzieLet2_4QVal_Int_5QNone_Int_1_argbuf_r;
  MyDTInt_Int_Int_t _14_d;
  logic _14_r;
  assign _14_r = 1'd1;
  MyDTInt_Int_Int_t lizzieLet2_4QVal_Int_6QVal_Int_d;
  logic lizzieLet2_4QVal_Int_6QVal_Int_r;
  MyDTInt_Int_Int_t _13_d;
  logic _13_r;
  assign _13_r = 1'd1;
  MyDTInt_Int_Int_t _12_d;
  logic _12_r;
  assign _12_r = 1'd1;
  MyDTInt_Int_Int_t lizzieLet2_4QVal_Int_6QVal_Int_1_argbuf_d;
  logic lizzieLet2_4QVal_Int_6QVal_Int_1_argbuf_r;
  TupMyDTInt_Int_Int___Int___Int_t applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_d;
  logic applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_r;
  Int_t _11_d;
  logic _11_r;
  assign _11_r = 1'd1;
  Int_t lizzieLet2_4QVal_Int_7QVal_Int_d;
  logic lizzieLet2_4QVal_Int_7QVal_Int_r;
  Int_t _10_d;
  logic _10_r;
  assign _10_r = 1'd1;
  Int_t _9_d;
  logic _9_r;
  assign _9_r = 1'd1;
  Int_t lizzieLet2_4QVal_Int_7QVal_Int_1_argbuf_d;
  logic lizzieLet2_4QVal_Int_7QVal_Int_1_argbuf_r;
  Pointer_CT$wmAdd_Int_t lizzieLet2_5QNone_Int_d;
  logic lizzieLet2_5QNone_Int_r;
  Pointer_CT$wmAdd_Int_t lizzieLet2_5QVal_Int_d;
  logic lizzieLet2_5QVal_Int_r;
  Pointer_CT$wmAdd_Int_t lizzieLet2_5QNode_Int_d;
  logic lizzieLet2_5QNode_Int_r;
  Pointer_CT$wmAdd_Int_t lizzieLet2_5QError_Int_d;
  logic lizzieLet2_5QError_Int_r;
  Pointer_CT$wmAdd_Int_t lizzieLet2_5QError_Int_1_argbuf_d;
  logic lizzieLet2_5QError_Int_1_argbuf_r;
  Pointer_CT$wmAdd_Int_t lizzieLet2_5QNone_Int_1_argbuf_d;
  logic lizzieLet2_5QNone_Int_1_argbuf_r;
  Pointer_QTree_Int_t _8_d;
  logic _8_r;
  assign _8_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet2_6QVal_Int_d;
  logic lizzieLet2_6QVal_Int_r;
  Pointer_QTree_Int_t lizzieLet2_6QNode_Int_d;
  logic lizzieLet2_6QNode_Int_r;
  Pointer_QTree_Int_t _7_d;
  logic _7_r;
  assign _7_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet2_7QNone_Int_d;
  logic lizzieLet2_7QNone_Int_r;
  Pointer_QTree_Int_t _6_d;
  logic _6_r;
  assign _6_r = 1'd1;
  Pointer_QTree_Int_t _5_d;
  logic _5_r;
  assign _5_r = 1'd1;
  Pointer_QTree_Int_t _4_d;
  logic _4_r;
  assign _4_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet2_7QNone_Int_1_argbuf_d;
  logic lizzieLet2_7QNone_Int_1_argbuf_r;
  MyDTInt_Int_Int_t _3_d;
  logic _3_r;
  assign _3_r = 1'd1;
  MyDTInt_Int_Int_t lizzieLet2_8QVal_Int_d;
  logic lizzieLet2_8QVal_Int_r;
  MyDTInt_Int_Int_t lizzieLet2_8QNode_Int_d;
  logic lizzieLet2_8QNode_Int_r;
  MyDTInt_Int_Int_t _2_d;
  logic _2_r;
  assign _2_r = 1'd1;
  Pointer_QTree_Int_t es_1_1_destruct_d;
  logic es_1_1_destruct_r;
  Pointer_QTree_Int_t es_2_2_destruct_d;
  logic es_2_2_destruct_r;
  Pointer_QTree_Int_t es_3_5_destruct_d;
  logic es_3_5_destruct_r;
  Pointer_CTmain_mask_Int_t sc_0_14_destruct_d;
  logic sc_0_14_destruct_r;
  Pointer_QTree_Int_t es_2_1_destruct_d;
  logic es_2_1_destruct_r;
  Pointer_QTree_Int_t es_3_4_destruct_d;
  logic es_3_4_destruct_r;
  Pointer_CTmain_mask_Int_t sc_0_13_destruct_d;
  logic sc_0_13_destruct_r;
  Pointer_QTree_Int_t t1a8x_3_destruct_d;
  logic t1a8x_3_destruct_r;
  Pointer_MaskQTree_t q1a8s_3_destruct_d;
  logic q1a8s_3_destruct_r;
  Pointer_QTree_Int_t es_3_3_destruct_d;
  logic es_3_3_destruct_r;
  Pointer_CTmain_mask_Int_t sc_0_12_destruct_d;
  logic sc_0_12_destruct_r;
  Pointer_QTree_Int_t t1a8x_2_destruct_d;
  logic t1a8x_2_destruct_r;
  Pointer_MaskQTree_t q1a8s_2_destruct_d;
  logic q1a8s_2_destruct_r;
  Pointer_QTree_Int_t t2a8y_2_destruct_d;
  logic t2a8y_2_destruct_r;
  Pointer_MaskQTree_t q2a8t_2_destruct_d;
  logic q2a8t_2_destruct_r;
  Pointer_CTmain_mask_Int_t sc_0_11_destruct_d;
  logic sc_0_11_destruct_r;
  Pointer_QTree_Int_t t1a8x_1_destruct_d;
  logic t1a8x_1_destruct_r;
  Pointer_MaskQTree_t q1a8s_1_destruct_d;
  logic q1a8s_1_destruct_r;
  Pointer_QTree_Int_t t2a8y_1_destruct_d;
  logic t2a8y_1_destruct_r;
  Pointer_MaskQTree_t q2a8t_1_destruct_d;
  logic q2a8t_1_destruct_r;
  Pointer_QTree_Int_t t3a8z_1_destruct_d;
  logic t3a8z_1_destruct_r;
  Pointer_MaskQTree_t q3a8u_1_destruct_d;
  logic q3a8u_1_destruct_r;
  CTmain_mask_Int_t _1_d;
  logic _1_r;
  assign _1_r = 1'd1;
  CTmain_mask_Int_t lizzieLet31_1Lcall_main_mask_Int3_d;
  logic lizzieLet31_1Lcall_main_mask_Int3_r;
  CTmain_mask_Int_t lizzieLet31_1Lcall_main_mask_Int2_d;
  logic lizzieLet31_1Lcall_main_mask_Int2_r;
  CTmain_mask_Int_t lizzieLet31_1Lcall_main_mask_Int1_d;
  logic lizzieLet31_1Lcall_main_mask_Int1_r;
  CTmain_mask_Int_t lizzieLet31_1Lcall_main_mask_Int0_d;
  logic lizzieLet31_1Lcall_main_mask_Int0_r;
  Go_t _0_d;
  logic _0_r;
  assign _0_r = 1'd1;
  Go_t lizzieLet31_3Lcall_main_mask_Int3_d;
  logic lizzieLet31_3Lcall_main_mask_Int3_r;
  Go_t lizzieLet31_3Lcall_main_mask_Int2_d;
  logic lizzieLet31_3Lcall_main_mask_Int2_r;
  Go_t lizzieLet31_3Lcall_main_mask_Int1_d;
  logic lizzieLet31_3Lcall_main_mask_Int1_r;
  Go_t lizzieLet31_3Lcall_main_mask_Int0_d;
  logic lizzieLet31_3Lcall_main_mask_Int0_r;
  Go_t lizzieLet31_3Lcall_main_mask_Int0_1_argbuf_d;
  logic lizzieLet31_3Lcall_main_mask_Int0_1_argbuf_r;
  Go_t lizzieLet31_3Lcall_main_mask_Int1_1_argbuf_d;
  logic lizzieLet31_3Lcall_main_mask_Int1_1_argbuf_r;
  Go_t lizzieLet31_3Lcall_main_mask_Int2_1_argbuf_d;
  logic lizzieLet31_3Lcall_main_mask_Int2_1_argbuf_r;
  Go_t lizzieLet31_3Lcall_main_mask_Int3_1_argbuf_d;
  logic lizzieLet31_3Lcall_main_mask_Int3_1_argbuf_r;
  Pointer_QTree_Int_t lizzieLet31_4Lmain_mask_Intsbos_d;
  logic lizzieLet31_4Lmain_mask_Intsbos_r;
  Pointer_QTree_Int_t lizzieLet31_4Lcall_main_mask_Int3_d;
  logic lizzieLet31_4Lcall_main_mask_Int3_r;
  Pointer_QTree_Int_t lizzieLet31_4Lcall_main_mask_Int2_d;
  logic lizzieLet31_4Lcall_main_mask_Int2_r;
  Pointer_QTree_Int_t lizzieLet31_4Lcall_main_mask_Int1_d;
  logic lizzieLet31_4Lcall_main_mask_Int1_r;
  Pointer_QTree_Int_t lizzieLet31_4Lcall_main_mask_Int0_d;
  logic lizzieLet31_4Lcall_main_mask_Int0_r;
  QTree_Int_t lizzieLet31_4Lcall_main_mask_Int0_1es_1_1_1es_2_2_1es_3_5_1QNode_Int_d;
  logic lizzieLet31_4Lcall_main_mask_Int0_1es_1_1_1es_2_2_1es_3_5_1QNode_Int_r;
  QTree_Int_t lizzieLet35_1_argbuf_d;
  logic lizzieLet35_1_argbuf_r;
  CTmain_mask_Int_t lizzieLet31_4Lcall_main_mask_Int1_1es_2_1_1es_3_4_1sc_0_13_1Lcall_main_mask_Int0_d;
  logic lizzieLet31_4Lcall_main_mask_Int1_1es_2_1_1es_3_4_1sc_0_13_1Lcall_main_mask_Int0_r;
  CTmain_mask_Int_t lizzieLet34_1_argbuf_d;
  logic lizzieLet34_1_argbuf_r;
  CTmain_mask_Int_t lizzieLet31_4Lcall_main_mask_Int2_1es_3_3_1sc_0_12_1t1a8x_2_1q1a8s_2_1Lcall_main_mask_Int1_d;
  logic lizzieLet31_4Lcall_main_mask_Int2_1es_3_3_1sc_0_12_1t1a8x_2_1q1a8s_2_1Lcall_main_mask_Int1_r;
  CTmain_mask_Int_t lizzieLet33_1_argbuf_d;
  logic lizzieLet33_1_argbuf_r;
  CTmain_mask_Int_t lizzieLet31_4Lcall_main_mask_Int3_1sc_0_11_1t1a8x_1_1q1a8s_1_1t2a8y_1_1q2a8t_1_1Lcall_main_mask_Int2_d;
  logic lizzieLet31_4Lcall_main_mask_Int3_1sc_0_11_1t1a8x_1_1q1a8s_1_1t2a8y_1_1q2a8t_1_1Lcall_main_mask_Int2_r;
  CTmain_mask_Int_t lizzieLet32_1_argbuf_d;
  logic lizzieLet32_1_argbuf_r;
  Pointer_QTree_Int_t lizzieLet31_4Lmain_mask_Intsbos_1_merge_merge_fork_1_d;
  logic lizzieLet31_4Lmain_mask_Intsbos_1_merge_merge_fork_1_r;
  Pointer_QTree_Int_t lizzieLet31_4Lmain_mask_Intsbos_1_merge_merge_fork_2_d;
  logic lizzieLet31_4Lmain_mask_Intsbos_1_merge_merge_fork_2_r;
  Go_t call_main_mask_Int_goConst_d;
  logic call_main_mask_Int_goConst_r;
  Pointer_QTree_Int_t main_mask_Int_resbuf_d;
  logic main_mask_Int_resbuf_r;
  Pointer_QTree_Int_t ma8q_1_argbuf_d;
  logic ma8q_1_argbuf_r;
  Pointer_QTree_Int_t ma8q_1_d;
  logic ma8q_1_r;
  Pointer_QTree_Int_t ma8q_2_d;
  logic ma8q_2_r;
  Go_t main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreego_9_d;
  logic main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreego_9_r;
  Pointer_QTree_Int_t main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreema8q_1_d;
  logic main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreema8q_1_r;
  Pointer_MaskQTree_t main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreemska8r_1_d;
  logic main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreemska8r_1_r;
  Go_t go_9_1_d;
  logic go_9_1_r;
  Go_t go_9_2_d;
  logic go_9_2_r;
  Pointer_QTree_Int_t ma8q_1_1_argbuf_d;
  logic ma8q_1_1_argbuf_r;
  Pointer_MaskQTree_t mska8r_1_1_argbuf_d;
  logic mska8r_1_1_argbuf_r;
  Pointer_QTree_Int_t es_0_1_argbuf_d;
  logic es_0_1_argbuf_r;
  Pointer_MaskQTree_t mska8r_1_argbuf_d;
  logic mska8r_1_argbuf_r;
  Pointer_QTree_Int_t q1a8C_1_argbuf_d;
  logic q1a8C_1_argbuf_r;
  Pointer_QTree_Int_t q1a8h_3_1_argbuf_d;
  logic q1a8h_3_1_argbuf_r;
  Pointer_MaskQTree_t q1a8s_3_1_argbuf_d;
  logic q1a8s_3_1_argbuf_r;
  Pointer_QTree_Int_t q2a8D_1_1_argbuf_d;
  logic q2a8D_1_1_argbuf_r;
  Pointer_QTree_Int_t q2a8i_2_1_argbuf_d;
  logic q2a8i_2_1_argbuf_r;
  Pointer_MaskQTree_t q2a8t_2_1_argbuf_d;
  logic q2a8t_2_1_argbuf_r;
  Pointer_QTree_Int_t q3a8E_2_1_argbuf_d;
  logic q3a8E_2_1_argbuf_r;
  Pointer_QTree_Int_t q3a8j_1_1_argbuf_d;
  logic q3a8j_1_1_argbuf_r;
  Pointer_MaskQTree_t q3a8u_1_1_argbuf_d;
  logic q3a8u_1_1_argbuf_r;
  Pointer_QTree_Int_t q4a8F_3_1_argbuf_d;
  logic q4a8F_3_1_argbuf_r;
  CT$wmAdd_Int_t readPointer_CT$wmAdd_Intscfarg_0_1_argbuf_rwb_d;
  logic readPointer_CT$wmAdd_Intscfarg_0_1_argbuf_rwb_r;
  CT$wmAdd_Int_t lizzieLet22_1_d;
  logic lizzieLet22_1_r;
  CT$wmAdd_Int_t lizzieLet22_2_d;
  logic lizzieLet22_2_r;
  CT$wmAdd_Int_t lizzieLet22_3_d;
  logic lizzieLet22_3_r;
  CT$wmAdd_Int_t lizzieLet22_4_d;
  logic lizzieLet22_4_r;
  CT$wnnz_Int_t readPointer_CT$wnnz_Intscfarg_0_1_1_argbuf_rwb_d;
  logic readPointer_CT$wnnz_Intscfarg_0_1_1_argbuf_rwb_r;
  CT$wnnz_Int_t lizzieLet27_1_d;
  logic lizzieLet27_1_r;
  CT$wnnz_Int_t lizzieLet27_2_d;
  logic lizzieLet27_2_r;
  CT$wnnz_Int_t lizzieLet27_3_d;
  logic lizzieLet27_3_r;
  CT$wnnz_Int_t lizzieLet27_4_d;
  logic lizzieLet27_4_r;
  CTmain_mask_Int_t readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf_rwb_d;
  logic readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf_rwb_r;
  CTmain_mask_Int_t lizzieLet31_1_d;
  logic lizzieLet31_1_r;
  CTmain_mask_Int_t lizzieLet31_2_d;
  logic lizzieLet31_2_r;
  CTmain_mask_Int_t lizzieLet31_3_d;
  logic lizzieLet31_3_r;
  CTmain_mask_Int_t lizzieLet31_4_d;
  logic lizzieLet31_4_r;
  MaskQTree_t readPointer_MaskQTreemska8r_1_argbuf_rwb_d;
  logic readPointer_MaskQTreemska8r_1_argbuf_rwb_r;
  MaskQTree_t lizzieLet14_1_1_d;
  logic lizzieLet14_1_1_r;
  MaskQTree_t lizzieLet14_1_2_d;
  logic lizzieLet14_1_2_r;
  MaskQTree_t lizzieLet14_1_3_d;
  logic lizzieLet14_1_3_r;
  MaskQTree_t lizzieLet14_1_4_d;
  logic lizzieLet14_1_4_r;
  MaskQTree_t lizzieLet14_1_5_d;
  logic lizzieLet14_1_5_r;
  MaskQTree_t lizzieLet14_1_6_d;
  logic lizzieLet14_1_6_r;
  QTree_Int_t readPointer_QTree_Intma8q_1_argbuf_rwb_d;
  logic readPointer_QTree_Intma8q_1_argbuf_rwb_r;
  QTree_Int_t readPointer_QTree_Intw1sif_1_1_argbuf_rwb_d;
  logic readPointer_QTree_Intw1sif_1_1_argbuf_rwb_r;
  QTree_Int_t lizzieLet2_1_d;
  logic lizzieLet2_1_r;
  QTree_Int_t lizzieLet2_2_d;
  logic lizzieLet2_2_r;
  QTree_Int_t lizzieLet2_3_d;
  logic lizzieLet2_3_r;
  QTree_Int_t lizzieLet2_4_d;
  logic lizzieLet2_4_r;
  QTree_Int_t lizzieLet2_5_d;
  logic lizzieLet2_5_r;
  QTree_Int_t lizzieLet2_6_d;
  logic lizzieLet2_6_r;
  QTree_Int_t lizzieLet2_7_d;
  logic lizzieLet2_7_r;
  QTree_Int_t lizzieLet2_8_d;
  logic lizzieLet2_8_r;
  QTree_Int_t readPointer_QTree_Intw2sig_1_1_argbuf_rwb_d;
  logic readPointer_QTree_Intw2sig_1_1_argbuf_rwb_r;
  QTree_Int_t readPointer_QTree_Intwsij_1_1_argbuf_rwb_d;
  logic readPointer_QTree_Intwsij_1_1_argbuf_rwb_r;
  QTree_Int_t lizzieLet12_1_1_d;
  logic lizzieLet12_1_1_r;
  QTree_Int_t lizzieLet12_1_2_d;
  logic lizzieLet12_1_2_r;
  QTree_Int_t lizzieLet12_1_3_d;
  logic lizzieLet12_1_3_r;
  QTree_Int_t lizzieLet12_1_4_d;
  logic lizzieLet12_1_4_r;
  Pointer_CT$wnnz_Int_t sc_0_10_1_argbuf_d;
  logic sc_0_10_1_argbuf_r;
  Pointer_CTmain_mask_Int_t sc_0_14_1_argbuf_d;
  logic sc_0_14_1_argbuf_r;
  Pointer_CT$wmAdd_Int_t sc_0_6_1_argbuf_d;
  logic sc_0_6_1_argbuf_r;
  Pointer_CT$wnnz_Int_t scfarg_0_1_1_argbuf_d;
  logic scfarg_0_1_1_argbuf_r;
  Pointer_CTmain_mask_Int_t scfarg_0_2_1_argbuf_d;
  logic scfarg_0_2_1_argbuf_r;
  Pointer_CT$wmAdd_Int_t scfarg_0_1_argbuf_d;
  logic scfarg_0_1_argbuf_r;
  Pointer_QTree_Int_t t1a8m_3_1_argbuf_d;
  logic t1a8m_3_1_argbuf_r;
  Pointer_QTree_Int_t t1a8x_3_1_argbuf_d;
  logic t1a8x_3_1_argbuf_r;
  Pointer_QTree_Int_t t2a8n_2_1_argbuf_d;
  logic t2a8n_2_1_argbuf_r;
  Pointer_QTree_Int_t t2a8y_2_1_argbuf_d;
  logic t2a8y_2_1_argbuf_r;
  Pointer_QTree_Int_t t3a8o_1_1_argbuf_d;
  logic t3a8o_1_1_argbuf_r;
  Pointer_QTree_Int_t t3a8z_1_1_argbuf_d;
  logic t3a8z_1_1_argbuf_r;
  Pointer_QTree_Int_t t4a8A_1_argbuf_d;
  logic t4a8A_1_argbuf_r;
  Pointer_QTree_Int_t t4a8p_1_argbuf_d;
  logic t4a8p_1_argbuf_r;
  Int_t va8c_1_argbuf_d;
  logic va8c_1_argbuf_r;
  Pointer_QTree_Int_t w1sif_1_1_argbuf_d;
  logic w1sif_1_1_argbuf_r;
  Pointer_QTree_Int_t w1sif_1_1_d;
  logic w1sif_1_1_r;
  Pointer_QTree_Int_t w1sif_1_2_d;
  logic w1sif_1_2_r;
  Pointer_QTree_Int_t w2sig_1_1_argbuf_d;
  logic w2sig_1_1_argbuf_r;
  Pointer_QTree_Int_t w2sig_1_1_d;
  logic w2sig_1_1_r;
  Pointer_QTree_Int_t w2sig_1_2_d;
  logic w2sig_1_2_r;
  Pointer_CT$wmAdd_Int_t writeCT$wmAdd_IntlizzieLet0_1_argbuf_rwb_d;
  logic writeCT$wmAdd_IntlizzieLet0_1_argbuf_rwb_r;
  Pointer_CT$wmAdd_Int_t lizzieLet14_1_argbuf_d;
  logic lizzieLet14_1_argbuf_r;
  Pointer_CT$wmAdd_Int_t writeCT$wmAdd_IntlizzieLet23_1_argbuf_rwb_d;
  logic writeCT$wmAdd_IntlizzieLet23_1_argbuf_rwb_r;
  Pointer_CT$wmAdd_Int_t sca2_1_argbuf_d;
  logic sca2_1_argbuf_r;
  Pointer_CT$wmAdd_Int_t writeCT$wmAdd_IntlizzieLet24_1_argbuf_rwb_d;
  logic writeCT$wmAdd_IntlizzieLet24_1_argbuf_rwb_r;
  Pointer_CT$wmAdd_Int_t sca1_1_argbuf_d;
  logic sca1_1_argbuf_r;
  Pointer_CT$wmAdd_Int_t writeCT$wmAdd_IntlizzieLet25_1_argbuf_rwb_d;
  logic writeCT$wmAdd_IntlizzieLet25_1_argbuf_rwb_r;
  Pointer_CT$wmAdd_Int_t sca0_1_argbuf_d;
  logic sca0_1_argbuf_r;
  Pointer_CT$wmAdd_Int_t writeCT$wmAdd_IntlizzieLet9_1_1_argbuf_rwb_d;
  logic writeCT$wmAdd_IntlizzieLet9_1_1_argbuf_rwb_r;
  Pointer_CT$wmAdd_Int_t sca3_1_argbuf_d;
  logic sca3_1_argbuf_r;
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet13_1_1_argbuf_rwb_d;
  logic writeCT$wnnz_IntlizzieLet13_1_1_argbuf_rwb_r;
  Pointer_CT$wnnz_Int_t sca3_1_1_argbuf_d;
  logic sca3_1_1_argbuf_r;
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet1_1_argbuf_rwb_d;
  logic writeCT$wnnz_IntlizzieLet1_1_argbuf_rwb_r;
  Pointer_CT$wnnz_Int_t lizzieLet7_1_argbuf_d;
  logic lizzieLet7_1_argbuf_r;
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet28_1_argbuf_rwb_d;
  logic writeCT$wnnz_IntlizzieLet28_1_argbuf_rwb_r;
  Pointer_CT$wnnz_Int_t sca2_1_1_argbuf_d;
  logic sca2_1_1_argbuf_r;
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet29_1_argbuf_rwb_d;
  logic writeCT$wnnz_IntlizzieLet29_1_argbuf_rwb_r;
  Pointer_CT$wnnz_Int_t sca1_1_1_argbuf_d;
  logic sca1_1_1_argbuf_r;
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet30_1_argbuf_rwb_d;
  logic writeCT$wnnz_IntlizzieLet30_1_argbuf_rwb_r;
  Pointer_CT$wnnz_Int_t sca0_1_1_argbuf_d;
  logic sca0_1_1_argbuf_r;
  Pointer_CTmain_mask_Int_t writeCTmain_mask_IntlizzieLet19_1_argbuf_rwb_d;
  logic writeCTmain_mask_IntlizzieLet19_1_argbuf_rwb_r;
  Pointer_CTmain_mask_Int_t sca3_2_1_argbuf_d;
  logic sca3_2_1_argbuf_r;
  Pointer_CTmain_mask_Int_t writeCTmain_mask_IntlizzieLet21_1_argbuf_rwb_d;
  logic writeCTmain_mask_IntlizzieLet21_1_argbuf_rwb_r;
  Pointer_CTmain_mask_Int_t lizzieLet4_1_1_argbuf_d;
  logic lizzieLet4_1_1_argbuf_r;
  Pointer_CTmain_mask_Int_t writeCTmain_mask_IntlizzieLet32_1_argbuf_rwb_d;
  logic writeCTmain_mask_IntlizzieLet32_1_argbuf_rwb_r;
  Pointer_CTmain_mask_Int_t sca2_2_1_argbuf_d;
  logic sca2_2_1_argbuf_r;
  Pointer_CTmain_mask_Int_t writeCTmain_mask_IntlizzieLet33_1_argbuf_rwb_d;
  logic writeCTmain_mask_IntlizzieLet33_1_argbuf_rwb_r;
  Pointer_CTmain_mask_Int_t sca1_2_1_argbuf_d;
  logic sca1_2_1_argbuf_r;
  Pointer_CTmain_mask_Int_t writeCTmain_mask_IntlizzieLet34_1_argbuf_rwb_d;
  logic writeCTmain_mask_IntlizzieLet34_1_argbuf_rwb_r;
  Pointer_CTmain_mask_Int_t sca0_2_1_argbuf_d;
  logic sca0_2_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet10_1_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet10_1_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet12_1_argbuf_d;
  logic lizzieLet12_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet11_1_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet11_1_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet13_1_argbuf_d;
  logic lizzieLet13_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet15_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet15_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet0_1_1_argbuf_d;
  logic lizzieLet0_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet17_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet17_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet1_1_1_argbuf_d;
  logic lizzieLet1_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet18_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet18_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet2_1_1_argbuf_d;
  logic lizzieLet2_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet20_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet20_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet3_1_1_argbuf_d;
  logic lizzieLet3_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet26_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet26_1_argbuf_rwb_r;
  Pointer_QTree_Int_t contRet_0_1_argbuf_d;
  logic contRet_0_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet35_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet35_1_argbuf_rwb_r;
  Pointer_QTree_Int_t contRet_0_2_1_argbuf_d;
  logic contRet_0_2_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet4_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet4_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet8_1_argbuf_d;
  logic lizzieLet8_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet5_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet5_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet9_1_argbuf_d;
  logic lizzieLet9_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet6_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet6_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet10_1_argbuf_d;
  logic lizzieLet10_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet8_1_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet8_1_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet11_1_argbuf_d;
  logic lizzieLet11_1_argbuf_r;
  MyDTInt_Int_Int_t wsie_2_2_argbuf_d;
  logic wsie_2_2_argbuf_r;
  MyDTInt_Int_Int_t wsie_2_1_d;
  logic wsie_2_1_r;
  MyDTInt_Int_Int_t wsie_2_2_d;
  logic wsie_2_2_r;
  MyDTInt_Int_Int_t wsie_3_2_argbuf_d;
  logic wsie_3_2_argbuf_r;
  MyDTInt_Int_Int_t wsie_3_1_d;
  logic wsie_3_1_r;
  MyDTInt_Int_Int_t wsie_3_2_d;
  logic wsie_3_2_r;
  MyDTInt_Int_Int_t wsie_4_1_argbuf_d;
  logic wsie_4_1_argbuf_r;
  Pointer_QTree_Int_t wsij_1_1_argbuf_d;
  logic wsij_1_1_argbuf_r;
  CT$wnnz_Int_t lizzieLet29_1_argbuf_d;
  logic lizzieLet29_1_argbuf_r;
  CT$wnnz_Int_t wwsim_2_1lizzieLet27_4Lcall_$wnnz_Int2_1sc_0_8_1q4a8F_2_1Lcall_$wnnz_Int1_d;
  logic wwsim_2_1lizzieLet27_4Lcall_$wnnz_Int2_1sc_0_8_1q4a8F_2_1Lcall_$wnnz_Int1_r;
  CT$wnnz_Int_t lizzieLet30_1_argbuf_d;
  logic lizzieLet30_1_argbuf_r;
  CT$wnnz_Int_t wwsim_3_1ww1XiS_1_1lizzieLet27_4Lcall_$wnnz_Int1_1sc_0_9_1Lcall_$wnnz_Int0_d;
  logic wwsim_3_1ww1XiS_1_1lizzieLet27_4Lcall_$wnnz_Int1_1sc_0_9_1Lcall_$wnnz_Int0_r;
  \Int#_t  es_6_1_1ww2XiV_1_1_Add32_d;
  logic es_6_1_1ww2XiV_1_1_Add32_r;
  \Int#_t  wwsim_4_1ww1XiS_2_1_Add32_d;
  logic wwsim_4_1ww1XiS_2_1_Add32_r;
  
  /* fork (Ty Go) : (sourceGo,Go) > [(go_1,Go),
                                (go_2,Go),
                                (go_3,Go),
                                (go_4,Go),
                                (go__5,Go),
                                (go__6,Go),
                                (go__7,Go),
                                (go__8,Go),
                                (go__9,Go),
                                (go__10,Go)] */
  logic [9:0] sourceGo_emitted;
  logic [9:0] sourceGo_done;
  assign go_1_d = (sourceGo_d[0] && (! sourceGo_emitted[0]));
  assign go_2_d = (sourceGo_d[0] && (! sourceGo_emitted[1]));
  assign go_3_d = (sourceGo_d[0] && (! sourceGo_emitted[2]));
  assign go_4_d = (sourceGo_d[0] && (! sourceGo_emitted[3]));
  assign go__5_d = (sourceGo_d[0] && (! sourceGo_emitted[4]));
  assign go__6_d = (sourceGo_d[0] && (! sourceGo_emitted[5]));
  assign go__7_d = (sourceGo_d[0] && (! sourceGo_emitted[6]));
  assign go__8_d = (sourceGo_d[0] && (! sourceGo_emitted[7]));
  assign go__9_d = (sourceGo_d[0] && (! sourceGo_emitted[8]));
  assign go__10_d = (sourceGo_d[0] && (! sourceGo_emitted[9]));
  assign sourceGo_done = (sourceGo_emitted | ({go__10_d[0],
                                               go__9_d[0],
                                               go__8_d[0],
                                               go__7_d[0],
                                               go__6_d[0],
                                               go__5_d[0],
                                               go_4_d[0],
                                               go_3_d[0],
                                               go_2_d[0],
                                               go_1_d[0]} & {go__10_r,
                                                             go__9_r,
                                                             go__8_r,
                                                             go__7_r,
                                                             go__6_r,
                                                             go__5_r,
                                                             go_4_r,
                                                             go_3_r,
                                                             go_2_r,
                                                             go_1_r}));
  assign sourceGo_r = (& sourceGo_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) sourceGo_emitted <= 10'd0;
    else
      sourceGo_emitted <= (sourceGo_r ? 10'd0 :
                           sourceGo_done);
  
  /* const (Ty Word16#,
       Lit 0) : (go__5,Go) > (initHP_CT$wmAdd_Int,Word16#) */
  assign initHP_CT$wmAdd_Int_d = {16'd0, go__5_d[0]};
  assign go__5_r = initHP_CT$wmAdd_Int_r;
  
  /* const (Ty Word16#,
       Lit 1) : (incrHP_CT$wmAdd_Int1,Go) > (incrHP_CT$wmAdd_Int,Word16#) */
  assign incrHP_CT$wmAdd_Int_d = {16'd1, incrHP_CT$wmAdd_Int1_d[0]};
  assign incrHP_CT$wmAdd_Int1_r = incrHP_CT$wmAdd_Int_r;
  
  /* merge (Ty Go) : [(go__6,Go),
                 (incrHP_CT$wmAdd_Int2,Go)] > (incrHP_mergeCT$wmAdd_Int,Go) */
  logic [1:0] incrHP_mergeCT$wmAdd_Int_selected;
  logic [1:0] incrHP_mergeCT$wmAdd_Int_select;
  always_comb
    begin
      incrHP_mergeCT$wmAdd_Int_selected = 2'd0;
      if ((| incrHP_mergeCT$wmAdd_Int_select))
        incrHP_mergeCT$wmAdd_Int_selected = incrHP_mergeCT$wmAdd_Int_select;
      else
        if (go__6_d[0]) incrHP_mergeCT$wmAdd_Int_selected[0] = 1'd1;
        else if (incrHP_CT$wmAdd_Int2_d[0])
          incrHP_mergeCT$wmAdd_Int_selected[1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeCT$wmAdd_Int_select <= 2'd0;
    else
      incrHP_mergeCT$wmAdd_Int_select <= (incrHP_mergeCT$wmAdd_Int_r ? 2'd0 :
                                          incrHP_mergeCT$wmAdd_Int_selected);
  always_comb
    if (incrHP_mergeCT$wmAdd_Int_selected[0])
      incrHP_mergeCT$wmAdd_Int_d = go__6_d;
    else if (incrHP_mergeCT$wmAdd_Int_selected[1])
      incrHP_mergeCT$wmAdd_Int_d = incrHP_CT$wmAdd_Int2_d;
    else incrHP_mergeCT$wmAdd_Int_d = 1'd0;
  assign {incrHP_CT$wmAdd_Int2_r,
          go__6_r} = (incrHP_mergeCT$wmAdd_Int_r ? incrHP_mergeCT$wmAdd_Int_selected :
                      2'd0);
  
  /* fork (Ty Go) : (incrHP_mergeCT$wmAdd_Int_buf,Go) > [(incrHP_CT$wmAdd_Int1,Go),
                                                    (incrHP_CT$wmAdd_Int2,Go)] */
  logic [1:0] incrHP_mergeCT$wmAdd_Int_buf_emitted;
  logic [1:0] incrHP_mergeCT$wmAdd_Int_buf_done;
  assign incrHP_CT$wmAdd_Int1_d = (incrHP_mergeCT$wmAdd_Int_buf_d[0] && (! incrHP_mergeCT$wmAdd_Int_buf_emitted[0]));
  assign incrHP_CT$wmAdd_Int2_d = (incrHP_mergeCT$wmAdd_Int_buf_d[0] && (! incrHP_mergeCT$wmAdd_Int_buf_emitted[1]));
  assign incrHP_mergeCT$wmAdd_Int_buf_done = (incrHP_mergeCT$wmAdd_Int_buf_emitted | ({incrHP_CT$wmAdd_Int2_d[0],
                                                                                       incrHP_CT$wmAdd_Int1_d[0]} & {incrHP_CT$wmAdd_Int2_r,
                                                                                                                     incrHP_CT$wmAdd_Int1_r}));
  assign incrHP_mergeCT$wmAdd_Int_buf_r = (& incrHP_mergeCT$wmAdd_Int_buf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeCT$wmAdd_Int_buf_emitted <= 2'd0;
    else
      incrHP_mergeCT$wmAdd_Int_buf_emitted <= (incrHP_mergeCT$wmAdd_Int_buf_r ? 2'd0 :
                                               incrHP_mergeCT$wmAdd_Int_buf_done);
  
  /* op_add (Ty Word16#) : (incrHP_CT$wmAdd_Int,Word16#) (forkHP1_CT$wmAdd_Int,Word16#) > (addHP_CT$wmAdd_Int,Word16#) */
  assign addHP_CT$wmAdd_Int_d = {(incrHP_CT$wmAdd_Int_d[16:1] + forkHP1_CT$wmAdd_Int_d[16:1]),
                                 (incrHP_CT$wmAdd_Int_d[0] && forkHP1_CT$wmAdd_Int_d[0])};
  assign {incrHP_CT$wmAdd_Int_r,
          forkHP1_CT$wmAdd_Int_r} = {2 {(addHP_CT$wmAdd_Int_r && addHP_CT$wmAdd_Int_d[0])}};
  
  /* merge (Ty Word16#) : [(initHP_CT$wmAdd_Int,Word16#),
                      (addHP_CT$wmAdd_Int,Word16#)] > (mergeHP_CT$wmAdd_Int,Word16#) */
  logic [1:0] mergeHP_CT$wmAdd_Int_selected;
  logic [1:0] mergeHP_CT$wmAdd_Int_select;
  always_comb
    begin
      mergeHP_CT$wmAdd_Int_selected = 2'd0;
      if ((| mergeHP_CT$wmAdd_Int_select))
        mergeHP_CT$wmAdd_Int_selected = mergeHP_CT$wmAdd_Int_select;
      else
        if (initHP_CT$wmAdd_Int_d[0])
          mergeHP_CT$wmAdd_Int_selected[0] = 1'd1;
        else if (addHP_CT$wmAdd_Int_d[0])
          mergeHP_CT$wmAdd_Int_selected[1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_CT$wmAdd_Int_select <= 2'd0;
    else
      mergeHP_CT$wmAdd_Int_select <= (mergeHP_CT$wmAdd_Int_r ? 2'd0 :
                                      mergeHP_CT$wmAdd_Int_selected);
  always_comb
    if (mergeHP_CT$wmAdd_Int_selected[0])
      mergeHP_CT$wmAdd_Int_d = initHP_CT$wmAdd_Int_d;
    else if (mergeHP_CT$wmAdd_Int_selected[1])
      mergeHP_CT$wmAdd_Int_d = addHP_CT$wmAdd_Int_d;
    else mergeHP_CT$wmAdd_Int_d = {16'd0, 1'd0};
  assign {addHP_CT$wmAdd_Int_r,
          initHP_CT$wmAdd_Int_r} = (mergeHP_CT$wmAdd_Int_r ? mergeHP_CT$wmAdd_Int_selected :
                                    2'd0);
  
  /* buf (Ty Go) : (incrHP_mergeCT$wmAdd_Int,Go) > (incrHP_mergeCT$wmAdd_Int_buf,Go) */
  Go_t incrHP_mergeCT$wmAdd_Int_bufchan_d;
  logic incrHP_mergeCT$wmAdd_Int_bufchan_r;
  assign incrHP_mergeCT$wmAdd_Int_r = ((! incrHP_mergeCT$wmAdd_Int_bufchan_d[0]) || incrHP_mergeCT$wmAdd_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeCT$wmAdd_Int_bufchan_d <= 1'd0;
    else
      if (incrHP_mergeCT$wmAdd_Int_r)
        incrHP_mergeCT$wmAdd_Int_bufchan_d <= incrHP_mergeCT$wmAdd_Int_d;
  Go_t incrHP_mergeCT$wmAdd_Int_bufchan_buf;
  assign incrHP_mergeCT$wmAdd_Int_bufchan_r = (! incrHP_mergeCT$wmAdd_Int_bufchan_buf[0]);
  assign incrHP_mergeCT$wmAdd_Int_buf_d = (incrHP_mergeCT$wmAdd_Int_bufchan_buf[0] ? incrHP_mergeCT$wmAdd_Int_bufchan_buf :
                                           incrHP_mergeCT$wmAdd_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeCT$wmAdd_Int_bufchan_buf <= 1'd0;
    else
      if ((incrHP_mergeCT$wmAdd_Int_buf_r && incrHP_mergeCT$wmAdd_Int_bufchan_buf[0]))
        incrHP_mergeCT$wmAdd_Int_bufchan_buf <= 1'd0;
      else if (((! incrHP_mergeCT$wmAdd_Int_buf_r) && (! incrHP_mergeCT$wmAdd_Int_bufchan_buf[0])))
        incrHP_mergeCT$wmAdd_Int_bufchan_buf <= incrHP_mergeCT$wmAdd_Int_bufchan_d;
  
  /* buf (Ty Word16#) : (mergeHP_CT$wmAdd_Int,Word16#) > (mergeHP_CT$wmAdd_Int_buf,Word16#) */
  \Word16#_t  mergeHP_CT$wmAdd_Int_bufchan_d;
  logic mergeHP_CT$wmAdd_Int_bufchan_r;
  assign mergeHP_CT$wmAdd_Int_r = ((! mergeHP_CT$wmAdd_Int_bufchan_d[0]) || mergeHP_CT$wmAdd_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      mergeHP_CT$wmAdd_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (mergeHP_CT$wmAdd_Int_r)
        mergeHP_CT$wmAdd_Int_bufchan_d <= mergeHP_CT$wmAdd_Int_d;
  \Word16#_t  mergeHP_CT$wmAdd_Int_bufchan_buf;
  assign mergeHP_CT$wmAdd_Int_bufchan_r = (! mergeHP_CT$wmAdd_Int_bufchan_buf[0]);
  assign mergeHP_CT$wmAdd_Int_buf_d = (mergeHP_CT$wmAdd_Int_bufchan_buf[0] ? mergeHP_CT$wmAdd_Int_bufchan_buf :
                                       mergeHP_CT$wmAdd_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      mergeHP_CT$wmAdd_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((mergeHP_CT$wmAdd_Int_buf_r && mergeHP_CT$wmAdd_Int_bufchan_buf[0]))
        mergeHP_CT$wmAdd_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! mergeHP_CT$wmAdd_Int_buf_r) && (! mergeHP_CT$wmAdd_Int_bufchan_buf[0])))
        mergeHP_CT$wmAdd_Int_bufchan_buf <= mergeHP_CT$wmAdd_Int_bufchan_d;
  
  /* fork (Ty Word16#) : (mergeHP_CT$wmAdd_Int_buf,Word16#) > [(forkHP1_CT$wmAdd_Int,Word16#),
                                                          (forkHP1_CT$wmAdd_In2,Word16#),
                                                          (forkHP1_CT$wmAdd_In3,Word16#)] */
  logic [2:0] mergeHP_CT$wmAdd_Int_buf_emitted;
  logic [2:0] mergeHP_CT$wmAdd_Int_buf_done;
  assign forkHP1_CT$wmAdd_Int_d = {mergeHP_CT$wmAdd_Int_buf_d[16:1],
                                   (mergeHP_CT$wmAdd_Int_buf_d[0] && (! mergeHP_CT$wmAdd_Int_buf_emitted[0]))};
  assign forkHP1_CT$wmAdd_In2_d = {mergeHP_CT$wmAdd_Int_buf_d[16:1],
                                   (mergeHP_CT$wmAdd_Int_buf_d[0] && (! mergeHP_CT$wmAdd_Int_buf_emitted[1]))};
  assign forkHP1_CT$wmAdd_In3_d = {mergeHP_CT$wmAdd_Int_buf_d[16:1],
                                   (mergeHP_CT$wmAdd_Int_buf_d[0] && (! mergeHP_CT$wmAdd_Int_buf_emitted[2]))};
  assign mergeHP_CT$wmAdd_Int_buf_done = (mergeHP_CT$wmAdd_Int_buf_emitted | ({forkHP1_CT$wmAdd_In3_d[0],
                                                                               forkHP1_CT$wmAdd_In2_d[0],
                                                                               forkHP1_CT$wmAdd_Int_d[0]} & {forkHP1_CT$wmAdd_In3_r,
                                                                                                             forkHP1_CT$wmAdd_In2_r,
                                                                                                             forkHP1_CT$wmAdd_Int_r}));
  assign mergeHP_CT$wmAdd_Int_buf_r = (& mergeHP_CT$wmAdd_Int_buf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_CT$wmAdd_Int_buf_emitted <= 3'd0;
    else
      mergeHP_CT$wmAdd_Int_buf_emitted <= (mergeHP_CT$wmAdd_Int_buf_r ? 3'd0 :
                                           mergeHP_CT$wmAdd_Int_buf_done);
  
  /* mergectrl (Ty C2,
           Ty MemIn_CT$wmAdd_Int) : [(dconReadIn_CT$wmAdd_Int,MemIn_CT$wmAdd_Int),
                                     (dconWriteIn_CT$wmAdd_Int,MemIn_CT$wmAdd_Int)] > (memMergeChoice_CT$wmAdd_Int,C2) (memMergeIn_CT$wmAdd_Int,MemIn_CT$wmAdd_Int) */
  logic [1:0] dconReadIn_CT$wmAdd_Int_select_d;
  assign dconReadIn_CT$wmAdd_Int_select_d = ((| dconReadIn_CT$wmAdd_Int_select_q) ? dconReadIn_CT$wmAdd_Int_select_q :
                                             (dconReadIn_CT$wmAdd_Int_d[0] ? 2'd1 :
                                              (dconWriteIn_CT$wmAdd_Int_d[0] ? 2'd2 :
                                               2'd0)));
  logic [1:0] dconReadIn_CT$wmAdd_Int_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) dconReadIn_CT$wmAdd_Int_select_q <= 2'd0;
    else
      dconReadIn_CT$wmAdd_Int_select_q <= (dconReadIn_CT$wmAdd_Int_done ? 2'd0 :
                                           dconReadIn_CT$wmAdd_Int_select_d);
  logic [1:0] dconReadIn_CT$wmAdd_Int_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) dconReadIn_CT$wmAdd_Int_emit_q <= 2'd0;
    else
      dconReadIn_CT$wmAdd_Int_emit_q <= (dconReadIn_CT$wmAdd_Int_done ? 2'd0 :
                                         dconReadIn_CT$wmAdd_Int_emit_d);
  logic [1:0] dconReadIn_CT$wmAdd_Int_emit_d;
  assign dconReadIn_CT$wmAdd_Int_emit_d = (dconReadIn_CT$wmAdd_Int_emit_q | ({memMergeChoice_CT$wmAdd_Int_d[0],
                                                                              memMergeIn_CT$wmAdd_Int_d[0]} & {memMergeChoice_CT$wmAdd_Int_r,
                                                                                                               memMergeIn_CT$wmAdd_Int_r}));
  logic dconReadIn_CT$wmAdd_Int_done;
  assign dconReadIn_CT$wmAdd_Int_done = (& dconReadIn_CT$wmAdd_Int_emit_d);
  assign {dconWriteIn_CT$wmAdd_Int_r,
          dconReadIn_CT$wmAdd_Int_r} = (dconReadIn_CT$wmAdd_Int_done ? dconReadIn_CT$wmAdd_Int_select_d :
                                        2'd0);
  assign memMergeIn_CT$wmAdd_Int_d = ((dconReadIn_CT$wmAdd_Int_select_d[0] && (! dconReadIn_CT$wmAdd_Int_emit_q[0])) ? dconReadIn_CT$wmAdd_Int_d :
                                      ((dconReadIn_CT$wmAdd_Int_select_d[1] && (! dconReadIn_CT$wmAdd_Int_emit_q[0])) ? dconWriteIn_CT$wmAdd_Int_d :
                                       {132'd0, 1'd0}));
  assign memMergeChoice_CT$wmAdd_Int_d = ((dconReadIn_CT$wmAdd_Int_select_d[0] && (! dconReadIn_CT$wmAdd_Int_emit_q[1])) ? C1_2_dc(1'd1) :
                                          ((dconReadIn_CT$wmAdd_Int_select_d[1] && (! dconReadIn_CT$wmAdd_Int_emit_q[1])) ? C2_2_dc(1'd1) :
                                           {1'd0, 1'd0}));
  
  /* bram (Ty MemIn_CT$wmAdd_Int,
      Ty MemOut_CT$wmAdd_Int) : (memMergeIn_CT$wmAdd_Int_dbuf,MemIn_CT$wmAdd_Int) > (memOut_CT$wmAdd_Int,MemOut_CT$wmAdd_Int) */
  logic [114:0] memMergeIn_CT$wmAdd_Int_dbuf_mem[65535:0];
  logic [15:0] memMergeIn_CT$wmAdd_Int_dbuf_address;
  logic [114:0] memMergeIn_CT$wmAdd_Int_dbuf_din;
  logic [114:0] memOut_CT$wmAdd_Int_q;
  logic memOut_CT$wmAdd_Int_valid;
  logic memMergeIn_CT$wmAdd_Int_dbuf_we;
  logic memOut_CT$wmAdd_Int_we;
  assign memMergeIn_CT$wmAdd_Int_dbuf_din = memMergeIn_CT$wmAdd_Int_dbuf_d[132:18];
  assign memMergeIn_CT$wmAdd_Int_dbuf_address = memMergeIn_CT$wmAdd_Int_dbuf_d[17:2];
  assign memMergeIn_CT$wmAdd_Int_dbuf_we = (memMergeIn_CT$wmAdd_Int_dbuf_d[1:1] && memMergeIn_CT$wmAdd_Int_dbuf_d[0]);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        memOut_CT$wmAdd_Int_we <= 1'd0;
        memOut_CT$wmAdd_Int_valid <= 1'd0;
      end
    else
      begin
        memOut_CT$wmAdd_Int_we <= memMergeIn_CT$wmAdd_Int_dbuf_we;
        memOut_CT$wmAdd_Int_valid <= memMergeIn_CT$wmAdd_Int_dbuf_d[0];
        if (memMergeIn_CT$wmAdd_Int_dbuf_we)
          begin
            memMergeIn_CT$wmAdd_Int_dbuf_mem[memMergeIn_CT$wmAdd_Int_dbuf_address] <= memMergeIn_CT$wmAdd_Int_dbuf_din;
            memOut_CT$wmAdd_Int_q <= memMergeIn_CT$wmAdd_Int_dbuf_din;
          end
        else
          memOut_CT$wmAdd_Int_q <= memMergeIn_CT$wmAdd_Int_dbuf_mem[memMergeIn_CT$wmAdd_Int_dbuf_address];
      end
  assign memOut_CT$wmAdd_Int_d = {memOut_CT$wmAdd_Int_q,
                                  memOut_CT$wmAdd_Int_we,
                                  memOut_CT$wmAdd_Int_valid};
  assign memMergeIn_CT$wmAdd_Int_dbuf_r = ((! memOut_CT$wmAdd_Int_valid) || memOut_CT$wmAdd_Int_r);
  
  /* demux (Ty C2,
       Ty MemOut_CT$wmAdd_Int) : (memMergeChoice_CT$wmAdd_Int,C2) (memOut_CT$wmAdd_Int_dbuf,MemOut_CT$wmAdd_Int) > [(memReadOut_CT$wmAdd_Int,MemOut_CT$wmAdd_Int),
                                                                                                                    (memWriteOut_CT$wmAdd_Int,MemOut_CT$wmAdd_Int)] */
  logic [1:0] memOut_CT$wmAdd_Int_dbuf_onehotd;
  always_comb
    if ((memMergeChoice_CT$wmAdd_Int_d[0] && memOut_CT$wmAdd_Int_dbuf_d[0]))
      unique case (memMergeChoice_CT$wmAdd_Int_d[1:1])
        1'd0: memOut_CT$wmAdd_Int_dbuf_onehotd = 2'd1;
        1'd1: memOut_CT$wmAdd_Int_dbuf_onehotd = 2'd2;
        default: memOut_CT$wmAdd_Int_dbuf_onehotd = 2'd0;
      endcase
    else memOut_CT$wmAdd_Int_dbuf_onehotd = 2'd0;
  assign memReadOut_CT$wmAdd_Int_d = {memOut_CT$wmAdd_Int_dbuf_d[116:1],
                                      memOut_CT$wmAdd_Int_dbuf_onehotd[0]};
  assign memWriteOut_CT$wmAdd_Int_d = {memOut_CT$wmAdd_Int_dbuf_d[116:1],
                                       memOut_CT$wmAdd_Int_dbuf_onehotd[1]};
  assign memOut_CT$wmAdd_Int_dbuf_r = (| (memOut_CT$wmAdd_Int_dbuf_onehotd & {memWriteOut_CT$wmAdd_Int_r,
                                                                              memReadOut_CT$wmAdd_Int_r}));
  assign memMergeChoice_CT$wmAdd_Int_r = memOut_CT$wmAdd_Int_dbuf_r;
  
  /* dbuf (Ty MemIn_CT$wmAdd_Int) : (memMergeIn_CT$wmAdd_Int_rbuf,MemIn_CT$wmAdd_Int) > (memMergeIn_CT$wmAdd_Int_dbuf,MemIn_CT$wmAdd_Int) */
  assign memMergeIn_CT$wmAdd_Int_rbuf_r = ((! memMergeIn_CT$wmAdd_Int_dbuf_d[0]) || memMergeIn_CT$wmAdd_Int_dbuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      memMergeIn_CT$wmAdd_Int_dbuf_d <= {132'd0, 1'd0};
    else
      if (memMergeIn_CT$wmAdd_Int_rbuf_r)
        memMergeIn_CT$wmAdd_Int_dbuf_d <= memMergeIn_CT$wmAdd_Int_rbuf_d;
  
  /* rbuf (Ty MemIn_CT$wmAdd_Int) : (memMergeIn_CT$wmAdd_Int,MemIn_CT$wmAdd_Int) > (memMergeIn_CT$wmAdd_Int_rbuf,MemIn_CT$wmAdd_Int) */
  MemIn_CT$wmAdd_Int_t memMergeIn_CT$wmAdd_Int_buf;
  assign memMergeIn_CT$wmAdd_Int_r = (! memMergeIn_CT$wmAdd_Int_buf[0]);
  assign memMergeIn_CT$wmAdd_Int_rbuf_d = (memMergeIn_CT$wmAdd_Int_buf[0] ? memMergeIn_CT$wmAdd_Int_buf :
                                           memMergeIn_CT$wmAdd_Int_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memMergeIn_CT$wmAdd_Int_buf <= {132'd0, 1'd0};
    else
      if ((memMergeIn_CT$wmAdd_Int_rbuf_r && memMergeIn_CT$wmAdd_Int_buf[0]))
        memMergeIn_CT$wmAdd_Int_buf <= {132'd0, 1'd0};
      else if (((! memMergeIn_CT$wmAdd_Int_rbuf_r) && (! memMergeIn_CT$wmAdd_Int_buf[0])))
        memMergeIn_CT$wmAdd_Int_buf <= memMergeIn_CT$wmAdd_Int_d;
  
  /* dbuf (Ty MemOut_CT$wmAdd_Int) : (memOut_CT$wmAdd_Int_rbuf,MemOut_CT$wmAdd_Int) > (memOut_CT$wmAdd_Int_dbuf,MemOut_CT$wmAdd_Int) */
  assign memOut_CT$wmAdd_Int_rbuf_r = ((! memOut_CT$wmAdd_Int_dbuf_d[0]) || memOut_CT$wmAdd_Int_dbuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memOut_CT$wmAdd_Int_dbuf_d <= {116'd0, 1'd0};
    else
      if (memOut_CT$wmAdd_Int_rbuf_r)
        memOut_CT$wmAdd_Int_dbuf_d <= memOut_CT$wmAdd_Int_rbuf_d;
  
  /* rbuf (Ty MemOut_CT$wmAdd_Int) : (memOut_CT$wmAdd_Int,MemOut_CT$wmAdd_Int) > (memOut_CT$wmAdd_Int_rbuf,MemOut_CT$wmAdd_Int) */
  MemOut_CT$wmAdd_Int_t memOut_CT$wmAdd_Int_buf;
  assign memOut_CT$wmAdd_Int_r = (! memOut_CT$wmAdd_Int_buf[0]);
  assign memOut_CT$wmAdd_Int_rbuf_d = (memOut_CT$wmAdd_Int_buf[0] ? memOut_CT$wmAdd_Int_buf :
                                       memOut_CT$wmAdd_Int_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memOut_CT$wmAdd_Int_buf <= {116'd0, 1'd0};
    else
      if ((memOut_CT$wmAdd_Int_rbuf_r && memOut_CT$wmAdd_Int_buf[0]))
        memOut_CT$wmAdd_Int_buf <= {116'd0, 1'd0};
      else if (((! memOut_CT$wmAdd_Int_rbuf_r) && (! memOut_CT$wmAdd_Int_buf[0])))
        memOut_CT$wmAdd_Int_buf <= memOut_CT$wmAdd_Int_d;
  
  /* destruct (Ty Pointer_CT$wmAdd_Int,
          Dcon Pointer_CT$wmAdd_Int) : (scfarg_0_1_argbuf,Pointer_CT$wmAdd_Int) > [(destructReadIn_CT$wmAdd_Int,Word16#)] */
  assign destructReadIn_CT$wmAdd_Int_d = {scfarg_0_1_argbuf_d[16:1],
                                          scfarg_0_1_argbuf_d[0]};
  assign scfarg_0_1_argbuf_r = destructReadIn_CT$wmAdd_Int_r;
  
  /* dcon (Ty MemIn_CT$wmAdd_Int,
      Dcon ReadIn_CT$wmAdd_Int) : [(destructReadIn_CT$wmAdd_Int,Word16#)] > (dconReadIn_CT$wmAdd_Int,MemIn_CT$wmAdd_Int) */
  assign dconReadIn_CT$wmAdd_Int_d = ReadIn_CT$wmAdd_Int_dc((& {destructReadIn_CT$wmAdd_Int_d[0]}), destructReadIn_CT$wmAdd_Int_d);
  assign {destructReadIn_CT$wmAdd_Int_r} = {1 {(dconReadIn_CT$wmAdd_Int_r && dconReadIn_CT$wmAdd_Int_d[0])}};
  
  /* destruct (Ty MemOut_CT$wmAdd_Int,
          Dcon ReadOut_CT$wmAdd_Int) : (memReadOut_CT$wmAdd_Int,MemOut_CT$wmAdd_Int) > [(readPointer_CT$wmAdd_Intscfarg_0_1_argbuf,CT$wmAdd_Int)] */
  assign readPointer_CT$wmAdd_Intscfarg_0_1_argbuf_d = {memReadOut_CT$wmAdd_Int_d[116:2],
                                                        memReadOut_CT$wmAdd_Int_d[0]};
  assign memReadOut_CT$wmAdd_Int_r = readPointer_CT$wmAdd_Intscfarg_0_1_argbuf_r;
  
  /* mergectrl (Ty C5,
           Ty CT$wmAdd_Int) : [(lizzieLet0_1_argbuf,CT$wmAdd_Int),
                               (lizzieLet23_1_argbuf,CT$wmAdd_Int),
                               (lizzieLet24_1_argbuf,CT$wmAdd_Int),
                               (lizzieLet25_1_argbuf,CT$wmAdd_Int),
                               (lizzieLet9_1_1_argbuf,CT$wmAdd_Int)] > (writeMerge_choice_CT$wmAdd_Int,C5) (writeMerge_data_CT$wmAdd_Int,CT$wmAdd_Int) */
  logic [4:0] lizzieLet0_1_argbuf_select_d;
  assign lizzieLet0_1_argbuf_select_d = ((| lizzieLet0_1_argbuf_select_q) ? lizzieLet0_1_argbuf_select_q :
                                         (lizzieLet0_1_argbuf_d[0] ? 5'd1 :
                                          (lizzieLet23_1_argbuf_d[0] ? 5'd2 :
                                           (lizzieLet24_1_argbuf_d[0] ? 5'd4 :
                                            (lizzieLet25_1_argbuf_d[0] ? 5'd8 :
                                             (lizzieLet9_1_1_argbuf_d[0] ? 5'd16 :
                                              5'd0))))));
  logic [4:0] lizzieLet0_1_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet0_1_argbuf_select_q <= 5'd0;
    else
      lizzieLet0_1_argbuf_select_q <= (lizzieLet0_1_argbuf_done ? 5'd0 :
                                       lizzieLet0_1_argbuf_select_d);
  logic [1:0] lizzieLet0_1_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet0_1_argbuf_emit_q <= 2'd0;
    else
      lizzieLet0_1_argbuf_emit_q <= (lizzieLet0_1_argbuf_done ? 2'd0 :
                                     lizzieLet0_1_argbuf_emit_d);
  logic [1:0] lizzieLet0_1_argbuf_emit_d;
  assign lizzieLet0_1_argbuf_emit_d = (lizzieLet0_1_argbuf_emit_q | ({writeMerge_choice_CT$wmAdd_Int_d[0],
                                                                      writeMerge_data_CT$wmAdd_Int_d[0]} & {writeMerge_choice_CT$wmAdd_Int_r,
                                                                                                            writeMerge_data_CT$wmAdd_Int_r}));
  logic lizzieLet0_1_argbuf_done;
  assign lizzieLet0_1_argbuf_done = (& lizzieLet0_1_argbuf_emit_d);
  assign {lizzieLet9_1_1_argbuf_r,
          lizzieLet25_1_argbuf_r,
          lizzieLet24_1_argbuf_r,
          lizzieLet23_1_argbuf_r,
          lizzieLet0_1_argbuf_r} = (lizzieLet0_1_argbuf_done ? lizzieLet0_1_argbuf_select_d :
                                    5'd0);
  assign writeMerge_data_CT$wmAdd_Int_d = ((lizzieLet0_1_argbuf_select_d[0] && (! lizzieLet0_1_argbuf_emit_q[0])) ? lizzieLet0_1_argbuf_d :
                                           ((lizzieLet0_1_argbuf_select_d[1] && (! lizzieLet0_1_argbuf_emit_q[0])) ? lizzieLet23_1_argbuf_d :
                                            ((lizzieLet0_1_argbuf_select_d[2] && (! lizzieLet0_1_argbuf_emit_q[0])) ? lizzieLet24_1_argbuf_d :
                                             ((lizzieLet0_1_argbuf_select_d[3] && (! lizzieLet0_1_argbuf_emit_q[0])) ? lizzieLet25_1_argbuf_d :
                                              ((lizzieLet0_1_argbuf_select_d[4] && (! lizzieLet0_1_argbuf_emit_q[0])) ? lizzieLet9_1_1_argbuf_d :
                                               {115'd0, 1'd0})))));
  assign writeMerge_choice_CT$wmAdd_Int_d = ((lizzieLet0_1_argbuf_select_d[0] && (! lizzieLet0_1_argbuf_emit_q[1])) ? C1_5_dc(1'd1) :
                                             ((lizzieLet0_1_argbuf_select_d[1] && (! lizzieLet0_1_argbuf_emit_q[1])) ? C2_5_dc(1'd1) :
                                              ((lizzieLet0_1_argbuf_select_d[2] && (! lizzieLet0_1_argbuf_emit_q[1])) ? C3_5_dc(1'd1) :
                                               ((lizzieLet0_1_argbuf_select_d[3] && (! lizzieLet0_1_argbuf_emit_q[1])) ? C4_5_dc(1'd1) :
                                                ((lizzieLet0_1_argbuf_select_d[4] && (! lizzieLet0_1_argbuf_emit_q[1])) ? C5_5_dc(1'd1) :
                                                 {3'd0, 1'd0})))));
  
  /* demux (Ty C5,
       Ty Pointer_CT$wmAdd_Int) : (writeMerge_choice_CT$wmAdd_Int,C5) (demuxWriteResult_CT$wmAdd_Int,Pointer_CT$wmAdd_Int) > [(writeCT$wmAdd_IntlizzieLet0_1_argbuf,Pointer_CT$wmAdd_Int),
                                                                                                                              (writeCT$wmAdd_IntlizzieLet23_1_argbuf,Pointer_CT$wmAdd_Int),
                                                                                                                              (writeCT$wmAdd_IntlizzieLet24_1_argbuf,Pointer_CT$wmAdd_Int),
                                                                                                                              (writeCT$wmAdd_IntlizzieLet25_1_argbuf,Pointer_CT$wmAdd_Int),
                                                                                                                              (writeCT$wmAdd_IntlizzieLet9_1_1_argbuf,Pointer_CT$wmAdd_Int)] */
  logic [4:0] demuxWriteResult_CT$wmAdd_Int_onehotd;
  always_comb
    if ((writeMerge_choice_CT$wmAdd_Int_d[0] && demuxWriteResult_CT$wmAdd_Int_d[0]))
      unique case (writeMerge_choice_CT$wmAdd_Int_d[3:1])
        3'd0: demuxWriteResult_CT$wmAdd_Int_onehotd = 5'd1;
        3'd1: demuxWriteResult_CT$wmAdd_Int_onehotd = 5'd2;
        3'd2: demuxWriteResult_CT$wmAdd_Int_onehotd = 5'd4;
        3'd3: demuxWriteResult_CT$wmAdd_Int_onehotd = 5'd8;
        3'd4: demuxWriteResult_CT$wmAdd_Int_onehotd = 5'd16;
        default: demuxWriteResult_CT$wmAdd_Int_onehotd = 5'd0;
      endcase
    else demuxWriteResult_CT$wmAdd_Int_onehotd = 5'd0;
  assign writeCT$wmAdd_IntlizzieLet0_1_argbuf_d = {demuxWriteResult_CT$wmAdd_Int_d[16:1],
                                                   demuxWriteResult_CT$wmAdd_Int_onehotd[0]};
  assign writeCT$wmAdd_IntlizzieLet23_1_argbuf_d = {demuxWriteResult_CT$wmAdd_Int_d[16:1],
                                                    demuxWriteResult_CT$wmAdd_Int_onehotd[1]};
  assign writeCT$wmAdd_IntlizzieLet24_1_argbuf_d = {demuxWriteResult_CT$wmAdd_Int_d[16:1],
                                                    demuxWriteResult_CT$wmAdd_Int_onehotd[2]};
  assign writeCT$wmAdd_IntlizzieLet25_1_argbuf_d = {demuxWriteResult_CT$wmAdd_Int_d[16:1],
                                                    demuxWriteResult_CT$wmAdd_Int_onehotd[3]};
  assign writeCT$wmAdd_IntlizzieLet9_1_1_argbuf_d = {demuxWriteResult_CT$wmAdd_Int_d[16:1],
                                                     demuxWriteResult_CT$wmAdd_Int_onehotd[4]};
  assign demuxWriteResult_CT$wmAdd_Int_r = (| (demuxWriteResult_CT$wmAdd_Int_onehotd & {writeCT$wmAdd_IntlizzieLet9_1_1_argbuf_r,
                                                                                        writeCT$wmAdd_IntlizzieLet25_1_argbuf_r,
                                                                                        writeCT$wmAdd_IntlizzieLet24_1_argbuf_r,
                                                                                        writeCT$wmAdd_IntlizzieLet23_1_argbuf_r,
                                                                                        writeCT$wmAdd_IntlizzieLet0_1_argbuf_r}));
  assign writeMerge_choice_CT$wmAdd_Int_r = demuxWriteResult_CT$wmAdd_Int_r;
  
  /* dcon (Ty MemIn_CT$wmAdd_Int,
      Dcon WriteIn_CT$wmAdd_Int) : [(forkHP1_CT$wmAdd_In2,Word16#),
                                    (writeMerge_data_CT$wmAdd_Int,CT$wmAdd_Int)] > (dconWriteIn_CT$wmAdd_Int,MemIn_CT$wmAdd_Int) */
  assign dconWriteIn_CT$wmAdd_Int_d = WriteIn_CT$wmAdd_Int_dc((& {forkHP1_CT$wmAdd_In2_d[0],
                                                                  writeMerge_data_CT$wmAdd_Int_d[0]}), forkHP1_CT$wmAdd_In2_d, writeMerge_data_CT$wmAdd_Int_d);
  assign {forkHP1_CT$wmAdd_In2_r,
          writeMerge_data_CT$wmAdd_Int_r} = {2 {(dconWriteIn_CT$wmAdd_Int_r && dconWriteIn_CT$wmAdd_Int_d[0])}};
  
  /* dcon (Ty Pointer_CT$wmAdd_Int,
      Dcon Pointer_CT$wmAdd_Int) : [(forkHP1_CT$wmAdd_In3,Word16#)] > (dconPtr_CT$wmAdd_Int,Pointer_CT$wmAdd_Int) */
  assign dconPtr_CT$wmAdd_Int_d = Pointer_CT$wmAdd_Int_dc((& {forkHP1_CT$wmAdd_In3_d[0]}), forkHP1_CT$wmAdd_In3_d);
  assign {forkHP1_CT$wmAdd_In3_r} = {1 {(dconPtr_CT$wmAdd_Int_r && dconPtr_CT$wmAdd_Int_d[0])}};
  
  /* demux (Ty MemOut_CT$wmAdd_Int,
       Ty Pointer_CT$wmAdd_Int) : (memWriteOut_CT$wmAdd_Int,MemOut_CT$wmAdd_Int) (dconPtr_CT$wmAdd_Int,Pointer_CT$wmAdd_Int) > [(_78,Pointer_CT$wmAdd_Int),
                                                                                                                                (demuxWriteResult_CT$wmAdd_Int,Pointer_CT$wmAdd_Int)] */
  logic [1:0] dconPtr_CT$wmAdd_Int_onehotd;
  always_comb
    if ((memWriteOut_CT$wmAdd_Int_d[0] && dconPtr_CT$wmAdd_Int_d[0]))
      unique case (memWriteOut_CT$wmAdd_Int_d[1:1])
        1'd0: dconPtr_CT$wmAdd_Int_onehotd = 2'd1;
        1'd1: dconPtr_CT$wmAdd_Int_onehotd = 2'd2;
        default: dconPtr_CT$wmAdd_Int_onehotd = 2'd0;
      endcase
    else dconPtr_CT$wmAdd_Int_onehotd = 2'd0;
  assign _78_d = {dconPtr_CT$wmAdd_Int_d[16:1],
                  dconPtr_CT$wmAdd_Int_onehotd[0]};
  assign demuxWriteResult_CT$wmAdd_Int_d = {dconPtr_CT$wmAdd_Int_d[16:1],
                                            dconPtr_CT$wmAdd_Int_onehotd[1]};
  assign dconPtr_CT$wmAdd_Int_r = (| (dconPtr_CT$wmAdd_Int_onehotd & {demuxWriteResult_CT$wmAdd_Int_r,
                                                                      _78_r}));
  assign memWriteOut_CT$wmAdd_Int_r = dconPtr_CT$wmAdd_Int_r;
  
  /* const (Ty Word16#,
       Lit 0) : (go_1_dummy_write_QTree_Int,Go) > (initHP_QTree_Int,Word16#) */
  assign initHP_QTree_Int_d = {16'd0,
                               go_1_dummy_write_QTree_Int_d[0]};
  assign go_1_dummy_write_QTree_Int_r = initHP_QTree_Int_r;
  
  /* const (Ty Word16#,
       Lit 1) : (incrHP_QTree_Int1,Go) > (incrHP_QTree_Int,Word16#) */
  assign incrHP_QTree_Int_d = {16'd1, incrHP_QTree_Int1_d[0]};
  assign incrHP_QTree_Int1_r = incrHP_QTree_Int_r;
  
  /* merge (Ty Go) : [(go_2_dummy_write_QTree_Int,Go),
                 (incrHP_QTree_Int2,Go)] > (incrHP_mergeQTree_Int,Go) */
  logic [1:0] incrHP_mergeQTree_Int_selected;
  logic [1:0] incrHP_mergeQTree_Int_select;
  always_comb
    begin
      incrHP_mergeQTree_Int_selected = 2'd0;
      if ((| incrHP_mergeQTree_Int_select))
        incrHP_mergeQTree_Int_selected = incrHP_mergeQTree_Int_select;
      else
        if (go_2_dummy_write_QTree_Int_d[0])
          incrHP_mergeQTree_Int_selected[0] = 1'd1;
        else if (incrHP_QTree_Int2_d[0])
          incrHP_mergeQTree_Int_selected[1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeQTree_Int_select <= 2'd0;
    else
      incrHP_mergeQTree_Int_select <= (incrHP_mergeQTree_Int_r ? 2'd0 :
                                       incrHP_mergeQTree_Int_selected);
  always_comb
    if (incrHP_mergeQTree_Int_selected[0])
      incrHP_mergeQTree_Int_d = go_2_dummy_write_QTree_Int_d;
    else if (incrHP_mergeQTree_Int_selected[1])
      incrHP_mergeQTree_Int_d = incrHP_QTree_Int2_d;
    else incrHP_mergeQTree_Int_d = 1'd0;
  assign {incrHP_QTree_Int2_r,
          go_2_dummy_write_QTree_Int_r} = (incrHP_mergeQTree_Int_r ? incrHP_mergeQTree_Int_selected :
                                           2'd0);
  
  /* fork (Ty Go) : (incrHP_mergeQTree_Int_buf,Go) > [(incrHP_QTree_Int1,Go),
                                                 (incrHP_QTree_Int2,Go)] */
  logic [1:0] incrHP_mergeQTree_Int_buf_emitted;
  logic [1:0] incrHP_mergeQTree_Int_buf_done;
  assign incrHP_QTree_Int1_d = (incrHP_mergeQTree_Int_buf_d[0] && (! incrHP_mergeQTree_Int_buf_emitted[0]));
  assign incrHP_QTree_Int2_d = (incrHP_mergeQTree_Int_buf_d[0] && (! incrHP_mergeQTree_Int_buf_emitted[1]));
  assign incrHP_mergeQTree_Int_buf_done = (incrHP_mergeQTree_Int_buf_emitted | ({incrHP_QTree_Int2_d[0],
                                                                                 incrHP_QTree_Int1_d[0]} & {incrHP_QTree_Int2_r,
                                                                                                            incrHP_QTree_Int1_r}));
  assign incrHP_mergeQTree_Int_buf_r = (& incrHP_mergeQTree_Int_buf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeQTree_Int_buf_emitted <= 2'd0;
    else
      incrHP_mergeQTree_Int_buf_emitted <= (incrHP_mergeQTree_Int_buf_r ? 2'd0 :
                                            incrHP_mergeQTree_Int_buf_done);
  
  /* op_add (Ty Word16#) : (incrHP_QTree_Int,Word16#) (forkHP1_QTree_Int,Word16#) > (addHP_QTree_Int,Word16#) */
  assign addHP_QTree_Int_d = {(incrHP_QTree_Int_d[16:1] + forkHP1_QTree_Int_d[16:1]),
                              (incrHP_QTree_Int_d[0] && forkHP1_QTree_Int_d[0])};
  assign {incrHP_QTree_Int_r,
          forkHP1_QTree_Int_r} = {2 {(addHP_QTree_Int_r && addHP_QTree_Int_d[0])}};
  
  /* merge (Ty Word16#) : [(initHP_QTree_Int,Word16#),
                      (addHP_QTree_Int,Word16#)] > (mergeHP_QTree_Int,Word16#) */
  logic [1:0] mergeHP_QTree_Int_selected;
  logic [1:0] mergeHP_QTree_Int_select;
  always_comb
    begin
      mergeHP_QTree_Int_selected = 2'd0;
      if ((| mergeHP_QTree_Int_select))
        mergeHP_QTree_Int_selected = mergeHP_QTree_Int_select;
      else
        if (initHP_QTree_Int_d[0]) mergeHP_QTree_Int_selected[0] = 1'd1;
        else if (addHP_QTree_Int_d[0])
          mergeHP_QTree_Int_selected[1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_QTree_Int_select <= 2'd0;
    else
      mergeHP_QTree_Int_select <= (mergeHP_QTree_Int_r ? 2'd0 :
                                   mergeHP_QTree_Int_selected);
  always_comb
    if (mergeHP_QTree_Int_selected[0])
      mergeHP_QTree_Int_d = initHP_QTree_Int_d;
    else if (mergeHP_QTree_Int_selected[1])
      mergeHP_QTree_Int_d = addHP_QTree_Int_d;
    else mergeHP_QTree_Int_d = {16'd0, 1'd0};
  assign {addHP_QTree_Int_r,
          initHP_QTree_Int_r} = (mergeHP_QTree_Int_r ? mergeHP_QTree_Int_selected :
                                 2'd0);
  
  /* buf (Ty Go) : (incrHP_mergeQTree_Int,Go) > (incrHP_mergeQTree_Int_buf,Go) */
  Go_t incrHP_mergeQTree_Int_bufchan_d;
  logic incrHP_mergeQTree_Int_bufchan_r;
  assign incrHP_mergeQTree_Int_r = ((! incrHP_mergeQTree_Int_bufchan_d[0]) || incrHP_mergeQTree_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeQTree_Int_bufchan_d <= 1'd0;
    else
      if (incrHP_mergeQTree_Int_r)
        incrHP_mergeQTree_Int_bufchan_d <= incrHP_mergeQTree_Int_d;
  Go_t incrHP_mergeQTree_Int_bufchan_buf;
  assign incrHP_mergeQTree_Int_bufchan_r = (! incrHP_mergeQTree_Int_bufchan_buf[0]);
  assign incrHP_mergeQTree_Int_buf_d = (incrHP_mergeQTree_Int_bufchan_buf[0] ? incrHP_mergeQTree_Int_bufchan_buf :
                                        incrHP_mergeQTree_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeQTree_Int_bufchan_buf <= 1'd0;
    else
      if ((incrHP_mergeQTree_Int_buf_r && incrHP_mergeQTree_Int_bufchan_buf[0]))
        incrHP_mergeQTree_Int_bufchan_buf <= 1'd0;
      else if (((! incrHP_mergeQTree_Int_buf_r) && (! incrHP_mergeQTree_Int_bufchan_buf[0])))
        incrHP_mergeQTree_Int_bufchan_buf <= incrHP_mergeQTree_Int_bufchan_d;
  
  /* buf (Ty Word16#) : (mergeHP_QTree_Int,Word16#) > (mergeHP_QTree_Int_buf,Word16#) */
  \Word16#_t  mergeHP_QTree_Int_bufchan_d;
  logic mergeHP_QTree_Int_bufchan_r;
  assign mergeHP_QTree_Int_r = ((! mergeHP_QTree_Int_bufchan_d[0]) || mergeHP_QTree_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_QTree_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (mergeHP_QTree_Int_r)
        mergeHP_QTree_Int_bufchan_d <= mergeHP_QTree_Int_d;
  \Word16#_t  mergeHP_QTree_Int_bufchan_buf;
  assign mergeHP_QTree_Int_bufchan_r = (! mergeHP_QTree_Int_bufchan_buf[0]);
  assign mergeHP_QTree_Int_buf_d = (mergeHP_QTree_Int_bufchan_buf[0] ? mergeHP_QTree_Int_bufchan_buf :
                                    mergeHP_QTree_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      mergeHP_QTree_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((mergeHP_QTree_Int_buf_r && mergeHP_QTree_Int_bufchan_buf[0]))
        mergeHP_QTree_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! mergeHP_QTree_Int_buf_r) && (! mergeHP_QTree_Int_bufchan_buf[0])))
        mergeHP_QTree_Int_bufchan_buf <= mergeHP_QTree_Int_bufchan_d;
  
  /* sink (Ty Word16#) : (forkHP1_QTree_Int_snk,Word16#) > */
  assign {forkHP1_QTree_Int_snk_r,
          forkHP1_QTree_Int_snk_dout} = {forkHP1_QTree_Int_snk_rout,
                                         forkHP1_QTree_Int_snk_d};
  
  /* source (Ty Go) : > (\QTree_Int_src,Go) */
  
  /* fork (Ty Go) : (\QTree_Int_src,Go) > [(go_1_dummy_write_QTree_Int,Go),
                                      (go_2_dummy_write_QTree_Int,Go)] */
  logic [1:0] \\QTree_Int_src_emitted ;
  logic [1:0] \\QTree_Int_src_done ;
  assign go_1_dummy_write_QTree_Int_d = (\\QTree_Int_src_d [0] && (! \\QTree_Int_src_emitted [0]));
  assign go_2_dummy_write_QTree_Int_d = (\\QTree_Int_src_d [0] && (! \\QTree_Int_src_emitted [1]));
  assign \\QTree_Int_src_done  = (\\QTree_Int_src_emitted  | ({go_2_dummy_write_QTree_Int_d[0],
                                                               go_1_dummy_write_QTree_Int_d[0]} & {go_2_dummy_write_QTree_Int_r,
                                                                                                   go_1_dummy_write_QTree_Int_r}));
  assign \\QTree_Int_src_r  = (& \\QTree_Int_src_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \\QTree_Int_src_emitted  <= 2'd0;
    else
      \\QTree_Int_src_emitted  <= (\\QTree_Int_src_r  ? 2'd0 :
                                   \\QTree_Int_src_done );
  
  /* source (Ty QTree_Int) : > (dummy_write_QTree_Int,QTree_Int) */
  
  /* sink (Ty Pointer_QTree_Int) : (dummy_write_QTree_Int_sink,Pointer_QTree_Int) > */
  assign {dummy_write_QTree_Int_sink_r,
          dummy_write_QTree_Int_sink_dout} = {dummy_write_QTree_Int_sink_rout,
                                              dummy_write_QTree_Int_sink_d};
  
  /* fork (Ty Word16#) : (mergeHP_QTree_Int_buf,Word16#) > [(forkHP1_QTree_Int,Word16#),
                                                       (forkHP1_QTree_Int_snk,Word16#),
                                                       (forkHP1_QTree_In3,Word16#),
                                                       (forkHP1_QTree_In4,Word16#)] */
  logic [3:0] mergeHP_QTree_Int_buf_emitted;
  logic [3:0] mergeHP_QTree_Int_buf_done;
  assign forkHP1_QTree_Int_d = {mergeHP_QTree_Int_buf_d[16:1],
                                (mergeHP_QTree_Int_buf_d[0] && (! mergeHP_QTree_Int_buf_emitted[0]))};
  assign forkHP1_QTree_Int_snk_d = {mergeHP_QTree_Int_buf_d[16:1],
                                    (mergeHP_QTree_Int_buf_d[0] && (! mergeHP_QTree_Int_buf_emitted[1]))};
  assign forkHP1_QTree_In3_d = {mergeHP_QTree_Int_buf_d[16:1],
                                (mergeHP_QTree_Int_buf_d[0] && (! mergeHP_QTree_Int_buf_emitted[2]))};
  assign forkHP1_QTree_In4_d = {mergeHP_QTree_Int_buf_d[16:1],
                                (mergeHP_QTree_Int_buf_d[0] && (! mergeHP_QTree_Int_buf_emitted[3]))};
  assign mergeHP_QTree_Int_buf_done = (mergeHP_QTree_Int_buf_emitted | ({forkHP1_QTree_In4_d[0],
                                                                         forkHP1_QTree_In3_d[0],
                                                                         forkHP1_QTree_Int_snk_d[0],
                                                                         forkHP1_QTree_Int_d[0]} & {forkHP1_QTree_In4_r,
                                                                                                    forkHP1_QTree_In3_r,
                                                                                                    forkHP1_QTree_Int_snk_r,
                                                                                                    forkHP1_QTree_Int_r}));
  assign mergeHP_QTree_Int_buf_r = (& mergeHP_QTree_Int_buf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_QTree_Int_buf_emitted <= 4'd0;
    else
      mergeHP_QTree_Int_buf_emitted <= (mergeHP_QTree_Int_buf_r ? 4'd0 :
                                        mergeHP_QTree_Int_buf_done);
  
  /* mergectrl (Ty C2,
           Ty MemIn_QTree_Int) : [(dconReadIn_QTree_Int,MemIn_QTree_Int),
                                  (dconWriteIn_QTree_Int,MemIn_QTree_Int)] > (memMergeChoice_QTree_Int,C2) (memMergeIn_QTree_Int,MemIn_QTree_Int) */
  logic [1:0] dconReadIn_QTree_Int_select_d;
  assign dconReadIn_QTree_Int_select_d = ((| dconReadIn_QTree_Int_select_q) ? dconReadIn_QTree_Int_select_q :
                                          (dconReadIn_QTree_Int_d[0] ? 2'd1 :
                                           (dconWriteIn_QTree_Int_d[0] ? 2'd2 :
                                            2'd0)));
  logic [1:0] dconReadIn_QTree_Int_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) dconReadIn_QTree_Int_select_q <= 2'd0;
    else
      dconReadIn_QTree_Int_select_q <= (dconReadIn_QTree_Int_done ? 2'd0 :
                                        dconReadIn_QTree_Int_select_d);
  logic [1:0] dconReadIn_QTree_Int_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) dconReadIn_QTree_Int_emit_q <= 2'd0;
    else
      dconReadIn_QTree_Int_emit_q <= (dconReadIn_QTree_Int_done ? 2'd0 :
                                      dconReadIn_QTree_Int_emit_d);
  logic [1:0] dconReadIn_QTree_Int_emit_d;
  assign dconReadIn_QTree_Int_emit_d = (dconReadIn_QTree_Int_emit_q | ({memMergeChoice_QTree_Int_d[0],
                                                                        memMergeIn_QTree_Int_d[0]} & {memMergeChoice_QTree_Int_r,
                                                                                                      memMergeIn_QTree_Int_r}));
  logic dconReadIn_QTree_Int_done;
  assign dconReadIn_QTree_Int_done = (& dconReadIn_QTree_Int_emit_d);
  assign {dconWriteIn_QTree_Int_r,
          dconReadIn_QTree_Int_r} = (dconReadIn_QTree_Int_done ? dconReadIn_QTree_Int_select_d :
                                     2'd0);
  assign memMergeIn_QTree_Int_d = ((dconReadIn_QTree_Int_select_d[0] && (! dconReadIn_QTree_Int_emit_q[0])) ? dconReadIn_QTree_Int_d :
                                   ((dconReadIn_QTree_Int_select_d[1] && (! dconReadIn_QTree_Int_emit_q[0])) ? dconWriteIn_QTree_Int_d :
                                    {83'd0, 1'd0}));
  assign memMergeChoice_QTree_Int_d = ((dconReadIn_QTree_Int_select_d[0] && (! dconReadIn_QTree_Int_emit_q[1])) ? C1_2_dc(1'd1) :
                                       ((dconReadIn_QTree_Int_select_d[1] && (! dconReadIn_QTree_Int_emit_q[1])) ? C2_2_dc(1'd1) :
                                        {1'd0, 1'd0}));
  
  /* bram (Ty MemIn_QTree_Int,
      Ty MemOut_QTree_Int) : (memMergeIn_QTree_Int_dbuf,MemIn_QTree_Int) > (memOut_QTree_Int,MemOut_QTree_Int) */
  logic [65:0] memMergeIn_QTree_Int_dbuf_mem[65535:0];
  logic [15:0] memMergeIn_QTree_Int_dbuf_address;
  logic [65:0] memMergeIn_QTree_Int_dbuf_din;
  logic [65:0] memOut_QTree_Int_q;
  logic memOut_QTree_Int_valid;
  logic memMergeIn_QTree_Int_dbuf_we;
  logic memOut_QTree_Int_we;
  assign memMergeIn_QTree_Int_dbuf_din = memMergeIn_QTree_Int_dbuf_d[83:18];
  assign memMergeIn_QTree_Int_dbuf_address = memMergeIn_QTree_Int_dbuf_d[17:2];
  assign memMergeIn_QTree_Int_dbuf_we = (memMergeIn_QTree_Int_dbuf_d[1:1] && memMergeIn_QTree_Int_dbuf_d[0]);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        memOut_QTree_Int_we <= 1'd0;
        memOut_QTree_Int_valid <= 1'd0;
      end
    else
      begin
        memOut_QTree_Int_we <= memMergeIn_QTree_Int_dbuf_we;
        memOut_QTree_Int_valid <= memMergeIn_QTree_Int_dbuf_d[0];
        if (memMergeIn_QTree_Int_dbuf_we)
          begin
            memMergeIn_QTree_Int_dbuf_mem[memMergeIn_QTree_Int_dbuf_address] <= memMergeIn_QTree_Int_dbuf_din;
            memOut_QTree_Int_q <= memMergeIn_QTree_Int_dbuf_din;
          end
        else
          memOut_QTree_Int_q <= memMergeIn_QTree_Int_dbuf_mem[memMergeIn_QTree_Int_dbuf_address];
      end
  assign memOut_QTree_Int_d = {memOut_QTree_Int_q,
                               memOut_QTree_Int_we,
                               memOut_QTree_Int_valid};
  assign memMergeIn_QTree_Int_dbuf_r = ((! memOut_QTree_Int_valid) || memOut_QTree_Int_r);
  
  /* demux (Ty C2,
       Ty MemOut_QTree_Int) : (memMergeChoice_QTree_Int,C2) (memOut_QTree_Int_dbuf,MemOut_QTree_Int) > [(memReadOut_QTree_Int,MemOut_QTree_Int),
                                                                                                        (memWriteOut_QTree_Int,MemOut_QTree_Int)] */
  logic [1:0] memOut_QTree_Int_dbuf_onehotd;
  always_comb
    if ((memMergeChoice_QTree_Int_d[0] && memOut_QTree_Int_dbuf_d[0]))
      unique case (memMergeChoice_QTree_Int_d[1:1])
        1'd0: memOut_QTree_Int_dbuf_onehotd = 2'd1;
        1'd1: memOut_QTree_Int_dbuf_onehotd = 2'd2;
        default: memOut_QTree_Int_dbuf_onehotd = 2'd0;
      endcase
    else memOut_QTree_Int_dbuf_onehotd = 2'd0;
  assign memReadOut_QTree_Int_d = {memOut_QTree_Int_dbuf_d[67:1],
                                   memOut_QTree_Int_dbuf_onehotd[0]};
  assign memWriteOut_QTree_Int_d = {memOut_QTree_Int_dbuf_d[67:1],
                                    memOut_QTree_Int_dbuf_onehotd[1]};
  assign memOut_QTree_Int_dbuf_r = (| (memOut_QTree_Int_dbuf_onehotd & {memWriteOut_QTree_Int_r,
                                                                        memReadOut_QTree_Int_r}));
  assign memMergeChoice_QTree_Int_r = memOut_QTree_Int_dbuf_r;
  
  /* dbuf (Ty MemIn_QTree_Int) : (memMergeIn_QTree_Int_rbuf,MemIn_QTree_Int) > (memMergeIn_QTree_Int_dbuf,MemIn_QTree_Int) */
  assign memMergeIn_QTree_Int_rbuf_r = ((! memMergeIn_QTree_Int_dbuf_d[0]) || memMergeIn_QTree_Int_dbuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memMergeIn_QTree_Int_dbuf_d <= {83'd0, 1'd0};
    else
      if (memMergeIn_QTree_Int_rbuf_r)
        memMergeIn_QTree_Int_dbuf_d <= memMergeIn_QTree_Int_rbuf_d;
  
  /* rbuf (Ty MemIn_QTree_Int) : (memMergeIn_QTree_Int,MemIn_QTree_Int) > (memMergeIn_QTree_Int_rbuf,MemIn_QTree_Int) */
  MemIn_QTree_Int_t memMergeIn_QTree_Int_buf;
  assign memMergeIn_QTree_Int_r = (! memMergeIn_QTree_Int_buf[0]);
  assign memMergeIn_QTree_Int_rbuf_d = (memMergeIn_QTree_Int_buf[0] ? memMergeIn_QTree_Int_buf :
                                        memMergeIn_QTree_Int_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memMergeIn_QTree_Int_buf <= {83'd0, 1'd0};
    else
      if ((memMergeIn_QTree_Int_rbuf_r && memMergeIn_QTree_Int_buf[0]))
        memMergeIn_QTree_Int_buf <= {83'd0, 1'd0};
      else if (((! memMergeIn_QTree_Int_rbuf_r) && (! memMergeIn_QTree_Int_buf[0])))
        memMergeIn_QTree_Int_buf <= memMergeIn_QTree_Int_d;
  
  /* dbuf (Ty MemOut_QTree_Int) : (memOut_QTree_Int_rbuf,MemOut_QTree_Int) > (memOut_QTree_Int_dbuf,MemOut_QTree_Int) */
  assign memOut_QTree_Int_rbuf_r = ((! memOut_QTree_Int_dbuf_d[0]) || memOut_QTree_Int_dbuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memOut_QTree_Int_dbuf_d <= {67'd0, 1'd0};
    else
      if (memOut_QTree_Int_rbuf_r)
        memOut_QTree_Int_dbuf_d <= memOut_QTree_Int_rbuf_d;
  
  /* rbuf (Ty MemOut_QTree_Int) : (memOut_QTree_Int,MemOut_QTree_Int) > (memOut_QTree_Int_rbuf,MemOut_QTree_Int) */
  MemOut_QTree_Int_t memOut_QTree_Int_buf;
  assign memOut_QTree_Int_r = (! memOut_QTree_Int_buf[0]);
  assign memOut_QTree_Int_rbuf_d = (memOut_QTree_Int_buf[0] ? memOut_QTree_Int_buf :
                                    memOut_QTree_Int_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memOut_QTree_Int_buf <= {67'd0, 1'd0};
    else
      if ((memOut_QTree_Int_rbuf_r && memOut_QTree_Int_buf[0]))
        memOut_QTree_Int_buf <= {67'd0, 1'd0};
      else if (((! memOut_QTree_Int_rbuf_r) && (! memOut_QTree_Int_buf[0])))
        memOut_QTree_Int_buf <= memOut_QTree_Int_d;
  
  /* mergectrl (Ty C4,
           Ty Pointer_QTree_Int) : [(ma8q_1_argbuf,Pointer_QTree_Int),
                                    (w1sif_1_1_argbuf,Pointer_QTree_Int),
                                    (w2sig_1_1_argbuf,Pointer_QTree_Int),
                                    (wsij_1_1_argbuf,Pointer_QTree_Int)] > (readMerge_choice_QTree_Int,C4) (readMerge_data_QTree_Int,Pointer_QTree_Int) */
  logic [3:0] ma8q_1_argbuf_select_d;
  assign ma8q_1_argbuf_select_d = ((| ma8q_1_argbuf_select_q) ? ma8q_1_argbuf_select_q :
                                   (ma8q_1_argbuf_d[0] ? 4'd1 :
                                    (w1sif_1_1_argbuf_d[0] ? 4'd2 :
                                     (w2sig_1_1_argbuf_d[0] ? 4'd4 :
                                      (wsij_1_1_argbuf_d[0] ? 4'd8 :
                                       4'd0)))));
  logic [3:0] ma8q_1_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) ma8q_1_argbuf_select_q <= 4'd0;
    else
      ma8q_1_argbuf_select_q <= (ma8q_1_argbuf_done ? 4'd0 :
                                 ma8q_1_argbuf_select_d);
  logic [1:0] ma8q_1_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) ma8q_1_argbuf_emit_q <= 2'd0;
    else
      ma8q_1_argbuf_emit_q <= (ma8q_1_argbuf_done ? 2'd0 :
                               ma8q_1_argbuf_emit_d);
  logic [1:0] ma8q_1_argbuf_emit_d;
  assign ma8q_1_argbuf_emit_d = (ma8q_1_argbuf_emit_q | ({readMerge_choice_QTree_Int_d[0],
                                                          readMerge_data_QTree_Int_d[0]} & {readMerge_choice_QTree_Int_r,
                                                                                            readMerge_data_QTree_Int_r}));
  logic ma8q_1_argbuf_done;
  assign ma8q_1_argbuf_done = (& ma8q_1_argbuf_emit_d);
  assign {wsij_1_1_argbuf_r,
          w2sig_1_1_argbuf_r,
          w1sif_1_1_argbuf_r,
          ma8q_1_argbuf_r} = (ma8q_1_argbuf_done ? ma8q_1_argbuf_select_d :
                              4'd0);
  assign readMerge_data_QTree_Int_d = ((ma8q_1_argbuf_select_d[0] && (! ma8q_1_argbuf_emit_q[0])) ? ma8q_1_argbuf_d :
                                       ((ma8q_1_argbuf_select_d[1] && (! ma8q_1_argbuf_emit_q[0])) ? w1sif_1_1_argbuf_d :
                                        ((ma8q_1_argbuf_select_d[2] && (! ma8q_1_argbuf_emit_q[0])) ? w2sig_1_1_argbuf_d :
                                         ((ma8q_1_argbuf_select_d[3] && (! ma8q_1_argbuf_emit_q[0])) ? wsij_1_1_argbuf_d :
                                          {16'd0, 1'd0}))));
  assign readMerge_choice_QTree_Int_d = ((ma8q_1_argbuf_select_d[0] && (! ma8q_1_argbuf_emit_q[1])) ? C1_4_dc(1'd1) :
                                         ((ma8q_1_argbuf_select_d[1] && (! ma8q_1_argbuf_emit_q[1])) ? C2_4_dc(1'd1) :
                                          ((ma8q_1_argbuf_select_d[2] && (! ma8q_1_argbuf_emit_q[1])) ? C3_4_dc(1'd1) :
                                           ((ma8q_1_argbuf_select_d[3] && (! ma8q_1_argbuf_emit_q[1])) ? C4_4_dc(1'd1) :
                                            {2'd0, 1'd0}))));
  
  /* demux (Ty C4,
       Ty QTree_Int) : (readMerge_choice_QTree_Int,C4) (destructReadOut_QTree_Int,QTree_Int) > [(readPointer_QTree_Intma8q_1_argbuf,QTree_Int),
                                                                                                (readPointer_QTree_Intw1sif_1_1_argbuf,QTree_Int),
                                                                                                (readPointer_QTree_Intw2sig_1_1_argbuf,QTree_Int),
                                                                                                (readPointer_QTree_Intwsij_1_1_argbuf,QTree_Int)] */
  logic [3:0] destructReadOut_QTree_Int_onehotd;
  always_comb
    if ((readMerge_choice_QTree_Int_d[0] && destructReadOut_QTree_Int_d[0]))
      unique case (readMerge_choice_QTree_Int_d[2:1])
        2'd0: destructReadOut_QTree_Int_onehotd = 4'd1;
        2'd1: destructReadOut_QTree_Int_onehotd = 4'd2;
        2'd2: destructReadOut_QTree_Int_onehotd = 4'd4;
        2'd3: destructReadOut_QTree_Int_onehotd = 4'd8;
        default: destructReadOut_QTree_Int_onehotd = 4'd0;
      endcase
    else destructReadOut_QTree_Int_onehotd = 4'd0;
  assign readPointer_QTree_Intma8q_1_argbuf_d = {destructReadOut_QTree_Int_d[66:1],
                                                 destructReadOut_QTree_Int_onehotd[0]};
  assign readPointer_QTree_Intw1sif_1_1_argbuf_d = {destructReadOut_QTree_Int_d[66:1],
                                                    destructReadOut_QTree_Int_onehotd[1]};
  assign readPointer_QTree_Intw2sig_1_1_argbuf_d = {destructReadOut_QTree_Int_d[66:1],
                                                    destructReadOut_QTree_Int_onehotd[2]};
  assign readPointer_QTree_Intwsij_1_1_argbuf_d = {destructReadOut_QTree_Int_d[66:1],
                                                   destructReadOut_QTree_Int_onehotd[3]};
  assign destructReadOut_QTree_Int_r = (| (destructReadOut_QTree_Int_onehotd & {readPointer_QTree_Intwsij_1_1_argbuf_r,
                                                                                readPointer_QTree_Intw2sig_1_1_argbuf_r,
                                                                                readPointer_QTree_Intw1sif_1_1_argbuf_r,
                                                                                readPointer_QTree_Intma8q_1_argbuf_r}));
  assign readMerge_choice_QTree_Int_r = destructReadOut_QTree_Int_r;
  
  /* destruct (Ty Pointer_QTree_Int,
          Dcon Pointer_QTree_Int) : (readMerge_data_QTree_Int,Pointer_QTree_Int) > [(destructReadIn_QTree_Int,Word16#)] */
  assign destructReadIn_QTree_Int_d = {readMerge_data_QTree_Int_d[16:1],
                                       readMerge_data_QTree_Int_d[0]};
  assign readMerge_data_QTree_Int_r = destructReadIn_QTree_Int_r;
  
  /* dcon (Ty MemIn_QTree_Int,
      Dcon ReadIn_QTree_Int) : [(destructReadIn_QTree_Int,Word16#)] > (dconReadIn_QTree_Int,MemIn_QTree_Int) */
  assign dconReadIn_QTree_Int_d = ReadIn_QTree_Int_dc((& {destructReadIn_QTree_Int_d[0]}), destructReadIn_QTree_Int_d);
  assign {destructReadIn_QTree_Int_r} = {1 {(dconReadIn_QTree_Int_r && dconReadIn_QTree_Int_d[0])}};
  
  /* destruct (Ty MemOut_QTree_Int,
          Dcon ReadOut_QTree_Int) : (memReadOut_QTree_Int,MemOut_QTree_Int) > [(destructReadOut_QTree_Int,QTree_Int)] */
  assign destructReadOut_QTree_Int_d = {memReadOut_QTree_Int_d[67:2],
                                        memReadOut_QTree_Int_d[0]};
  assign memReadOut_QTree_Int_r = destructReadOut_QTree_Int_r;
  
  /* mergectrl (Ty C13,
           Ty QTree_Int) : [(lizzieLet10_1_1_argbuf,QTree_Int),
                            (lizzieLet11_1_1_argbuf,QTree_Int),
                            (lizzieLet15_1_argbuf,QTree_Int),
                            (lizzieLet17_1_argbuf,QTree_Int),
                            (lizzieLet18_1_argbuf,QTree_Int),
                            (lizzieLet20_1_argbuf,QTree_Int),
                            (lizzieLet26_1_argbuf,QTree_Int),
                            (lizzieLet35_1_argbuf,QTree_Int),
                            (lizzieLet4_1_argbuf,QTree_Int),
                            (lizzieLet5_1_argbuf,QTree_Int),
                            (lizzieLet6_1_argbuf,QTree_Int),
                            (lizzieLet8_1_1_argbuf,QTree_Int),
                            (dummy_write_QTree_Int,QTree_Int)] > (writeMerge_choice_QTree_Int,C13) (writeMerge_data_QTree_Int,QTree_Int) */
  logic [12:0] lizzieLet10_1_1_argbuf_select_d;
  assign lizzieLet10_1_1_argbuf_select_d = ((| lizzieLet10_1_1_argbuf_select_q) ? lizzieLet10_1_1_argbuf_select_q :
                                            (lizzieLet10_1_1_argbuf_d[0] ? 13'd1 :
                                             (lizzieLet11_1_1_argbuf_d[0] ? 13'd2 :
                                              (lizzieLet15_1_argbuf_d[0] ? 13'd4 :
                                               (lizzieLet17_1_argbuf_d[0] ? 13'd8 :
                                                (lizzieLet18_1_argbuf_d[0] ? 13'd16 :
                                                 (lizzieLet20_1_argbuf_d[0] ? 13'd32 :
                                                  (lizzieLet26_1_argbuf_d[0] ? 13'd64 :
                                                   (lizzieLet35_1_argbuf_d[0] ? 13'd128 :
                                                    (lizzieLet4_1_argbuf_d[0] ? 13'd256 :
                                                     (lizzieLet5_1_argbuf_d[0] ? 13'd512 :
                                                      (lizzieLet6_1_argbuf_d[0] ? 13'd1024 :
                                                       (lizzieLet8_1_1_argbuf_d[0] ? 13'd2048 :
                                                        (dummy_write_QTree_Int_d[0] ? 13'd4096 :
                                                         13'd0))))))))))))));
  logic [12:0] lizzieLet10_1_1_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet10_1_1_argbuf_select_q <= 13'd0;
    else
      lizzieLet10_1_1_argbuf_select_q <= (lizzieLet10_1_1_argbuf_done ? 13'd0 :
                                          lizzieLet10_1_1_argbuf_select_d);
  logic [1:0] lizzieLet10_1_1_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet10_1_1_argbuf_emit_q <= 2'd0;
    else
      lizzieLet10_1_1_argbuf_emit_q <= (lizzieLet10_1_1_argbuf_done ? 2'd0 :
                                        lizzieLet10_1_1_argbuf_emit_d);
  logic [1:0] lizzieLet10_1_1_argbuf_emit_d;
  assign lizzieLet10_1_1_argbuf_emit_d = (lizzieLet10_1_1_argbuf_emit_q | ({writeMerge_choice_QTree_Int_d[0],
                                                                            writeMerge_data_QTree_Int_d[0]} & {writeMerge_choice_QTree_Int_r,
                                                                                                               writeMerge_data_QTree_Int_r}));
  logic lizzieLet10_1_1_argbuf_done;
  assign lizzieLet10_1_1_argbuf_done = (& lizzieLet10_1_1_argbuf_emit_d);
  assign {dummy_write_QTree_Int_r,
          lizzieLet8_1_1_argbuf_r,
          lizzieLet6_1_argbuf_r,
          lizzieLet5_1_argbuf_r,
          lizzieLet4_1_argbuf_r,
          lizzieLet35_1_argbuf_r,
          lizzieLet26_1_argbuf_r,
          lizzieLet20_1_argbuf_r,
          lizzieLet18_1_argbuf_r,
          lizzieLet17_1_argbuf_r,
          lizzieLet15_1_argbuf_r,
          lizzieLet11_1_1_argbuf_r,
          lizzieLet10_1_1_argbuf_r} = (lizzieLet10_1_1_argbuf_done ? lizzieLet10_1_1_argbuf_select_d :
                                       13'd0);
  assign writeMerge_data_QTree_Int_d = ((lizzieLet10_1_1_argbuf_select_d[0] && (! lizzieLet10_1_1_argbuf_emit_q[0])) ? lizzieLet10_1_1_argbuf_d :
                                        ((lizzieLet10_1_1_argbuf_select_d[1] && (! lizzieLet10_1_1_argbuf_emit_q[0])) ? lizzieLet11_1_1_argbuf_d :
                                         ((lizzieLet10_1_1_argbuf_select_d[2] && (! lizzieLet10_1_1_argbuf_emit_q[0])) ? lizzieLet15_1_argbuf_d :
                                          ((lizzieLet10_1_1_argbuf_select_d[3] && (! lizzieLet10_1_1_argbuf_emit_q[0])) ? lizzieLet17_1_argbuf_d :
                                           ((lizzieLet10_1_1_argbuf_select_d[4] && (! lizzieLet10_1_1_argbuf_emit_q[0])) ? lizzieLet18_1_argbuf_d :
                                            ((lizzieLet10_1_1_argbuf_select_d[5] && (! lizzieLet10_1_1_argbuf_emit_q[0])) ? lizzieLet20_1_argbuf_d :
                                             ((lizzieLet10_1_1_argbuf_select_d[6] && (! lizzieLet10_1_1_argbuf_emit_q[0])) ? lizzieLet26_1_argbuf_d :
                                              ((lizzieLet10_1_1_argbuf_select_d[7] && (! lizzieLet10_1_1_argbuf_emit_q[0])) ? lizzieLet35_1_argbuf_d :
                                               ((lizzieLet10_1_1_argbuf_select_d[8] && (! lizzieLet10_1_1_argbuf_emit_q[0])) ? lizzieLet4_1_argbuf_d :
                                                ((lizzieLet10_1_1_argbuf_select_d[9] && (! lizzieLet10_1_1_argbuf_emit_q[0])) ? lizzieLet5_1_argbuf_d :
                                                 ((lizzieLet10_1_1_argbuf_select_d[10] && (! lizzieLet10_1_1_argbuf_emit_q[0])) ? lizzieLet6_1_argbuf_d :
                                                  ((lizzieLet10_1_1_argbuf_select_d[11] && (! lizzieLet10_1_1_argbuf_emit_q[0])) ? lizzieLet8_1_1_argbuf_d :
                                                   ((lizzieLet10_1_1_argbuf_select_d[12] && (! lizzieLet10_1_1_argbuf_emit_q[0])) ? dummy_write_QTree_Int_d :
                                                    {66'd0, 1'd0})))))))))))));
  assign writeMerge_choice_QTree_Int_d = ((lizzieLet10_1_1_argbuf_select_d[0] && (! lizzieLet10_1_1_argbuf_emit_q[1])) ? C1_13_dc(1'd1) :
                                          ((lizzieLet10_1_1_argbuf_select_d[1] && (! lizzieLet10_1_1_argbuf_emit_q[1])) ? C2_13_dc(1'd1) :
                                           ((lizzieLet10_1_1_argbuf_select_d[2] && (! lizzieLet10_1_1_argbuf_emit_q[1])) ? C3_13_dc(1'd1) :
                                            ((lizzieLet10_1_1_argbuf_select_d[3] && (! lizzieLet10_1_1_argbuf_emit_q[1])) ? C4_13_dc(1'd1) :
                                             ((lizzieLet10_1_1_argbuf_select_d[4] && (! lizzieLet10_1_1_argbuf_emit_q[1])) ? C5_13_dc(1'd1) :
                                              ((lizzieLet10_1_1_argbuf_select_d[5] && (! lizzieLet10_1_1_argbuf_emit_q[1])) ? C6_13_dc(1'd1) :
                                               ((lizzieLet10_1_1_argbuf_select_d[6] && (! lizzieLet10_1_1_argbuf_emit_q[1])) ? C7_13_dc(1'd1) :
                                                ((lizzieLet10_1_1_argbuf_select_d[7] && (! lizzieLet10_1_1_argbuf_emit_q[1])) ? C8_13_dc(1'd1) :
                                                 ((lizzieLet10_1_1_argbuf_select_d[8] && (! lizzieLet10_1_1_argbuf_emit_q[1])) ? C9_13_dc(1'd1) :
                                                  ((lizzieLet10_1_1_argbuf_select_d[9] && (! lizzieLet10_1_1_argbuf_emit_q[1])) ? C10_13_dc(1'd1) :
                                                   ((lizzieLet10_1_1_argbuf_select_d[10] && (! lizzieLet10_1_1_argbuf_emit_q[1])) ? C11_13_dc(1'd1) :
                                                    ((lizzieLet10_1_1_argbuf_select_d[11] && (! lizzieLet10_1_1_argbuf_emit_q[1])) ? C12_13_dc(1'd1) :
                                                     ((lizzieLet10_1_1_argbuf_select_d[12] && (! lizzieLet10_1_1_argbuf_emit_q[1])) ? C13_13_dc(1'd1) :
                                                      {4'd0, 1'd0})))))))))))));
  
  /* demux (Ty C13,
       Ty Pointer_QTree_Int) : (writeMerge_choice_QTree_Int,C13) (demuxWriteResult_QTree_Int,Pointer_QTree_Int) > [(writeQTree_IntlizzieLet10_1_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet11_1_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet15_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet17_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet18_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet20_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet26_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet35_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet4_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet5_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet6_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet8_1_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (dummy_write_QTree_Int_sink,Pointer_QTree_Int)] */
  logic [12:0] demuxWriteResult_QTree_Int_onehotd;
  always_comb
    if ((writeMerge_choice_QTree_Int_d[0] && demuxWriteResult_QTree_Int_d[0]))
      unique case (writeMerge_choice_QTree_Int_d[4:1])
        4'd0: demuxWriteResult_QTree_Int_onehotd = 13'd1;
        4'd1: demuxWriteResult_QTree_Int_onehotd = 13'd2;
        4'd2: demuxWriteResult_QTree_Int_onehotd = 13'd4;
        4'd3: demuxWriteResult_QTree_Int_onehotd = 13'd8;
        4'd4: demuxWriteResult_QTree_Int_onehotd = 13'd16;
        4'd5: demuxWriteResult_QTree_Int_onehotd = 13'd32;
        4'd6: demuxWriteResult_QTree_Int_onehotd = 13'd64;
        4'd7: demuxWriteResult_QTree_Int_onehotd = 13'd128;
        4'd8: demuxWriteResult_QTree_Int_onehotd = 13'd256;
        4'd9: demuxWriteResult_QTree_Int_onehotd = 13'd512;
        4'd10: demuxWriteResult_QTree_Int_onehotd = 13'd1024;
        4'd11: demuxWriteResult_QTree_Int_onehotd = 13'd2048;
        4'd12: demuxWriteResult_QTree_Int_onehotd = 13'd4096;
        default: demuxWriteResult_QTree_Int_onehotd = 13'd0;
      endcase
    else demuxWriteResult_QTree_Int_onehotd = 13'd0;
  assign writeQTree_IntlizzieLet10_1_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                   demuxWriteResult_QTree_Int_onehotd[0]};
  assign writeQTree_IntlizzieLet11_1_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                   demuxWriteResult_QTree_Int_onehotd[1]};
  assign writeQTree_IntlizzieLet15_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                 demuxWriteResult_QTree_Int_onehotd[2]};
  assign writeQTree_IntlizzieLet17_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                 demuxWriteResult_QTree_Int_onehotd[3]};
  assign writeQTree_IntlizzieLet18_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                 demuxWriteResult_QTree_Int_onehotd[4]};
  assign writeQTree_IntlizzieLet20_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                 demuxWriteResult_QTree_Int_onehotd[5]};
  assign writeQTree_IntlizzieLet26_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                 demuxWriteResult_QTree_Int_onehotd[6]};
  assign writeQTree_IntlizzieLet35_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                 demuxWriteResult_QTree_Int_onehotd[7]};
  assign writeQTree_IntlizzieLet4_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                demuxWriteResult_QTree_Int_onehotd[8]};
  assign writeQTree_IntlizzieLet5_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                demuxWriteResult_QTree_Int_onehotd[9]};
  assign writeQTree_IntlizzieLet6_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                demuxWriteResult_QTree_Int_onehotd[10]};
  assign writeQTree_IntlizzieLet8_1_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                  demuxWriteResult_QTree_Int_onehotd[11]};
  assign dummy_write_QTree_Int_sink_d = {demuxWriteResult_QTree_Int_d[16:1],
                                         demuxWriteResult_QTree_Int_onehotd[12]};
  assign demuxWriteResult_QTree_Int_r = (| (demuxWriteResult_QTree_Int_onehotd & {dummy_write_QTree_Int_sink_r,
                                                                                  writeQTree_IntlizzieLet8_1_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet6_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet5_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet4_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet35_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet26_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet20_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet18_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet17_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet15_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet11_1_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet10_1_1_argbuf_r}));
  assign writeMerge_choice_QTree_Int_r = demuxWriteResult_QTree_Int_r;
  
  /* dcon (Ty MemIn_QTree_Int,
      Dcon WriteIn_QTree_Int) : [(forkHP1_QTree_In3,Word16#),
                                 (writeMerge_data_QTree_Int,QTree_Int)] > (dconWriteIn_QTree_Int,MemIn_QTree_Int) */
  assign dconWriteIn_QTree_Int_d = WriteIn_QTree_Int_dc((& {forkHP1_QTree_In3_d[0],
                                                            writeMerge_data_QTree_Int_d[0]}), forkHP1_QTree_In3_d, writeMerge_data_QTree_Int_d);
  assign {forkHP1_QTree_In3_r,
          writeMerge_data_QTree_Int_r} = {2 {(dconWriteIn_QTree_Int_r && dconWriteIn_QTree_Int_d[0])}};
  
  /* dcon (Ty Pointer_QTree_Int,
      Dcon Pointer_QTree_Int) : [(forkHP1_QTree_In4,Word16#)] > (dconPtr_QTree_Int,Pointer_QTree_Int) */
  assign dconPtr_QTree_Int_d = Pointer_QTree_Int_dc((& {forkHP1_QTree_In4_d[0]}), forkHP1_QTree_In4_d);
  assign {forkHP1_QTree_In4_r} = {1 {(dconPtr_QTree_Int_r && dconPtr_QTree_Int_d[0])}};
  
  /* demux (Ty MemOut_QTree_Int,
       Ty Pointer_QTree_Int) : (memWriteOut_QTree_Int,MemOut_QTree_Int) (dconPtr_QTree_Int,Pointer_QTree_Int) > [(_77,Pointer_QTree_Int),
                                                                                                                 (demuxWriteResult_QTree_Int,Pointer_QTree_Int)] */
  logic [1:0] dconPtr_QTree_Int_onehotd;
  always_comb
    if ((memWriteOut_QTree_Int_d[0] && dconPtr_QTree_Int_d[0]))
      unique case (memWriteOut_QTree_Int_d[1:1])
        1'd0: dconPtr_QTree_Int_onehotd = 2'd1;
        1'd1: dconPtr_QTree_Int_onehotd = 2'd2;
        default: dconPtr_QTree_Int_onehotd = 2'd0;
      endcase
    else dconPtr_QTree_Int_onehotd = 2'd0;
  assign _77_d = {dconPtr_QTree_Int_d[16:1],
                  dconPtr_QTree_Int_onehotd[0]};
  assign demuxWriteResult_QTree_Int_d = {dconPtr_QTree_Int_d[16:1],
                                         dconPtr_QTree_Int_onehotd[1]};
  assign dconPtr_QTree_Int_r = (| (dconPtr_QTree_Int_onehotd & {demuxWriteResult_QTree_Int_r,
                                                                _77_r}));
  assign memWriteOut_QTree_Int_r = dconPtr_QTree_Int_r;
  
  /* const (Ty Word16#,
       Lit 0) : (go__7,Go) > (initHP_CT$wnnz_Int,Word16#) */
  assign initHP_CT$wnnz_Int_d = {16'd0, go__7_d[0]};
  assign go__7_r = initHP_CT$wnnz_Int_r;
  
  /* const (Ty Word16#,
       Lit 1) : (incrHP_CT$wnnz_Int1,Go) > (incrHP_CT$wnnz_Int,Word16#) */
  assign incrHP_CT$wnnz_Int_d = {16'd1, incrHP_CT$wnnz_Int1_d[0]};
  assign incrHP_CT$wnnz_Int1_r = incrHP_CT$wnnz_Int_r;
  
  /* merge (Ty Go) : [(go__8,Go),
                 (incrHP_CT$wnnz_Int2,Go)] > (incrHP_mergeCT$wnnz_Int,Go) */
  logic [1:0] incrHP_mergeCT$wnnz_Int_selected;
  logic [1:0] incrHP_mergeCT$wnnz_Int_select;
  always_comb
    begin
      incrHP_mergeCT$wnnz_Int_selected = 2'd0;
      if ((| incrHP_mergeCT$wnnz_Int_select))
        incrHP_mergeCT$wnnz_Int_selected = incrHP_mergeCT$wnnz_Int_select;
      else
        if (go__8_d[0]) incrHP_mergeCT$wnnz_Int_selected[0] = 1'd1;
        else if (incrHP_CT$wnnz_Int2_d[0])
          incrHP_mergeCT$wnnz_Int_selected[1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeCT$wnnz_Int_select <= 2'd0;
    else
      incrHP_mergeCT$wnnz_Int_select <= (incrHP_mergeCT$wnnz_Int_r ? 2'd0 :
                                         incrHP_mergeCT$wnnz_Int_selected);
  always_comb
    if (incrHP_mergeCT$wnnz_Int_selected[0])
      incrHP_mergeCT$wnnz_Int_d = go__8_d;
    else if (incrHP_mergeCT$wnnz_Int_selected[1])
      incrHP_mergeCT$wnnz_Int_d = incrHP_CT$wnnz_Int2_d;
    else incrHP_mergeCT$wnnz_Int_d = 1'd0;
  assign {incrHP_CT$wnnz_Int2_r,
          go__8_r} = (incrHP_mergeCT$wnnz_Int_r ? incrHP_mergeCT$wnnz_Int_selected :
                      2'd0);
  
  /* fork (Ty Go) : (incrHP_mergeCT$wnnz_Int_buf,Go) > [(incrHP_CT$wnnz_Int1,Go),
                                                   (incrHP_CT$wnnz_Int2,Go)] */
  logic [1:0] incrHP_mergeCT$wnnz_Int_buf_emitted;
  logic [1:0] incrHP_mergeCT$wnnz_Int_buf_done;
  assign incrHP_CT$wnnz_Int1_d = (incrHP_mergeCT$wnnz_Int_buf_d[0] && (! incrHP_mergeCT$wnnz_Int_buf_emitted[0]));
  assign incrHP_CT$wnnz_Int2_d = (incrHP_mergeCT$wnnz_Int_buf_d[0] && (! incrHP_mergeCT$wnnz_Int_buf_emitted[1]));
  assign incrHP_mergeCT$wnnz_Int_buf_done = (incrHP_mergeCT$wnnz_Int_buf_emitted | ({incrHP_CT$wnnz_Int2_d[0],
                                                                                     incrHP_CT$wnnz_Int1_d[0]} & {incrHP_CT$wnnz_Int2_r,
                                                                                                                  incrHP_CT$wnnz_Int1_r}));
  assign incrHP_mergeCT$wnnz_Int_buf_r = (& incrHP_mergeCT$wnnz_Int_buf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeCT$wnnz_Int_buf_emitted <= 2'd0;
    else
      incrHP_mergeCT$wnnz_Int_buf_emitted <= (incrHP_mergeCT$wnnz_Int_buf_r ? 2'd0 :
                                              incrHP_mergeCT$wnnz_Int_buf_done);
  
  /* op_add (Ty Word16#) : (incrHP_CT$wnnz_Int,Word16#) (forkHP1_CT$wnnz_Int,Word16#) > (addHP_CT$wnnz_Int,Word16#) */
  assign addHP_CT$wnnz_Int_d = {(incrHP_CT$wnnz_Int_d[16:1] + forkHP1_CT$wnnz_Int_d[16:1]),
                                (incrHP_CT$wnnz_Int_d[0] && forkHP1_CT$wnnz_Int_d[0])};
  assign {incrHP_CT$wnnz_Int_r,
          forkHP1_CT$wnnz_Int_r} = {2 {(addHP_CT$wnnz_Int_r && addHP_CT$wnnz_Int_d[0])}};
  
  /* merge (Ty Word16#) : [(initHP_CT$wnnz_Int,Word16#),
                      (addHP_CT$wnnz_Int,Word16#)] > (mergeHP_CT$wnnz_Int,Word16#) */
  logic [1:0] mergeHP_CT$wnnz_Int_selected;
  logic [1:0] mergeHP_CT$wnnz_Int_select;
  always_comb
    begin
      mergeHP_CT$wnnz_Int_selected = 2'd0;
      if ((| mergeHP_CT$wnnz_Int_select))
        mergeHP_CT$wnnz_Int_selected = mergeHP_CT$wnnz_Int_select;
      else
        if (initHP_CT$wnnz_Int_d[0])
          mergeHP_CT$wnnz_Int_selected[0] = 1'd1;
        else if (addHP_CT$wnnz_Int_d[0])
          mergeHP_CT$wnnz_Int_selected[1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_CT$wnnz_Int_select <= 2'd0;
    else
      mergeHP_CT$wnnz_Int_select <= (mergeHP_CT$wnnz_Int_r ? 2'd0 :
                                     mergeHP_CT$wnnz_Int_selected);
  always_comb
    if (mergeHP_CT$wnnz_Int_selected[0])
      mergeHP_CT$wnnz_Int_d = initHP_CT$wnnz_Int_d;
    else if (mergeHP_CT$wnnz_Int_selected[1])
      mergeHP_CT$wnnz_Int_d = addHP_CT$wnnz_Int_d;
    else mergeHP_CT$wnnz_Int_d = {16'd0, 1'd0};
  assign {addHP_CT$wnnz_Int_r,
          initHP_CT$wnnz_Int_r} = (mergeHP_CT$wnnz_Int_r ? mergeHP_CT$wnnz_Int_selected :
                                   2'd0);
  
  /* buf (Ty Go) : (incrHP_mergeCT$wnnz_Int,Go) > (incrHP_mergeCT$wnnz_Int_buf,Go) */
  Go_t incrHP_mergeCT$wnnz_Int_bufchan_d;
  logic incrHP_mergeCT$wnnz_Int_bufchan_r;
  assign incrHP_mergeCT$wnnz_Int_r = ((! incrHP_mergeCT$wnnz_Int_bufchan_d[0]) || incrHP_mergeCT$wnnz_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeCT$wnnz_Int_bufchan_d <= 1'd0;
    else
      if (incrHP_mergeCT$wnnz_Int_r)
        incrHP_mergeCT$wnnz_Int_bufchan_d <= incrHP_mergeCT$wnnz_Int_d;
  Go_t incrHP_mergeCT$wnnz_Int_bufchan_buf;
  assign incrHP_mergeCT$wnnz_Int_bufchan_r = (! incrHP_mergeCT$wnnz_Int_bufchan_buf[0]);
  assign incrHP_mergeCT$wnnz_Int_buf_d = (incrHP_mergeCT$wnnz_Int_bufchan_buf[0] ? incrHP_mergeCT$wnnz_Int_bufchan_buf :
                                          incrHP_mergeCT$wnnz_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeCT$wnnz_Int_bufchan_buf <= 1'd0;
    else
      if ((incrHP_mergeCT$wnnz_Int_buf_r && incrHP_mergeCT$wnnz_Int_bufchan_buf[0]))
        incrHP_mergeCT$wnnz_Int_bufchan_buf <= 1'd0;
      else if (((! incrHP_mergeCT$wnnz_Int_buf_r) && (! incrHP_mergeCT$wnnz_Int_bufchan_buf[0])))
        incrHP_mergeCT$wnnz_Int_bufchan_buf <= incrHP_mergeCT$wnnz_Int_bufchan_d;
  
  /* buf (Ty Word16#) : (mergeHP_CT$wnnz_Int,Word16#) > (mergeHP_CT$wnnz_Int_buf,Word16#) */
  \Word16#_t  mergeHP_CT$wnnz_Int_bufchan_d;
  logic mergeHP_CT$wnnz_Int_bufchan_r;
  assign mergeHP_CT$wnnz_Int_r = ((! mergeHP_CT$wnnz_Int_bufchan_d[0]) || mergeHP_CT$wnnz_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      mergeHP_CT$wnnz_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (mergeHP_CT$wnnz_Int_r)
        mergeHP_CT$wnnz_Int_bufchan_d <= mergeHP_CT$wnnz_Int_d;
  \Word16#_t  mergeHP_CT$wnnz_Int_bufchan_buf;
  assign mergeHP_CT$wnnz_Int_bufchan_r = (! mergeHP_CT$wnnz_Int_bufchan_buf[0]);
  assign mergeHP_CT$wnnz_Int_buf_d = (mergeHP_CT$wnnz_Int_bufchan_buf[0] ? mergeHP_CT$wnnz_Int_bufchan_buf :
                                      mergeHP_CT$wnnz_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      mergeHP_CT$wnnz_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((mergeHP_CT$wnnz_Int_buf_r && mergeHP_CT$wnnz_Int_bufchan_buf[0]))
        mergeHP_CT$wnnz_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! mergeHP_CT$wnnz_Int_buf_r) && (! mergeHP_CT$wnnz_Int_bufchan_buf[0])))
        mergeHP_CT$wnnz_Int_bufchan_buf <= mergeHP_CT$wnnz_Int_bufchan_d;
  
  /* fork (Ty Word16#) : (mergeHP_CT$wnnz_Int_buf,Word16#) > [(forkHP1_CT$wnnz_Int,Word16#),
                                                         (forkHP1_CT$wnnz_In2,Word16#),
                                                         (forkHP1_CT$wnnz_In3,Word16#)] */
  logic [2:0] mergeHP_CT$wnnz_Int_buf_emitted;
  logic [2:0] mergeHP_CT$wnnz_Int_buf_done;
  assign forkHP1_CT$wnnz_Int_d = {mergeHP_CT$wnnz_Int_buf_d[16:1],
                                  (mergeHP_CT$wnnz_Int_buf_d[0] && (! mergeHP_CT$wnnz_Int_buf_emitted[0]))};
  assign forkHP1_CT$wnnz_In2_d = {mergeHP_CT$wnnz_Int_buf_d[16:1],
                                  (mergeHP_CT$wnnz_Int_buf_d[0] && (! mergeHP_CT$wnnz_Int_buf_emitted[1]))};
  assign forkHP1_CT$wnnz_In3_d = {mergeHP_CT$wnnz_Int_buf_d[16:1],
                                  (mergeHP_CT$wnnz_Int_buf_d[0] && (! mergeHP_CT$wnnz_Int_buf_emitted[2]))};
  assign mergeHP_CT$wnnz_Int_buf_done = (mergeHP_CT$wnnz_Int_buf_emitted | ({forkHP1_CT$wnnz_In3_d[0],
                                                                             forkHP1_CT$wnnz_In2_d[0],
                                                                             forkHP1_CT$wnnz_Int_d[0]} & {forkHP1_CT$wnnz_In3_r,
                                                                                                          forkHP1_CT$wnnz_In2_r,
                                                                                                          forkHP1_CT$wnnz_Int_r}));
  assign mergeHP_CT$wnnz_Int_buf_r = (& mergeHP_CT$wnnz_Int_buf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_CT$wnnz_Int_buf_emitted <= 3'd0;
    else
      mergeHP_CT$wnnz_Int_buf_emitted <= (mergeHP_CT$wnnz_Int_buf_r ? 3'd0 :
                                          mergeHP_CT$wnnz_Int_buf_done);
  
  /* mergectrl (Ty C2,
           Ty MemIn_CT$wnnz_Int) : [(dconReadIn_CT$wnnz_Int,MemIn_CT$wnnz_Int),
                                    (dconWriteIn_CT$wnnz_Int,MemIn_CT$wnnz_Int)] > (memMergeChoice_CT$wnnz_Int,C2) (memMergeIn_CT$wnnz_Int,MemIn_CT$wnnz_Int) */
  logic [1:0] dconReadIn_CT$wnnz_Int_select_d;
  assign dconReadIn_CT$wnnz_Int_select_d = ((| dconReadIn_CT$wnnz_Int_select_q) ? dconReadIn_CT$wnnz_Int_select_q :
                                            (dconReadIn_CT$wnnz_Int_d[0] ? 2'd1 :
                                             (dconWriteIn_CT$wnnz_Int_d[0] ? 2'd2 :
                                              2'd0)));
  logic [1:0] dconReadIn_CT$wnnz_Int_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) dconReadIn_CT$wnnz_Int_select_q <= 2'd0;
    else
      dconReadIn_CT$wnnz_Int_select_q <= (dconReadIn_CT$wnnz_Int_done ? 2'd0 :
                                          dconReadIn_CT$wnnz_Int_select_d);
  logic [1:0] dconReadIn_CT$wnnz_Int_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) dconReadIn_CT$wnnz_Int_emit_q <= 2'd0;
    else
      dconReadIn_CT$wnnz_Int_emit_q <= (dconReadIn_CT$wnnz_Int_done ? 2'd0 :
                                        dconReadIn_CT$wnnz_Int_emit_d);
  logic [1:0] dconReadIn_CT$wnnz_Int_emit_d;
  assign dconReadIn_CT$wnnz_Int_emit_d = (dconReadIn_CT$wnnz_Int_emit_q | ({memMergeChoice_CT$wnnz_Int_d[0],
                                                                            memMergeIn_CT$wnnz_Int_d[0]} & {memMergeChoice_CT$wnnz_Int_r,
                                                                                                            memMergeIn_CT$wnnz_Int_r}));
  logic dconReadIn_CT$wnnz_Int_done;
  assign dconReadIn_CT$wnnz_Int_done = (& dconReadIn_CT$wnnz_Int_emit_d);
  assign {dconWriteIn_CT$wnnz_Int_r,
          dconReadIn_CT$wnnz_Int_r} = (dconReadIn_CT$wnnz_Int_done ? dconReadIn_CT$wnnz_Int_select_d :
                                       2'd0);
  assign memMergeIn_CT$wnnz_Int_d = ((dconReadIn_CT$wnnz_Int_select_d[0] && (! dconReadIn_CT$wnnz_Int_emit_q[0])) ? dconReadIn_CT$wnnz_Int_d :
                                     ((dconReadIn_CT$wnnz_Int_select_d[1] && (! dconReadIn_CT$wnnz_Int_emit_q[0])) ? dconWriteIn_CT$wnnz_Int_d :
                                      {132'd0, 1'd0}));
  assign memMergeChoice_CT$wnnz_Int_d = ((dconReadIn_CT$wnnz_Int_select_d[0] && (! dconReadIn_CT$wnnz_Int_emit_q[1])) ? C1_2_dc(1'd1) :
                                         ((dconReadIn_CT$wnnz_Int_select_d[1] && (! dconReadIn_CT$wnnz_Int_emit_q[1])) ? C2_2_dc(1'd1) :
                                          {1'd0, 1'd0}));
  
  /* bram (Ty MemIn_CT$wnnz_Int,
      Ty MemOut_CT$wnnz_Int) : (memMergeIn_CT$wnnz_Int_dbuf,MemIn_CT$wnnz_Int) > (memOut_CT$wnnz_Int,MemOut_CT$wnnz_Int) */
  logic [114:0] memMergeIn_CT$wnnz_Int_dbuf_mem[65535:0];
  logic [15:0] memMergeIn_CT$wnnz_Int_dbuf_address;
  logic [114:0] memMergeIn_CT$wnnz_Int_dbuf_din;
  logic [114:0] memOut_CT$wnnz_Int_q;
  logic memOut_CT$wnnz_Int_valid;
  logic memMergeIn_CT$wnnz_Int_dbuf_we;
  logic memOut_CT$wnnz_Int_we;
  assign memMergeIn_CT$wnnz_Int_dbuf_din = memMergeIn_CT$wnnz_Int_dbuf_d[132:18];
  assign memMergeIn_CT$wnnz_Int_dbuf_address = memMergeIn_CT$wnnz_Int_dbuf_d[17:2];
  assign memMergeIn_CT$wnnz_Int_dbuf_we = (memMergeIn_CT$wnnz_Int_dbuf_d[1:1] && memMergeIn_CT$wnnz_Int_dbuf_d[0]);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        memOut_CT$wnnz_Int_we <= 1'd0;
        memOut_CT$wnnz_Int_valid <= 1'd0;
      end
    else
      begin
        memOut_CT$wnnz_Int_we <= memMergeIn_CT$wnnz_Int_dbuf_we;
        memOut_CT$wnnz_Int_valid <= memMergeIn_CT$wnnz_Int_dbuf_d[0];
        if (memMergeIn_CT$wnnz_Int_dbuf_we)
          begin
            memMergeIn_CT$wnnz_Int_dbuf_mem[memMergeIn_CT$wnnz_Int_dbuf_address] <= memMergeIn_CT$wnnz_Int_dbuf_din;
            memOut_CT$wnnz_Int_q <= memMergeIn_CT$wnnz_Int_dbuf_din;
          end
        else
          memOut_CT$wnnz_Int_q <= memMergeIn_CT$wnnz_Int_dbuf_mem[memMergeIn_CT$wnnz_Int_dbuf_address];
      end
  assign memOut_CT$wnnz_Int_d = {memOut_CT$wnnz_Int_q,
                                 memOut_CT$wnnz_Int_we,
                                 memOut_CT$wnnz_Int_valid};
  assign memMergeIn_CT$wnnz_Int_dbuf_r = ((! memOut_CT$wnnz_Int_valid) || memOut_CT$wnnz_Int_r);
  
  /* demux (Ty C2,
       Ty MemOut_CT$wnnz_Int) : (memMergeChoice_CT$wnnz_Int,C2) (memOut_CT$wnnz_Int_dbuf,MemOut_CT$wnnz_Int) > [(memReadOut_CT$wnnz_Int,MemOut_CT$wnnz_Int),
                                                                                                                (memWriteOut_CT$wnnz_Int,MemOut_CT$wnnz_Int)] */
  logic [1:0] memOut_CT$wnnz_Int_dbuf_onehotd;
  always_comb
    if ((memMergeChoice_CT$wnnz_Int_d[0] && memOut_CT$wnnz_Int_dbuf_d[0]))
      unique case (memMergeChoice_CT$wnnz_Int_d[1:1])
        1'd0: memOut_CT$wnnz_Int_dbuf_onehotd = 2'd1;
        1'd1: memOut_CT$wnnz_Int_dbuf_onehotd = 2'd2;
        default: memOut_CT$wnnz_Int_dbuf_onehotd = 2'd0;
      endcase
    else memOut_CT$wnnz_Int_dbuf_onehotd = 2'd0;
  assign memReadOut_CT$wnnz_Int_d = {memOut_CT$wnnz_Int_dbuf_d[116:1],
                                     memOut_CT$wnnz_Int_dbuf_onehotd[0]};
  assign memWriteOut_CT$wnnz_Int_d = {memOut_CT$wnnz_Int_dbuf_d[116:1],
                                      memOut_CT$wnnz_Int_dbuf_onehotd[1]};
  assign memOut_CT$wnnz_Int_dbuf_r = (| (memOut_CT$wnnz_Int_dbuf_onehotd & {memWriteOut_CT$wnnz_Int_r,
                                                                            memReadOut_CT$wnnz_Int_r}));
  assign memMergeChoice_CT$wnnz_Int_r = memOut_CT$wnnz_Int_dbuf_r;
  
  /* dbuf (Ty MemIn_CT$wnnz_Int) : (memMergeIn_CT$wnnz_Int_rbuf,MemIn_CT$wnnz_Int) > (memMergeIn_CT$wnnz_Int_dbuf,MemIn_CT$wnnz_Int) */
  assign memMergeIn_CT$wnnz_Int_rbuf_r = ((! memMergeIn_CT$wnnz_Int_dbuf_d[0]) || memMergeIn_CT$wnnz_Int_dbuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      memMergeIn_CT$wnnz_Int_dbuf_d <= {132'd0, 1'd0};
    else
      if (memMergeIn_CT$wnnz_Int_rbuf_r)
        memMergeIn_CT$wnnz_Int_dbuf_d <= memMergeIn_CT$wnnz_Int_rbuf_d;
  
  /* rbuf (Ty MemIn_CT$wnnz_Int) : (memMergeIn_CT$wnnz_Int,MemIn_CT$wnnz_Int) > (memMergeIn_CT$wnnz_Int_rbuf,MemIn_CT$wnnz_Int) */
  MemIn_CT$wnnz_Int_t memMergeIn_CT$wnnz_Int_buf;
  assign memMergeIn_CT$wnnz_Int_r = (! memMergeIn_CT$wnnz_Int_buf[0]);
  assign memMergeIn_CT$wnnz_Int_rbuf_d = (memMergeIn_CT$wnnz_Int_buf[0] ? memMergeIn_CT$wnnz_Int_buf :
                                          memMergeIn_CT$wnnz_Int_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memMergeIn_CT$wnnz_Int_buf <= {132'd0, 1'd0};
    else
      if ((memMergeIn_CT$wnnz_Int_rbuf_r && memMergeIn_CT$wnnz_Int_buf[0]))
        memMergeIn_CT$wnnz_Int_buf <= {132'd0, 1'd0};
      else if (((! memMergeIn_CT$wnnz_Int_rbuf_r) && (! memMergeIn_CT$wnnz_Int_buf[0])))
        memMergeIn_CT$wnnz_Int_buf <= memMergeIn_CT$wnnz_Int_d;
  
  /* dbuf (Ty MemOut_CT$wnnz_Int) : (memOut_CT$wnnz_Int_rbuf,MemOut_CT$wnnz_Int) > (memOut_CT$wnnz_Int_dbuf,MemOut_CT$wnnz_Int) */
  assign memOut_CT$wnnz_Int_rbuf_r = ((! memOut_CT$wnnz_Int_dbuf_d[0]) || memOut_CT$wnnz_Int_dbuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memOut_CT$wnnz_Int_dbuf_d <= {116'd0, 1'd0};
    else
      if (memOut_CT$wnnz_Int_rbuf_r)
        memOut_CT$wnnz_Int_dbuf_d <= memOut_CT$wnnz_Int_rbuf_d;
  
  /* rbuf (Ty MemOut_CT$wnnz_Int) : (memOut_CT$wnnz_Int,MemOut_CT$wnnz_Int) > (memOut_CT$wnnz_Int_rbuf,MemOut_CT$wnnz_Int) */
  MemOut_CT$wnnz_Int_t memOut_CT$wnnz_Int_buf;
  assign memOut_CT$wnnz_Int_r = (! memOut_CT$wnnz_Int_buf[0]);
  assign memOut_CT$wnnz_Int_rbuf_d = (memOut_CT$wnnz_Int_buf[0] ? memOut_CT$wnnz_Int_buf :
                                      memOut_CT$wnnz_Int_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memOut_CT$wnnz_Int_buf <= {116'd0, 1'd0};
    else
      if ((memOut_CT$wnnz_Int_rbuf_r && memOut_CT$wnnz_Int_buf[0]))
        memOut_CT$wnnz_Int_buf <= {116'd0, 1'd0};
      else if (((! memOut_CT$wnnz_Int_rbuf_r) && (! memOut_CT$wnnz_Int_buf[0])))
        memOut_CT$wnnz_Int_buf <= memOut_CT$wnnz_Int_d;
  
  /* destruct (Ty Pointer_CT$wnnz_Int,
          Dcon Pointer_CT$wnnz_Int) : (scfarg_0_1_1_argbuf,Pointer_CT$wnnz_Int) > [(destructReadIn_CT$wnnz_Int,Word16#)] */
  assign destructReadIn_CT$wnnz_Int_d = {scfarg_0_1_1_argbuf_d[16:1],
                                         scfarg_0_1_1_argbuf_d[0]};
  assign scfarg_0_1_1_argbuf_r = destructReadIn_CT$wnnz_Int_r;
  
  /* dcon (Ty MemIn_CT$wnnz_Int,
      Dcon ReadIn_CT$wnnz_Int) : [(destructReadIn_CT$wnnz_Int,Word16#)] > (dconReadIn_CT$wnnz_Int,MemIn_CT$wnnz_Int) */
  assign dconReadIn_CT$wnnz_Int_d = ReadIn_CT$wnnz_Int_dc((& {destructReadIn_CT$wnnz_Int_d[0]}), destructReadIn_CT$wnnz_Int_d);
  assign {destructReadIn_CT$wnnz_Int_r} = {1 {(dconReadIn_CT$wnnz_Int_r && dconReadIn_CT$wnnz_Int_d[0])}};
  
  /* destruct (Ty MemOut_CT$wnnz_Int,
          Dcon ReadOut_CT$wnnz_Int) : (memReadOut_CT$wnnz_Int,MemOut_CT$wnnz_Int) > [(readPointer_CT$wnnz_Intscfarg_0_1_1_argbuf,CT$wnnz_Int)] */
  assign readPointer_CT$wnnz_Intscfarg_0_1_1_argbuf_d = {memReadOut_CT$wnnz_Int_d[116:2],
                                                         memReadOut_CT$wnnz_Int_d[0]};
  assign memReadOut_CT$wnnz_Int_r = readPointer_CT$wnnz_Intscfarg_0_1_1_argbuf_r;
  
  /* mergectrl (Ty C5,
           Ty CT$wnnz_Int) : [(lizzieLet13_1_1_argbuf,CT$wnnz_Int),
                              (lizzieLet1_1_argbuf,CT$wnnz_Int),
                              (lizzieLet28_1_argbuf,CT$wnnz_Int),
                              (lizzieLet29_1_argbuf,CT$wnnz_Int),
                              (lizzieLet30_1_argbuf,CT$wnnz_Int)] > (writeMerge_choice_CT$wnnz_Int,C5) (writeMerge_data_CT$wnnz_Int,CT$wnnz_Int) */
  logic [4:0] lizzieLet13_1_1_argbuf_select_d;
  assign lizzieLet13_1_1_argbuf_select_d = ((| lizzieLet13_1_1_argbuf_select_q) ? lizzieLet13_1_1_argbuf_select_q :
                                            (lizzieLet13_1_1_argbuf_d[0] ? 5'd1 :
                                             (lizzieLet1_1_argbuf_d[0] ? 5'd2 :
                                              (lizzieLet28_1_argbuf_d[0] ? 5'd4 :
                                               (lizzieLet29_1_argbuf_d[0] ? 5'd8 :
                                                (lizzieLet30_1_argbuf_d[0] ? 5'd16 :
                                                 5'd0))))));
  logic [4:0] lizzieLet13_1_1_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet13_1_1_argbuf_select_q <= 5'd0;
    else
      lizzieLet13_1_1_argbuf_select_q <= (lizzieLet13_1_1_argbuf_done ? 5'd0 :
                                          lizzieLet13_1_1_argbuf_select_d);
  logic [1:0] lizzieLet13_1_1_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet13_1_1_argbuf_emit_q <= 2'd0;
    else
      lizzieLet13_1_1_argbuf_emit_q <= (lizzieLet13_1_1_argbuf_done ? 2'd0 :
                                        lizzieLet13_1_1_argbuf_emit_d);
  logic [1:0] lizzieLet13_1_1_argbuf_emit_d;
  assign lizzieLet13_1_1_argbuf_emit_d = (lizzieLet13_1_1_argbuf_emit_q | ({writeMerge_choice_CT$wnnz_Int_d[0],
                                                                            writeMerge_data_CT$wnnz_Int_d[0]} & {writeMerge_choice_CT$wnnz_Int_r,
                                                                                                                 writeMerge_data_CT$wnnz_Int_r}));
  logic lizzieLet13_1_1_argbuf_done;
  assign lizzieLet13_1_1_argbuf_done = (& lizzieLet13_1_1_argbuf_emit_d);
  assign {lizzieLet30_1_argbuf_r,
          lizzieLet29_1_argbuf_r,
          lizzieLet28_1_argbuf_r,
          lizzieLet1_1_argbuf_r,
          lizzieLet13_1_1_argbuf_r} = (lizzieLet13_1_1_argbuf_done ? lizzieLet13_1_1_argbuf_select_d :
                                       5'd0);
  assign writeMerge_data_CT$wnnz_Int_d = ((lizzieLet13_1_1_argbuf_select_d[0] && (! lizzieLet13_1_1_argbuf_emit_q[0])) ? lizzieLet13_1_1_argbuf_d :
                                          ((lizzieLet13_1_1_argbuf_select_d[1] && (! lizzieLet13_1_1_argbuf_emit_q[0])) ? lizzieLet1_1_argbuf_d :
                                           ((lizzieLet13_1_1_argbuf_select_d[2] && (! lizzieLet13_1_1_argbuf_emit_q[0])) ? lizzieLet28_1_argbuf_d :
                                            ((lizzieLet13_1_1_argbuf_select_d[3] && (! lizzieLet13_1_1_argbuf_emit_q[0])) ? lizzieLet29_1_argbuf_d :
                                             ((lizzieLet13_1_1_argbuf_select_d[4] && (! lizzieLet13_1_1_argbuf_emit_q[0])) ? lizzieLet30_1_argbuf_d :
                                              {115'd0, 1'd0})))));
  assign writeMerge_choice_CT$wnnz_Int_d = ((lizzieLet13_1_1_argbuf_select_d[0] && (! lizzieLet13_1_1_argbuf_emit_q[1])) ? C1_5_dc(1'd1) :
                                            ((lizzieLet13_1_1_argbuf_select_d[1] && (! lizzieLet13_1_1_argbuf_emit_q[1])) ? C2_5_dc(1'd1) :
                                             ((lizzieLet13_1_1_argbuf_select_d[2] && (! lizzieLet13_1_1_argbuf_emit_q[1])) ? C3_5_dc(1'd1) :
                                              ((lizzieLet13_1_1_argbuf_select_d[3] && (! lizzieLet13_1_1_argbuf_emit_q[1])) ? C4_5_dc(1'd1) :
                                               ((lizzieLet13_1_1_argbuf_select_d[4] && (! lizzieLet13_1_1_argbuf_emit_q[1])) ? C5_5_dc(1'd1) :
                                                {3'd0, 1'd0})))));
  
  /* demux (Ty C5,
       Ty Pointer_CT$wnnz_Int) : (writeMerge_choice_CT$wnnz_Int,C5) (demuxWriteResult_CT$wnnz_Int,Pointer_CT$wnnz_Int) > [(writeCT$wnnz_IntlizzieLet13_1_1_argbuf,Pointer_CT$wnnz_Int),
                                                                                                                          (writeCT$wnnz_IntlizzieLet1_1_argbuf,Pointer_CT$wnnz_Int),
                                                                                                                          (writeCT$wnnz_IntlizzieLet28_1_argbuf,Pointer_CT$wnnz_Int),
                                                                                                                          (writeCT$wnnz_IntlizzieLet29_1_argbuf,Pointer_CT$wnnz_Int),
                                                                                                                          (writeCT$wnnz_IntlizzieLet30_1_argbuf,Pointer_CT$wnnz_Int)] */
  logic [4:0] demuxWriteResult_CT$wnnz_Int_onehotd;
  always_comb
    if ((writeMerge_choice_CT$wnnz_Int_d[0] && demuxWriteResult_CT$wnnz_Int_d[0]))
      unique case (writeMerge_choice_CT$wnnz_Int_d[3:1])
        3'd0: demuxWriteResult_CT$wnnz_Int_onehotd = 5'd1;
        3'd1: demuxWriteResult_CT$wnnz_Int_onehotd = 5'd2;
        3'd2: demuxWriteResult_CT$wnnz_Int_onehotd = 5'd4;
        3'd3: demuxWriteResult_CT$wnnz_Int_onehotd = 5'd8;
        3'd4: demuxWriteResult_CT$wnnz_Int_onehotd = 5'd16;
        default: demuxWriteResult_CT$wnnz_Int_onehotd = 5'd0;
      endcase
    else demuxWriteResult_CT$wnnz_Int_onehotd = 5'd0;
  assign writeCT$wnnz_IntlizzieLet13_1_1_argbuf_d = {demuxWriteResult_CT$wnnz_Int_d[16:1],
                                                     demuxWriteResult_CT$wnnz_Int_onehotd[0]};
  assign writeCT$wnnz_IntlizzieLet1_1_argbuf_d = {demuxWriteResult_CT$wnnz_Int_d[16:1],
                                                  demuxWriteResult_CT$wnnz_Int_onehotd[1]};
  assign writeCT$wnnz_IntlizzieLet28_1_argbuf_d = {demuxWriteResult_CT$wnnz_Int_d[16:1],
                                                   demuxWriteResult_CT$wnnz_Int_onehotd[2]};
  assign writeCT$wnnz_IntlizzieLet29_1_argbuf_d = {demuxWriteResult_CT$wnnz_Int_d[16:1],
                                                   demuxWriteResult_CT$wnnz_Int_onehotd[3]};
  assign writeCT$wnnz_IntlizzieLet30_1_argbuf_d = {demuxWriteResult_CT$wnnz_Int_d[16:1],
                                                   demuxWriteResult_CT$wnnz_Int_onehotd[4]};
  assign demuxWriteResult_CT$wnnz_Int_r = (| (demuxWriteResult_CT$wnnz_Int_onehotd & {writeCT$wnnz_IntlizzieLet30_1_argbuf_r,
                                                                                      writeCT$wnnz_IntlizzieLet29_1_argbuf_r,
                                                                                      writeCT$wnnz_IntlizzieLet28_1_argbuf_r,
                                                                                      writeCT$wnnz_IntlizzieLet1_1_argbuf_r,
                                                                                      writeCT$wnnz_IntlizzieLet13_1_1_argbuf_r}));
  assign writeMerge_choice_CT$wnnz_Int_r = demuxWriteResult_CT$wnnz_Int_r;
  
  /* dcon (Ty MemIn_CT$wnnz_Int,
      Dcon WriteIn_CT$wnnz_Int) : [(forkHP1_CT$wnnz_In2,Word16#),
                                   (writeMerge_data_CT$wnnz_Int,CT$wnnz_Int)] > (dconWriteIn_CT$wnnz_Int,MemIn_CT$wnnz_Int) */
  assign dconWriteIn_CT$wnnz_Int_d = WriteIn_CT$wnnz_Int_dc((& {forkHP1_CT$wnnz_In2_d[0],
                                                                writeMerge_data_CT$wnnz_Int_d[0]}), forkHP1_CT$wnnz_In2_d, writeMerge_data_CT$wnnz_Int_d);
  assign {forkHP1_CT$wnnz_In2_r,
          writeMerge_data_CT$wnnz_Int_r} = {2 {(dconWriteIn_CT$wnnz_Int_r && dconWriteIn_CT$wnnz_Int_d[0])}};
  
  /* dcon (Ty Pointer_CT$wnnz_Int,
      Dcon Pointer_CT$wnnz_Int) : [(forkHP1_CT$wnnz_In3,Word16#)] > (dconPtr_CT$wnnz_Int,Pointer_CT$wnnz_Int) */
  assign dconPtr_CT$wnnz_Int_d = Pointer_CT$wnnz_Int_dc((& {forkHP1_CT$wnnz_In3_d[0]}), forkHP1_CT$wnnz_In3_d);
  assign {forkHP1_CT$wnnz_In3_r} = {1 {(dconPtr_CT$wnnz_Int_r && dconPtr_CT$wnnz_Int_d[0])}};
  
  /* demux (Ty MemOut_CT$wnnz_Int,
       Ty Pointer_CT$wnnz_Int) : (memWriteOut_CT$wnnz_Int,MemOut_CT$wnnz_Int) (dconPtr_CT$wnnz_Int,Pointer_CT$wnnz_Int) > [(_76,Pointer_CT$wnnz_Int),
                                                                                                                           (demuxWriteResult_CT$wnnz_Int,Pointer_CT$wnnz_Int)] */
  logic [1:0] dconPtr_CT$wnnz_Int_onehotd;
  always_comb
    if ((memWriteOut_CT$wnnz_Int_d[0] && dconPtr_CT$wnnz_Int_d[0]))
      unique case (memWriteOut_CT$wnnz_Int_d[1:1])
        1'd0: dconPtr_CT$wnnz_Int_onehotd = 2'd1;
        1'd1: dconPtr_CT$wnnz_Int_onehotd = 2'd2;
        default: dconPtr_CT$wnnz_Int_onehotd = 2'd0;
      endcase
    else dconPtr_CT$wnnz_Int_onehotd = 2'd0;
  assign _76_d = {dconPtr_CT$wnnz_Int_d[16:1],
                  dconPtr_CT$wnnz_Int_onehotd[0]};
  assign demuxWriteResult_CT$wnnz_Int_d = {dconPtr_CT$wnnz_Int_d[16:1],
                                           dconPtr_CT$wnnz_Int_onehotd[1]};
  assign dconPtr_CT$wnnz_Int_r = (| (dconPtr_CT$wnnz_Int_onehotd & {demuxWriteResult_CT$wnnz_Int_r,
                                                                    _76_r}));
  assign memWriteOut_CT$wnnz_Int_r = dconPtr_CT$wnnz_Int_r;
  
  /* const (Ty Word16#,
       Lit 0) : (go__9,Go) > (initHP_CTmain_mask_Int,Word16#) */
  assign initHP_CTmain_mask_Int_d = {16'd0, go__9_d[0]};
  assign go__9_r = initHP_CTmain_mask_Int_r;
  
  /* const (Ty Word16#,
       Lit 1) : (incrHP_CTmain_mask_Int1,Go) > (incrHP_CTmain_mask_Int,Word16#) */
  assign incrHP_CTmain_mask_Int_d = {16'd1,
                                     incrHP_CTmain_mask_Int1_d[0]};
  assign incrHP_CTmain_mask_Int1_r = incrHP_CTmain_mask_Int_r;
  
  /* merge (Ty Go) : [(go__10,Go),
                 (incrHP_CTmain_mask_Int2,Go)] > (incrHP_mergeCTmain_mask_Int,Go) */
  logic [1:0] incrHP_mergeCTmain_mask_Int_selected;
  logic [1:0] incrHP_mergeCTmain_mask_Int_select;
  always_comb
    begin
      incrHP_mergeCTmain_mask_Int_selected = 2'd0;
      if ((| incrHP_mergeCTmain_mask_Int_select))
        incrHP_mergeCTmain_mask_Int_selected = incrHP_mergeCTmain_mask_Int_select;
      else
        if (go__10_d[0]) incrHP_mergeCTmain_mask_Int_selected[0] = 1'd1;
        else if (incrHP_CTmain_mask_Int2_d[0])
          incrHP_mergeCTmain_mask_Int_selected[1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeCTmain_mask_Int_select <= 2'd0;
    else
      incrHP_mergeCTmain_mask_Int_select <= (incrHP_mergeCTmain_mask_Int_r ? 2'd0 :
                                             incrHP_mergeCTmain_mask_Int_selected);
  always_comb
    if (incrHP_mergeCTmain_mask_Int_selected[0])
      incrHP_mergeCTmain_mask_Int_d = go__10_d;
    else if (incrHP_mergeCTmain_mask_Int_selected[1])
      incrHP_mergeCTmain_mask_Int_d = incrHP_CTmain_mask_Int2_d;
    else incrHP_mergeCTmain_mask_Int_d = 1'd0;
  assign {incrHP_CTmain_mask_Int2_r,
          go__10_r} = (incrHP_mergeCTmain_mask_Int_r ? incrHP_mergeCTmain_mask_Int_selected :
                       2'd0);
  
  /* fork (Ty Go) : (incrHP_mergeCTmain_mask_Int_buf,Go) > [(incrHP_CTmain_mask_Int1,Go),
                                                       (incrHP_CTmain_mask_Int2,Go)] */
  logic [1:0] incrHP_mergeCTmain_mask_Int_buf_emitted;
  logic [1:0] incrHP_mergeCTmain_mask_Int_buf_done;
  assign incrHP_CTmain_mask_Int1_d = (incrHP_mergeCTmain_mask_Int_buf_d[0] && (! incrHP_mergeCTmain_mask_Int_buf_emitted[0]));
  assign incrHP_CTmain_mask_Int2_d = (incrHP_mergeCTmain_mask_Int_buf_d[0] && (! incrHP_mergeCTmain_mask_Int_buf_emitted[1]));
  assign incrHP_mergeCTmain_mask_Int_buf_done = (incrHP_mergeCTmain_mask_Int_buf_emitted | ({incrHP_CTmain_mask_Int2_d[0],
                                                                                             incrHP_CTmain_mask_Int1_d[0]} & {incrHP_CTmain_mask_Int2_r,
                                                                                                                              incrHP_CTmain_mask_Int1_r}));
  assign incrHP_mergeCTmain_mask_Int_buf_r = (& incrHP_mergeCTmain_mask_Int_buf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      incrHP_mergeCTmain_mask_Int_buf_emitted <= 2'd0;
    else
      incrHP_mergeCTmain_mask_Int_buf_emitted <= (incrHP_mergeCTmain_mask_Int_buf_r ? 2'd0 :
                                                  incrHP_mergeCTmain_mask_Int_buf_done);
  
  /* op_add (Ty Word16#) : (incrHP_CTmain_mask_Int,Word16#) (forkHP1_CTmain_mask_Int,Word16#) > (addHP_CTmain_mask_Int,Word16#) */
  assign addHP_CTmain_mask_Int_d = {(incrHP_CTmain_mask_Int_d[16:1] + forkHP1_CTmain_mask_Int_d[16:1]),
                                    (incrHP_CTmain_mask_Int_d[0] && forkHP1_CTmain_mask_Int_d[0])};
  assign {incrHP_CTmain_mask_Int_r,
          forkHP1_CTmain_mask_Int_r} = {2 {(addHP_CTmain_mask_Int_r && addHP_CTmain_mask_Int_d[0])}};
  
  /* merge (Ty Word16#) : [(initHP_CTmain_mask_Int,Word16#),
                      (addHP_CTmain_mask_Int,Word16#)] > (mergeHP_CTmain_mask_Int,Word16#) */
  logic [1:0] mergeHP_CTmain_mask_Int_selected;
  logic [1:0] mergeHP_CTmain_mask_Int_select;
  always_comb
    begin
      mergeHP_CTmain_mask_Int_selected = 2'd0;
      if ((| mergeHP_CTmain_mask_Int_select))
        mergeHP_CTmain_mask_Int_selected = mergeHP_CTmain_mask_Int_select;
      else
        if (initHP_CTmain_mask_Int_d[0])
          mergeHP_CTmain_mask_Int_selected[0] = 1'd1;
        else if (addHP_CTmain_mask_Int_d[0])
          mergeHP_CTmain_mask_Int_selected[1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_CTmain_mask_Int_select <= 2'd0;
    else
      mergeHP_CTmain_mask_Int_select <= (mergeHP_CTmain_mask_Int_r ? 2'd0 :
                                         mergeHP_CTmain_mask_Int_selected);
  always_comb
    if (mergeHP_CTmain_mask_Int_selected[0])
      mergeHP_CTmain_mask_Int_d = initHP_CTmain_mask_Int_d;
    else if (mergeHP_CTmain_mask_Int_selected[1])
      mergeHP_CTmain_mask_Int_d = addHP_CTmain_mask_Int_d;
    else mergeHP_CTmain_mask_Int_d = {16'd0, 1'd0};
  assign {addHP_CTmain_mask_Int_r,
          initHP_CTmain_mask_Int_r} = (mergeHP_CTmain_mask_Int_r ? mergeHP_CTmain_mask_Int_selected :
                                       2'd0);
  
  /* buf (Ty Go) : (incrHP_mergeCTmain_mask_Int,Go) > (incrHP_mergeCTmain_mask_Int_buf,Go) */
  Go_t incrHP_mergeCTmain_mask_Int_bufchan_d;
  logic incrHP_mergeCTmain_mask_Int_bufchan_r;
  assign incrHP_mergeCTmain_mask_Int_r = ((! incrHP_mergeCTmain_mask_Int_bufchan_d[0]) || incrHP_mergeCTmain_mask_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeCTmain_mask_Int_bufchan_d <= 1'd0;
    else
      if (incrHP_mergeCTmain_mask_Int_r)
        incrHP_mergeCTmain_mask_Int_bufchan_d <= incrHP_mergeCTmain_mask_Int_d;
  Go_t incrHP_mergeCTmain_mask_Int_bufchan_buf;
  assign incrHP_mergeCTmain_mask_Int_bufchan_r = (! incrHP_mergeCTmain_mask_Int_bufchan_buf[0]);
  assign incrHP_mergeCTmain_mask_Int_buf_d = (incrHP_mergeCTmain_mask_Int_bufchan_buf[0] ? incrHP_mergeCTmain_mask_Int_bufchan_buf :
                                              incrHP_mergeCTmain_mask_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      incrHP_mergeCTmain_mask_Int_bufchan_buf <= 1'd0;
    else
      if ((incrHP_mergeCTmain_mask_Int_buf_r && incrHP_mergeCTmain_mask_Int_bufchan_buf[0]))
        incrHP_mergeCTmain_mask_Int_bufchan_buf <= 1'd0;
      else if (((! incrHP_mergeCTmain_mask_Int_buf_r) && (! incrHP_mergeCTmain_mask_Int_bufchan_buf[0])))
        incrHP_mergeCTmain_mask_Int_bufchan_buf <= incrHP_mergeCTmain_mask_Int_bufchan_d;
  
  /* buf (Ty Word16#) : (mergeHP_CTmain_mask_Int,Word16#) > (mergeHP_CTmain_mask_Int_buf,Word16#) */
  \Word16#_t  mergeHP_CTmain_mask_Int_bufchan_d;
  logic mergeHP_CTmain_mask_Int_bufchan_r;
  assign mergeHP_CTmain_mask_Int_r = ((! mergeHP_CTmain_mask_Int_bufchan_d[0]) || mergeHP_CTmain_mask_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      mergeHP_CTmain_mask_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (mergeHP_CTmain_mask_Int_r)
        mergeHP_CTmain_mask_Int_bufchan_d <= mergeHP_CTmain_mask_Int_d;
  \Word16#_t  mergeHP_CTmain_mask_Int_bufchan_buf;
  assign mergeHP_CTmain_mask_Int_bufchan_r = (! mergeHP_CTmain_mask_Int_bufchan_buf[0]);
  assign mergeHP_CTmain_mask_Int_buf_d = (mergeHP_CTmain_mask_Int_bufchan_buf[0] ? mergeHP_CTmain_mask_Int_bufchan_buf :
                                          mergeHP_CTmain_mask_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      mergeHP_CTmain_mask_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((mergeHP_CTmain_mask_Int_buf_r && mergeHP_CTmain_mask_Int_bufchan_buf[0]))
        mergeHP_CTmain_mask_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! mergeHP_CTmain_mask_Int_buf_r) && (! mergeHP_CTmain_mask_Int_bufchan_buf[0])))
        mergeHP_CTmain_mask_Int_bufchan_buf <= mergeHP_CTmain_mask_Int_bufchan_d;
  
  /* fork (Ty Word16#) : (mergeHP_CTmain_mask_Int_buf,Word16#) > [(forkHP1_CTmain_mask_Int,Word16#),
                                                             (forkHP1_CTmain_mask_In2,Word16#),
                                                             (forkHP1_CTmain_mask_In3,Word16#)] */
  logic [2:0] mergeHP_CTmain_mask_Int_buf_emitted;
  logic [2:0] mergeHP_CTmain_mask_Int_buf_done;
  assign forkHP1_CTmain_mask_Int_d = {mergeHP_CTmain_mask_Int_buf_d[16:1],
                                      (mergeHP_CTmain_mask_Int_buf_d[0] && (! mergeHP_CTmain_mask_Int_buf_emitted[0]))};
  assign forkHP1_CTmain_mask_In2_d = {mergeHP_CTmain_mask_Int_buf_d[16:1],
                                      (mergeHP_CTmain_mask_Int_buf_d[0] && (! mergeHP_CTmain_mask_Int_buf_emitted[1]))};
  assign forkHP1_CTmain_mask_In3_d = {mergeHP_CTmain_mask_Int_buf_d[16:1],
                                      (mergeHP_CTmain_mask_Int_buf_d[0] && (! mergeHP_CTmain_mask_Int_buf_emitted[2]))};
  assign mergeHP_CTmain_mask_Int_buf_done = (mergeHP_CTmain_mask_Int_buf_emitted | ({forkHP1_CTmain_mask_In3_d[0],
                                                                                     forkHP1_CTmain_mask_In2_d[0],
                                                                                     forkHP1_CTmain_mask_Int_d[0]} & {forkHP1_CTmain_mask_In3_r,
                                                                                                                      forkHP1_CTmain_mask_In2_r,
                                                                                                                      forkHP1_CTmain_mask_Int_r}));
  assign mergeHP_CTmain_mask_Int_buf_r = (& mergeHP_CTmain_mask_Int_buf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_CTmain_mask_Int_buf_emitted <= 3'd0;
    else
      mergeHP_CTmain_mask_Int_buf_emitted <= (mergeHP_CTmain_mask_Int_buf_r ? 3'd0 :
                                              mergeHP_CTmain_mask_Int_buf_done);
  
  /* mergectrl (Ty C2,
           Ty MemIn_CTmain_mask_Int) : [(dconReadIn_CTmain_mask_Int,MemIn_CTmain_mask_Int),
                                        (dconWriteIn_CTmain_mask_Int,MemIn_CTmain_mask_Int)] > (memMergeChoice_CTmain_mask_Int,C2) (memMergeIn_CTmain_mask_Int,MemIn_CTmain_mask_Int) */
  logic [1:0] dconReadIn_CTmain_mask_Int_select_d;
  assign dconReadIn_CTmain_mask_Int_select_d = ((| dconReadIn_CTmain_mask_Int_select_q) ? dconReadIn_CTmain_mask_Int_select_q :
                                                (dconReadIn_CTmain_mask_Int_d[0] ? 2'd1 :
                                                 (dconWriteIn_CTmain_mask_Int_d[0] ? 2'd2 :
                                                  2'd0)));
  logic [1:0] dconReadIn_CTmain_mask_Int_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) dconReadIn_CTmain_mask_Int_select_q <= 2'd0;
    else
      dconReadIn_CTmain_mask_Int_select_q <= (dconReadIn_CTmain_mask_Int_done ? 2'd0 :
                                              dconReadIn_CTmain_mask_Int_select_d);
  logic [1:0] dconReadIn_CTmain_mask_Int_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) dconReadIn_CTmain_mask_Int_emit_q <= 2'd0;
    else
      dconReadIn_CTmain_mask_Int_emit_q <= (dconReadIn_CTmain_mask_Int_done ? 2'd0 :
                                            dconReadIn_CTmain_mask_Int_emit_d);
  logic [1:0] dconReadIn_CTmain_mask_Int_emit_d;
  assign dconReadIn_CTmain_mask_Int_emit_d = (dconReadIn_CTmain_mask_Int_emit_q | ({memMergeChoice_CTmain_mask_Int_d[0],
                                                                                    memMergeIn_CTmain_mask_Int_d[0]} & {memMergeChoice_CTmain_mask_Int_r,
                                                                                                                        memMergeIn_CTmain_mask_Int_r}));
  logic dconReadIn_CTmain_mask_Int_done;
  assign dconReadIn_CTmain_mask_Int_done = (& dconReadIn_CTmain_mask_Int_emit_d);
  assign {dconWriteIn_CTmain_mask_Int_r,
          dconReadIn_CTmain_mask_Int_r} = (dconReadIn_CTmain_mask_Int_done ? dconReadIn_CTmain_mask_Int_select_d :
                                           2'd0);
  assign memMergeIn_CTmain_mask_Int_d = ((dconReadIn_CTmain_mask_Int_select_d[0] && (! dconReadIn_CTmain_mask_Int_emit_q[0])) ? dconReadIn_CTmain_mask_Int_d :
                                         ((dconReadIn_CTmain_mask_Int_select_d[1] && (! dconReadIn_CTmain_mask_Int_emit_q[0])) ? dconWriteIn_CTmain_mask_Int_d :
                                          {132'd0, 1'd0}));
  assign memMergeChoice_CTmain_mask_Int_d = ((dconReadIn_CTmain_mask_Int_select_d[0] && (! dconReadIn_CTmain_mask_Int_emit_q[1])) ? C1_2_dc(1'd1) :
                                             ((dconReadIn_CTmain_mask_Int_select_d[1] && (! dconReadIn_CTmain_mask_Int_emit_q[1])) ? C2_2_dc(1'd1) :
                                              {1'd0, 1'd0}));
  
  /* bram (Ty MemIn_CTmain_mask_Int,
      Ty MemOut_CTmain_mask_Int) : (memMergeIn_CTmain_mask_Int_dbuf,MemIn_CTmain_mask_Int) > (memOut_CTmain_mask_Int,MemOut_CTmain_mask_Int) */
  logic [114:0] memMergeIn_CTmain_mask_Int_dbuf_mem[65535:0];
  logic [15:0] memMergeIn_CTmain_mask_Int_dbuf_address;
  logic [114:0] memMergeIn_CTmain_mask_Int_dbuf_din;
  logic [114:0] memOut_CTmain_mask_Int_q;
  logic memOut_CTmain_mask_Int_valid;
  logic memMergeIn_CTmain_mask_Int_dbuf_we;
  logic memOut_CTmain_mask_Int_we;
  assign memMergeIn_CTmain_mask_Int_dbuf_din = memMergeIn_CTmain_mask_Int_dbuf_d[132:18];
  assign memMergeIn_CTmain_mask_Int_dbuf_address = memMergeIn_CTmain_mask_Int_dbuf_d[17:2];
  assign memMergeIn_CTmain_mask_Int_dbuf_we = (memMergeIn_CTmain_mask_Int_dbuf_d[1:1] && memMergeIn_CTmain_mask_Int_dbuf_d[0]);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        memOut_CTmain_mask_Int_we <= 1'd0;
        memOut_CTmain_mask_Int_valid <= 1'd0;
      end
    else
      begin
        memOut_CTmain_mask_Int_we <= memMergeIn_CTmain_mask_Int_dbuf_we;
        memOut_CTmain_mask_Int_valid <= memMergeIn_CTmain_mask_Int_dbuf_d[0];
        if (memMergeIn_CTmain_mask_Int_dbuf_we)
          begin
            memMergeIn_CTmain_mask_Int_dbuf_mem[memMergeIn_CTmain_mask_Int_dbuf_address] <= memMergeIn_CTmain_mask_Int_dbuf_din;
            memOut_CTmain_mask_Int_q <= memMergeIn_CTmain_mask_Int_dbuf_din;
          end
        else
          memOut_CTmain_mask_Int_q <= memMergeIn_CTmain_mask_Int_dbuf_mem[memMergeIn_CTmain_mask_Int_dbuf_address];
      end
  assign memOut_CTmain_mask_Int_d = {memOut_CTmain_mask_Int_q,
                                     memOut_CTmain_mask_Int_we,
                                     memOut_CTmain_mask_Int_valid};
  assign memMergeIn_CTmain_mask_Int_dbuf_r = ((! memOut_CTmain_mask_Int_valid) || memOut_CTmain_mask_Int_r);
  
  /* demux (Ty C2,
       Ty MemOut_CTmain_mask_Int) : (memMergeChoice_CTmain_mask_Int,C2) (memOut_CTmain_mask_Int_dbuf,MemOut_CTmain_mask_Int) > [(memReadOut_CTmain_mask_Int,MemOut_CTmain_mask_Int),
                                                                                                                                (memWriteOut_CTmain_mask_Int,MemOut_CTmain_mask_Int)] */
  logic [1:0] memOut_CTmain_mask_Int_dbuf_onehotd;
  always_comb
    if ((memMergeChoice_CTmain_mask_Int_d[0] && memOut_CTmain_mask_Int_dbuf_d[0]))
      unique case (memMergeChoice_CTmain_mask_Int_d[1:1])
        1'd0: memOut_CTmain_mask_Int_dbuf_onehotd = 2'd1;
        1'd1: memOut_CTmain_mask_Int_dbuf_onehotd = 2'd2;
        default: memOut_CTmain_mask_Int_dbuf_onehotd = 2'd0;
      endcase
    else memOut_CTmain_mask_Int_dbuf_onehotd = 2'd0;
  assign memReadOut_CTmain_mask_Int_d = {memOut_CTmain_mask_Int_dbuf_d[116:1],
                                         memOut_CTmain_mask_Int_dbuf_onehotd[0]};
  assign memWriteOut_CTmain_mask_Int_d = {memOut_CTmain_mask_Int_dbuf_d[116:1],
                                          memOut_CTmain_mask_Int_dbuf_onehotd[1]};
  assign memOut_CTmain_mask_Int_dbuf_r = (| (memOut_CTmain_mask_Int_dbuf_onehotd & {memWriteOut_CTmain_mask_Int_r,
                                                                                    memReadOut_CTmain_mask_Int_r}));
  assign memMergeChoice_CTmain_mask_Int_r = memOut_CTmain_mask_Int_dbuf_r;
  
  /* dbuf (Ty MemIn_CTmain_mask_Int) : (memMergeIn_CTmain_mask_Int_rbuf,MemIn_CTmain_mask_Int) > (memMergeIn_CTmain_mask_Int_dbuf,MemIn_CTmain_mask_Int) */
  assign memMergeIn_CTmain_mask_Int_rbuf_r = ((! memMergeIn_CTmain_mask_Int_dbuf_d[0]) || memMergeIn_CTmain_mask_Int_dbuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      memMergeIn_CTmain_mask_Int_dbuf_d <= {132'd0, 1'd0};
    else
      if (memMergeIn_CTmain_mask_Int_rbuf_r)
        memMergeIn_CTmain_mask_Int_dbuf_d <= memMergeIn_CTmain_mask_Int_rbuf_d;
  
  /* rbuf (Ty MemIn_CTmain_mask_Int) : (memMergeIn_CTmain_mask_Int,MemIn_CTmain_mask_Int) > (memMergeIn_CTmain_mask_Int_rbuf,MemIn_CTmain_mask_Int) */
  MemIn_CTmain_mask_Int_t memMergeIn_CTmain_mask_Int_buf;
  assign memMergeIn_CTmain_mask_Int_r = (! memMergeIn_CTmain_mask_Int_buf[0]);
  assign memMergeIn_CTmain_mask_Int_rbuf_d = (memMergeIn_CTmain_mask_Int_buf[0] ? memMergeIn_CTmain_mask_Int_buf :
                                              memMergeIn_CTmain_mask_Int_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      memMergeIn_CTmain_mask_Int_buf <= {132'd0, 1'd0};
    else
      if ((memMergeIn_CTmain_mask_Int_rbuf_r && memMergeIn_CTmain_mask_Int_buf[0]))
        memMergeIn_CTmain_mask_Int_buf <= {132'd0, 1'd0};
      else if (((! memMergeIn_CTmain_mask_Int_rbuf_r) && (! memMergeIn_CTmain_mask_Int_buf[0])))
        memMergeIn_CTmain_mask_Int_buf <= memMergeIn_CTmain_mask_Int_d;
  
  /* dbuf (Ty MemOut_CTmain_mask_Int) : (memOut_CTmain_mask_Int_rbuf,MemOut_CTmain_mask_Int) > (memOut_CTmain_mask_Int_dbuf,MemOut_CTmain_mask_Int) */
  assign memOut_CTmain_mask_Int_rbuf_r = ((! memOut_CTmain_mask_Int_dbuf_d[0]) || memOut_CTmain_mask_Int_dbuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      memOut_CTmain_mask_Int_dbuf_d <= {116'd0, 1'd0};
    else
      if (memOut_CTmain_mask_Int_rbuf_r)
        memOut_CTmain_mask_Int_dbuf_d <= memOut_CTmain_mask_Int_rbuf_d;
  
  /* rbuf (Ty MemOut_CTmain_mask_Int) : (memOut_CTmain_mask_Int,MemOut_CTmain_mask_Int) > (memOut_CTmain_mask_Int_rbuf,MemOut_CTmain_mask_Int) */
  MemOut_CTmain_mask_Int_t memOut_CTmain_mask_Int_buf;
  assign memOut_CTmain_mask_Int_r = (! memOut_CTmain_mask_Int_buf[0]);
  assign memOut_CTmain_mask_Int_rbuf_d = (memOut_CTmain_mask_Int_buf[0] ? memOut_CTmain_mask_Int_buf :
                                          memOut_CTmain_mask_Int_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memOut_CTmain_mask_Int_buf <= {116'd0, 1'd0};
    else
      if ((memOut_CTmain_mask_Int_rbuf_r && memOut_CTmain_mask_Int_buf[0]))
        memOut_CTmain_mask_Int_buf <= {116'd0, 1'd0};
      else if (((! memOut_CTmain_mask_Int_rbuf_r) && (! memOut_CTmain_mask_Int_buf[0])))
        memOut_CTmain_mask_Int_buf <= memOut_CTmain_mask_Int_d;
  
  /* destruct (Ty Pointer_CTmain_mask_Int,
          Dcon Pointer_CTmain_mask_Int) : (scfarg_0_2_1_argbuf,Pointer_CTmain_mask_Int) > [(destructReadIn_CTmain_mask_Int,Word16#)] */
  assign destructReadIn_CTmain_mask_Int_d = {scfarg_0_2_1_argbuf_d[16:1],
                                             scfarg_0_2_1_argbuf_d[0]};
  assign scfarg_0_2_1_argbuf_r = destructReadIn_CTmain_mask_Int_r;
  
  /* dcon (Ty MemIn_CTmain_mask_Int,
      Dcon ReadIn_CTmain_mask_Int) : [(destructReadIn_CTmain_mask_Int,Word16#)] > (dconReadIn_CTmain_mask_Int,MemIn_CTmain_mask_Int) */
  assign dconReadIn_CTmain_mask_Int_d = ReadIn_CTmain_mask_Int_dc((& {destructReadIn_CTmain_mask_Int_d[0]}), destructReadIn_CTmain_mask_Int_d);
  assign {destructReadIn_CTmain_mask_Int_r} = {1 {(dconReadIn_CTmain_mask_Int_r && dconReadIn_CTmain_mask_Int_d[0])}};
  
  /* destruct (Ty MemOut_CTmain_mask_Int,
          Dcon ReadOut_CTmain_mask_Int) : (memReadOut_CTmain_mask_Int,MemOut_CTmain_mask_Int) > [(readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf,CTmain_mask_Int)] */
  assign readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf_d = {memReadOut_CTmain_mask_Int_d[116:2],
                                                             memReadOut_CTmain_mask_Int_d[0]};
  assign memReadOut_CTmain_mask_Int_r = readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf_r;
  
  /* mergectrl (Ty C5,
           Ty CTmain_mask_Int) : [(lizzieLet19_1_argbuf,CTmain_mask_Int),
                                  (lizzieLet21_1_argbuf,CTmain_mask_Int),
                                  (lizzieLet32_1_argbuf,CTmain_mask_Int),
                                  (lizzieLet33_1_argbuf,CTmain_mask_Int),
                                  (lizzieLet34_1_argbuf,CTmain_mask_Int)] > (writeMerge_choice_CTmain_mask_Int,C5) (writeMerge_data_CTmain_mask_Int,CTmain_mask_Int) */
  logic [4:0] lizzieLet19_1_argbuf_select_d;
  assign lizzieLet19_1_argbuf_select_d = ((| lizzieLet19_1_argbuf_select_q) ? lizzieLet19_1_argbuf_select_q :
                                          (lizzieLet19_1_argbuf_d[0] ? 5'd1 :
                                           (lizzieLet21_1_argbuf_d[0] ? 5'd2 :
                                            (lizzieLet32_1_argbuf_d[0] ? 5'd4 :
                                             (lizzieLet33_1_argbuf_d[0] ? 5'd8 :
                                              (lizzieLet34_1_argbuf_d[0] ? 5'd16 :
                                               5'd0))))));
  logic [4:0] lizzieLet19_1_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet19_1_argbuf_select_q <= 5'd0;
    else
      lizzieLet19_1_argbuf_select_q <= (lizzieLet19_1_argbuf_done ? 5'd0 :
                                        lizzieLet19_1_argbuf_select_d);
  logic [1:0] lizzieLet19_1_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet19_1_argbuf_emit_q <= 2'd0;
    else
      lizzieLet19_1_argbuf_emit_q <= (lizzieLet19_1_argbuf_done ? 2'd0 :
                                      lizzieLet19_1_argbuf_emit_d);
  logic [1:0] lizzieLet19_1_argbuf_emit_d;
  assign lizzieLet19_1_argbuf_emit_d = (lizzieLet19_1_argbuf_emit_q | ({writeMerge_choice_CTmain_mask_Int_d[0],
                                                                        writeMerge_data_CTmain_mask_Int_d[0]} & {writeMerge_choice_CTmain_mask_Int_r,
                                                                                                                 writeMerge_data_CTmain_mask_Int_r}));
  logic lizzieLet19_1_argbuf_done;
  assign lizzieLet19_1_argbuf_done = (& lizzieLet19_1_argbuf_emit_d);
  assign {lizzieLet34_1_argbuf_r,
          lizzieLet33_1_argbuf_r,
          lizzieLet32_1_argbuf_r,
          lizzieLet21_1_argbuf_r,
          lizzieLet19_1_argbuf_r} = (lizzieLet19_1_argbuf_done ? lizzieLet19_1_argbuf_select_d :
                                     5'd0);
  assign writeMerge_data_CTmain_mask_Int_d = ((lizzieLet19_1_argbuf_select_d[0] && (! lizzieLet19_1_argbuf_emit_q[0])) ? lizzieLet19_1_argbuf_d :
                                              ((lizzieLet19_1_argbuf_select_d[1] && (! lizzieLet19_1_argbuf_emit_q[0])) ? lizzieLet21_1_argbuf_d :
                                               ((lizzieLet19_1_argbuf_select_d[2] && (! lizzieLet19_1_argbuf_emit_q[0])) ? lizzieLet32_1_argbuf_d :
                                                ((lizzieLet19_1_argbuf_select_d[3] && (! lizzieLet19_1_argbuf_emit_q[0])) ? lizzieLet33_1_argbuf_d :
                                                 ((lizzieLet19_1_argbuf_select_d[4] && (! lizzieLet19_1_argbuf_emit_q[0])) ? lizzieLet34_1_argbuf_d :
                                                  {115'd0, 1'd0})))));
  assign writeMerge_choice_CTmain_mask_Int_d = ((lizzieLet19_1_argbuf_select_d[0] && (! lizzieLet19_1_argbuf_emit_q[1])) ? C1_5_dc(1'd1) :
                                                ((lizzieLet19_1_argbuf_select_d[1] && (! lizzieLet19_1_argbuf_emit_q[1])) ? C2_5_dc(1'd1) :
                                                 ((lizzieLet19_1_argbuf_select_d[2] && (! lizzieLet19_1_argbuf_emit_q[1])) ? C3_5_dc(1'd1) :
                                                  ((lizzieLet19_1_argbuf_select_d[3] && (! lizzieLet19_1_argbuf_emit_q[1])) ? C4_5_dc(1'd1) :
                                                   ((lizzieLet19_1_argbuf_select_d[4] && (! lizzieLet19_1_argbuf_emit_q[1])) ? C5_5_dc(1'd1) :
                                                    {3'd0, 1'd0})))));
  
  /* demux (Ty C5,
       Ty Pointer_CTmain_mask_Int) : (writeMerge_choice_CTmain_mask_Int,C5) (demuxWriteResult_CTmain_mask_Int,Pointer_CTmain_mask_Int) > [(writeCTmain_mask_IntlizzieLet19_1_argbuf,Pointer_CTmain_mask_Int),
                                                                                                                                          (writeCTmain_mask_IntlizzieLet21_1_argbuf,Pointer_CTmain_mask_Int),
                                                                                                                                          (writeCTmain_mask_IntlizzieLet32_1_argbuf,Pointer_CTmain_mask_Int),
                                                                                                                                          (writeCTmain_mask_IntlizzieLet33_1_argbuf,Pointer_CTmain_mask_Int),
                                                                                                                                          (writeCTmain_mask_IntlizzieLet34_1_argbuf,Pointer_CTmain_mask_Int)] */
  logic [4:0] demuxWriteResult_CTmain_mask_Int_onehotd;
  always_comb
    if ((writeMerge_choice_CTmain_mask_Int_d[0] && demuxWriteResult_CTmain_mask_Int_d[0]))
      unique case (writeMerge_choice_CTmain_mask_Int_d[3:1])
        3'd0: demuxWriteResult_CTmain_mask_Int_onehotd = 5'd1;
        3'd1: demuxWriteResult_CTmain_mask_Int_onehotd = 5'd2;
        3'd2: demuxWriteResult_CTmain_mask_Int_onehotd = 5'd4;
        3'd3: demuxWriteResult_CTmain_mask_Int_onehotd = 5'd8;
        3'd4: demuxWriteResult_CTmain_mask_Int_onehotd = 5'd16;
        default: demuxWriteResult_CTmain_mask_Int_onehotd = 5'd0;
      endcase
    else demuxWriteResult_CTmain_mask_Int_onehotd = 5'd0;
  assign writeCTmain_mask_IntlizzieLet19_1_argbuf_d = {demuxWriteResult_CTmain_mask_Int_d[16:1],
                                                       demuxWriteResult_CTmain_mask_Int_onehotd[0]};
  assign writeCTmain_mask_IntlizzieLet21_1_argbuf_d = {demuxWriteResult_CTmain_mask_Int_d[16:1],
                                                       demuxWriteResult_CTmain_mask_Int_onehotd[1]};
  assign writeCTmain_mask_IntlizzieLet32_1_argbuf_d = {demuxWriteResult_CTmain_mask_Int_d[16:1],
                                                       demuxWriteResult_CTmain_mask_Int_onehotd[2]};
  assign writeCTmain_mask_IntlizzieLet33_1_argbuf_d = {demuxWriteResult_CTmain_mask_Int_d[16:1],
                                                       demuxWriteResult_CTmain_mask_Int_onehotd[3]};
  assign writeCTmain_mask_IntlizzieLet34_1_argbuf_d = {demuxWriteResult_CTmain_mask_Int_d[16:1],
                                                       demuxWriteResult_CTmain_mask_Int_onehotd[4]};
  assign demuxWriteResult_CTmain_mask_Int_r = (| (demuxWriteResult_CTmain_mask_Int_onehotd & {writeCTmain_mask_IntlizzieLet34_1_argbuf_r,
                                                                                              writeCTmain_mask_IntlizzieLet33_1_argbuf_r,
                                                                                              writeCTmain_mask_IntlizzieLet32_1_argbuf_r,
                                                                                              writeCTmain_mask_IntlizzieLet21_1_argbuf_r,
                                                                                              writeCTmain_mask_IntlizzieLet19_1_argbuf_r}));
  assign writeMerge_choice_CTmain_mask_Int_r = demuxWriteResult_CTmain_mask_Int_r;
  
  /* dcon (Ty MemIn_CTmain_mask_Int,
      Dcon WriteIn_CTmain_mask_Int) : [(forkHP1_CTmain_mask_In2,Word16#),
                                       (writeMerge_data_CTmain_mask_Int,CTmain_mask_Int)] > (dconWriteIn_CTmain_mask_Int,MemIn_CTmain_mask_Int) */
  assign dconWriteIn_CTmain_mask_Int_d = WriteIn_CTmain_mask_Int_dc((& {forkHP1_CTmain_mask_In2_d[0],
                                                                        writeMerge_data_CTmain_mask_Int_d[0]}), forkHP1_CTmain_mask_In2_d, writeMerge_data_CTmain_mask_Int_d);
  assign {forkHP1_CTmain_mask_In2_r,
          writeMerge_data_CTmain_mask_Int_r} = {2 {(dconWriteIn_CTmain_mask_Int_r && dconWriteIn_CTmain_mask_Int_d[0])}};
  
  /* dcon (Ty Pointer_CTmain_mask_Int,
      Dcon Pointer_CTmain_mask_Int) : [(forkHP1_CTmain_mask_In3,Word16#)] > (dconPtr_CTmain_mask_Int,Pointer_CTmain_mask_Int) */
  assign dconPtr_CTmain_mask_Int_d = Pointer_CTmain_mask_Int_dc((& {forkHP1_CTmain_mask_In3_d[0]}), forkHP1_CTmain_mask_In3_d);
  assign {forkHP1_CTmain_mask_In3_r} = {1 {(dconPtr_CTmain_mask_Int_r && dconPtr_CTmain_mask_Int_d[0])}};
  
  /* demux (Ty MemOut_CTmain_mask_Int,
       Ty Pointer_CTmain_mask_Int) : (memWriteOut_CTmain_mask_Int,MemOut_CTmain_mask_Int) (dconPtr_CTmain_mask_Int,Pointer_CTmain_mask_Int) > [(_75,Pointer_CTmain_mask_Int),
                                                                                                                                               (demuxWriteResult_CTmain_mask_Int,Pointer_CTmain_mask_Int)] */
  logic [1:0] dconPtr_CTmain_mask_Int_onehotd;
  always_comb
    if ((memWriteOut_CTmain_mask_Int_d[0] && dconPtr_CTmain_mask_Int_d[0]))
      unique case (memWriteOut_CTmain_mask_Int_d[1:1])
        1'd0: dconPtr_CTmain_mask_Int_onehotd = 2'd1;
        1'd1: dconPtr_CTmain_mask_Int_onehotd = 2'd2;
        default: dconPtr_CTmain_mask_Int_onehotd = 2'd0;
      endcase
    else dconPtr_CTmain_mask_Int_onehotd = 2'd0;
  assign _75_d = {dconPtr_CTmain_mask_Int_d[16:1],
                  dconPtr_CTmain_mask_Int_onehotd[0]};
  assign demuxWriteResult_CTmain_mask_Int_d = {dconPtr_CTmain_mask_Int_d[16:1],
                                               dconPtr_CTmain_mask_Int_onehotd[1]};
  assign dconPtr_CTmain_mask_Int_r = (| (dconPtr_CTmain_mask_Int_onehotd & {demuxWriteResult_CTmain_mask_Int_r,
                                                                            _75_r}));
  assign memWriteOut_CTmain_mask_Int_r = dconPtr_CTmain_mask_Int_r;
  
  /* const (Ty Word16#,
       Lit 0) : (go_1_dummy_write_MaskQTree,Go) > (initHP_MaskQTree,Word16#) */
  assign initHP_MaskQTree_d = {16'd0,
                               go_1_dummy_write_MaskQTree_d[0]};
  assign go_1_dummy_write_MaskQTree_r = initHP_MaskQTree_r;
  
  /* const (Ty Word16#,
       Lit 1) : (incrHP_MaskQTree1,Go) > (incrHP_MaskQTree,Word16#) */
  assign incrHP_MaskQTree_d = {16'd1, incrHP_MaskQTree1_d[0]};
  assign incrHP_MaskQTree1_r = incrHP_MaskQTree_r;
  
  /* merge (Ty Go) : [(go_2_dummy_write_MaskQTree,Go),
                 (incrHP_MaskQTree2,Go)] > (incrHP_mergeMaskQTree,Go) */
  logic [1:0] incrHP_mergeMaskQTree_selected;
  logic [1:0] incrHP_mergeMaskQTree_select;
  always_comb
    begin
      incrHP_mergeMaskQTree_selected = 2'd0;
      if ((| incrHP_mergeMaskQTree_select))
        incrHP_mergeMaskQTree_selected = incrHP_mergeMaskQTree_select;
      else
        if (go_2_dummy_write_MaskQTree_d[0])
          incrHP_mergeMaskQTree_selected[0] = 1'd1;
        else if (incrHP_MaskQTree2_d[0])
          incrHP_mergeMaskQTree_selected[1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeMaskQTree_select <= 2'd0;
    else
      incrHP_mergeMaskQTree_select <= (incrHP_mergeMaskQTree_r ? 2'd0 :
                                       incrHP_mergeMaskQTree_selected);
  always_comb
    if (incrHP_mergeMaskQTree_selected[0])
      incrHP_mergeMaskQTree_d = go_2_dummy_write_MaskQTree_d;
    else if (incrHP_mergeMaskQTree_selected[1])
      incrHP_mergeMaskQTree_d = incrHP_MaskQTree2_d;
    else incrHP_mergeMaskQTree_d = 1'd0;
  assign {incrHP_MaskQTree2_r,
          go_2_dummy_write_MaskQTree_r} = (incrHP_mergeMaskQTree_r ? incrHP_mergeMaskQTree_selected :
                                           2'd0);
  
  /* fork (Ty Go) : (incrHP_mergeMaskQTree_buf,Go) > [(incrHP_MaskQTree1,Go),
                                                 (incrHP_MaskQTree2,Go)] */
  logic [1:0] incrHP_mergeMaskQTree_buf_emitted;
  logic [1:0] incrHP_mergeMaskQTree_buf_done;
  assign incrHP_MaskQTree1_d = (incrHP_mergeMaskQTree_buf_d[0] && (! incrHP_mergeMaskQTree_buf_emitted[0]));
  assign incrHP_MaskQTree2_d = (incrHP_mergeMaskQTree_buf_d[0] && (! incrHP_mergeMaskQTree_buf_emitted[1]));
  assign incrHP_mergeMaskQTree_buf_done = (incrHP_mergeMaskQTree_buf_emitted | ({incrHP_MaskQTree2_d[0],
                                                                                 incrHP_MaskQTree1_d[0]} & {incrHP_MaskQTree2_r,
                                                                                                            incrHP_MaskQTree1_r}));
  assign incrHP_mergeMaskQTree_buf_r = (& incrHP_mergeMaskQTree_buf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeMaskQTree_buf_emitted <= 2'd0;
    else
      incrHP_mergeMaskQTree_buf_emitted <= (incrHP_mergeMaskQTree_buf_r ? 2'd0 :
                                            incrHP_mergeMaskQTree_buf_done);
  
  /* op_add (Ty Word16#) : (incrHP_MaskQTree,Word16#) (forkHP1_MaskQTree,Word16#) > (addHP_MaskQTree,Word16#) */
  assign addHP_MaskQTree_d = {(incrHP_MaskQTree_d[16:1] + forkHP1_MaskQTree_d[16:1]),
                              (incrHP_MaskQTree_d[0] && forkHP1_MaskQTree_d[0])};
  assign {incrHP_MaskQTree_r,
          forkHP1_MaskQTree_r} = {2 {(addHP_MaskQTree_r && addHP_MaskQTree_d[0])}};
  
  /* merge (Ty Word16#) : [(initHP_MaskQTree,Word16#),
                      (addHP_MaskQTree,Word16#)] > (mergeHP_MaskQTree,Word16#) */
  logic [1:0] mergeHP_MaskQTree_selected;
  logic [1:0] mergeHP_MaskQTree_select;
  always_comb
    begin
      mergeHP_MaskQTree_selected = 2'd0;
      if ((| mergeHP_MaskQTree_select))
        mergeHP_MaskQTree_selected = mergeHP_MaskQTree_select;
      else
        if (initHP_MaskQTree_d[0]) mergeHP_MaskQTree_selected[0] = 1'd1;
        else if (addHP_MaskQTree_d[0])
          mergeHP_MaskQTree_selected[1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_MaskQTree_select <= 2'd0;
    else
      mergeHP_MaskQTree_select <= (mergeHP_MaskQTree_r ? 2'd0 :
                                   mergeHP_MaskQTree_selected);
  always_comb
    if (mergeHP_MaskQTree_selected[0])
      mergeHP_MaskQTree_d = initHP_MaskQTree_d;
    else if (mergeHP_MaskQTree_selected[1])
      mergeHP_MaskQTree_d = addHP_MaskQTree_d;
    else mergeHP_MaskQTree_d = {16'd0, 1'd0};
  assign {addHP_MaskQTree_r,
          initHP_MaskQTree_r} = (mergeHP_MaskQTree_r ? mergeHP_MaskQTree_selected :
                                 2'd0);
  
  /* buf (Ty Go) : (incrHP_mergeMaskQTree,Go) > (incrHP_mergeMaskQTree_buf,Go) */
  Go_t incrHP_mergeMaskQTree_bufchan_d;
  logic incrHP_mergeMaskQTree_bufchan_r;
  assign incrHP_mergeMaskQTree_r = ((! incrHP_mergeMaskQTree_bufchan_d[0]) || incrHP_mergeMaskQTree_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeMaskQTree_bufchan_d <= 1'd0;
    else
      if (incrHP_mergeMaskQTree_r)
        incrHP_mergeMaskQTree_bufchan_d <= incrHP_mergeMaskQTree_d;
  Go_t incrHP_mergeMaskQTree_bufchan_buf;
  assign incrHP_mergeMaskQTree_bufchan_r = (! incrHP_mergeMaskQTree_bufchan_buf[0]);
  assign incrHP_mergeMaskQTree_buf_d = (incrHP_mergeMaskQTree_bufchan_buf[0] ? incrHP_mergeMaskQTree_bufchan_buf :
                                        incrHP_mergeMaskQTree_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeMaskQTree_bufchan_buf <= 1'd0;
    else
      if ((incrHP_mergeMaskQTree_buf_r && incrHP_mergeMaskQTree_bufchan_buf[0]))
        incrHP_mergeMaskQTree_bufchan_buf <= 1'd0;
      else if (((! incrHP_mergeMaskQTree_buf_r) && (! incrHP_mergeMaskQTree_bufchan_buf[0])))
        incrHP_mergeMaskQTree_bufchan_buf <= incrHP_mergeMaskQTree_bufchan_d;
  
  /* buf (Ty Word16#) : (mergeHP_MaskQTree,Word16#) > (mergeHP_MaskQTree_buf,Word16#) */
  \Word16#_t  mergeHP_MaskQTree_bufchan_d;
  logic mergeHP_MaskQTree_bufchan_r;
  assign mergeHP_MaskQTree_r = ((! mergeHP_MaskQTree_bufchan_d[0]) || mergeHP_MaskQTree_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_MaskQTree_bufchan_d <= {16'd0, 1'd0};
    else
      if (mergeHP_MaskQTree_r)
        mergeHP_MaskQTree_bufchan_d <= mergeHP_MaskQTree_d;
  \Word16#_t  mergeHP_MaskQTree_bufchan_buf;
  assign mergeHP_MaskQTree_bufchan_r = (! mergeHP_MaskQTree_bufchan_buf[0]);
  assign mergeHP_MaskQTree_buf_d = (mergeHP_MaskQTree_bufchan_buf[0] ? mergeHP_MaskQTree_bufchan_buf :
                                    mergeHP_MaskQTree_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      mergeHP_MaskQTree_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((mergeHP_MaskQTree_buf_r && mergeHP_MaskQTree_bufchan_buf[0]))
        mergeHP_MaskQTree_bufchan_buf <= {16'd0, 1'd0};
      else if (((! mergeHP_MaskQTree_buf_r) && (! mergeHP_MaskQTree_bufchan_buf[0])))
        mergeHP_MaskQTree_bufchan_buf <= mergeHP_MaskQTree_bufchan_d;
  
  /* sink (Ty Word16#) : (forkHP1_MaskQTree_snk,Word16#) > */
  assign {forkHP1_MaskQTree_snk_r,
          forkHP1_MaskQTree_snk_dout} = {forkHP1_MaskQTree_snk_rout,
                                         forkHP1_MaskQTree_snk_d};
  
  /* source (Ty Go) : > (\MaskQTree_src,Go) */
  
  /* fork (Ty Go) : (\MaskQTree_src,Go) > [(go_1_dummy_write_MaskQTree,Go),
                                      (go_2_dummy_write_MaskQTree,Go)] */
  logic [1:0] \\MaskQTree_src_emitted ;
  logic [1:0] \\MaskQTree_src_done ;
  assign go_1_dummy_write_MaskQTree_d = (\\MaskQTree_src_d [0] && (! \\MaskQTree_src_emitted [0]));
  assign go_2_dummy_write_MaskQTree_d = (\\MaskQTree_src_d [0] && (! \\MaskQTree_src_emitted [1]));
  assign \\MaskQTree_src_done  = (\\MaskQTree_src_emitted  | ({go_2_dummy_write_MaskQTree_d[0],
                                                               go_1_dummy_write_MaskQTree_d[0]} & {go_2_dummy_write_MaskQTree_r,
                                                                                                   go_1_dummy_write_MaskQTree_r}));
  assign \\MaskQTree_src_r  = (& \\MaskQTree_src_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \\MaskQTree_src_emitted  <= 2'd0;
    else
      \\MaskQTree_src_emitted  <= (\\MaskQTree_src_r  ? 2'd0 :
                                   \\MaskQTree_src_done );
  
  /* source (Ty MaskQTree) : > (dummy_write_MaskQTree,MaskQTree) */
  
  /* sink (Ty Pointer_MaskQTree) : (dummy_write_MaskQTree_sink,Pointer_MaskQTree) > */
  assign {dummy_write_MaskQTree_sink_r,
          dummy_write_MaskQTree_sink_dout} = {dummy_write_MaskQTree_sink_rout,
                                              dummy_write_MaskQTree_sink_d};
  
  /* fork (Ty Word16#) : (mergeHP_MaskQTree_buf,Word16#) > [(forkHP1_MaskQTree,Word16#),
                                                       (forkHP1_MaskQTree_snk,Word16#),
                                                       (forkHP1_MaskQTre3,Word16#),
                                                       (forkHP1_MaskQTre4,Word16#)] */
  logic [3:0] mergeHP_MaskQTree_buf_emitted;
  logic [3:0] mergeHP_MaskQTree_buf_done;
  assign forkHP1_MaskQTree_d = {mergeHP_MaskQTree_buf_d[16:1],
                                (mergeHP_MaskQTree_buf_d[0] && (! mergeHP_MaskQTree_buf_emitted[0]))};
  assign forkHP1_MaskQTree_snk_d = {mergeHP_MaskQTree_buf_d[16:1],
                                    (mergeHP_MaskQTree_buf_d[0] && (! mergeHP_MaskQTree_buf_emitted[1]))};
  assign forkHP1_MaskQTre3_d = {mergeHP_MaskQTree_buf_d[16:1],
                                (mergeHP_MaskQTree_buf_d[0] && (! mergeHP_MaskQTree_buf_emitted[2]))};
  assign forkHP1_MaskQTre4_d = {mergeHP_MaskQTree_buf_d[16:1],
                                (mergeHP_MaskQTree_buf_d[0] && (! mergeHP_MaskQTree_buf_emitted[3]))};
  assign mergeHP_MaskQTree_buf_done = (mergeHP_MaskQTree_buf_emitted | ({forkHP1_MaskQTre4_d[0],
                                                                         forkHP1_MaskQTre3_d[0],
                                                                         forkHP1_MaskQTree_snk_d[0],
                                                                         forkHP1_MaskQTree_d[0]} & {forkHP1_MaskQTre4_r,
                                                                                                    forkHP1_MaskQTre3_r,
                                                                                                    forkHP1_MaskQTree_snk_r,
                                                                                                    forkHP1_MaskQTree_r}));
  assign mergeHP_MaskQTree_buf_r = (& mergeHP_MaskQTree_buf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_MaskQTree_buf_emitted <= 4'd0;
    else
      mergeHP_MaskQTree_buf_emitted <= (mergeHP_MaskQTree_buf_r ? 4'd0 :
                                        mergeHP_MaskQTree_buf_done);
  
  /* mergectrl (Ty C2,
           Ty MemIn_MaskQTree) : [(dconReadIn_MaskQTree,MemIn_MaskQTree),
                                  (dconWriteIn_MaskQTree,MemIn_MaskQTree)] > (memMergeChoice_MaskQTree,C2) (memMergeIn_MaskQTree,MemIn_MaskQTree) */
  logic [1:0] dconReadIn_MaskQTree_select_d;
  assign dconReadIn_MaskQTree_select_d = ((| dconReadIn_MaskQTree_select_q) ? dconReadIn_MaskQTree_select_q :
                                          (dconReadIn_MaskQTree_d[0] ? 2'd1 :
                                           (dconWriteIn_MaskQTree_d[0] ? 2'd2 :
                                            2'd0)));
  logic [1:0] dconReadIn_MaskQTree_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) dconReadIn_MaskQTree_select_q <= 2'd0;
    else
      dconReadIn_MaskQTree_select_q <= (dconReadIn_MaskQTree_done ? 2'd0 :
                                        dconReadIn_MaskQTree_select_d);
  logic [1:0] dconReadIn_MaskQTree_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) dconReadIn_MaskQTree_emit_q <= 2'd0;
    else
      dconReadIn_MaskQTree_emit_q <= (dconReadIn_MaskQTree_done ? 2'd0 :
                                      dconReadIn_MaskQTree_emit_d);
  logic [1:0] dconReadIn_MaskQTree_emit_d;
  assign dconReadIn_MaskQTree_emit_d = (dconReadIn_MaskQTree_emit_q | ({memMergeChoice_MaskQTree_d[0],
                                                                        memMergeIn_MaskQTree_d[0]} & {memMergeChoice_MaskQTree_r,
                                                                                                      memMergeIn_MaskQTree_r}));
  logic dconReadIn_MaskQTree_done;
  assign dconReadIn_MaskQTree_done = (& dconReadIn_MaskQTree_emit_d);
  assign {dconWriteIn_MaskQTree_r,
          dconReadIn_MaskQTree_r} = (dconReadIn_MaskQTree_done ? dconReadIn_MaskQTree_select_d :
                                     2'd0);
  assign memMergeIn_MaskQTree_d = ((dconReadIn_MaskQTree_select_d[0] && (! dconReadIn_MaskQTree_emit_q[0])) ? dconReadIn_MaskQTree_d :
                                   ((dconReadIn_MaskQTree_select_d[1] && (! dconReadIn_MaskQTree_emit_q[0])) ? dconWriteIn_MaskQTree_d :
                                    {83'd0, 1'd0}));
  assign memMergeChoice_MaskQTree_d = ((dconReadIn_MaskQTree_select_d[0] && (! dconReadIn_MaskQTree_emit_q[1])) ? C1_2_dc(1'd1) :
                                       ((dconReadIn_MaskQTree_select_d[1] && (! dconReadIn_MaskQTree_emit_q[1])) ? C2_2_dc(1'd1) :
                                        {1'd0, 1'd0}));
  
  /* bram (Ty MemIn_MaskQTree,
      Ty MemOut_MaskQTree) : (memMergeIn_MaskQTree_dbuf,MemIn_MaskQTree) > (memOut_MaskQTree,MemOut_MaskQTree) */
  logic [65:0] memMergeIn_MaskQTree_dbuf_mem[65535:0];
  logic [15:0] memMergeIn_MaskQTree_dbuf_address;
  logic [65:0] memMergeIn_MaskQTree_dbuf_din;
  logic [65:0] memOut_MaskQTree_q;
  logic memOut_MaskQTree_valid;
  logic memMergeIn_MaskQTree_dbuf_we;
  logic memOut_MaskQTree_we;
  assign memMergeIn_MaskQTree_dbuf_din = memMergeIn_MaskQTree_dbuf_d[83:18];
  assign memMergeIn_MaskQTree_dbuf_address = memMergeIn_MaskQTree_dbuf_d[17:2];
  assign memMergeIn_MaskQTree_dbuf_we = (memMergeIn_MaskQTree_dbuf_d[1:1] && memMergeIn_MaskQTree_dbuf_d[0]);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        memOut_MaskQTree_we <= 1'd0;
        memOut_MaskQTree_valid <= 1'd0;
      end
    else
      begin
        memOut_MaskQTree_we <= memMergeIn_MaskQTree_dbuf_we;
        memOut_MaskQTree_valid <= memMergeIn_MaskQTree_dbuf_d[0];
        if (memMergeIn_MaskQTree_dbuf_we)
          begin
            memMergeIn_MaskQTree_dbuf_mem[memMergeIn_MaskQTree_dbuf_address] <= memMergeIn_MaskQTree_dbuf_din;
            memOut_MaskQTree_q <= memMergeIn_MaskQTree_dbuf_din;
          end
        else
          memOut_MaskQTree_q <= memMergeIn_MaskQTree_dbuf_mem[memMergeIn_MaskQTree_dbuf_address];
      end
  assign memOut_MaskQTree_d = {memOut_MaskQTree_q,
                               memOut_MaskQTree_we,
                               memOut_MaskQTree_valid};
  assign memMergeIn_MaskQTree_dbuf_r = ((! memOut_MaskQTree_valid) || memOut_MaskQTree_r);
  
  /* demux (Ty C2,
       Ty MemOut_MaskQTree) : (memMergeChoice_MaskQTree,C2) (memOut_MaskQTree_dbuf,MemOut_MaskQTree) > [(memReadOut_MaskQTree,MemOut_MaskQTree),
                                                                                                        (memWriteOut_MaskQTree,MemOut_MaskQTree)] */
  logic [1:0] memOut_MaskQTree_dbuf_onehotd;
  always_comb
    if ((memMergeChoice_MaskQTree_d[0] && memOut_MaskQTree_dbuf_d[0]))
      unique case (memMergeChoice_MaskQTree_d[1:1])
        1'd0: memOut_MaskQTree_dbuf_onehotd = 2'd1;
        1'd1: memOut_MaskQTree_dbuf_onehotd = 2'd2;
        default: memOut_MaskQTree_dbuf_onehotd = 2'd0;
      endcase
    else memOut_MaskQTree_dbuf_onehotd = 2'd0;
  assign memReadOut_MaskQTree_d = {memOut_MaskQTree_dbuf_d[67:1],
                                   memOut_MaskQTree_dbuf_onehotd[0]};
  assign memWriteOut_MaskQTree_d = {memOut_MaskQTree_dbuf_d[67:1],
                                    memOut_MaskQTree_dbuf_onehotd[1]};
  assign memOut_MaskQTree_dbuf_r = (| (memOut_MaskQTree_dbuf_onehotd & {memWriteOut_MaskQTree_r,
                                                                        memReadOut_MaskQTree_r}));
  assign memMergeChoice_MaskQTree_r = memOut_MaskQTree_dbuf_r;
  
  /* dbuf (Ty MemIn_MaskQTree) : (memMergeIn_MaskQTree_rbuf,MemIn_MaskQTree) > (memMergeIn_MaskQTree_dbuf,MemIn_MaskQTree) */
  assign memMergeIn_MaskQTree_rbuf_r = ((! memMergeIn_MaskQTree_dbuf_d[0]) || memMergeIn_MaskQTree_dbuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memMergeIn_MaskQTree_dbuf_d <= {83'd0, 1'd0};
    else
      if (memMergeIn_MaskQTree_rbuf_r)
        memMergeIn_MaskQTree_dbuf_d <= memMergeIn_MaskQTree_rbuf_d;
  
  /* rbuf (Ty MemIn_MaskQTree) : (memMergeIn_MaskQTree,MemIn_MaskQTree) > (memMergeIn_MaskQTree_rbuf,MemIn_MaskQTree) */
  MemIn_MaskQTree_t memMergeIn_MaskQTree_buf;
  assign memMergeIn_MaskQTree_r = (! memMergeIn_MaskQTree_buf[0]);
  assign memMergeIn_MaskQTree_rbuf_d = (memMergeIn_MaskQTree_buf[0] ? memMergeIn_MaskQTree_buf :
                                        memMergeIn_MaskQTree_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memMergeIn_MaskQTree_buf <= {83'd0, 1'd0};
    else
      if ((memMergeIn_MaskQTree_rbuf_r && memMergeIn_MaskQTree_buf[0]))
        memMergeIn_MaskQTree_buf <= {83'd0, 1'd0};
      else if (((! memMergeIn_MaskQTree_rbuf_r) && (! memMergeIn_MaskQTree_buf[0])))
        memMergeIn_MaskQTree_buf <= memMergeIn_MaskQTree_d;
  
  /* dbuf (Ty MemOut_MaskQTree) : (memOut_MaskQTree_rbuf,MemOut_MaskQTree) > (memOut_MaskQTree_dbuf,MemOut_MaskQTree) */
  assign memOut_MaskQTree_rbuf_r = ((! memOut_MaskQTree_dbuf_d[0]) || memOut_MaskQTree_dbuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memOut_MaskQTree_dbuf_d <= {67'd0, 1'd0};
    else
      if (memOut_MaskQTree_rbuf_r)
        memOut_MaskQTree_dbuf_d <= memOut_MaskQTree_rbuf_d;
  
  /* rbuf (Ty MemOut_MaskQTree) : (memOut_MaskQTree,MemOut_MaskQTree) > (memOut_MaskQTree_rbuf,MemOut_MaskQTree) */
  MemOut_MaskQTree_t memOut_MaskQTree_buf;
  assign memOut_MaskQTree_r = (! memOut_MaskQTree_buf[0]);
  assign memOut_MaskQTree_rbuf_d = (memOut_MaskQTree_buf[0] ? memOut_MaskQTree_buf :
                                    memOut_MaskQTree_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memOut_MaskQTree_buf <= {67'd0, 1'd0};
    else
      if ((memOut_MaskQTree_rbuf_r && memOut_MaskQTree_buf[0]))
        memOut_MaskQTree_buf <= {67'd0, 1'd0};
      else if (((! memOut_MaskQTree_rbuf_r) && (! memOut_MaskQTree_buf[0])))
        memOut_MaskQTree_buf <= memOut_MaskQTree_d;
  
  /* destruct (Ty Pointer_MaskQTree,
          Dcon Pointer_MaskQTree) : (mska8r_1_argbuf,Pointer_MaskQTree) > [(destructReadIn_MaskQTree,Word16#)] */
  assign destructReadIn_MaskQTree_d = {mska8r_1_argbuf_d[16:1],
                                       mska8r_1_argbuf_d[0]};
  assign mska8r_1_argbuf_r = destructReadIn_MaskQTree_r;
  
  /* dcon (Ty MemIn_MaskQTree,
      Dcon ReadIn_MaskQTree) : [(destructReadIn_MaskQTree,Word16#)] > (dconReadIn_MaskQTree,MemIn_MaskQTree) */
  assign dconReadIn_MaskQTree_d = ReadIn_MaskQTree_dc((& {destructReadIn_MaskQTree_d[0]}), destructReadIn_MaskQTree_d);
  assign {destructReadIn_MaskQTree_r} = {1 {(dconReadIn_MaskQTree_r && dconReadIn_MaskQTree_d[0])}};
  
  /* destruct (Ty MemOut_MaskQTree,
          Dcon ReadOut_MaskQTree) : (memReadOut_MaskQTree,MemOut_MaskQTree) > [(readPointer_MaskQTreemska8r_1_argbuf,MaskQTree)] */
  assign readPointer_MaskQTreemska8r_1_argbuf_d = {memReadOut_MaskQTree_d[67:2],
                                                   memReadOut_MaskQTree_d[0]};
  assign memReadOut_MaskQTree_r = readPointer_MaskQTreemska8r_1_argbuf_r;
  
  /* dcon (Ty MemIn_MaskQTree,
      Dcon WriteIn_MaskQTree) : [(forkHP1_MaskQTre3,Word16#),
                                 (dummy_write_MaskQTree,MaskQTree)] > (dconWriteIn_MaskQTree,MemIn_MaskQTree) */
  assign dconWriteIn_MaskQTree_d = WriteIn_MaskQTree_dc((& {forkHP1_MaskQTre3_d[0],
                                                            dummy_write_MaskQTree_d[0]}), forkHP1_MaskQTre3_d, dummy_write_MaskQTree_d);
  assign {forkHP1_MaskQTre3_r,
          dummy_write_MaskQTree_r} = {2 {(dconWriteIn_MaskQTree_r && dconWriteIn_MaskQTree_d[0])}};
  
  /* dcon (Ty Pointer_MaskQTree,
      Dcon Pointer_MaskQTree) : [(forkHP1_MaskQTre4,Word16#)] > (dconPtr_MaskQTree,Pointer_MaskQTree) */
  assign dconPtr_MaskQTree_d = Pointer_MaskQTree_dc((& {forkHP1_MaskQTre4_d[0]}), forkHP1_MaskQTre4_d);
  assign {forkHP1_MaskQTre4_r} = {1 {(dconPtr_MaskQTree_r && dconPtr_MaskQTree_d[0])}};
  
  /* demux (Ty MemOut_MaskQTree,
       Ty Pointer_MaskQTree) : (memWriteOut_MaskQTree,MemOut_MaskQTree) (dconPtr_MaskQTree,Pointer_MaskQTree) > [(_74,Pointer_MaskQTree),
                                                                                                                 (dummy_write_MaskQTree_sink,Pointer_MaskQTree)] */
  logic [1:0] dconPtr_MaskQTree_onehotd;
  always_comb
    if ((memWriteOut_MaskQTree_d[0] && dconPtr_MaskQTree_d[0]))
      unique case (memWriteOut_MaskQTree_d[1:1])
        1'd0: dconPtr_MaskQTree_onehotd = 2'd1;
        1'd1: dconPtr_MaskQTree_onehotd = 2'd2;
        default: dconPtr_MaskQTree_onehotd = 2'd0;
      endcase
    else dconPtr_MaskQTree_onehotd = 2'd0;
  assign _74_d = {dconPtr_MaskQTree_d[16:1],
                  dconPtr_MaskQTree_onehotd[0]};
  assign dummy_write_MaskQTree_sink_d = {dconPtr_MaskQTree_d[16:1],
                                         dconPtr_MaskQTree_onehotd[1]};
  assign dconPtr_MaskQTree_r = (| (dconPtr_MaskQTree_onehotd & {dummy_write_MaskQTree_sink_r,
                                                                _74_r}));
  assign memWriteOut_MaskQTree_r = dconPtr_MaskQTree_r;
  
  /* source (Ty Go) : > (sourceGo,Go) */
  
  /* source (Ty Pointer_MaskQTree) : > (m1a92_0,Pointer_MaskQTree) */
  
  /* source (Ty Pointer_QTree_Int) : > (m2a93_1,Pointer_QTree_Int) */
  
  /* source (Ty Pointer_QTree_Int) : > (m3a94_2,Pointer_QTree_Int) */
  
  /* destruct (Ty TupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int,
          Dcon TupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int) : ($wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1,TupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int) > [($wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgo_4,Go),
                                                                                                                                                                                                                                   ($wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intwsie,MyDTInt_Int_Int),
                                                                                                                                                                                                                                   ($wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw1sif,Pointer_QTree_Int),
                                                                                                                                                                                                                                   ($wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw2sig,Pointer_QTree_Int)] */
  logic [3:0] \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1_emitted ;
  logic [3:0] \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1_done ;
  assign \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgo_4_d  = (\$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1_d [0] && (! \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1_emitted [0]));
  assign \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intwsie_d  = (\$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1_d [0] && (! \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1_emitted [1]));
  assign \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw1sif_d  = {\$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1_d [16:1],
                                                                                               (\$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1_d [0] && (! \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1_emitted [2]))};
  assign \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw2sig_d  = {\$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1_d [32:17],
                                                                                               (\$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1_d [0] && (! \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1_emitted [3]))};
  assign \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1_done  = (\$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1_emitted  | ({\$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw2sig_d [0],
                                                                                                                                                                                         \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw1sif_d [0],
                                                                                                                                                                                         \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intwsie_d [0],
                                                                                                                                                                                         \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgo_4_d [0]} & {\$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw2sig_r ,
                                                                                                                                                                                                                                                                                  \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw1sif_r ,
                                                                                                                                                                                                                                                                                  \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intwsie_r ,
                                                                                                                                                                                                                                                                                  \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgo_4_r }));
  assign \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1_r  = (& \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1_emitted  <= 4'd0;
    else
      \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1_emitted  <= (\$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1_r  ? 4'd0 :
                                                                                                \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1_done );
  
  /* fork (Ty Go) : ($wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgo_4,Go) > [(go_4_1,Go),
                                                                                                     (go_4_2,Go)] */
  logic [1:0] \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgo_4_emitted ;
  logic [1:0] \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgo_4_done ;
  assign go_4_1_d = (\$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgo_4_d [0] && (! \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgo_4_emitted [0]));
  assign go_4_2_d = (\$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgo_4_d [0] && (! \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgo_4_emitted [1]));
  assign \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgo_4_done  = (\$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgo_4_emitted  | ({go_4_2_d[0],
                                                                                                                                                                                             go_4_1_d[0]} & {go_4_2_r,
                                                                                                                                                                                                             go_4_1_r}));
  assign \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgo_4_r  = (& \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgo_4_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgo_4_emitted  <= 2'd0;
    else
      \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgo_4_emitted  <= (\$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgo_4_r  ? 2'd0 :
                                                                                                  \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgo_4_done );
  
  /* buf (Ty Pointer_QTree_Int) : ($wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw1sif,Pointer_QTree_Int) > (w1sif_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw1sif_bufchan_d ;
  logic \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw1sif_bufchan_r ;
  assign \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw1sif_r  = ((! \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw1sif_bufchan_d [0]) || \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw1sif_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw1sif_bufchan_d  <= {16'd0,
                                                                                                     1'd0};
    else
      if (\$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw1sif_r )
        \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw1sif_bufchan_d  <= \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw1sif_d ;
  Pointer_QTree_Int_t \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw1sif_bufchan_buf ;
  assign \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw1sif_bufchan_r  = (! \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw1sif_bufchan_buf [0]);
  assign w1sif_1_argbuf_d = (\$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw1sif_bufchan_buf [0] ? \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw1sif_bufchan_buf  :
                             \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw1sif_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw1sif_bufchan_buf  <= {16'd0,
                                                                                                       1'd0};
    else
      if ((w1sif_1_argbuf_r && \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw1sif_bufchan_buf [0]))
        \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw1sif_bufchan_buf  <= {16'd0,
                                                                                                         1'd0};
      else if (((! w1sif_1_argbuf_r) && (! \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw1sif_bufchan_buf [0])))
        \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw1sif_bufchan_buf  <= \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw1sif_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Int) : ($wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw2sig,Pointer_QTree_Int) > (w2sig_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw2sig_bufchan_d ;
  logic \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw2sig_bufchan_r ;
  assign \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw2sig_r  = ((! \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw2sig_bufchan_d [0]) || \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw2sig_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw2sig_bufchan_d  <= {16'd0,
                                                                                                     1'd0};
    else
      if (\$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw2sig_r )
        \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw2sig_bufchan_d  <= \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw2sig_d ;
  Pointer_QTree_Int_t \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw2sig_bufchan_buf ;
  assign \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw2sig_bufchan_r  = (! \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw2sig_bufchan_buf [0]);
  assign w2sig_1_argbuf_d = (\$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw2sig_bufchan_buf [0] ? \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw2sig_bufchan_buf  :
                             \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw2sig_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw2sig_bufchan_buf  <= {16'd0,
                                                                                                       1'd0};
    else
      if ((w2sig_1_argbuf_r && \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw2sig_bufchan_buf [0]))
        \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw2sig_bufchan_buf  <= {16'd0,
                                                                                                         1'd0};
      else if (((! w2sig_1_argbuf_r) && (! \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw2sig_bufchan_buf [0])))
        \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw2sig_bufchan_buf  <= \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw2sig_bufchan_d ;
  
  /* buf (Ty MyDTInt_Int_Int) : ($wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intwsie,MyDTInt_Int_Int) > (wsie_1_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intwsie_bufchan_d ;
  logic \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intwsie_bufchan_r ;
  assign \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intwsie_r  = ((! \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intwsie_bufchan_d [0]) || \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intwsie_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intwsie_bufchan_d  <= 1'd0;
    else
      if (\$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intwsie_r )
        \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intwsie_bufchan_d  <= \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intwsie_d ;
  MyDTInt_Int_Int_t \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intwsie_bufchan_buf ;
  assign \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intwsie_bufchan_r  = (! \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intwsie_bufchan_buf [0]);
  assign wsie_1_argbuf_d = (\$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intwsie_bufchan_buf [0] ? \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intwsie_bufchan_buf  :
                            \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intwsie_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intwsie_bufchan_buf  <= 1'd0;
    else
      if ((wsie_1_argbuf_r && \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intwsie_bufchan_buf [0]))
        \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intwsie_bufchan_buf  <= 1'd0;
      else if (((! wsie_1_argbuf_r) && (! \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intwsie_bufchan_buf [0])))
        \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intwsie_bufchan_buf  <= \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intwsie_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Int) : ($wmAdd_Int_resbuf,Pointer_QTree_Int) > (es_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t \$wmAdd_Int_resbuf_bufchan_d ;
  logic \$wmAdd_Int_resbuf_bufchan_r ;
  assign \$wmAdd_Int_resbuf_r  = ((! \$wmAdd_Int_resbuf_bufchan_d [0]) || \$wmAdd_Int_resbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \$wmAdd_Int_resbuf_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\$wmAdd_Int_resbuf_r )
        \$wmAdd_Int_resbuf_bufchan_d  <= \$wmAdd_Int_resbuf_d ;
  Pointer_QTree_Int_t \$wmAdd_Int_resbuf_bufchan_buf ;
  assign \$wmAdd_Int_resbuf_bufchan_r  = (! \$wmAdd_Int_resbuf_bufchan_buf [0]);
  assign es_1_1_argbuf_d = (\$wmAdd_Int_resbuf_bufchan_buf [0] ? \$wmAdd_Int_resbuf_bufchan_buf  :
                            \$wmAdd_Int_resbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \$wmAdd_Int_resbuf_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((es_1_1_argbuf_r && \$wmAdd_Int_resbuf_bufchan_buf [0]))
        \$wmAdd_Int_resbuf_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! es_1_1_argbuf_r) && (! \$wmAdd_Int_resbuf_bufchan_buf [0])))
        \$wmAdd_Int_resbuf_bufchan_buf  <= \$wmAdd_Int_resbuf_bufchan_d ;
  
  /* destruct (Ty TupGo___Pointer_QTree_Int,
          Dcon TupGo___Pointer_QTree_Int) : ($wnnz_IntTupGo___Pointer_QTree_Int_1,TupGo___Pointer_QTree_Int) > [($wnnz_IntTupGo___Pointer_QTree_Intgo_5,Go),
                                                                                                                ($wnnz_IntTupGo___Pointer_QTree_Intwsij,Pointer_QTree_Int)] */
  logic [1:0] \$wnnz_IntTupGo___Pointer_QTree_Int_1_emitted ;
  logic [1:0] \$wnnz_IntTupGo___Pointer_QTree_Int_1_done ;
  assign \$wnnz_IntTupGo___Pointer_QTree_Intgo_5_d  = (\$wnnz_IntTupGo___Pointer_QTree_Int_1_d [0] && (! \$wnnz_IntTupGo___Pointer_QTree_Int_1_emitted [0]));
  assign \$wnnz_IntTupGo___Pointer_QTree_Intwsij_d  = {\$wnnz_IntTupGo___Pointer_QTree_Int_1_d [16:1],
                                                       (\$wnnz_IntTupGo___Pointer_QTree_Int_1_d [0] && (! \$wnnz_IntTupGo___Pointer_QTree_Int_1_emitted [1]))};
  assign \$wnnz_IntTupGo___Pointer_QTree_Int_1_done  = (\$wnnz_IntTupGo___Pointer_QTree_Int_1_emitted  | ({\$wnnz_IntTupGo___Pointer_QTree_Intwsij_d [0],
                                                                                                           \$wnnz_IntTupGo___Pointer_QTree_Intgo_5_d [0]} & {\$wnnz_IntTupGo___Pointer_QTree_Intwsij_r ,
                                                                                                                                                             \$wnnz_IntTupGo___Pointer_QTree_Intgo_5_r }));
  assign \$wnnz_IntTupGo___Pointer_QTree_Int_1_r  = (& \$wnnz_IntTupGo___Pointer_QTree_Int_1_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \$wnnz_IntTupGo___Pointer_QTree_Int_1_emitted  <= 2'd0;
    else
      \$wnnz_IntTupGo___Pointer_QTree_Int_1_emitted  <= (\$wnnz_IntTupGo___Pointer_QTree_Int_1_r  ? 2'd0 :
                                                         \$wnnz_IntTupGo___Pointer_QTree_Int_1_done );
  
  /* fork (Ty Go) : ($wnnz_IntTupGo___Pointer_QTree_Intgo_5,Go) > [(go_5_1,Go),
                                                              (go_5_2,Go)] */
  logic [1:0] \$wnnz_IntTupGo___Pointer_QTree_Intgo_5_emitted ;
  logic [1:0] \$wnnz_IntTupGo___Pointer_QTree_Intgo_5_done ;
  assign go_5_1_d = (\$wnnz_IntTupGo___Pointer_QTree_Intgo_5_d [0] && (! \$wnnz_IntTupGo___Pointer_QTree_Intgo_5_emitted [0]));
  assign go_5_2_d = (\$wnnz_IntTupGo___Pointer_QTree_Intgo_5_d [0] && (! \$wnnz_IntTupGo___Pointer_QTree_Intgo_5_emitted [1]));
  assign \$wnnz_IntTupGo___Pointer_QTree_Intgo_5_done  = (\$wnnz_IntTupGo___Pointer_QTree_Intgo_5_emitted  | ({go_5_2_d[0],
                                                                                                               go_5_1_d[0]} & {go_5_2_r,
                                                                                                                               go_5_1_r}));
  assign \$wnnz_IntTupGo___Pointer_QTree_Intgo_5_r  = (& \$wnnz_IntTupGo___Pointer_QTree_Intgo_5_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \$wnnz_IntTupGo___Pointer_QTree_Intgo_5_emitted  <= 2'd0;
    else
      \$wnnz_IntTupGo___Pointer_QTree_Intgo_5_emitted  <= (\$wnnz_IntTupGo___Pointer_QTree_Intgo_5_r  ? 2'd0 :
                                                           \$wnnz_IntTupGo___Pointer_QTree_Intgo_5_done );
  
  /* buf (Ty Pointer_QTree_Int) : ($wnnz_IntTupGo___Pointer_QTree_Intwsij,Pointer_QTree_Int) > (wsij_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t \$wnnz_IntTupGo___Pointer_QTree_Intwsij_bufchan_d ;
  logic \$wnnz_IntTupGo___Pointer_QTree_Intwsij_bufchan_r ;
  assign \$wnnz_IntTupGo___Pointer_QTree_Intwsij_r  = ((! \$wnnz_IntTupGo___Pointer_QTree_Intwsij_bufchan_d [0]) || \$wnnz_IntTupGo___Pointer_QTree_Intwsij_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \$wnnz_IntTupGo___Pointer_QTree_Intwsij_bufchan_d  <= {16'd0,
                                                             1'd0};
    else
      if (\$wnnz_IntTupGo___Pointer_QTree_Intwsij_r )
        \$wnnz_IntTupGo___Pointer_QTree_Intwsij_bufchan_d  <= \$wnnz_IntTupGo___Pointer_QTree_Intwsij_d ;
  Pointer_QTree_Int_t \$wnnz_IntTupGo___Pointer_QTree_Intwsij_bufchan_buf ;
  assign \$wnnz_IntTupGo___Pointer_QTree_Intwsij_bufchan_r  = (! \$wnnz_IntTupGo___Pointer_QTree_Intwsij_bufchan_buf [0]);
  assign wsij_1_argbuf_d = (\$wnnz_IntTupGo___Pointer_QTree_Intwsij_bufchan_buf [0] ? \$wnnz_IntTupGo___Pointer_QTree_Intwsij_bufchan_buf  :
                            \$wnnz_IntTupGo___Pointer_QTree_Intwsij_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \$wnnz_IntTupGo___Pointer_QTree_Intwsij_bufchan_buf  <= {16'd0,
                                                               1'd0};
    else
      if ((wsij_1_argbuf_r && \$wnnz_IntTupGo___Pointer_QTree_Intwsij_bufchan_buf [0]))
        \$wnnz_IntTupGo___Pointer_QTree_Intwsij_bufchan_buf  <= {16'd0,
                                                                 1'd0};
      else if (((! wsij_1_argbuf_r) && (! \$wnnz_IntTupGo___Pointer_QTree_Intwsij_bufchan_buf [0])))
        \$wnnz_IntTupGo___Pointer_QTree_Intwsij_bufchan_buf  <= \$wnnz_IntTupGo___Pointer_QTree_Intwsij_bufchan_d ;
  
  /* dcon (Ty Int,Dcon I#) : [($wnnz_Int_resbuf,Int#)] > (es_6_1I#,Int) */
  assign \es_6_1I#_d  = \I#_dc ((& {\$wnnz_Int_resbuf_d [0]}), \$wnnz_Int_resbuf_d );
  assign {\$wnnz_Int_resbuf_r } = {1 {(\es_6_1I#_r  && \es_6_1I#_d [0])}};
  
  /* destruct (Ty TupMyDTInt_Int_Int___Int___Int,
          Dcon TupMyDTInt_Int_Int___Int___Int) : (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1,TupMyDTInt_Int_Int___Int___Int) > [(applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0,MyDTInt_Int_Int),
                                                                                                                                          (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg2,Int),
                                                                                                                                          (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg1,Int)] */
  logic [2:0] applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_emitted;
  logic [2:0] applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_done;
  assign applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_d = (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_d[0] && (! applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_emitted[0]));
  assign applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg2_d = {applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_d[32:1],
                                                                     (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_d[0] && (! applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_emitted[1]))};
  assign applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg1_d = {applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_d[64:33],
                                                                     (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_d[0] && (! applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_emitted[2]))};
  assign applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_done = (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_emitted | ({applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg1_d[0],
                                                                                                                                       applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg2_d[0],
                                                                                                                                       applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_d[0]} & {applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg1_r,
                                                                                                                                                                                                       applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg2_r,
                                                                                                                                                                                                       applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_r}));
  assign applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_r = (& applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_emitted <= 3'd0;
    else
      applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_emitted <= (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_r ? 3'd0 :
                                                                       applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_done);
  
  /* fork (Ty MyDTInt_Int_Int) : (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0,MyDTInt_Int_Int) > [(arg0_1,MyDTInt_Int_Int),
                                                                                                        (arg0_2,MyDTInt_Int_Int),
                                                                                                        (arg0_3,MyDTInt_Int_Int)] */
  logic [2:0] applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_emitted;
  logic [2:0] applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_done;
  assign arg0_1_d = (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_d[0] && (! applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_emitted[0]));
  assign arg0_2_d = (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_d[0] && (! applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_emitted[1]));
  assign arg0_3_d = (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_d[0] && (! applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_emitted[2]));
  assign applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_done = (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_emitted | ({arg0_3_d[0],
                                                                                                                                           arg0_2_d[0],
                                                                                                                                           arg0_1_d[0]} & {arg0_3_r,
                                                                                                                                                           arg0_2_r,
                                                                                                                                                           arg0_1_r}));
  assign applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_r = (& applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_emitted <= 3'd0;
    else
      applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_emitted <= (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_r ? 3'd0 :
                                                                         applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_done);
  
  /* dcon (Ty QTree_Int,
      Dcon QVal_Int) : [(applyfnInt_Int_Int_5_resbuf,Int)] > (es_0_2_1QVal_Int,QTree_Int) */
  assign es_0_2_1QVal_Int_d = QVal_Int_dc((& {applyfnInt_Int_Int_5_resbuf_d[0]}), applyfnInt_Int_Int_5_resbuf_d);
  assign {applyfnInt_Int_Int_5_resbuf_r} = {1 {(es_0_2_1QVal_Int_r && es_0_2_1QVal_Int_d[0])}};
  
  /* demux (Ty MyDTInt_Int_Int,
       Ty Int) : (arg0_1,MyDTInt_Int_Int) (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg1,Int) > [(arg0_1Dcon_$fNumInt_$c+,Int)] */
  assign \arg0_1Dcon_$fNumInt_$c+_d  = {applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg1_d[32:1],
                                        (arg0_1_d[0] && applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg1_d[0])};
  assign applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg1_r = (\arg0_1Dcon_$fNumInt_$c+_r  && (arg0_1_d[0] && applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg1_d[0]));
  assign arg0_1_r = (\arg0_1Dcon_$fNumInt_$c+_r  && (arg0_1_d[0] && applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg1_d[0]));
  
  /* demux (Ty MyDTInt_Int_Int,
       Ty Int) : (arg0_2,MyDTInt_Int_Int) (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg2,Int) > [(arg0_2Dcon_$fNumInt_$c+,Int)] */
  assign \arg0_2Dcon_$fNumInt_$c+_d  = {applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg2_d[32:1],
                                        (arg0_2_d[0] && applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg2_d[0])};
  assign applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg2_r = (\arg0_2Dcon_$fNumInt_$c+_r  && (arg0_2_d[0] && applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg2_d[0]));
  assign arg0_2_r = (\arg0_2Dcon_$fNumInt_$c+_r  && (arg0_2_d[0] && applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg2_d[0]));
  
  /* fork (Ty Int) : (arg0_2Dcon_$fNumInt_$c+,Int) > [(arg0_2Dcon_$fNumInt_$c+_1,Int),
                                                 (arg0_2Dcon_$fNumInt_$c+_2,Int),
                                                 (arg0_2Dcon_$fNumInt_$c+_3,Int),
                                                 (arg0_2Dcon_$fNumInt_$c+_4,Int)] */
  logic [3:0] \arg0_2Dcon_$fNumInt_$c+_emitted ;
  logic [3:0] \arg0_2Dcon_$fNumInt_$c+_done ;
  assign \arg0_2Dcon_$fNumInt_$c+_1_d  = {\arg0_2Dcon_$fNumInt_$c+_d [32:1],
                                          (\arg0_2Dcon_$fNumInt_$c+_d [0] && (! \arg0_2Dcon_$fNumInt_$c+_emitted [0]))};
  assign \arg0_2Dcon_$fNumInt_$c+_2_d  = {\arg0_2Dcon_$fNumInt_$c+_d [32:1],
                                          (\arg0_2Dcon_$fNumInt_$c+_d [0] && (! \arg0_2Dcon_$fNumInt_$c+_emitted [1]))};
  assign \arg0_2Dcon_$fNumInt_$c+_3_d  = {\arg0_2Dcon_$fNumInt_$c+_d [32:1],
                                          (\arg0_2Dcon_$fNumInt_$c+_d [0] && (! \arg0_2Dcon_$fNumInt_$c+_emitted [2]))};
  assign \arg0_2Dcon_$fNumInt_$c+_4_d  = {\arg0_2Dcon_$fNumInt_$c+_d [32:1],
                                          (\arg0_2Dcon_$fNumInt_$c+_d [0] && (! \arg0_2Dcon_$fNumInt_$c+_emitted [3]))};
  assign \arg0_2Dcon_$fNumInt_$c+_done  = (\arg0_2Dcon_$fNumInt_$c+_emitted  | ({\arg0_2Dcon_$fNumInt_$c+_4_d [0],
                                                                                 \arg0_2Dcon_$fNumInt_$c+_3_d [0],
                                                                                 \arg0_2Dcon_$fNumInt_$c+_2_d [0],
                                                                                 \arg0_2Dcon_$fNumInt_$c+_1_d [0]} & {\arg0_2Dcon_$fNumInt_$c+_4_r ,
                                                                                                                      \arg0_2Dcon_$fNumInt_$c+_3_r ,
                                                                                                                      \arg0_2Dcon_$fNumInt_$c+_2_r ,
                                                                                                                      \arg0_2Dcon_$fNumInt_$c+_1_r }));
  assign \arg0_2Dcon_$fNumInt_$c+_r  = (& \arg0_2Dcon_$fNumInt_$c+_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \arg0_2Dcon_$fNumInt_$c+_emitted  <= 4'd0;
    else
      \arg0_2Dcon_$fNumInt_$c+_emitted  <= (\arg0_2Dcon_$fNumInt_$c+_r  ? 4'd0 :
                                            \arg0_2Dcon_$fNumInt_$c+_done );
  
  /* destruct (Ty Int,
          Dcon I#) : (arg0_2Dcon_$fNumInt_$c+_1I#,Int) > [(xa1lV_destruct,Int#)] */
  assign xa1lV_destruct_d = {\arg0_2Dcon_$fNumInt_$c+_1I#_d [32:1],
                             \arg0_2Dcon_$fNumInt_$c+_1I#_d [0]};
  assign \arg0_2Dcon_$fNumInt_$c+_1I#_r  = xa1lV_destruct_r;
  
  /* demux (Ty Int,
       Ty Int) : (arg0_2Dcon_$fNumInt_$c+_2,Int) (arg0_2Dcon_$fNumInt_$c+_1,Int) > [(arg0_2Dcon_$fNumInt_$c+_1I#,Int)] */
  assign \arg0_2Dcon_$fNumInt_$c+_1I#_d  = {\arg0_2Dcon_$fNumInt_$c+_1_d [32:1],
                                            (\arg0_2Dcon_$fNumInt_$c+_2_d [0] && \arg0_2Dcon_$fNumInt_$c+_1_d [0])};
  assign \arg0_2Dcon_$fNumInt_$c+_1_r  = (\arg0_2Dcon_$fNumInt_$c+_1I#_r  && (\arg0_2Dcon_$fNumInt_$c+_2_d [0] && \arg0_2Dcon_$fNumInt_$c+_1_d [0]));
  assign \arg0_2Dcon_$fNumInt_$c+_2_r  = (\arg0_2Dcon_$fNumInt_$c+_1I#_r  && (\arg0_2Dcon_$fNumInt_$c+_2_d [0] && \arg0_2Dcon_$fNumInt_$c+_1_d [0]));
  
  /* demux (Ty Int,
       Ty Int) : (arg0_2Dcon_$fNumInt_$c+_3,Int) (arg0_1Dcon_$fNumInt_$c+,Int) > [(arg0_2Dcon_$fNumInt_$c+_3I#,Int)] */
  assign \arg0_2Dcon_$fNumInt_$c+_3I#_d  = {\arg0_1Dcon_$fNumInt_$c+_d [32:1],
                                            (\arg0_2Dcon_$fNumInt_$c+_3_d [0] && \arg0_1Dcon_$fNumInt_$c+_d [0])};
  assign \arg0_1Dcon_$fNumInt_$c+_r  = (\arg0_2Dcon_$fNumInt_$c+_3I#_r  && (\arg0_2Dcon_$fNumInt_$c+_3_d [0] && \arg0_1Dcon_$fNumInt_$c+_d [0]));
  assign \arg0_2Dcon_$fNumInt_$c+_3_r  = (\arg0_2Dcon_$fNumInt_$c+_3I#_r  && (\arg0_2Dcon_$fNumInt_$c+_3_d [0] && \arg0_1Dcon_$fNumInt_$c+_d [0]));
  
  /* fork (Ty Int) : (arg0_2Dcon_$fNumInt_$c+_3I#,Int) > [(arg0_2Dcon_$fNumInt_$c+_3I#_1,Int),
                                                     (arg0_2Dcon_$fNumInt_$c+_3I#_2,Int),
                                                     (arg0_2Dcon_$fNumInt_$c+_3I#_3,Int),
                                                     (arg0_2Dcon_$fNumInt_$c+_3I#_4,Int)] */
  logic [3:0] \arg0_2Dcon_$fNumInt_$c+_3I#_emitted ;
  logic [3:0] \arg0_2Dcon_$fNumInt_$c+_3I#_done ;
  assign \arg0_2Dcon_$fNumInt_$c+_3I#_1_d  = {\arg0_2Dcon_$fNumInt_$c+_3I#_d [32:1],
                                              (\arg0_2Dcon_$fNumInt_$c+_3I#_d [0] && (! \arg0_2Dcon_$fNumInt_$c+_3I#_emitted [0]))};
  assign \arg0_2Dcon_$fNumInt_$c+_3I#_2_d  = {\arg0_2Dcon_$fNumInt_$c+_3I#_d [32:1],
                                              (\arg0_2Dcon_$fNumInt_$c+_3I#_d [0] && (! \arg0_2Dcon_$fNumInt_$c+_3I#_emitted [1]))};
  assign \arg0_2Dcon_$fNumInt_$c+_3I#_3_d  = {\arg0_2Dcon_$fNumInt_$c+_3I#_d [32:1],
                                              (\arg0_2Dcon_$fNumInt_$c+_3I#_d [0] && (! \arg0_2Dcon_$fNumInt_$c+_3I#_emitted [2]))};
  assign \arg0_2Dcon_$fNumInt_$c+_3I#_4_d  = {\arg0_2Dcon_$fNumInt_$c+_3I#_d [32:1],
                                              (\arg0_2Dcon_$fNumInt_$c+_3I#_d [0] && (! \arg0_2Dcon_$fNumInt_$c+_3I#_emitted [3]))};
  assign \arg0_2Dcon_$fNumInt_$c+_3I#_done  = (\arg0_2Dcon_$fNumInt_$c+_3I#_emitted  | ({\arg0_2Dcon_$fNumInt_$c+_3I#_4_d [0],
                                                                                         \arg0_2Dcon_$fNumInt_$c+_3I#_3_d [0],
                                                                                         \arg0_2Dcon_$fNumInt_$c+_3I#_2_d [0],
                                                                                         \arg0_2Dcon_$fNumInt_$c+_3I#_1_d [0]} & {\arg0_2Dcon_$fNumInt_$c+_3I#_4_r ,
                                                                                                                                  \arg0_2Dcon_$fNumInt_$c+_3I#_3_r ,
                                                                                                                                  \arg0_2Dcon_$fNumInt_$c+_3I#_2_r ,
                                                                                                                                  \arg0_2Dcon_$fNumInt_$c+_3I#_1_r }));
  assign \arg0_2Dcon_$fNumInt_$c+_3I#_r  = (& \arg0_2Dcon_$fNumInt_$c+_3I#_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \arg0_2Dcon_$fNumInt_$c+_3I#_emitted  <= 4'd0;
    else
      \arg0_2Dcon_$fNumInt_$c+_3I#_emitted  <= (\arg0_2Dcon_$fNumInt_$c+_3I#_r  ? 4'd0 :
                                                \arg0_2Dcon_$fNumInt_$c+_3I#_done );
  
  /* destruct (Ty Int,
          Dcon I#) : (arg0_2Dcon_$fNumInt_$c+_3I#_1I#,Int) > [(ya1lW_destruct,Int#)] */
  assign ya1lW_destruct_d = {\arg0_2Dcon_$fNumInt_$c+_3I#_1I#_d [32:1],
                             \arg0_2Dcon_$fNumInt_$c+_3I#_1I#_d [0]};
  assign \arg0_2Dcon_$fNumInt_$c+_3I#_1I#_r  = ya1lW_destruct_r;
  
  /* demux (Ty Int,
       Ty Int) : (arg0_2Dcon_$fNumInt_$c+_3I#_2,Int) (arg0_2Dcon_$fNumInt_$c+_3I#_1,Int) > [(arg0_2Dcon_$fNumInt_$c+_3I#_1I#,Int)] */
  assign \arg0_2Dcon_$fNumInt_$c+_3I#_1I#_d  = {\arg0_2Dcon_$fNumInt_$c+_3I#_1_d [32:1],
                                                (\arg0_2Dcon_$fNumInt_$c+_3I#_2_d [0] && \arg0_2Dcon_$fNumInt_$c+_3I#_1_d [0])};
  assign \arg0_2Dcon_$fNumInt_$c+_3I#_1_r  = (\arg0_2Dcon_$fNumInt_$c+_3I#_1I#_r  && (\arg0_2Dcon_$fNumInt_$c+_3I#_2_d [0] && \arg0_2Dcon_$fNumInt_$c+_3I#_1_d [0]));
  assign \arg0_2Dcon_$fNumInt_$c+_3I#_2_r  = (\arg0_2Dcon_$fNumInt_$c+_3I#_1I#_r  && (\arg0_2Dcon_$fNumInt_$c+_3I#_2_d [0] && \arg0_2Dcon_$fNumInt_$c+_3I#_1_d [0]));
  
  /* demux (Ty Int,
       Ty Int#) : (arg0_2Dcon_$fNumInt_$c+_3I#_3,Int) (xa1lV_destruct,Int#) > [(arg0_2Dcon_$fNumInt_$c+_3I#_3I#,Int#)] */
  assign \arg0_2Dcon_$fNumInt_$c+_3I#_3I#_d  = {xa1lV_destruct_d[32:1],
                                                (\arg0_2Dcon_$fNumInt_$c+_3I#_3_d [0] && xa1lV_destruct_d[0])};
  assign xa1lV_destruct_r = (\arg0_2Dcon_$fNumInt_$c+_3I#_3I#_r  && (\arg0_2Dcon_$fNumInt_$c+_3I#_3_d [0] && xa1lV_destruct_d[0]));
  assign \arg0_2Dcon_$fNumInt_$c+_3I#_3_r  = (\arg0_2Dcon_$fNumInt_$c+_3I#_3I#_r  && (\arg0_2Dcon_$fNumInt_$c+_3I#_3_d [0] && xa1lV_destruct_d[0]));
  
  /* op_add (Ty Int#) : (arg0_2Dcon_$fNumInt_$c+_3I#_3I#,Int#) (ya1lW_destruct,Int#) > (arg0_2Dcon_$fNumInt_$c+_3I#_3I#_1ya1lW_1_Add32,Int#) */
  assign \arg0_2Dcon_$fNumInt_$c+_3I#_3I#_1ya1lW_1_Add32_d  = {(\arg0_2Dcon_$fNumInt_$c+_3I#_3I#_d [32:1] + ya1lW_destruct_d[32:1]),
                                                               (\arg0_2Dcon_$fNumInt_$c+_3I#_3I#_d [0] && ya1lW_destruct_d[0])};
  assign {\arg0_2Dcon_$fNumInt_$c+_3I#_3I#_r ,
          ya1lW_destruct_r} = {2 {(\arg0_2Dcon_$fNumInt_$c+_3I#_3I#_1ya1lW_1_Add32_r  && \arg0_2Dcon_$fNumInt_$c+_3I#_3I#_1ya1lW_1_Add32_d [0])}};
  
  /* dcon (Ty Int,
      Dcon I#) : [(arg0_2Dcon_$fNumInt_$c+_3I#_3I#_1ya1lW_1_Add32,Int#)] > (es_0_1_1I#,Int) */
  assign \es_0_1_1I#_d  = \I#_dc ((& {\arg0_2Dcon_$fNumInt_$c+_3I#_3I#_1ya1lW_1_Add32_d [0]}), \arg0_2Dcon_$fNumInt_$c+_3I#_3I#_1ya1lW_1_Add32_d );
  assign {\arg0_2Dcon_$fNumInt_$c+_3I#_3I#_1ya1lW_1_Add32_r } = {1 {(\es_0_1_1I#_r  && \es_0_1_1I#_d [0])}};
  
  /* mux (Ty Int,
     Ty Int) : (arg0_2Dcon_$fNumInt_$c+_3I#_4,Int) [(es_0_1_1I#,Int)] > (es_0_1_1I#_mux,Int) */
  assign \es_0_1_1I#_mux_d  = {\es_0_1_1I#_d [32:1],
                               (\arg0_2Dcon_$fNumInt_$c+_3I#_4_d [0] && \es_0_1_1I#_d [0])};
  assign \es_0_1_1I#_r  = (\es_0_1_1I#_mux_r  && (\arg0_2Dcon_$fNumInt_$c+_3I#_4_d [0] && \es_0_1_1I#_d [0]));
  assign \arg0_2Dcon_$fNumInt_$c+_3I#_4_r  = (\es_0_1_1I#_mux_r  && (\arg0_2Dcon_$fNumInt_$c+_3I#_4_d [0] && \es_0_1_1I#_d [0]));
  
  /* mux (Ty Int,
     Ty Int) : (arg0_2Dcon_$fNumInt_$c+_4,Int) [(es_0_1_1I#_mux,Int)] > (es_0_1_1I#_mux_mux,Int) */
  assign \es_0_1_1I#_mux_mux_d  = {\es_0_1_1I#_mux_d [32:1],
                                   (\arg0_2Dcon_$fNumInt_$c+_4_d [0] && \es_0_1_1I#_mux_d [0])};
  assign \es_0_1_1I#_mux_r  = (\es_0_1_1I#_mux_mux_r  && (\arg0_2Dcon_$fNumInt_$c+_4_d [0] && \es_0_1_1I#_mux_d [0]));
  assign \arg0_2Dcon_$fNumInt_$c+_4_r  = (\es_0_1_1I#_mux_mux_r  && (\arg0_2Dcon_$fNumInt_$c+_4_d [0] && \es_0_1_1I#_mux_d [0]));
  
  /* mux (Ty MyDTInt_Int_Int,
     Ty Int) : (arg0_3,MyDTInt_Int_Int) [(es_0_1_1I#_mux_mux,Int)] > (es_0_1_1I#_mux_mux_mux,Int) */
  assign \es_0_1_1I#_mux_mux_mux_d  = {\es_0_1_1I#_mux_mux_d [32:1],
                                       (arg0_3_d[0] && \es_0_1_1I#_mux_mux_d [0])};
  assign \es_0_1_1I#_mux_mux_r  = (\es_0_1_1I#_mux_mux_mux_r  && (arg0_3_d[0] && \es_0_1_1I#_mux_mux_d [0]));
  assign arg0_3_r = (\es_0_1_1I#_mux_mux_mux_r  && (arg0_3_d[0] && \es_0_1_1I#_mux_mux_d [0]));
  
  /* destruct (Ty TupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Int,
          Dcon TupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Int) : (call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Int_1,TupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Int) > [(call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Intgo_6,Go),
                                                                                                                                                                                                                                                                                                             (call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Intwsie_1,MyDTInt_Int_Int),
                                                                                                                                                                                                                                                                                                             (call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Intw1sif_1,Pointer_QTree_Int),
                                                                                                                                                                                                                                                                                                             (call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Intw2sig_1,Pointer_QTree_Int),
                                                                                                                                                                                                                                                                                                             (call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Intsc_0,Pointer_CT$wmAdd_Int)] */
  logic [4:0] call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Int_1_emitted;
  logic [4:0] call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Int_1_done;
  assign call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Intgo_6_d = (call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Int_1_d[0] && (! call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Int_1_emitted[0]));
  assign call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Intwsie_1_d = (call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Int_1_d[0] && (! call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Int_1_emitted[1]));
  assign call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Intw1sif_1_d = {call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Int_1_d[16:1],
                                                                                                                           (call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Int_1_d[0] && (! call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Int_1_emitted[2]))};
  assign call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Intw2sig_1_d = {call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Int_1_d[32:17],
                                                                                                                           (call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Int_1_d[0] && (! call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Int_1_emitted[3]))};
  assign call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Intsc_0_d = {call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Int_1_d[48:33],
                                                                                                                        (call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Int_1_d[0] && (! call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Int_1_emitted[4]))};
  assign call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Int_1_done = (call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Int_1_emitted | ({call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Intsc_0_d[0],
                                                                                                                                                                                                                                             call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Intw2sig_1_d[0],
                                                                                                                                                                                                                                             call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Intw1sif_1_d[0],
                                                                                                                                                                                                                                             call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Intwsie_1_d[0],
                                                                                                                                                                                                                                             call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Intgo_6_d[0]} & {call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Intsc_0_r,
                                                                                                                                                                                                                                                                                                                                                                call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Intw2sig_1_r,
                                                                                                                                                                                                                                                                                                                                                                call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Intw1sif_1_r,
                                                                                                                                                                                                                                                                                                                                                                call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Intwsie_1_r,
                                                                                                                                                                                                                                                                                                                                                                call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Intgo_6_r}));
  assign call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Int_1_r = (& call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Int_1_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Int_1_emitted <= 5'd0;
    else
      call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Int_1_emitted <= (call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Int_1_r ? 5'd0 :
                                                                                                                          call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Int_1_done);
  
  /* rbuf (Ty Go) : (call_$wmAdd_Int_goConst,Go) > (call_$wmAdd_Int_initBufi,Go) */
  Go_t call_$wmAdd_Int_goConst_buf;
  assign call_$wmAdd_Int_goConst_r = (! call_$wmAdd_Int_goConst_buf[0]);
  assign call_$wmAdd_Int_initBufi_d = (call_$wmAdd_Int_goConst_buf[0] ? call_$wmAdd_Int_goConst_buf :
                                       call_$wmAdd_Int_goConst_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_$wmAdd_Int_goConst_buf <= 1'd0;
    else
      if ((call_$wmAdd_Int_initBufi_r && call_$wmAdd_Int_goConst_buf[0]))
        call_$wmAdd_Int_goConst_buf <= 1'd0;
      else if (((! call_$wmAdd_Int_initBufi_r) && (! call_$wmAdd_Int_goConst_buf[0])))
        call_$wmAdd_Int_goConst_buf <= call_$wmAdd_Int_goConst_d;
  
  /* mergectrl (Ty C5,Ty Go) : [(call_$wmAdd_Int_goMux1,Go),
                           (lizzieLet22_3Lcall_$wmAdd_Int3_1_argbuf,Go),
                           (lizzieLet22_3Lcall_$wmAdd_Int2_1_argbuf,Go),
                           (lizzieLet22_3Lcall_$wmAdd_Int1_1_argbuf,Go),
                           (lizzieLet2_4QNode_Int_3QNode_Int_1_argbuf,Go)] > (go_6_goMux_choice,C5) (go_6_goMux_data,Go) */
  logic [4:0] call_$wmAdd_Int_goMux1_select_d;
  assign call_$wmAdd_Int_goMux1_select_d = ((| call_$wmAdd_Int_goMux1_select_q) ? call_$wmAdd_Int_goMux1_select_q :
                                            (call_$wmAdd_Int_goMux1_d[0] ? 5'd1 :
                                             (lizzieLet22_3Lcall_$wmAdd_Int3_1_argbuf_d[0] ? 5'd2 :
                                              (lizzieLet22_3Lcall_$wmAdd_Int2_1_argbuf_d[0] ? 5'd4 :
                                               (lizzieLet22_3Lcall_$wmAdd_Int1_1_argbuf_d[0] ? 5'd8 :
                                                (lizzieLet2_4QNode_Int_3QNode_Int_1_argbuf_d[0] ? 5'd16 :
                                                 5'd0))))));
  logic [4:0] call_$wmAdd_Int_goMux1_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_$wmAdd_Int_goMux1_select_q <= 5'd0;
    else
      call_$wmAdd_Int_goMux1_select_q <= (call_$wmAdd_Int_goMux1_done ? 5'd0 :
                                          call_$wmAdd_Int_goMux1_select_d);
  logic [1:0] call_$wmAdd_Int_goMux1_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_$wmAdd_Int_goMux1_emit_q <= 2'd0;
    else
      call_$wmAdd_Int_goMux1_emit_q <= (call_$wmAdd_Int_goMux1_done ? 2'd0 :
                                        call_$wmAdd_Int_goMux1_emit_d);
  logic [1:0] call_$wmAdd_Int_goMux1_emit_d;
  assign call_$wmAdd_Int_goMux1_emit_d = (call_$wmAdd_Int_goMux1_emit_q | ({go_6_goMux_choice_d[0],
                                                                            go_6_goMux_data_d[0]} & {go_6_goMux_choice_r,
                                                                                                     go_6_goMux_data_r}));
  logic call_$wmAdd_Int_goMux1_done;
  assign call_$wmAdd_Int_goMux1_done = (& call_$wmAdd_Int_goMux1_emit_d);
  assign {lizzieLet2_4QNode_Int_3QNode_Int_1_argbuf_r,
          lizzieLet22_3Lcall_$wmAdd_Int1_1_argbuf_r,
          lizzieLet22_3Lcall_$wmAdd_Int2_1_argbuf_r,
          lizzieLet22_3Lcall_$wmAdd_Int3_1_argbuf_r,
          call_$wmAdd_Int_goMux1_r} = (call_$wmAdd_Int_goMux1_done ? call_$wmAdd_Int_goMux1_select_d :
                                       5'd0);
  assign go_6_goMux_data_d = ((call_$wmAdd_Int_goMux1_select_d[0] && (! call_$wmAdd_Int_goMux1_emit_q[0])) ? call_$wmAdd_Int_goMux1_d :
                              ((call_$wmAdd_Int_goMux1_select_d[1] && (! call_$wmAdd_Int_goMux1_emit_q[0])) ? lizzieLet22_3Lcall_$wmAdd_Int3_1_argbuf_d :
                               ((call_$wmAdd_Int_goMux1_select_d[2] && (! call_$wmAdd_Int_goMux1_emit_q[0])) ? lizzieLet22_3Lcall_$wmAdd_Int2_1_argbuf_d :
                                ((call_$wmAdd_Int_goMux1_select_d[3] && (! call_$wmAdd_Int_goMux1_emit_q[0])) ? lizzieLet22_3Lcall_$wmAdd_Int1_1_argbuf_d :
                                 ((call_$wmAdd_Int_goMux1_select_d[4] && (! call_$wmAdd_Int_goMux1_emit_q[0])) ? lizzieLet2_4QNode_Int_3QNode_Int_1_argbuf_d :
                                  1'd0)))));
  assign go_6_goMux_choice_d = ((call_$wmAdd_Int_goMux1_select_d[0] && (! call_$wmAdd_Int_goMux1_emit_q[1])) ? C1_5_dc(1'd1) :
                                ((call_$wmAdd_Int_goMux1_select_d[1] && (! call_$wmAdd_Int_goMux1_emit_q[1])) ? C2_5_dc(1'd1) :
                                 ((call_$wmAdd_Int_goMux1_select_d[2] && (! call_$wmAdd_Int_goMux1_emit_q[1])) ? C3_5_dc(1'd1) :
                                  ((call_$wmAdd_Int_goMux1_select_d[3] && (! call_$wmAdd_Int_goMux1_emit_q[1])) ? C4_5_dc(1'd1) :
                                   ((call_$wmAdd_Int_goMux1_select_d[4] && (! call_$wmAdd_Int_goMux1_emit_q[1])) ? C5_5_dc(1'd1) :
                                    {3'd0, 1'd0})))));
  
  /* fork (Ty Go) : (call_$wmAdd_Int_initBuf,Go) > [(call_$wmAdd_Int_unlockFork1,Go),
                                               (call_$wmAdd_Int_unlockFork2,Go),
                                               (call_$wmAdd_Int_unlockFork3,Go),
                                               (call_$wmAdd_Int_unlockFork4,Go),
                                               (call_$wmAdd_Int_unlockFork5,Go)] */
  logic [4:0] call_$wmAdd_Int_initBuf_emitted;
  logic [4:0] call_$wmAdd_Int_initBuf_done;
  assign call_$wmAdd_Int_unlockFork1_d = (call_$wmAdd_Int_initBuf_d[0] && (! call_$wmAdd_Int_initBuf_emitted[0]));
  assign call_$wmAdd_Int_unlockFork2_d = (call_$wmAdd_Int_initBuf_d[0] && (! call_$wmAdd_Int_initBuf_emitted[1]));
  assign call_$wmAdd_Int_unlockFork3_d = (call_$wmAdd_Int_initBuf_d[0] && (! call_$wmAdd_Int_initBuf_emitted[2]));
  assign call_$wmAdd_Int_unlockFork4_d = (call_$wmAdd_Int_initBuf_d[0] && (! call_$wmAdd_Int_initBuf_emitted[3]));
  assign call_$wmAdd_Int_unlockFork5_d = (call_$wmAdd_Int_initBuf_d[0] && (! call_$wmAdd_Int_initBuf_emitted[4]));
  assign call_$wmAdd_Int_initBuf_done = (call_$wmAdd_Int_initBuf_emitted | ({call_$wmAdd_Int_unlockFork5_d[0],
                                                                             call_$wmAdd_Int_unlockFork4_d[0],
                                                                             call_$wmAdd_Int_unlockFork3_d[0],
                                                                             call_$wmAdd_Int_unlockFork2_d[0],
                                                                             call_$wmAdd_Int_unlockFork1_d[0]} & {call_$wmAdd_Int_unlockFork5_r,
                                                                                                                  call_$wmAdd_Int_unlockFork4_r,
                                                                                                                  call_$wmAdd_Int_unlockFork3_r,
                                                                                                                  call_$wmAdd_Int_unlockFork2_r,
                                                                                                                  call_$wmAdd_Int_unlockFork1_r}));
  assign call_$wmAdd_Int_initBuf_r = (& call_$wmAdd_Int_initBuf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_$wmAdd_Int_initBuf_emitted <= 5'd0;
    else
      call_$wmAdd_Int_initBuf_emitted <= (call_$wmAdd_Int_initBuf_r ? 5'd0 :
                                          call_$wmAdd_Int_initBuf_done);
  
  /* initbuf (Ty Go,
         Dcon Go) : (call_$wmAdd_Int_initBufi,Go) > (call_$wmAdd_Int_initBuf,Go) */
  assign call_$wmAdd_Int_initBufi_r = ((! call_$wmAdd_Int_initBuf_d[0]) || call_$wmAdd_Int_initBuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_$wmAdd_Int_initBuf_d <= Go_dc(1'd1);
    else
      if (call_$wmAdd_Int_initBufi_r)
        call_$wmAdd_Int_initBuf_d <= call_$wmAdd_Int_initBufi_d;
  
  /* mux (Ty Go,
     Ty Go) : (call_$wmAdd_Int_unlockFork1,Go) [(call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Intgo_6,Go)] > (call_$wmAdd_Int_goMux1,Go) */
  assign call_$wmAdd_Int_goMux1_d = (call_$wmAdd_Int_unlockFork1_d[0] && call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Intgo_6_d[0]);
  assign call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Intgo_6_r = (call_$wmAdd_Int_goMux1_r && (call_$wmAdd_Int_unlockFork1_d[0] && call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Intgo_6_d[0]));
  assign call_$wmAdd_Int_unlockFork1_r = (call_$wmAdd_Int_goMux1_r && (call_$wmAdd_Int_unlockFork1_d[0] && call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Intgo_6_d[0]));
  
  /* mux (Ty Go,
     Ty MyDTInt_Int_Int) : (call_$wmAdd_Int_unlockFork2,Go) [(call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Intwsie_1,MyDTInt_Int_Int)] > (call_$wmAdd_Int_goMux2,MyDTInt_Int_Int) */
  assign call_$wmAdd_Int_goMux2_d = (call_$wmAdd_Int_unlockFork2_d[0] && call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Intwsie_1_d[0]);
  assign call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Intwsie_1_r = (call_$wmAdd_Int_goMux2_r && (call_$wmAdd_Int_unlockFork2_d[0] && call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Intwsie_1_d[0]));
  assign call_$wmAdd_Int_unlockFork2_r = (call_$wmAdd_Int_goMux2_r && (call_$wmAdd_Int_unlockFork2_d[0] && call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Intwsie_1_d[0]));
  
  /* mux (Ty Go,
     Ty Pointer_QTree_Int) : (call_$wmAdd_Int_unlockFork3,Go) [(call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Intw1sif_1,Pointer_QTree_Int)] > (call_$wmAdd_Int_goMux3,Pointer_QTree_Int) */
  assign call_$wmAdd_Int_goMux3_d = {call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Intw1sif_1_d[16:1],
                                     (call_$wmAdd_Int_unlockFork3_d[0] && call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Intw1sif_1_d[0])};
  assign call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Intw1sif_1_r = (call_$wmAdd_Int_goMux3_r && (call_$wmAdd_Int_unlockFork3_d[0] && call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Intw1sif_1_d[0]));
  assign call_$wmAdd_Int_unlockFork3_r = (call_$wmAdd_Int_goMux3_r && (call_$wmAdd_Int_unlockFork3_d[0] && call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Intw1sif_1_d[0]));
  
  /* mux (Ty Go,
     Ty Pointer_QTree_Int) : (call_$wmAdd_Int_unlockFork4,Go) [(call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Intw2sig_1,Pointer_QTree_Int)] > (call_$wmAdd_Int_goMux4,Pointer_QTree_Int) */
  assign call_$wmAdd_Int_goMux4_d = {call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Intw2sig_1_d[16:1],
                                     (call_$wmAdd_Int_unlockFork4_d[0] && call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Intw2sig_1_d[0])};
  assign call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Intw2sig_1_r = (call_$wmAdd_Int_goMux4_r && (call_$wmAdd_Int_unlockFork4_d[0] && call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Intw2sig_1_d[0]));
  assign call_$wmAdd_Int_unlockFork4_r = (call_$wmAdd_Int_goMux4_r && (call_$wmAdd_Int_unlockFork4_d[0] && call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Intw2sig_1_d[0]));
  
  /* mux (Ty Go,
     Ty Pointer_CT$wmAdd_Int) : (call_$wmAdd_Int_unlockFork5,Go) [(call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Intsc_0,Pointer_CT$wmAdd_Int)] > (call_$wmAdd_Int_goMux5,Pointer_CT$wmAdd_Int) */
  assign call_$wmAdd_Int_goMux5_d = {call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Intsc_0_d[16:1],
                                     (call_$wmAdd_Int_unlockFork5_d[0] && call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Intsc_0_d[0])};
  assign call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Intsc_0_r = (call_$wmAdd_Int_goMux5_r && (call_$wmAdd_Int_unlockFork5_d[0] && call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Intsc_0_d[0]));
  assign call_$wmAdd_Int_unlockFork5_r = (call_$wmAdd_Int_goMux5_r && (call_$wmAdd_Int_unlockFork5_d[0] && call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Intsc_0_d[0]));
  
  /* destruct (Ty TupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int,
          Dcon TupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int) : (call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1,TupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int) > [(call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intgo_7,Go),
                                                                                                                                                                                       (call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intwsij_1,Pointer_QTree_Int),
                                                                                                                                                                                       (call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intsc_0_1,Pointer_CT$wnnz_Int)] */
  logic [2:0] call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_emitted;
  logic [2:0] call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_done;
  assign call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intgo_7_d = (call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_d[0] && (! call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_emitted[0]));
  assign call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intwsij_1_d = {call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_d[16:1],
                                                                                  (call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_d[0] && (! call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_emitted[1]))};
  assign call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intsc_0_1_d = {call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_d[32:17],
                                                                                  (call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_d[0] && (! call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_emitted[2]))};
  assign call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_done = (call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_emitted | ({call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intsc_0_1_d[0],
                                                                                                                                                             call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intwsij_1_d[0],
                                                                                                                                                             call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intgo_7_d[0]} & {call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intsc_0_1_r,
                                                                                                                                                                                                                                        call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intwsij_1_r,
                                                                                                                                                                                                                                        call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intgo_7_r}));
  assign call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_r = (& call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_emitted <= 3'd0;
    else
      call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_emitted <= (call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_r ? 3'd0 :
                                                                                  call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_done);
  
  /* rbuf (Ty Go) : (call_$wnnz_Int_goConst,Go) > (call_$wnnz_Int_initBufi,Go) */
  Go_t call_$wnnz_Int_goConst_buf;
  assign call_$wnnz_Int_goConst_r = (! call_$wnnz_Int_goConst_buf[0]);
  assign call_$wnnz_Int_initBufi_d = (call_$wnnz_Int_goConst_buf[0] ? call_$wnnz_Int_goConst_buf :
                                      call_$wnnz_Int_goConst_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_$wnnz_Int_goConst_buf <= 1'd0;
    else
      if ((call_$wnnz_Int_initBufi_r && call_$wnnz_Int_goConst_buf[0]))
        call_$wnnz_Int_goConst_buf <= 1'd0;
      else if (((! call_$wnnz_Int_initBufi_r) && (! call_$wnnz_Int_goConst_buf[0])))
        call_$wnnz_Int_goConst_buf <= call_$wnnz_Int_goConst_d;
  
  /* mergectrl (Ty C5,Ty Go) : [(call_$wnnz_Int_goMux1,Go),
                           (lizzieLet27_3Lcall_$wnnz_Int3_1_argbuf,Go),
                           (lizzieLet27_3Lcall_$wnnz_Int2_1_argbuf,Go),
                           (lizzieLet27_3Lcall_$wnnz_Int1_1_argbuf,Go),
                           (lizzieLet12_1_3QNode_Int_1_argbuf,Go)] > (go_7_goMux_choice,C5) (go_7_goMux_data,Go) */
  logic [4:0] call_$wnnz_Int_goMux1_select_d;
  assign call_$wnnz_Int_goMux1_select_d = ((| call_$wnnz_Int_goMux1_select_q) ? call_$wnnz_Int_goMux1_select_q :
                                           (call_$wnnz_Int_goMux1_d[0] ? 5'd1 :
                                            (lizzieLet27_3Lcall_$wnnz_Int3_1_argbuf_d[0] ? 5'd2 :
                                             (lizzieLet27_3Lcall_$wnnz_Int2_1_argbuf_d[0] ? 5'd4 :
                                              (lizzieLet27_3Lcall_$wnnz_Int1_1_argbuf_d[0] ? 5'd8 :
                                               (lizzieLet12_1_3QNode_Int_1_argbuf_d[0] ? 5'd16 :
                                                5'd0))))));
  logic [4:0] call_$wnnz_Int_goMux1_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_$wnnz_Int_goMux1_select_q <= 5'd0;
    else
      call_$wnnz_Int_goMux1_select_q <= (call_$wnnz_Int_goMux1_done ? 5'd0 :
                                         call_$wnnz_Int_goMux1_select_d);
  logic [1:0] call_$wnnz_Int_goMux1_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_$wnnz_Int_goMux1_emit_q <= 2'd0;
    else
      call_$wnnz_Int_goMux1_emit_q <= (call_$wnnz_Int_goMux1_done ? 2'd0 :
                                       call_$wnnz_Int_goMux1_emit_d);
  logic [1:0] call_$wnnz_Int_goMux1_emit_d;
  assign call_$wnnz_Int_goMux1_emit_d = (call_$wnnz_Int_goMux1_emit_q | ({go_7_goMux_choice_d[0],
                                                                          go_7_goMux_data_d[0]} & {go_7_goMux_choice_r,
                                                                                                   go_7_goMux_data_r}));
  logic call_$wnnz_Int_goMux1_done;
  assign call_$wnnz_Int_goMux1_done = (& call_$wnnz_Int_goMux1_emit_d);
  assign {lizzieLet12_1_3QNode_Int_1_argbuf_r,
          lizzieLet27_3Lcall_$wnnz_Int1_1_argbuf_r,
          lizzieLet27_3Lcall_$wnnz_Int2_1_argbuf_r,
          lizzieLet27_3Lcall_$wnnz_Int3_1_argbuf_r,
          call_$wnnz_Int_goMux1_r} = (call_$wnnz_Int_goMux1_done ? call_$wnnz_Int_goMux1_select_d :
                                      5'd0);
  assign go_7_goMux_data_d = ((call_$wnnz_Int_goMux1_select_d[0] && (! call_$wnnz_Int_goMux1_emit_q[0])) ? call_$wnnz_Int_goMux1_d :
                              ((call_$wnnz_Int_goMux1_select_d[1] && (! call_$wnnz_Int_goMux1_emit_q[0])) ? lizzieLet27_3Lcall_$wnnz_Int3_1_argbuf_d :
                               ((call_$wnnz_Int_goMux1_select_d[2] && (! call_$wnnz_Int_goMux1_emit_q[0])) ? lizzieLet27_3Lcall_$wnnz_Int2_1_argbuf_d :
                                ((call_$wnnz_Int_goMux1_select_d[3] && (! call_$wnnz_Int_goMux1_emit_q[0])) ? lizzieLet27_3Lcall_$wnnz_Int1_1_argbuf_d :
                                 ((call_$wnnz_Int_goMux1_select_d[4] && (! call_$wnnz_Int_goMux1_emit_q[0])) ? lizzieLet12_1_3QNode_Int_1_argbuf_d :
                                  1'd0)))));
  assign go_7_goMux_choice_d = ((call_$wnnz_Int_goMux1_select_d[0] && (! call_$wnnz_Int_goMux1_emit_q[1])) ? C1_5_dc(1'd1) :
                                ((call_$wnnz_Int_goMux1_select_d[1] && (! call_$wnnz_Int_goMux1_emit_q[1])) ? C2_5_dc(1'd1) :
                                 ((call_$wnnz_Int_goMux1_select_d[2] && (! call_$wnnz_Int_goMux1_emit_q[1])) ? C3_5_dc(1'd1) :
                                  ((call_$wnnz_Int_goMux1_select_d[3] && (! call_$wnnz_Int_goMux1_emit_q[1])) ? C4_5_dc(1'd1) :
                                   ((call_$wnnz_Int_goMux1_select_d[4] && (! call_$wnnz_Int_goMux1_emit_q[1])) ? C5_5_dc(1'd1) :
                                    {3'd0, 1'd0})))));
  
  /* fork (Ty Go) : (call_$wnnz_Int_initBuf,Go) > [(call_$wnnz_Int_unlockFork1,Go),
                                              (call_$wnnz_Int_unlockFork2,Go),
                                              (call_$wnnz_Int_unlockFork3,Go)] */
  logic [2:0] call_$wnnz_Int_initBuf_emitted;
  logic [2:0] call_$wnnz_Int_initBuf_done;
  assign call_$wnnz_Int_unlockFork1_d = (call_$wnnz_Int_initBuf_d[0] && (! call_$wnnz_Int_initBuf_emitted[0]));
  assign call_$wnnz_Int_unlockFork2_d = (call_$wnnz_Int_initBuf_d[0] && (! call_$wnnz_Int_initBuf_emitted[1]));
  assign call_$wnnz_Int_unlockFork3_d = (call_$wnnz_Int_initBuf_d[0] && (! call_$wnnz_Int_initBuf_emitted[2]));
  assign call_$wnnz_Int_initBuf_done = (call_$wnnz_Int_initBuf_emitted | ({call_$wnnz_Int_unlockFork3_d[0],
                                                                           call_$wnnz_Int_unlockFork2_d[0],
                                                                           call_$wnnz_Int_unlockFork1_d[0]} & {call_$wnnz_Int_unlockFork3_r,
                                                                                                               call_$wnnz_Int_unlockFork2_r,
                                                                                                               call_$wnnz_Int_unlockFork1_r}));
  assign call_$wnnz_Int_initBuf_r = (& call_$wnnz_Int_initBuf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_$wnnz_Int_initBuf_emitted <= 3'd0;
    else
      call_$wnnz_Int_initBuf_emitted <= (call_$wnnz_Int_initBuf_r ? 3'd0 :
                                         call_$wnnz_Int_initBuf_done);
  
  /* initbuf (Ty Go,
         Dcon Go) : (call_$wnnz_Int_initBufi,Go) > (call_$wnnz_Int_initBuf,Go) */
  assign call_$wnnz_Int_initBufi_r = ((! call_$wnnz_Int_initBuf_d[0]) || call_$wnnz_Int_initBuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_$wnnz_Int_initBuf_d <= Go_dc(1'd1);
    else
      if (call_$wnnz_Int_initBufi_r)
        call_$wnnz_Int_initBuf_d <= call_$wnnz_Int_initBufi_d;
  
  /* mux (Ty Go,
     Ty Go) : (call_$wnnz_Int_unlockFork1,Go) [(call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intgo_7,Go)] > (call_$wnnz_Int_goMux1,Go) */
  assign call_$wnnz_Int_goMux1_d = (call_$wnnz_Int_unlockFork1_d[0] && call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intgo_7_d[0]);
  assign call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intgo_7_r = (call_$wnnz_Int_goMux1_r && (call_$wnnz_Int_unlockFork1_d[0] && call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intgo_7_d[0]));
  assign call_$wnnz_Int_unlockFork1_r = (call_$wnnz_Int_goMux1_r && (call_$wnnz_Int_unlockFork1_d[0] && call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intgo_7_d[0]));
  
  /* mux (Ty Go,
     Ty Pointer_QTree_Int) : (call_$wnnz_Int_unlockFork2,Go) [(call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intwsij_1,Pointer_QTree_Int)] > (call_$wnnz_Int_goMux2,Pointer_QTree_Int) */
  assign call_$wnnz_Int_goMux2_d = {call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intwsij_1_d[16:1],
                                    (call_$wnnz_Int_unlockFork2_d[0] && call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intwsij_1_d[0])};
  assign call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intwsij_1_r = (call_$wnnz_Int_goMux2_r && (call_$wnnz_Int_unlockFork2_d[0] && call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intwsij_1_d[0]));
  assign call_$wnnz_Int_unlockFork2_r = (call_$wnnz_Int_goMux2_r && (call_$wnnz_Int_unlockFork2_d[0] && call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intwsij_1_d[0]));
  
  /* mux (Ty Go,
     Ty Pointer_CT$wnnz_Int) : (call_$wnnz_Int_unlockFork3,Go) [(call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intsc_0_1,Pointer_CT$wnnz_Int)] > (call_$wnnz_Int_goMux3,Pointer_CT$wnnz_Int) */
  assign call_$wnnz_Int_goMux3_d = {call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intsc_0_1_d[16:1],
                                    (call_$wnnz_Int_unlockFork3_d[0] && call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intsc_0_1_d[0])};
  assign call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intsc_0_1_r = (call_$wnnz_Int_goMux3_r && (call_$wnnz_Int_unlockFork3_d[0] && call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intsc_0_1_d[0]));
  assign call_$wnnz_Int_unlockFork3_r = (call_$wnnz_Int_goMux3_r && (call_$wnnz_Int_unlockFork3_d[0] && call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intsc_0_1_d[0]));
  
  /* destruct (Ty TupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Int,
          Dcon TupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Int) : (call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Int_1,TupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Int) > [(call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Intgo_8,Go),
                                                                                                                                                                                                                                                                   (call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Intma8q,Pointer_QTree_Int),
                                                                                                                                                                                                                                                                   (call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Intmska8r,Pointer_MaskQTree),
                                                                                                                                                                                                                                                                   (call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Intsc_0_2,Pointer_CTmain_mask_Int)] */
  logic [3:0] call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Int_1_emitted;
  logic [3:0] call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Int_1_done;
  assign call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Intgo_8_d = (call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Int_1_d[0] && (! call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Int_1_emitted[0]));
  assign call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Intma8q_d = {call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Int_1_d[16:1],
                                                                                                            (call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Int_1_d[0] && (! call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Int_1_emitted[1]))};
  assign call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Intmska8r_d = {call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Int_1_d[32:17],
                                                                                                              (call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Int_1_d[0] && (! call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Int_1_emitted[2]))};
  assign call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Intsc_0_2_d = {call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Int_1_d[48:33],
                                                                                                              (call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Int_1_d[0] && (! call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Int_1_emitted[3]))};
  assign call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Int_1_done = (call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Int_1_emitted | ({call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Intsc_0_2_d[0],
                                                                                                                                                                                                                     call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Intmska8r_d[0],
                                                                                                                                                                                                                     call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Intma8q_d[0],
                                                                                                                                                                                                                     call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Intgo_8_d[0]} & {call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Intsc_0_2_r,
                                                                                                                                                                                                                                                                                                                            call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Intmska8r_r,
                                                                                                                                                                                                                                                                                                                            call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Intma8q_r,
                                                                                                                                                                                                                                                                                                                            call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Intgo_8_r}));
  assign call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Int_1_r = (& call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Int_1_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Int_1_emitted <= 4'd0;
    else
      call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Int_1_emitted <= (call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Int_1_r ? 4'd0 :
                                                                                                              call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Int_1_done);
  
  /* rbuf (Ty Go) : (call_main_mask_Int_goConst,Go) > (call_main_mask_Int_initBufi,Go) */
  Go_t call_main_mask_Int_goConst_buf;
  assign call_main_mask_Int_goConst_r = (! call_main_mask_Int_goConst_buf[0]);
  assign call_main_mask_Int_initBufi_d = (call_main_mask_Int_goConst_buf[0] ? call_main_mask_Int_goConst_buf :
                                          call_main_mask_Int_goConst_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_main_mask_Int_goConst_buf <= 1'd0;
    else
      if ((call_main_mask_Int_initBufi_r && call_main_mask_Int_goConst_buf[0]))
        call_main_mask_Int_goConst_buf <= 1'd0;
      else if (((! call_main_mask_Int_initBufi_r) && (! call_main_mask_Int_goConst_buf[0])))
        call_main_mask_Int_goConst_buf <= call_main_mask_Int_goConst_d;
  
  /* mergectrl (Ty C5,Ty Go) : [(call_main_mask_Int_goMux1,Go),
                           (lizzieLet31_3Lcall_main_mask_Int3_1_argbuf,Go),
                           (lizzieLet31_3Lcall_main_mask_Int2_1_argbuf,Go),
                           (lizzieLet31_3Lcall_main_mask_Int1_1_argbuf,Go),
                           (lizzieLet14_1_4MQNode_3QNode_Int_1_argbuf,Go)] > (go_8_goMux_choice,C5) (go_8_goMux_data,Go) */
  logic [4:0] call_main_mask_Int_goMux1_select_d;
  assign call_main_mask_Int_goMux1_select_d = ((| call_main_mask_Int_goMux1_select_q) ? call_main_mask_Int_goMux1_select_q :
                                               (call_main_mask_Int_goMux1_d[0] ? 5'd1 :
                                                (lizzieLet31_3Lcall_main_mask_Int3_1_argbuf_d[0] ? 5'd2 :
                                                 (lizzieLet31_3Lcall_main_mask_Int2_1_argbuf_d[0] ? 5'd4 :
                                                  (lizzieLet31_3Lcall_main_mask_Int1_1_argbuf_d[0] ? 5'd8 :
                                                   (lizzieLet14_1_4MQNode_3QNode_Int_1_argbuf_d[0] ? 5'd16 :
                                                    5'd0))))));
  logic [4:0] call_main_mask_Int_goMux1_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_main_mask_Int_goMux1_select_q <= 5'd0;
    else
      call_main_mask_Int_goMux1_select_q <= (call_main_mask_Int_goMux1_done ? 5'd0 :
                                             call_main_mask_Int_goMux1_select_d);
  logic [1:0] call_main_mask_Int_goMux1_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_main_mask_Int_goMux1_emit_q <= 2'd0;
    else
      call_main_mask_Int_goMux1_emit_q <= (call_main_mask_Int_goMux1_done ? 2'd0 :
                                           call_main_mask_Int_goMux1_emit_d);
  logic [1:0] call_main_mask_Int_goMux1_emit_d;
  assign call_main_mask_Int_goMux1_emit_d = (call_main_mask_Int_goMux1_emit_q | ({go_8_goMux_choice_d[0],
                                                                                  go_8_goMux_data_d[0]} & {go_8_goMux_choice_r,
                                                                                                           go_8_goMux_data_r}));
  logic call_main_mask_Int_goMux1_done;
  assign call_main_mask_Int_goMux1_done = (& call_main_mask_Int_goMux1_emit_d);
  assign {lizzieLet14_1_4MQNode_3QNode_Int_1_argbuf_r,
          lizzieLet31_3Lcall_main_mask_Int1_1_argbuf_r,
          lizzieLet31_3Lcall_main_mask_Int2_1_argbuf_r,
          lizzieLet31_3Lcall_main_mask_Int3_1_argbuf_r,
          call_main_mask_Int_goMux1_r} = (call_main_mask_Int_goMux1_done ? call_main_mask_Int_goMux1_select_d :
                                          5'd0);
  assign go_8_goMux_data_d = ((call_main_mask_Int_goMux1_select_d[0] && (! call_main_mask_Int_goMux1_emit_q[0])) ? call_main_mask_Int_goMux1_d :
                              ((call_main_mask_Int_goMux1_select_d[1] && (! call_main_mask_Int_goMux1_emit_q[0])) ? lizzieLet31_3Lcall_main_mask_Int3_1_argbuf_d :
                               ((call_main_mask_Int_goMux1_select_d[2] && (! call_main_mask_Int_goMux1_emit_q[0])) ? lizzieLet31_3Lcall_main_mask_Int2_1_argbuf_d :
                                ((call_main_mask_Int_goMux1_select_d[3] && (! call_main_mask_Int_goMux1_emit_q[0])) ? lizzieLet31_3Lcall_main_mask_Int1_1_argbuf_d :
                                 ((call_main_mask_Int_goMux1_select_d[4] && (! call_main_mask_Int_goMux1_emit_q[0])) ? lizzieLet14_1_4MQNode_3QNode_Int_1_argbuf_d :
                                  1'd0)))));
  assign go_8_goMux_choice_d = ((call_main_mask_Int_goMux1_select_d[0] && (! call_main_mask_Int_goMux1_emit_q[1])) ? C1_5_dc(1'd1) :
                                ((call_main_mask_Int_goMux1_select_d[1] && (! call_main_mask_Int_goMux1_emit_q[1])) ? C2_5_dc(1'd1) :
                                 ((call_main_mask_Int_goMux1_select_d[2] && (! call_main_mask_Int_goMux1_emit_q[1])) ? C3_5_dc(1'd1) :
                                  ((call_main_mask_Int_goMux1_select_d[3] && (! call_main_mask_Int_goMux1_emit_q[1])) ? C4_5_dc(1'd1) :
                                   ((call_main_mask_Int_goMux1_select_d[4] && (! call_main_mask_Int_goMux1_emit_q[1])) ? C5_5_dc(1'd1) :
                                    {3'd0, 1'd0})))));
  
  /* fork (Ty Go) : (call_main_mask_Int_initBuf,Go) > [(call_main_mask_Int_unlockFork1,Go),
                                                  (call_main_mask_Int_unlockFork2,Go),
                                                  (call_main_mask_Int_unlockFork3,Go),
                                                  (call_main_mask_Int_unlockFork4,Go)] */
  logic [3:0] call_main_mask_Int_initBuf_emitted;
  logic [3:0] call_main_mask_Int_initBuf_done;
  assign call_main_mask_Int_unlockFork1_d = (call_main_mask_Int_initBuf_d[0] && (! call_main_mask_Int_initBuf_emitted[0]));
  assign call_main_mask_Int_unlockFork2_d = (call_main_mask_Int_initBuf_d[0] && (! call_main_mask_Int_initBuf_emitted[1]));
  assign call_main_mask_Int_unlockFork3_d = (call_main_mask_Int_initBuf_d[0] && (! call_main_mask_Int_initBuf_emitted[2]));
  assign call_main_mask_Int_unlockFork4_d = (call_main_mask_Int_initBuf_d[0] && (! call_main_mask_Int_initBuf_emitted[3]));
  assign call_main_mask_Int_initBuf_done = (call_main_mask_Int_initBuf_emitted | ({call_main_mask_Int_unlockFork4_d[0],
                                                                                   call_main_mask_Int_unlockFork3_d[0],
                                                                                   call_main_mask_Int_unlockFork2_d[0],
                                                                                   call_main_mask_Int_unlockFork1_d[0]} & {call_main_mask_Int_unlockFork4_r,
                                                                                                                           call_main_mask_Int_unlockFork3_r,
                                                                                                                           call_main_mask_Int_unlockFork2_r,
                                                                                                                           call_main_mask_Int_unlockFork1_r}));
  assign call_main_mask_Int_initBuf_r = (& call_main_mask_Int_initBuf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_main_mask_Int_initBuf_emitted <= 4'd0;
    else
      call_main_mask_Int_initBuf_emitted <= (call_main_mask_Int_initBuf_r ? 4'd0 :
                                             call_main_mask_Int_initBuf_done);
  
  /* initbuf (Ty Go,
         Dcon Go) : (call_main_mask_Int_initBufi,Go) > (call_main_mask_Int_initBuf,Go) */
  assign call_main_mask_Int_initBufi_r = ((! call_main_mask_Int_initBuf_d[0]) || call_main_mask_Int_initBuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_main_mask_Int_initBuf_d <= Go_dc(1'd1);
    else
      if (call_main_mask_Int_initBufi_r)
        call_main_mask_Int_initBuf_d <= call_main_mask_Int_initBufi_d;
  
  /* mux (Ty Go,
     Ty Go) : (call_main_mask_Int_unlockFork1,Go) [(call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Intgo_8,Go)] > (call_main_mask_Int_goMux1,Go) */
  assign call_main_mask_Int_goMux1_d = (call_main_mask_Int_unlockFork1_d[0] && call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Intgo_8_d[0]);
  assign call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Intgo_8_r = (call_main_mask_Int_goMux1_r && (call_main_mask_Int_unlockFork1_d[0] && call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Intgo_8_d[0]));
  assign call_main_mask_Int_unlockFork1_r = (call_main_mask_Int_goMux1_r && (call_main_mask_Int_unlockFork1_d[0] && call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Intgo_8_d[0]));
  
  /* mux (Ty Go,
     Ty Pointer_QTree_Int) : (call_main_mask_Int_unlockFork2,Go) [(call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Intma8q,Pointer_QTree_Int)] > (call_main_mask_Int_goMux2,Pointer_QTree_Int) */
  assign call_main_mask_Int_goMux2_d = {call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Intma8q_d[16:1],
                                        (call_main_mask_Int_unlockFork2_d[0] && call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Intma8q_d[0])};
  assign call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Intma8q_r = (call_main_mask_Int_goMux2_r && (call_main_mask_Int_unlockFork2_d[0] && call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Intma8q_d[0]));
  assign call_main_mask_Int_unlockFork2_r = (call_main_mask_Int_goMux2_r && (call_main_mask_Int_unlockFork2_d[0] && call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Intma8q_d[0]));
  
  /* mux (Ty Go,
     Ty Pointer_MaskQTree) : (call_main_mask_Int_unlockFork3,Go) [(call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Intmska8r,Pointer_MaskQTree)] > (call_main_mask_Int_goMux3,Pointer_MaskQTree) */
  assign call_main_mask_Int_goMux3_d = {call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Intmska8r_d[16:1],
                                        (call_main_mask_Int_unlockFork3_d[0] && call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Intmska8r_d[0])};
  assign call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Intmska8r_r = (call_main_mask_Int_goMux3_r && (call_main_mask_Int_unlockFork3_d[0] && call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Intmska8r_d[0]));
  assign call_main_mask_Int_unlockFork3_r = (call_main_mask_Int_goMux3_r && (call_main_mask_Int_unlockFork3_d[0] && call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Intmska8r_d[0]));
  
  /* mux (Ty Go,
     Ty Pointer_CTmain_mask_Int) : (call_main_mask_Int_unlockFork4,Go) [(call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Intsc_0_2,Pointer_CTmain_mask_Int)] > (call_main_mask_Int_goMux4,Pointer_CTmain_mask_Int) */
  assign call_main_mask_Int_goMux4_d = {call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Intsc_0_2_d[16:1],
                                        (call_main_mask_Int_unlockFork4_d[0] && call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Intsc_0_2_d[0])};
  assign call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Intsc_0_2_r = (call_main_mask_Int_goMux4_r && (call_main_mask_Int_unlockFork4_d[0] && call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Intsc_0_2_d[0]));
  assign call_main_mask_Int_unlockFork4_r = (call_main_mask_Int_goMux4_r && (call_main_mask_Int_unlockFork4_d[0] && call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Intsc_0_2_d[0]));
  
  /* buf (Ty Int) : (es_0_1_1I#_mux_mux_mux,Int) > (applyfnInt_Int_Int_5_resbuf,Int) */
  Int_t \es_0_1_1I#_mux_mux_mux_bufchan_d ;
  logic \es_0_1_1I#_mux_mux_mux_bufchan_r ;
  assign \es_0_1_1I#_mux_mux_mux_r  = ((! \es_0_1_1I#_mux_mux_mux_bufchan_d [0]) || \es_0_1_1I#_mux_mux_mux_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \es_0_1_1I#_mux_mux_mux_bufchan_d  <= {32'd0, 1'd0};
    else
      if (\es_0_1_1I#_mux_mux_mux_r )
        \es_0_1_1I#_mux_mux_mux_bufchan_d  <= \es_0_1_1I#_mux_mux_mux_d ;
  Int_t \es_0_1_1I#_mux_mux_mux_bufchan_buf ;
  assign \es_0_1_1I#_mux_mux_mux_bufchan_r  = (! \es_0_1_1I#_mux_mux_mux_bufchan_buf [0]);
  assign applyfnInt_Int_Int_5_resbuf_d = (\es_0_1_1I#_mux_mux_mux_bufchan_buf [0] ? \es_0_1_1I#_mux_mux_mux_bufchan_buf  :
                                          \es_0_1_1I#_mux_mux_mux_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \es_0_1_1I#_mux_mux_mux_bufchan_buf  <= {32'd0, 1'd0};
    else
      if ((applyfnInt_Int_Int_5_resbuf_r && \es_0_1_1I#_mux_mux_mux_bufchan_buf [0]))
        \es_0_1_1I#_mux_mux_mux_bufchan_buf  <= {32'd0, 1'd0};
      else if (((! applyfnInt_Int_Int_5_resbuf_r) && (! \es_0_1_1I#_mux_mux_mux_bufchan_buf [0])))
        \es_0_1_1I#_mux_mux_mux_bufchan_buf  <= \es_0_1_1I#_mux_mux_mux_bufchan_d ;
  
  /* buf (Ty QTree_Int) : (es_0_2_1QVal_Int,QTree_Int) > (lizzieLet4_1_argbuf,QTree_Int) */
  QTree_Int_t es_0_2_1QVal_Int_bufchan_d;
  logic es_0_2_1QVal_Int_bufchan_r;
  assign es_0_2_1QVal_Int_r = ((! es_0_2_1QVal_Int_bufchan_d[0]) || es_0_2_1QVal_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_0_2_1QVal_Int_bufchan_d <= {66'd0, 1'd0};
    else
      if (es_0_2_1QVal_Int_r)
        es_0_2_1QVal_Int_bufchan_d <= es_0_2_1QVal_Int_d;
  QTree_Int_t es_0_2_1QVal_Int_bufchan_buf;
  assign es_0_2_1QVal_Int_bufchan_r = (! es_0_2_1QVal_Int_bufchan_buf[0]);
  assign lizzieLet4_1_argbuf_d = (es_0_2_1QVal_Int_bufchan_buf[0] ? es_0_2_1QVal_Int_bufchan_buf :
                                  es_0_2_1QVal_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_0_2_1QVal_Int_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((lizzieLet4_1_argbuf_r && es_0_2_1QVal_Int_bufchan_buf[0]))
        es_0_2_1QVal_Int_bufchan_buf <= {66'd0, 1'd0};
      else if (((! lizzieLet4_1_argbuf_r) && (! es_0_2_1QVal_Int_bufchan_buf[0])))
        es_0_2_1QVal_Int_bufchan_buf <= es_0_2_1QVal_Int_bufchan_d;
  
  /* buf (Ty Int#) : (es_4_3_1lizzieLet27_4Lcall_$wnnz_Int0_1_Add32,Int#) > (contRet_0_1_1_argbuf,Int#) */
  \Int#_t  es_4_3_1lizzieLet27_4Lcall_$wnnz_Int0_1_Add32_bufchan_d;
  logic es_4_3_1lizzieLet27_4Lcall_$wnnz_Int0_1_Add32_bufchan_r;
  assign es_4_3_1lizzieLet27_4Lcall_$wnnz_Int0_1_Add32_r = ((! es_4_3_1lizzieLet27_4Lcall_$wnnz_Int0_1_Add32_bufchan_d[0]) || es_4_3_1lizzieLet27_4Lcall_$wnnz_Int0_1_Add32_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_4_3_1lizzieLet27_4Lcall_$wnnz_Int0_1_Add32_bufchan_d <= {32'd0,
                                                                  1'd0};
    else
      if (es_4_3_1lizzieLet27_4Lcall_$wnnz_Int0_1_Add32_r)
        es_4_3_1lizzieLet27_4Lcall_$wnnz_Int0_1_Add32_bufchan_d <= es_4_3_1lizzieLet27_4Lcall_$wnnz_Int0_1_Add32_d;
  \Int#_t  es_4_3_1lizzieLet27_4Lcall_$wnnz_Int0_1_Add32_bufchan_buf;
  assign es_4_3_1lizzieLet27_4Lcall_$wnnz_Int0_1_Add32_bufchan_r = (! es_4_3_1lizzieLet27_4Lcall_$wnnz_Int0_1_Add32_bufchan_buf[0]);
  assign contRet_0_1_1_argbuf_d = (es_4_3_1lizzieLet27_4Lcall_$wnnz_Int0_1_Add32_bufchan_buf[0] ? es_4_3_1lizzieLet27_4Lcall_$wnnz_Int0_1_Add32_bufchan_buf :
                                   es_4_3_1lizzieLet27_4Lcall_$wnnz_Int0_1_Add32_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_4_3_1lizzieLet27_4Lcall_$wnnz_Int0_1_Add32_bufchan_buf <= {32'd0,
                                                                    1'd0};
    else
      if ((contRet_0_1_1_argbuf_r && es_4_3_1lizzieLet27_4Lcall_$wnnz_Int0_1_Add32_bufchan_buf[0]))
        es_4_3_1lizzieLet27_4Lcall_$wnnz_Int0_1_Add32_bufchan_buf <= {32'd0,
                                                                      1'd0};
      else if (((! contRet_0_1_1_argbuf_r) && (! es_4_3_1lizzieLet27_4Lcall_$wnnz_Int0_1_Add32_bufchan_buf[0])))
        es_4_3_1lizzieLet27_4Lcall_$wnnz_Int0_1_Add32_bufchan_buf <= es_4_3_1lizzieLet27_4Lcall_$wnnz_Int0_1_Add32_bufchan_d;
  
  /* sink (Ty Int) : (es_6_1I#,Int) > */
  assign {\es_6_1I#_r , \es_6_1I#_dout } = {\es_6_1I#_rout ,
                                            \es_6_1I#_d };
  
  /* op_add (Ty Int#) : (es_6_1_1ww2XiV_1_1_Add32,Int#) (lizzieLet27_4Lcall_$wnnz_Int0,Int#) > (es_4_3_1lizzieLet27_4Lcall_$wnnz_Int0_1_Add32,Int#) */
  assign es_4_3_1lizzieLet27_4Lcall_$wnnz_Int0_1_Add32_d = {(es_6_1_1ww2XiV_1_1_Add32_d[32:1] + lizzieLet27_4Lcall_$wnnz_Int0_d[32:1]),
                                                            (es_6_1_1ww2XiV_1_1_Add32_d[0] && lizzieLet27_4Lcall_$wnnz_Int0_d[0])};
  assign {es_6_1_1ww2XiV_1_1_Add32_r,
          lizzieLet27_4Lcall_$wnnz_Int0_r} = {2 {(es_4_3_1lizzieLet27_4Lcall_$wnnz_Int0_1_Add32_r && es_4_3_1lizzieLet27_4Lcall_$wnnz_Int0_1_Add32_d[0])}};
  
  /* dcon (Ty MyDTInt_Int_Int,
      Dcon Dcon_$fNumInt_$c+) : [(go_1,Go)] > (go_1Dcon_$fNumInt_$c+,MyDTInt_Int_Int) */
  assign \go_1Dcon_$fNumInt_$c+_d  = \Dcon_$fNumInt_$c+_dc ((& {go_1_d[0]}), go_1_d);
  assign {go_1_r} = {1 {(\go_1Dcon_$fNumInt_$c+_r  && \go_1Dcon_$fNumInt_$c+_d [0])}};
  
  /* fork (Ty C10) : (go_10_goMux_choice,C10) > [(go_10_goMux_choice_1,C10),
                                            (go_10_goMux_choice_2,C10)] */
  logic [1:0] go_10_goMux_choice_emitted;
  logic [1:0] go_10_goMux_choice_done;
  assign go_10_goMux_choice_1_d = {go_10_goMux_choice_d[4:1],
                                   (go_10_goMux_choice_d[0] && (! go_10_goMux_choice_emitted[0]))};
  assign go_10_goMux_choice_2_d = {go_10_goMux_choice_d[4:1],
                                   (go_10_goMux_choice_d[0] && (! go_10_goMux_choice_emitted[1]))};
  assign go_10_goMux_choice_done = (go_10_goMux_choice_emitted | ({go_10_goMux_choice_2_d[0],
                                                                   go_10_goMux_choice_1_d[0]} & {go_10_goMux_choice_2_r,
                                                                                                 go_10_goMux_choice_1_r}));
  assign go_10_goMux_choice_r = (& go_10_goMux_choice_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_10_goMux_choice_emitted <= 2'd0;
    else
      go_10_goMux_choice_emitted <= (go_10_goMux_choice_r ? 2'd0 :
                                     go_10_goMux_choice_done);
  
  /* mux (Ty C10,
     Ty Pointer_QTree_Int) : (go_10_goMux_choice_1,C10) [(lizzieLet2_7QNone_Int_1_argbuf,Pointer_QTree_Int),
                                                         (contRet_0_1_argbuf,Pointer_QTree_Int),
                                                         (lizzieLet2_4QVal_Int_5QNone_Int_1_argbuf,Pointer_QTree_Int),
                                                         (lizzieLet8_1_argbuf,Pointer_QTree_Int),
                                                         (lizzieLet9_1_argbuf,Pointer_QTree_Int),
                                                         (lizzieLet10_1_argbuf,Pointer_QTree_Int),
                                                         (lizzieLet2_4QNode_Int_5QNone_Int_1_argbuf,Pointer_QTree_Int),
                                                         (lizzieLet11_1_argbuf,Pointer_QTree_Int),
                                                         (lizzieLet12_1_argbuf,Pointer_QTree_Int),
                                                         (lizzieLet13_1_argbuf,Pointer_QTree_Int)] > (srtarg_0_goMux_mux,Pointer_QTree_Int) */
  logic [16:0] srtarg_0_goMux_mux_mux;
  logic [9:0] srtarg_0_goMux_mux_onehot;
  always_comb
    unique case (go_10_goMux_choice_1_d[4:1])
      4'd0:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {10'd1,
                                                               lizzieLet2_7QNone_Int_1_argbuf_d};
      4'd1:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {10'd2,
                                                               contRet_0_1_argbuf_d};
      4'd2:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {10'd4,
                                                               lizzieLet2_4QVal_Int_5QNone_Int_1_argbuf_d};
      4'd3:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {10'd8,
                                                               lizzieLet8_1_argbuf_d};
      4'd4:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {10'd16,
                                                               lizzieLet9_1_argbuf_d};
      4'd5:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {10'd32,
                                                               lizzieLet10_1_argbuf_d};
      4'd6:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {10'd64,
                                                               lizzieLet2_4QNode_Int_5QNone_Int_1_argbuf_d};
      4'd7:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {10'd128,
                                                               lizzieLet11_1_argbuf_d};
      4'd8:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {10'd256,
                                                               lizzieLet12_1_argbuf_d};
      4'd9:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {10'd512,
                                                               lizzieLet13_1_argbuf_d};
      default:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {10'd0,
                                                               {16'd0, 1'd0}};
    endcase
  assign srtarg_0_goMux_mux_d = {srtarg_0_goMux_mux_mux[16:1],
                                 (srtarg_0_goMux_mux_mux[0] && go_10_goMux_choice_1_d[0])};
  assign go_10_goMux_choice_1_r = (srtarg_0_goMux_mux_d[0] && srtarg_0_goMux_mux_r);
  assign {lizzieLet13_1_argbuf_r,
          lizzieLet12_1_argbuf_r,
          lizzieLet11_1_argbuf_r,
          lizzieLet2_4QNode_Int_5QNone_Int_1_argbuf_r,
          lizzieLet10_1_argbuf_r,
          lizzieLet9_1_argbuf_r,
          lizzieLet8_1_argbuf_r,
          lizzieLet2_4QVal_Int_5QNone_Int_1_argbuf_r,
          contRet_0_1_argbuf_r,
          lizzieLet2_7QNone_Int_1_argbuf_r} = (go_10_goMux_choice_1_r ? srtarg_0_goMux_mux_onehot :
                                               10'd0);
  
  /* mux (Ty C10,
     Ty Pointer_CT$wmAdd_Int) : (go_10_goMux_choice_2,C10) [(lizzieLet2_5QNone_Int_1_argbuf,Pointer_CT$wmAdd_Int),
                                                            (sc_0_6_1_argbuf,Pointer_CT$wmAdd_Int),
                                                            (lizzieLet2_4QVal_Int_4QNone_Int_1_argbuf,Pointer_CT$wmAdd_Int),
                                                            (lizzieLet2_4QVal_Int_4QVal_Int_1_argbuf,Pointer_CT$wmAdd_Int),
                                                            (lizzieLet2_4QVal_Int_4QNode_Int_1_argbuf,Pointer_CT$wmAdd_Int),
                                                            (lizzieLet2_4QVal_Int_4QError_Int_1_argbuf,Pointer_CT$wmAdd_Int),
                                                            (lizzieLet2_4QNode_Int_4QNone_Int_1_argbuf,Pointer_CT$wmAdd_Int),
                                                            (lizzieLet2_4QNode_Int_4QVal_Int_1_argbuf,Pointer_CT$wmAdd_Int),
                                                            (lizzieLet2_4QNode_Int_4QError_Int_1_argbuf,Pointer_CT$wmAdd_Int),
                                                            (lizzieLet2_5QError_Int_1_argbuf,Pointer_CT$wmAdd_Int)] > (scfarg_0_goMux_mux,Pointer_CT$wmAdd_Int) */
  logic [16:0] scfarg_0_goMux_mux_mux;
  logic [9:0] scfarg_0_goMux_mux_onehot;
  always_comb
    unique case (go_10_goMux_choice_2_d[4:1])
      4'd0:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {10'd1,
                                                               lizzieLet2_5QNone_Int_1_argbuf_d};
      4'd1:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {10'd2,
                                                               sc_0_6_1_argbuf_d};
      4'd2:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {10'd4,
                                                               lizzieLet2_4QVal_Int_4QNone_Int_1_argbuf_d};
      4'd3:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {10'd8,
                                                               lizzieLet2_4QVal_Int_4QVal_Int_1_argbuf_d};
      4'd4:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {10'd16,
                                                               lizzieLet2_4QVal_Int_4QNode_Int_1_argbuf_d};
      4'd5:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {10'd32,
                                                               lizzieLet2_4QVal_Int_4QError_Int_1_argbuf_d};
      4'd6:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {10'd64,
                                                               lizzieLet2_4QNode_Int_4QNone_Int_1_argbuf_d};
      4'd7:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {10'd128,
                                                               lizzieLet2_4QNode_Int_4QVal_Int_1_argbuf_d};
      4'd8:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {10'd256,
                                                               lizzieLet2_4QNode_Int_4QError_Int_1_argbuf_d};
      4'd9:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {10'd512,
                                                               lizzieLet2_5QError_Int_1_argbuf_d};
      default:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {10'd0,
                                                               {16'd0, 1'd0}};
    endcase
  assign scfarg_0_goMux_mux_d = {scfarg_0_goMux_mux_mux[16:1],
                                 (scfarg_0_goMux_mux_mux[0] && go_10_goMux_choice_2_d[0])};
  assign go_10_goMux_choice_2_r = (scfarg_0_goMux_mux_d[0] && scfarg_0_goMux_mux_r);
  assign {lizzieLet2_5QError_Int_1_argbuf_r,
          lizzieLet2_4QNode_Int_4QError_Int_1_argbuf_r,
          lizzieLet2_4QNode_Int_4QVal_Int_1_argbuf_r,
          lizzieLet2_4QNode_Int_4QNone_Int_1_argbuf_r,
          lizzieLet2_4QVal_Int_4QError_Int_1_argbuf_r,
          lizzieLet2_4QVal_Int_4QNode_Int_1_argbuf_r,
          lizzieLet2_4QVal_Int_4QVal_Int_1_argbuf_r,
          lizzieLet2_4QVal_Int_4QNone_Int_1_argbuf_r,
          sc_0_6_1_argbuf_r,
          lizzieLet2_5QNone_Int_1_argbuf_r} = (go_10_goMux_choice_2_r ? scfarg_0_goMux_mux_onehot :
                                               10'd0);
  
  /* fork (Ty C4) : (go_11_goMux_choice,C4) > [(go_11_goMux_choice_1,C4),
                                          (go_11_goMux_choice_2,C4)] */
  logic [1:0] go_11_goMux_choice_emitted;
  logic [1:0] go_11_goMux_choice_done;
  assign go_11_goMux_choice_1_d = {go_11_goMux_choice_d[2:1],
                                   (go_11_goMux_choice_d[0] && (! go_11_goMux_choice_emitted[0]))};
  assign go_11_goMux_choice_2_d = {go_11_goMux_choice_d[2:1],
                                   (go_11_goMux_choice_d[0] && (! go_11_goMux_choice_emitted[1]))};
  assign go_11_goMux_choice_done = (go_11_goMux_choice_emitted | ({go_11_goMux_choice_2_d[0],
                                                                   go_11_goMux_choice_1_d[0]} & {go_11_goMux_choice_2_r,
                                                                                                 go_11_goMux_choice_1_r}));
  assign go_11_goMux_choice_r = (& go_11_goMux_choice_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_11_goMux_choice_emitted <= 2'd0;
    else
      go_11_goMux_choice_emitted <= (go_11_goMux_choice_r ? 2'd0 :
                                     go_11_goMux_choice_done);
  
  /* mux (Ty C4,
     Ty Int#) : (go_11_goMux_choice_1,C4) [(lizzieLet5_1_1_argbuf,Int#),
                                           (contRet_0_1_1_argbuf,Int#),
                                           (lizzieLet6_1_1_argbuf,Int#),
                                           (lizzieLet5_2_1_argbuf,Int#)] > (srtarg_0_1_goMux_mux,Int#) */
  logic [32:0] srtarg_0_1_goMux_mux_mux;
  logic [3:0] srtarg_0_1_goMux_mux_onehot;
  always_comb
    unique case (go_11_goMux_choice_1_d[2:1])
      2'd0:
        {srtarg_0_1_goMux_mux_onehot, srtarg_0_1_goMux_mux_mux} = {4'd1,
                                                                   lizzieLet5_1_1_argbuf_d};
      2'd1:
        {srtarg_0_1_goMux_mux_onehot, srtarg_0_1_goMux_mux_mux} = {4'd2,
                                                                   contRet_0_1_1_argbuf_d};
      2'd2:
        {srtarg_0_1_goMux_mux_onehot, srtarg_0_1_goMux_mux_mux} = {4'd4,
                                                                   lizzieLet6_1_1_argbuf_d};
      2'd3:
        {srtarg_0_1_goMux_mux_onehot, srtarg_0_1_goMux_mux_mux} = {4'd8,
                                                                   lizzieLet5_2_1_argbuf_d};
      default:
        {srtarg_0_1_goMux_mux_onehot, srtarg_0_1_goMux_mux_mux} = {4'd0,
                                                                   {32'd0, 1'd0}};
    endcase
  assign srtarg_0_1_goMux_mux_d = {srtarg_0_1_goMux_mux_mux[32:1],
                                   (srtarg_0_1_goMux_mux_mux[0] && go_11_goMux_choice_1_d[0])};
  assign go_11_goMux_choice_1_r = (srtarg_0_1_goMux_mux_d[0] && srtarg_0_1_goMux_mux_r);
  assign {lizzieLet5_2_1_argbuf_r,
          lizzieLet6_1_1_argbuf_r,
          contRet_0_1_1_argbuf_r,
          lizzieLet5_1_1_argbuf_r} = (go_11_goMux_choice_1_r ? srtarg_0_1_goMux_mux_onehot :
                                      4'd0);
  
  /* mux (Ty C4,
     Ty Pointer_CT$wnnz_Int) : (go_11_goMux_choice_2,C4) [(lizzieLet12_1_4QNone_Int_1_argbuf,Pointer_CT$wnnz_Int),
                                                          (sc_0_10_1_argbuf,Pointer_CT$wnnz_Int),
                                                          (lizzieLet12_1_4QVal_Int_1_argbuf,Pointer_CT$wnnz_Int),
                                                          (lizzieLet12_1_4QError_Int_1_argbuf,Pointer_CT$wnnz_Int)] > (scfarg_0_1_goMux_mux,Pointer_CT$wnnz_Int) */
  logic [16:0] scfarg_0_1_goMux_mux_mux;
  logic [3:0] scfarg_0_1_goMux_mux_onehot;
  always_comb
    unique case (go_11_goMux_choice_2_d[2:1])
      2'd0:
        {scfarg_0_1_goMux_mux_onehot, scfarg_0_1_goMux_mux_mux} = {4'd1,
                                                                   lizzieLet12_1_4QNone_Int_1_argbuf_d};
      2'd1:
        {scfarg_0_1_goMux_mux_onehot, scfarg_0_1_goMux_mux_mux} = {4'd2,
                                                                   sc_0_10_1_argbuf_d};
      2'd2:
        {scfarg_0_1_goMux_mux_onehot, scfarg_0_1_goMux_mux_mux} = {4'd4,
                                                                   lizzieLet12_1_4QVal_Int_1_argbuf_d};
      2'd3:
        {scfarg_0_1_goMux_mux_onehot, scfarg_0_1_goMux_mux_mux} = {4'd8,
                                                                   lizzieLet12_1_4QError_Int_1_argbuf_d};
      default:
        {scfarg_0_1_goMux_mux_onehot, scfarg_0_1_goMux_mux_mux} = {4'd0,
                                                                   {16'd0, 1'd0}};
    endcase
  assign scfarg_0_1_goMux_mux_d = {scfarg_0_1_goMux_mux_mux[16:1],
                                   (scfarg_0_1_goMux_mux_mux[0] && go_11_goMux_choice_2_d[0])};
  assign go_11_goMux_choice_2_r = (scfarg_0_1_goMux_mux_d[0] && scfarg_0_1_goMux_mux_r);
  assign {lizzieLet12_1_4QError_Int_1_argbuf_r,
          lizzieLet12_1_4QVal_Int_1_argbuf_r,
          sc_0_10_1_argbuf_r,
          lizzieLet12_1_4QNone_Int_1_argbuf_r} = (go_11_goMux_choice_2_r ? scfarg_0_1_goMux_mux_onehot :
                                                  4'd0);
  
  /* fork (Ty C6) : (go_12_goMux_choice,C6) > [(go_12_goMux_choice_1,C6),
                                          (go_12_goMux_choice_2,C6)] */
  logic [1:0] go_12_goMux_choice_emitted;
  logic [1:0] go_12_goMux_choice_done;
  assign go_12_goMux_choice_1_d = {go_12_goMux_choice_d[3:1],
                                   (go_12_goMux_choice_d[0] && (! go_12_goMux_choice_emitted[0]))};
  assign go_12_goMux_choice_2_d = {go_12_goMux_choice_d[3:1],
                                   (go_12_goMux_choice_d[0] && (! go_12_goMux_choice_emitted[1]))};
  assign go_12_goMux_choice_done = (go_12_goMux_choice_emitted | ({go_12_goMux_choice_2_d[0],
                                                                   go_12_goMux_choice_1_d[0]} & {go_12_goMux_choice_2_r,
                                                                                                 go_12_goMux_choice_1_r}));
  assign go_12_goMux_choice_r = (& go_12_goMux_choice_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_12_goMux_choice_emitted <= 2'd0;
    else
      go_12_goMux_choice_emitted <= (go_12_goMux_choice_r ? 2'd0 :
                                     go_12_goMux_choice_done);
  
  /* mux (Ty C6,
     Ty Pointer_QTree_Int) : (go_12_goMux_choice_1,C6) [(lizzieLet0_1_1_argbuf,Pointer_QTree_Int),
                                                        (contRet_0_2_1_argbuf,Pointer_QTree_Int),
                                                        (lizzieLet14_1_5MQVal_1_argbuf,Pointer_QTree_Int),
                                                        (lizzieLet1_1_1_argbuf,Pointer_QTree_Int),
                                                        (lizzieLet2_1_1_argbuf,Pointer_QTree_Int),
                                                        (lizzieLet3_1_1_argbuf,Pointer_QTree_Int)] > (srtarg_0_2_goMux_mux,Pointer_QTree_Int) */
  logic [16:0] srtarg_0_2_goMux_mux_mux;
  logic [5:0] srtarg_0_2_goMux_mux_onehot;
  always_comb
    unique case (go_12_goMux_choice_1_d[3:1])
      3'd0:
        {srtarg_0_2_goMux_mux_onehot, srtarg_0_2_goMux_mux_mux} = {6'd1,
                                                                   lizzieLet0_1_1_argbuf_d};
      3'd1:
        {srtarg_0_2_goMux_mux_onehot, srtarg_0_2_goMux_mux_mux} = {6'd2,
                                                                   contRet_0_2_1_argbuf_d};
      3'd2:
        {srtarg_0_2_goMux_mux_onehot, srtarg_0_2_goMux_mux_mux} = {6'd4,
                                                                   lizzieLet14_1_5MQVal_1_argbuf_d};
      3'd3:
        {srtarg_0_2_goMux_mux_onehot, srtarg_0_2_goMux_mux_mux} = {6'd8,
                                                                   lizzieLet1_1_1_argbuf_d};
      3'd4:
        {srtarg_0_2_goMux_mux_onehot, srtarg_0_2_goMux_mux_mux} = {6'd16,
                                                                   lizzieLet2_1_1_argbuf_d};
      3'd5:
        {srtarg_0_2_goMux_mux_onehot, srtarg_0_2_goMux_mux_mux} = {6'd32,
                                                                   lizzieLet3_1_1_argbuf_d};
      default:
        {srtarg_0_2_goMux_mux_onehot, srtarg_0_2_goMux_mux_mux} = {6'd0,
                                                                   {16'd0, 1'd0}};
    endcase
  assign srtarg_0_2_goMux_mux_d = {srtarg_0_2_goMux_mux_mux[16:1],
                                   (srtarg_0_2_goMux_mux_mux[0] && go_12_goMux_choice_1_d[0])};
  assign go_12_goMux_choice_1_r = (srtarg_0_2_goMux_mux_d[0] && srtarg_0_2_goMux_mux_r);
  assign {lizzieLet3_1_1_argbuf_r,
          lizzieLet2_1_1_argbuf_r,
          lizzieLet1_1_1_argbuf_r,
          lizzieLet14_1_5MQVal_1_argbuf_r,
          contRet_0_2_1_argbuf_r,
          lizzieLet0_1_1_argbuf_r} = (go_12_goMux_choice_1_r ? srtarg_0_2_goMux_mux_onehot :
                                      6'd0);
  
  /* mux (Ty C6,
     Ty Pointer_CTmain_mask_Int) : (go_12_goMux_choice_2,C6) [(lizzieLet14_1_6MQNone_1_argbuf,Pointer_CTmain_mask_Int),
                                                              (sc_0_14_1_argbuf,Pointer_CTmain_mask_Int),
                                                              (lizzieLet14_1_6MQVal_1_argbuf,Pointer_CTmain_mask_Int),
                                                              (lizzieLet14_1_4MQNode_4QNone_Int_1_argbuf,Pointer_CTmain_mask_Int),
                                                              (lizzieLet14_1_4MQNode_4QVal_Int_1_argbuf,Pointer_CTmain_mask_Int),
                                                              (lizzieLet14_1_4MQNode_4QError_Int_1_argbuf,Pointer_CTmain_mask_Int)] > (scfarg_0_2_goMux_mux,Pointer_CTmain_mask_Int) */
  logic [16:0] scfarg_0_2_goMux_mux_mux;
  logic [5:0] scfarg_0_2_goMux_mux_onehot;
  always_comb
    unique case (go_12_goMux_choice_2_d[3:1])
      3'd0:
        {scfarg_0_2_goMux_mux_onehot, scfarg_0_2_goMux_mux_mux} = {6'd1,
                                                                   lizzieLet14_1_6MQNone_1_argbuf_d};
      3'd1:
        {scfarg_0_2_goMux_mux_onehot, scfarg_0_2_goMux_mux_mux} = {6'd2,
                                                                   sc_0_14_1_argbuf_d};
      3'd2:
        {scfarg_0_2_goMux_mux_onehot, scfarg_0_2_goMux_mux_mux} = {6'd4,
                                                                   lizzieLet14_1_6MQVal_1_argbuf_d};
      3'd3:
        {scfarg_0_2_goMux_mux_onehot, scfarg_0_2_goMux_mux_mux} = {6'd8,
                                                                   lizzieLet14_1_4MQNode_4QNone_Int_1_argbuf_d};
      3'd4:
        {scfarg_0_2_goMux_mux_onehot, scfarg_0_2_goMux_mux_mux} = {6'd16,
                                                                   lizzieLet14_1_4MQNode_4QVal_Int_1_argbuf_d};
      3'd5:
        {scfarg_0_2_goMux_mux_onehot, scfarg_0_2_goMux_mux_mux} = {6'd32,
                                                                   lizzieLet14_1_4MQNode_4QError_Int_1_argbuf_d};
      default:
        {scfarg_0_2_goMux_mux_onehot, scfarg_0_2_goMux_mux_mux} = {6'd0,
                                                                   {16'd0, 1'd0}};
    endcase
  assign scfarg_0_2_goMux_mux_d = {scfarg_0_2_goMux_mux_mux[16:1],
                                   (scfarg_0_2_goMux_mux_mux[0] && go_12_goMux_choice_2_d[0])};
  assign go_12_goMux_choice_2_r = (scfarg_0_2_goMux_mux_d[0] && scfarg_0_2_goMux_mux_r);
  assign {lizzieLet14_1_4MQNode_4QError_Int_1_argbuf_r,
          lizzieLet14_1_4MQNode_4QVal_Int_1_argbuf_r,
          lizzieLet14_1_4MQNode_4QNone_Int_1_argbuf_r,
          lizzieLet14_1_6MQVal_1_argbuf_r,
          sc_0_14_1_argbuf_r,
          lizzieLet14_1_6MQNone_1_argbuf_r} = (go_12_goMux_choice_2_r ? scfarg_0_2_goMux_mux_onehot :
                                               6'd0);
  
  /* buf (Ty MyDTInt_Int_Int) : (go_1Dcon_$fNumInt_$c+,MyDTInt_Int_Int) > (es_3_1_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t \go_1Dcon_$fNumInt_$c+_bufchan_d ;
  logic \go_1Dcon_$fNumInt_$c+_bufchan_r ;
  assign \go_1Dcon_$fNumInt_$c+_r  = ((! \go_1Dcon_$fNumInt_$c+_bufchan_d [0]) || \go_1Dcon_$fNumInt_$c+_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \go_1Dcon_$fNumInt_$c+_bufchan_d  <= 1'd0;
    else
      if (\go_1Dcon_$fNumInt_$c+_r )
        \go_1Dcon_$fNumInt_$c+_bufchan_d  <= \go_1Dcon_$fNumInt_$c+_d ;
  MyDTInt_Int_Int_t \go_1Dcon_$fNumInt_$c+_bufchan_buf ;
  assign \go_1Dcon_$fNumInt_$c+_bufchan_r  = (! \go_1Dcon_$fNumInt_$c+_bufchan_buf [0]);
  assign es_3_1_argbuf_d = (\go_1Dcon_$fNumInt_$c+_bufchan_buf [0] ? \go_1Dcon_$fNumInt_$c+_bufchan_buf  :
                            \go_1Dcon_$fNumInt_$c+_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \go_1Dcon_$fNumInt_$c+_bufchan_buf  <= 1'd0;
    else
      if ((es_3_1_argbuf_r && \go_1Dcon_$fNumInt_$c+_bufchan_buf [0]))
        \go_1Dcon_$fNumInt_$c+_bufchan_buf  <= 1'd0;
      else if (((! es_3_1_argbuf_r) && (! \go_1Dcon_$fNumInt_$c+_bufchan_buf [0])))
        \go_1Dcon_$fNumInt_$c+_bufchan_buf  <= \go_1Dcon_$fNumInt_$c+_bufchan_d ;
  
  /* buf (Ty Go) : (go_2,Go) > (go_2_argbuf,Go) */
  Go_t go_2_bufchan_d;
  logic go_2_bufchan_r;
  assign go_2_r = ((! go_2_bufchan_d[0]) || go_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_2_bufchan_d <= 1'd0;
    else if (go_2_r) go_2_bufchan_d <= go_2_d;
  Go_t go_2_bufchan_buf;
  assign go_2_bufchan_r = (! go_2_bufchan_buf[0]);
  assign go_2_argbuf_d = (go_2_bufchan_buf[0] ? go_2_bufchan_buf :
                          go_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_2_bufchan_buf <= 1'd0;
    else
      if ((go_2_argbuf_r && go_2_bufchan_buf[0]))
        go_2_bufchan_buf <= 1'd0;
      else if (((! go_2_argbuf_r) && (! go_2_bufchan_buf[0])))
        go_2_bufchan_buf <= go_2_bufchan_d;
  
  /* dcon (Ty TupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int,
      Dcon TupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int) : [(go_2_argbuf,Go),
                                                                               (es_3_1_argbuf,MyDTInt_Int_Int),
                                                                               (m2a93_1,Pointer_QTree_Int),
                                                                               (m3a94_2,Pointer_QTree_Int)] > ($wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1,TupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int) */
  assign \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1_d  = TupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_dc((& {go_2_argbuf_d[0],
                                                                                                                                                                  es_3_1_argbuf_d[0],
                                                                                                                                                                  m2a93_1_d[0],
                                                                                                                                                                  m3a94_2_d[0]}), go_2_argbuf_d, es_3_1_argbuf_d, m2a93_1_d, m3a94_2_d);
  assign {go_2_argbuf_r,
          es_3_1_argbuf_r,
          m2a93_1_r,
          m3a94_2_r} = {4 {(\$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1_r  && \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1_d [0])}};
  
  /* buf (Ty Go) : (go_3,Go) > (go_3_argbuf,Go) */
  Go_t go_3_bufchan_d;
  logic go_3_bufchan_r;
  assign go_3_r = ((! go_3_bufchan_d[0]) || go_3_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_3_bufchan_d <= 1'd0;
    else if (go_3_r) go_3_bufchan_d <= go_3_d;
  Go_t go_3_bufchan_buf;
  assign go_3_bufchan_r = (! go_3_bufchan_buf[0]);
  assign go_3_argbuf_d = (go_3_bufchan_buf[0] ? go_3_bufchan_buf :
                          go_3_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_3_bufchan_buf <= 1'd0;
    else
      if ((go_3_argbuf_r && go_3_bufchan_buf[0]))
        go_3_bufchan_buf <= 1'd0;
      else if (((! go_3_argbuf_r) && (! go_3_bufchan_buf[0])))
        go_3_bufchan_buf <= go_3_bufchan_d;
  
  /* dcon (Ty TupGo___Pointer_QTree_Int___Pointer_MaskQTree,
      Dcon TupGo___Pointer_QTree_Int___Pointer_MaskQTree) : [(go_3_argbuf,Go),
                                                             (es_1_1_argbuf,Pointer_QTree_Int),
                                                             (m1a92_0,Pointer_MaskQTree)] > (main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree_1,TupGo___Pointer_QTree_Int___Pointer_MaskQTree) */
  assign main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree_1_d = TupGo___Pointer_QTree_Int___Pointer_MaskQTree_dc((& {go_3_argbuf_d[0],
                                                                                                                               es_1_1_argbuf_d[0],
                                                                                                                               m1a92_0_d[0]}), go_3_argbuf_d, es_1_1_argbuf_d, m1a92_0_d);
  assign {go_3_argbuf_r,
          es_1_1_argbuf_r,
          m1a92_0_r} = {3 {(main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree_1_r && main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree_1_d[0])}};
  
  /* buf (Ty Go) : (go_4,Go) > (go_4_argbuf,Go) */
  Go_t go_4_bufchan_d;
  logic go_4_bufchan_r;
  assign go_4_r = ((! go_4_bufchan_d[0]) || go_4_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_4_bufchan_d <= 1'd0;
    else if (go_4_r) go_4_bufchan_d <= go_4_d;
  Go_t go_4_bufchan_buf;
  assign go_4_bufchan_r = (! go_4_bufchan_buf[0]);
  assign go_4_argbuf_d = (go_4_bufchan_buf[0] ? go_4_bufchan_buf :
                          go_4_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_4_bufchan_buf <= 1'd0;
    else
      if ((go_4_argbuf_r && go_4_bufchan_buf[0]))
        go_4_bufchan_buf <= 1'd0;
      else if (((! go_4_argbuf_r) && (! go_4_bufchan_buf[0])))
        go_4_bufchan_buf <= go_4_bufchan_d;
  
  /* dcon (Ty CT$wmAdd_Int,
      Dcon L$wmAdd_Intsbos) : [(go_4_1,Go)] > (go_4_1L$wmAdd_Intsbos,CT$wmAdd_Int) */
  assign go_4_1L$wmAdd_Intsbos_d = L$wmAdd_Intsbos_dc((& {go_4_1_d[0]}), go_4_1_d);
  assign {go_4_1_r} = {1 {(go_4_1L$wmAdd_Intsbos_r && go_4_1L$wmAdd_Intsbos_d[0])}};
  
  /* buf (Ty CT$wmAdd_Int) : (go_4_1L$wmAdd_Intsbos,CT$wmAdd_Int) > (lizzieLet0_1_argbuf,CT$wmAdd_Int) */
  CT$wmAdd_Int_t go_4_1L$wmAdd_Intsbos_bufchan_d;
  logic go_4_1L$wmAdd_Intsbos_bufchan_r;
  assign go_4_1L$wmAdd_Intsbos_r = ((! go_4_1L$wmAdd_Intsbos_bufchan_d[0]) || go_4_1L$wmAdd_Intsbos_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      go_4_1L$wmAdd_Intsbos_bufchan_d <= {115'd0, 1'd0};
    else
      if (go_4_1L$wmAdd_Intsbos_r)
        go_4_1L$wmAdd_Intsbos_bufchan_d <= go_4_1L$wmAdd_Intsbos_d;
  CT$wmAdd_Int_t go_4_1L$wmAdd_Intsbos_bufchan_buf;
  assign go_4_1L$wmAdd_Intsbos_bufchan_r = (! go_4_1L$wmAdd_Intsbos_bufchan_buf[0]);
  assign lizzieLet0_1_argbuf_d = (go_4_1L$wmAdd_Intsbos_bufchan_buf[0] ? go_4_1L$wmAdd_Intsbos_bufchan_buf :
                                  go_4_1L$wmAdd_Intsbos_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      go_4_1L$wmAdd_Intsbos_bufchan_buf <= {115'd0, 1'd0};
    else
      if ((lizzieLet0_1_argbuf_r && go_4_1L$wmAdd_Intsbos_bufchan_buf[0]))
        go_4_1L$wmAdd_Intsbos_bufchan_buf <= {115'd0, 1'd0};
      else if (((! lizzieLet0_1_argbuf_r) && (! go_4_1L$wmAdd_Intsbos_bufchan_buf[0])))
        go_4_1L$wmAdd_Intsbos_bufchan_buf <= go_4_1L$wmAdd_Intsbos_bufchan_d;
  
  /* buf (Ty Go) : (go_4_2,Go) > (go_4_2_argbuf,Go) */
  Go_t go_4_2_bufchan_d;
  logic go_4_2_bufchan_r;
  assign go_4_2_r = ((! go_4_2_bufchan_d[0]) || go_4_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_4_2_bufchan_d <= 1'd0;
    else if (go_4_2_r) go_4_2_bufchan_d <= go_4_2_d;
  Go_t go_4_2_bufchan_buf;
  assign go_4_2_bufchan_r = (! go_4_2_bufchan_buf[0]);
  assign go_4_2_argbuf_d = (go_4_2_bufchan_buf[0] ? go_4_2_bufchan_buf :
                            go_4_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_4_2_bufchan_buf <= 1'd0;
    else
      if ((go_4_2_argbuf_r && go_4_2_bufchan_buf[0]))
        go_4_2_bufchan_buf <= 1'd0;
      else if (((! go_4_2_argbuf_r) && (! go_4_2_bufchan_buf[0])))
        go_4_2_bufchan_buf <= go_4_2_bufchan_d;
  
  /* dcon (Ty TupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Int,
      Dcon TupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Int) : [(go_4_2_argbuf,Go),
                                                                                                      (wsie_1_argbuf,MyDTInt_Int_Int),
                                                                                                      (w1sif_1_argbuf,Pointer_QTree_Int),
                                                                                                      (w2sig_1_argbuf,Pointer_QTree_Int),
                                                                                                      (lizzieLet14_1_argbuf,Pointer_CT$wmAdd_Int)] > (call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Int_1,TupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Int) */
  assign call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Int_1_d = TupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Int_dc((& {go_4_2_argbuf_d[0],
                                                                                                                                                                                                                   wsie_1_argbuf_d[0],
                                                                                                                                                                                                                   w1sif_1_argbuf_d[0],
                                                                                                                                                                                                                   w2sig_1_argbuf_d[0],
                                                                                                                                                                                                                   lizzieLet14_1_argbuf_d[0]}), go_4_2_argbuf_d, wsie_1_argbuf_d, w1sif_1_argbuf_d, w2sig_1_argbuf_d, lizzieLet14_1_argbuf_d);
  assign {go_4_2_argbuf_r,
          wsie_1_argbuf_r,
          w1sif_1_argbuf_r,
          w2sig_1_argbuf_r,
          lizzieLet14_1_argbuf_r} = {5 {(call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Int_1_r && call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Int_1_d[0])}};
  
  /* dcon (Ty TupGo___Pointer_QTree_Int,
      Dcon TupGo___Pointer_QTree_Int) : [(go_4_argbuf,Go),
                                         (es_0_1_argbuf,Pointer_QTree_Int)] > ($wnnz_IntTupGo___Pointer_QTree_Int_1,TupGo___Pointer_QTree_Int) */
  assign \$wnnz_IntTupGo___Pointer_QTree_Int_1_d  = TupGo___Pointer_QTree_Int_dc((& {go_4_argbuf_d[0],
                                                                                     es_0_1_argbuf_d[0]}), go_4_argbuf_d, es_0_1_argbuf_d);
  assign {go_4_argbuf_r,
          es_0_1_argbuf_r} = {2 {(\$wnnz_IntTupGo___Pointer_QTree_Int_1_r  && \$wnnz_IntTupGo___Pointer_QTree_Int_1_d [0])}};
  
  /* dcon (Ty CT$wnnz_Int,
      Dcon L$wnnz_Intsbos) : [(go_5_1,Go)] > (go_5_1L$wnnz_Intsbos,CT$wnnz_Int) */
  assign go_5_1L$wnnz_Intsbos_d = L$wnnz_Intsbos_dc((& {go_5_1_d[0]}), go_5_1_d);
  assign {go_5_1_r} = {1 {(go_5_1L$wnnz_Intsbos_r && go_5_1L$wnnz_Intsbos_d[0])}};
  
  /* buf (Ty CT$wnnz_Int) : (go_5_1L$wnnz_Intsbos,CT$wnnz_Int) > (lizzieLet1_1_argbuf,CT$wnnz_Int) */
  CT$wnnz_Int_t go_5_1L$wnnz_Intsbos_bufchan_d;
  logic go_5_1L$wnnz_Intsbos_bufchan_r;
  assign go_5_1L$wnnz_Intsbos_r = ((! go_5_1L$wnnz_Intsbos_bufchan_d[0]) || go_5_1L$wnnz_Intsbos_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      go_5_1L$wnnz_Intsbos_bufchan_d <= {115'd0, 1'd0};
    else
      if (go_5_1L$wnnz_Intsbos_r)
        go_5_1L$wnnz_Intsbos_bufchan_d <= go_5_1L$wnnz_Intsbos_d;
  CT$wnnz_Int_t go_5_1L$wnnz_Intsbos_bufchan_buf;
  assign go_5_1L$wnnz_Intsbos_bufchan_r = (! go_5_1L$wnnz_Intsbos_bufchan_buf[0]);
  assign lizzieLet1_1_argbuf_d = (go_5_1L$wnnz_Intsbos_bufchan_buf[0] ? go_5_1L$wnnz_Intsbos_bufchan_buf :
                                  go_5_1L$wnnz_Intsbos_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      go_5_1L$wnnz_Intsbos_bufchan_buf <= {115'd0, 1'd0};
    else
      if ((lizzieLet1_1_argbuf_r && go_5_1L$wnnz_Intsbos_bufchan_buf[0]))
        go_5_1L$wnnz_Intsbos_bufchan_buf <= {115'd0, 1'd0};
      else if (((! lizzieLet1_1_argbuf_r) && (! go_5_1L$wnnz_Intsbos_bufchan_buf[0])))
        go_5_1L$wnnz_Intsbos_bufchan_buf <= go_5_1L$wnnz_Intsbos_bufchan_d;
  
  /* buf (Ty Go) : (go_5_2,Go) > (go_5_2_argbuf,Go) */
  Go_t go_5_2_bufchan_d;
  logic go_5_2_bufchan_r;
  assign go_5_2_r = ((! go_5_2_bufchan_d[0]) || go_5_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_5_2_bufchan_d <= 1'd0;
    else if (go_5_2_r) go_5_2_bufchan_d <= go_5_2_d;
  Go_t go_5_2_bufchan_buf;
  assign go_5_2_bufchan_r = (! go_5_2_bufchan_buf[0]);
  assign go_5_2_argbuf_d = (go_5_2_bufchan_buf[0] ? go_5_2_bufchan_buf :
                            go_5_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_5_2_bufchan_buf <= 1'd0;
    else
      if ((go_5_2_argbuf_r && go_5_2_bufchan_buf[0]))
        go_5_2_bufchan_buf <= 1'd0;
      else if (((! go_5_2_argbuf_r) && (! go_5_2_bufchan_buf[0])))
        go_5_2_bufchan_buf <= go_5_2_bufchan_d;
  
  /* dcon (Ty TupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int,
      Dcon TupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int) : [(go_5_2_argbuf,Go),
                                                               (wsij_1_argbuf,Pointer_QTree_Int),
                                                               (lizzieLet7_1_argbuf,Pointer_CT$wnnz_Int)] > (call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1,TupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int) */
  assign call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_d = TupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_dc((& {go_5_2_argbuf_d[0],
                                                                                                                                    wsij_1_argbuf_d[0],
                                                                                                                                    lizzieLet7_1_argbuf_d[0]}), go_5_2_argbuf_d, wsij_1_argbuf_d, lizzieLet7_1_argbuf_d);
  assign {go_5_2_argbuf_r,
          wsij_1_argbuf_r,
          lizzieLet7_1_argbuf_r} = {3 {(call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_r && call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_d[0])}};
  
  /* fork (Ty C5) : (go_6_goMux_choice,C5) > [(go_6_goMux_choice_1,C5),
                                         (go_6_goMux_choice_2,C5),
                                         (go_6_goMux_choice_3,C5),
                                         (go_6_goMux_choice_4,C5)] */
  logic [3:0] go_6_goMux_choice_emitted;
  logic [3:0] go_6_goMux_choice_done;
  assign go_6_goMux_choice_1_d = {go_6_goMux_choice_d[3:1],
                                  (go_6_goMux_choice_d[0] && (! go_6_goMux_choice_emitted[0]))};
  assign go_6_goMux_choice_2_d = {go_6_goMux_choice_d[3:1],
                                  (go_6_goMux_choice_d[0] && (! go_6_goMux_choice_emitted[1]))};
  assign go_6_goMux_choice_3_d = {go_6_goMux_choice_d[3:1],
                                  (go_6_goMux_choice_d[0] && (! go_6_goMux_choice_emitted[2]))};
  assign go_6_goMux_choice_4_d = {go_6_goMux_choice_d[3:1],
                                  (go_6_goMux_choice_d[0] && (! go_6_goMux_choice_emitted[3]))};
  assign go_6_goMux_choice_done = (go_6_goMux_choice_emitted | ({go_6_goMux_choice_4_d[0],
                                                                 go_6_goMux_choice_3_d[0],
                                                                 go_6_goMux_choice_2_d[0],
                                                                 go_6_goMux_choice_1_d[0]} & {go_6_goMux_choice_4_r,
                                                                                              go_6_goMux_choice_3_r,
                                                                                              go_6_goMux_choice_2_r,
                                                                                              go_6_goMux_choice_1_r}));
  assign go_6_goMux_choice_r = (& go_6_goMux_choice_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_6_goMux_choice_emitted <= 4'd0;
    else
      go_6_goMux_choice_emitted <= (go_6_goMux_choice_r ? 4'd0 :
                                    go_6_goMux_choice_done);
  
  /* mux (Ty C5,
     Ty MyDTInt_Int_Int) : (go_6_goMux_choice_1,C5) [(call_$wmAdd_Int_goMux2,MyDTInt_Int_Int),
                                                     (wsie_2_2_argbuf,MyDTInt_Int_Int),
                                                     (wsie_3_2_argbuf,MyDTInt_Int_Int),
                                                     (wsie_4_1_argbuf,MyDTInt_Int_Int),
                                                     (lizzieLet2_4QNode_Int_6QNode_Int_2_argbuf,MyDTInt_Int_Int)] > (wsie_1_goMux_mux,MyDTInt_Int_Int) */
  logic [0:0] wsie_1_goMux_mux_mux;
  logic [4:0] wsie_1_goMux_mux_onehot;
  always_comb
    unique case (go_6_goMux_choice_1_d[3:1])
      3'd0:
        {wsie_1_goMux_mux_onehot, wsie_1_goMux_mux_mux} = {5'd1,
                                                           call_$wmAdd_Int_goMux2_d};
      3'd1:
        {wsie_1_goMux_mux_onehot, wsie_1_goMux_mux_mux} = {5'd2,
                                                           wsie_2_2_argbuf_d};
      3'd2:
        {wsie_1_goMux_mux_onehot, wsie_1_goMux_mux_mux} = {5'd4,
                                                           wsie_3_2_argbuf_d};
      3'd3:
        {wsie_1_goMux_mux_onehot, wsie_1_goMux_mux_mux} = {5'd8,
                                                           wsie_4_1_argbuf_d};
      3'd4:
        {wsie_1_goMux_mux_onehot, wsie_1_goMux_mux_mux} = {5'd16,
                                                           lizzieLet2_4QNode_Int_6QNode_Int_2_argbuf_d};
      default:
        {wsie_1_goMux_mux_onehot, wsie_1_goMux_mux_mux} = {5'd0, 1'd0};
    endcase
  assign wsie_1_goMux_mux_d = (wsie_1_goMux_mux_mux[0] && go_6_goMux_choice_1_d[0]);
  assign go_6_goMux_choice_1_r = (wsie_1_goMux_mux_d[0] && wsie_1_goMux_mux_r);
  assign {lizzieLet2_4QNode_Int_6QNode_Int_2_argbuf_r,
          wsie_4_1_argbuf_r,
          wsie_3_2_argbuf_r,
          wsie_2_2_argbuf_r,
          call_$wmAdd_Int_goMux2_r} = (go_6_goMux_choice_1_r ? wsie_1_goMux_mux_onehot :
                                       5'd0);
  
  /* mux (Ty C5,
     Ty Pointer_QTree_Int) : (go_6_goMux_choice_2,C5) [(call_$wmAdd_Int_goMux3,Pointer_QTree_Int),
                                                       (q3a8j_1_1_argbuf,Pointer_QTree_Int),
                                                       (q2a8i_2_1_argbuf,Pointer_QTree_Int),
                                                       (q1a8h_3_1_argbuf,Pointer_QTree_Int),
                                                       (lizzieLet2_4QNode_Int_10QNode_Int_1_argbuf,Pointer_QTree_Int)] > (w1sif_1_goMux_mux,Pointer_QTree_Int) */
  logic [16:0] w1sif_1_goMux_mux_mux;
  logic [4:0] w1sif_1_goMux_mux_onehot;
  always_comb
    unique case (go_6_goMux_choice_2_d[3:1])
      3'd0:
        {w1sif_1_goMux_mux_onehot, w1sif_1_goMux_mux_mux} = {5'd1,
                                                             call_$wmAdd_Int_goMux3_d};
      3'd1:
        {w1sif_1_goMux_mux_onehot, w1sif_1_goMux_mux_mux} = {5'd2,
                                                             q3a8j_1_1_argbuf_d};
      3'd2:
        {w1sif_1_goMux_mux_onehot, w1sif_1_goMux_mux_mux} = {5'd4,
                                                             q2a8i_2_1_argbuf_d};
      3'd3:
        {w1sif_1_goMux_mux_onehot, w1sif_1_goMux_mux_mux} = {5'd8,
                                                             q1a8h_3_1_argbuf_d};
      3'd4:
        {w1sif_1_goMux_mux_onehot, w1sif_1_goMux_mux_mux} = {5'd16,
                                                             lizzieLet2_4QNode_Int_10QNode_Int_1_argbuf_d};
      default:
        {w1sif_1_goMux_mux_onehot, w1sif_1_goMux_mux_mux} = {5'd0,
                                                             {16'd0, 1'd0}};
    endcase
  assign w1sif_1_goMux_mux_d = {w1sif_1_goMux_mux_mux[16:1],
                                (w1sif_1_goMux_mux_mux[0] && go_6_goMux_choice_2_d[0])};
  assign go_6_goMux_choice_2_r = (w1sif_1_goMux_mux_d[0] && w1sif_1_goMux_mux_r);
  assign {lizzieLet2_4QNode_Int_10QNode_Int_1_argbuf_r,
          q1a8h_3_1_argbuf_r,
          q2a8i_2_1_argbuf_r,
          q3a8j_1_1_argbuf_r,
          call_$wmAdd_Int_goMux3_r} = (go_6_goMux_choice_2_r ? w1sif_1_goMux_mux_onehot :
                                       5'd0);
  
  /* mux (Ty C5,
     Ty Pointer_QTree_Int) : (go_6_goMux_choice_3,C5) [(call_$wmAdd_Int_goMux4,Pointer_QTree_Int),
                                                       (t3a8o_1_1_argbuf,Pointer_QTree_Int),
                                                       (t2a8n_2_1_argbuf,Pointer_QTree_Int),
                                                       (t1a8m_3_1_argbuf,Pointer_QTree_Int),
                                                       (t4a8p_1_argbuf,Pointer_QTree_Int)] > (w2sig_1_goMux_mux,Pointer_QTree_Int) */
  logic [16:0] w2sig_1_goMux_mux_mux;
  logic [4:0] w2sig_1_goMux_mux_onehot;
  always_comb
    unique case (go_6_goMux_choice_3_d[3:1])
      3'd0:
        {w2sig_1_goMux_mux_onehot, w2sig_1_goMux_mux_mux} = {5'd1,
                                                             call_$wmAdd_Int_goMux4_d};
      3'd1:
        {w2sig_1_goMux_mux_onehot, w2sig_1_goMux_mux_mux} = {5'd2,
                                                             t3a8o_1_1_argbuf_d};
      3'd2:
        {w2sig_1_goMux_mux_onehot, w2sig_1_goMux_mux_mux} = {5'd4,
                                                             t2a8n_2_1_argbuf_d};
      3'd3:
        {w2sig_1_goMux_mux_onehot, w2sig_1_goMux_mux_mux} = {5'd8,
                                                             t1a8m_3_1_argbuf_d};
      3'd4:
        {w2sig_1_goMux_mux_onehot, w2sig_1_goMux_mux_mux} = {5'd16,
                                                             t4a8p_1_argbuf_d};
      default:
        {w2sig_1_goMux_mux_onehot, w2sig_1_goMux_mux_mux} = {5'd0,
                                                             {16'd0, 1'd0}};
    endcase
  assign w2sig_1_goMux_mux_d = {w2sig_1_goMux_mux_mux[16:1],
                                (w2sig_1_goMux_mux_mux[0] && go_6_goMux_choice_3_d[0])};
  assign go_6_goMux_choice_3_r = (w2sig_1_goMux_mux_d[0] && w2sig_1_goMux_mux_r);
  assign {t4a8p_1_argbuf_r,
          t1a8m_3_1_argbuf_r,
          t2a8n_2_1_argbuf_r,
          t3a8o_1_1_argbuf_r,
          call_$wmAdd_Int_goMux4_r} = (go_6_goMux_choice_3_r ? w2sig_1_goMux_mux_onehot :
                                       5'd0);
  
  /* mux (Ty C5,
     Ty Pointer_CT$wmAdd_Int) : (go_6_goMux_choice_4,C5) [(call_$wmAdd_Int_goMux5,Pointer_CT$wmAdd_Int),
                                                          (sca2_1_argbuf,Pointer_CT$wmAdd_Int),
                                                          (sca1_1_argbuf,Pointer_CT$wmAdd_Int),
                                                          (sca0_1_argbuf,Pointer_CT$wmAdd_Int),
                                                          (sca3_1_argbuf,Pointer_CT$wmAdd_Int)] > (sc_0_goMux_mux,Pointer_CT$wmAdd_Int) */
  logic [16:0] sc_0_goMux_mux_mux;
  logic [4:0] sc_0_goMux_mux_onehot;
  always_comb
    unique case (go_6_goMux_choice_4_d[3:1])
      3'd0:
        {sc_0_goMux_mux_onehot, sc_0_goMux_mux_mux} = {5'd1,
                                                       call_$wmAdd_Int_goMux5_d};
      3'd1:
        {sc_0_goMux_mux_onehot, sc_0_goMux_mux_mux} = {5'd2,
                                                       sca2_1_argbuf_d};
      3'd2:
        {sc_0_goMux_mux_onehot, sc_0_goMux_mux_mux} = {5'd4,
                                                       sca1_1_argbuf_d};
      3'd3:
        {sc_0_goMux_mux_onehot, sc_0_goMux_mux_mux} = {5'd8,
                                                       sca0_1_argbuf_d};
      3'd4:
        {sc_0_goMux_mux_onehot, sc_0_goMux_mux_mux} = {5'd16,
                                                       sca3_1_argbuf_d};
      default:
        {sc_0_goMux_mux_onehot, sc_0_goMux_mux_mux} = {5'd0,
                                                       {16'd0, 1'd0}};
    endcase
  assign sc_0_goMux_mux_d = {sc_0_goMux_mux_mux[16:1],
                             (sc_0_goMux_mux_mux[0] && go_6_goMux_choice_4_d[0])};
  assign go_6_goMux_choice_4_r = (sc_0_goMux_mux_d[0] && sc_0_goMux_mux_r);
  assign {sca3_1_argbuf_r,
          sca0_1_argbuf_r,
          sca1_1_argbuf_r,
          sca2_1_argbuf_r,
          call_$wmAdd_Int_goMux5_r} = (go_6_goMux_choice_4_r ? sc_0_goMux_mux_onehot :
                                       5'd0);
  
  /* fork (Ty C5) : (go_7_goMux_choice,C5) > [(go_7_goMux_choice_1,C5),
                                         (go_7_goMux_choice_2,C5)] */
  logic [1:0] go_7_goMux_choice_emitted;
  logic [1:0] go_7_goMux_choice_done;
  assign go_7_goMux_choice_1_d = {go_7_goMux_choice_d[3:1],
                                  (go_7_goMux_choice_d[0] && (! go_7_goMux_choice_emitted[0]))};
  assign go_7_goMux_choice_2_d = {go_7_goMux_choice_d[3:1],
                                  (go_7_goMux_choice_d[0] && (! go_7_goMux_choice_emitted[1]))};
  assign go_7_goMux_choice_done = (go_7_goMux_choice_emitted | ({go_7_goMux_choice_2_d[0],
                                                                 go_7_goMux_choice_1_d[0]} & {go_7_goMux_choice_2_r,
                                                                                              go_7_goMux_choice_1_r}));
  assign go_7_goMux_choice_r = (& go_7_goMux_choice_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_7_goMux_choice_emitted <= 2'd0;
    else
      go_7_goMux_choice_emitted <= (go_7_goMux_choice_r ? 2'd0 :
                                    go_7_goMux_choice_done);
  
  /* mux (Ty C5,
     Ty Pointer_QTree_Int) : (go_7_goMux_choice_1,C5) [(call_$wnnz_Int_goMux2,Pointer_QTree_Int),
                                                       (q2a8D_1_1_argbuf,Pointer_QTree_Int),
                                                       (q3a8E_2_1_argbuf,Pointer_QTree_Int),
                                                       (q4a8F_3_1_argbuf,Pointer_QTree_Int),
                                                       (q1a8C_1_argbuf,Pointer_QTree_Int)] > (wsij_1_goMux_mux,Pointer_QTree_Int) */
  logic [16:0] wsij_1_goMux_mux_mux;
  logic [4:0] wsij_1_goMux_mux_onehot;
  always_comb
    unique case (go_7_goMux_choice_1_d[3:1])
      3'd0:
        {wsij_1_goMux_mux_onehot, wsij_1_goMux_mux_mux} = {5'd1,
                                                           call_$wnnz_Int_goMux2_d};
      3'd1:
        {wsij_1_goMux_mux_onehot, wsij_1_goMux_mux_mux} = {5'd2,
                                                           q2a8D_1_1_argbuf_d};
      3'd2:
        {wsij_1_goMux_mux_onehot, wsij_1_goMux_mux_mux} = {5'd4,
                                                           q3a8E_2_1_argbuf_d};
      3'd3:
        {wsij_1_goMux_mux_onehot, wsij_1_goMux_mux_mux} = {5'd8,
                                                           q4a8F_3_1_argbuf_d};
      3'd4:
        {wsij_1_goMux_mux_onehot, wsij_1_goMux_mux_mux} = {5'd16,
                                                           q1a8C_1_argbuf_d};
      default:
        {wsij_1_goMux_mux_onehot, wsij_1_goMux_mux_mux} = {5'd0,
                                                           {16'd0, 1'd0}};
    endcase
  assign wsij_1_goMux_mux_d = {wsij_1_goMux_mux_mux[16:1],
                               (wsij_1_goMux_mux_mux[0] && go_7_goMux_choice_1_d[0])};
  assign go_7_goMux_choice_1_r = (wsij_1_goMux_mux_d[0] && wsij_1_goMux_mux_r);
  assign {q1a8C_1_argbuf_r,
          q4a8F_3_1_argbuf_r,
          q3a8E_2_1_argbuf_r,
          q2a8D_1_1_argbuf_r,
          call_$wnnz_Int_goMux2_r} = (go_7_goMux_choice_1_r ? wsij_1_goMux_mux_onehot :
                                      5'd0);
  
  /* mux (Ty C5,
     Ty Pointer_CT$wnnz_Int) : (go_7_goMux_choice_2,C5) [(call_$wnnz_Int_goMux3,Pointer_CT$wnnz_Int),
                                                         (sca2_1_1_argbuf,Pointer_CT$wnnz_Int),
                                                         (sca1_1_1_argbuf,Pointer_CT$wnnz_Int),
                                                         (sca0_1_1_argbuf,Pointer_CT$wnnz_Int),
                                                         (sca3_1_1_argbuf,Pointer_CT$wnnz_Int)] > (sc_0_1_goMux_mux,Pointer_CT$wnnz_Int) */
  logic [16:0] sc_0_1_goMux_mux_mux;
  logic [4:0] sc_0_1_goMux_mux_onehot;
  always_comb
    unique case (go_7_goMux_choice_2_d[3:1])
      3'd0:
        {sc_0_1_goMux_mux_onehot, sc_0_1_goMux_mux_mux} = {5'd1,
                                                           call_$wnnz_Int_goMux3_d};
      3'd1:
        {sc_0_1_goMux_mux_onehot, sc_0_1_goMux_mux_mux} = {5'd2,
                                                           sca2_1_1_argbuf_d};
      3'd2:
        {sc_0_1_goMux_mux_onehot, sc_0_1_goMux_mux_mux} = {5'd4,
                                                           sca1_1_1_argbuf_d};
      3'd3:
        {sc_0_1_goMux_mux_onehot, sc_0_1_goMux_mux_mux} = {5'd8,
                                                           sca0_1_1_argbuf_d};
      3'd4:
        {sc_0_1_goMux_mux_onehot, sc_0_1_goMux_mux_mux} = {5'd16,
                                                           sca3_1_1_argbuf_d};
      default:
        {sc_0_1_goMux_mux_onehot, sc_0_1_goMux_mux_mux} = {5'd0,
                                                           {16'd0, 1'd0}};
    endcase
  assign sc_0_1_goMux_mux_d = {sc_0_1_goMux_mux_mux[16:1],
                               (sc_0_1_goMux_mux_mux[0] && go_7_goMux_choice_2_d[0])};
  assign go_7_goMux_choice_2_r = (sc_0_1_goMux_mux_d[0] && sc_0_1_goMux_mux_r);
  assign {sca3_1_1_argbuf_r,
          sca0_1_1_argbuf_r,
          sca1_1_1_argbuf_r,
          sca2_1_1_argbuf_r,
          call_$wnnz_Int_goMux3_r} = (go_7_goMux_choice_2_r ? sc_0_1_goMux_mux_onehot :
                                      5'd0);
  
  /* fork (Ty C5) : (go_8_goMux_choice,C5) > [(go_8_goMux_choice_1,C5),
                                         (go_8_goMux_choice_2,C5),
                                         (go_8_goMux_choice_3,C5)] */
  logic [2:0] go_8_goMux_choice_emitted;
  logic [2:0] go_8_goMux_choice_done;
  assign go_8_goMux_choice_1_d = {go_8_goMux_choice_d[3:1],
                                  (go_8_goMux_choice_d[0] && (! go_8_goMux_choice_emitted[0]))};
  assign go_8_goMux_choice_2_d = {go_8_goMux_choice_d[3:1],
                                  (go_8_goMux_choice_d[0] && (! go_8_goMux_choice_emitted[1]))};
  assign go_8_goMux_choice_3_d = {go_8_goMux_choice_d[3:1],
                                  (go_8_goMux_choice_d[0] && (! go_8_goMux_choice_emitted[2]))};
  assign go_8_goMux_choice_done = (go_8_goMux_choice_emitted | ({go_8_goMux_choice_3_d[0],
                                                                 go_8_goMux_choice_2_d[0],
                                                                 go_8_goMux_choice_1_d[0]} & {go_8_goMux_choice_3_r,
                                                                                              go_8_goMux_choice_2_r,
                                                                                              go_8_goMux_choice_1_r}));
  assign go_8_goMux_choice_r = (& go_8_goMux_choice_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_8_goMux_choice_emitted <= 3'd0;
    else
      go_8_goMux_choice_emitted <= (go_8_goMux_choice_r ? 3'd0 :
                                    go_8_goMux_choice_done);
  
  /* mux (Ty C5,
     Ty Pointer_QTree_Int) : (go_8_goMux_choice_1,C5) [(call_main_mask_Int_goMux2,Pointer_QTree_Int),
                                                       (t3a8z_1_1_argbuf,Pointer_QTree_Int),
                                                       (t2a8y_2_1_argbuf,Pointer_QTree_Int),
                                                       (t1a8x_3_1_argbuf,Pointer_QTree_Int),
                                                       (t4a8A_1_argbuf,Pointer_QTree_Int)] > (ma8q_goMux_mux,Pointer_QTree_Int) */
  logic [16:0] ma8q_goMux_mux_mux;
  logic [4:0] ma8q_goMux_mux_onehot;
  always_comb
    unique case (go_8_goMux_choice_1_d[3:1])
      3'd0:
        {ma8q_goMux_mux_onehot, ma8q_goMux_mux_mux} = {5'd1,
                                                       call_main_mask_Int_goMux2_d};
      3'd1:
        {ma8q_goMux_mux_onehot, ma8q_goMux_mux_mux} = {5'd2,
                                                       t3a8z_1_1_argbuf_d};
      3'd2:
        {ma8q_goMux_mux_onehot, ma8q_goMux_mux_mux} = {5'd4,
                                                       t2a8y_2_1_argbuf_d};
      3'd3:
        {ma8q_goMux_mux_onehot, ma8q_goMux_mux_mux} = {5'd8,
                                                       t1a8x_3_1_argbuf_d};
      3'd4:
        {ma8q_goMux_mux_onehot, ma8q_goMux_mux_mux} = {5'd16,
                                                       t4a8A_1_argbuf_d};
      default:
        {ma8q_goMux_mux_onehot, ma8q_goMux_mux_mux} = {5'd0,
                                                       {16'd0, 1'd0}};
    endcase
  assign ma8q_goMux_mux_d = {ma8q_goMux_mux_mux[16:1],
                             (ma8q_goMux_mux_mux[0] && go_8_goMux_choice_1_d[0])};
  assign go_8_goMux_choice_1_r = (ma8q_goMux_mux_d[0] && ma8q_goMux_mux_r);
  assign {t4a8A_1_argbuf_r,
          t1a8x_3_1_argbuf_r,
          t2a8y_2_1_argbuf_r,
          t3a8z_1_1_argbuf_r,
          call_main_mask_Int_goMux2_r} = (go_8_goMux_choice_1_r ? ma8q_goMux_mux_onehot :
                                          5'd0);
  
  /* mux (Ty C5,
     Ty Pointer_MaskQTree) : (go_8_goMux_choice_2,C5) [(call_main_mask_Int_goMux3,Pointer_MaskQTree),
                                                       (q3a8u_1_1_argbuf,Pointer_MaskQTree),
                                                       (q2a8t_2_1_argbuf,Pointer_MaskQTree),
                                                       (q1a8s_3_1_argbuf,Pointer_MaskQTree),
                                                       (lizzieLet14_1_4MQNode_8QNode_Int_1_argbuf,Pointer_MaskQTree)] > (mska8r_goMux_mux,Pointer_MaskQTree) */
  logic [16:0] mska8r_goMux_mux_mux;
  logic [4:0] mska8r_goMux_mux_onehot;
  always_comb
    unique case (go_8_goMux_choice_2_d[3:1])
      3'd0:
        {mska8r_goMux_mux_onehot, mska8r_goMux_mux_mux} = {5'd1,
                                                           call_main_mask_Int_goMux3_d};
      3'd1:
        {mska8r_goMux_mux_onehot, mska8r_goMux_mux_mux} = {5'd2,
                                                           q3a8u_1_1_argbuf_d};
      3'd2:
        {mska8r_goMux_mux_onehot, mska8r_goMux_mux_mux} = {5'd4,
                                                           q2a8t_2_1_argbuf_d};
      3'd3:
        {mska8r_goMux_mux_onehot, mska8r_goMux_mux_mux} = {5'd8,
                                                           q1a8s_3_1_argbuf_d};
      3'd4:
        {mska8r_goMux_mux_onehot, mska8r_goMux_mux_mux} = {5'd16,
                                                           lizzieLet14_1_4MQNode_8QNode_Int_1_argbuf_d};
      default:
        {mska8r_goMux_mux_onehot, mska8r_goMux_mux_mux} = {5'd0,
                                                           {16'd0, 1'd0}};
    endcase
  assign mska8r_goMux_mux_d = {mska8r_goMux_mux_mux[16:1],
                               (mska8r_goMux_mux_mux[0] && go_8_goMux_choice_2_d[0])};
  assign go_8_goMux_choice_2_r = (mska8r_goMux_mux_d[0] && mska8r_goMux_mux_r);
  assign {lizzieLet14_1_4MQNode_8QNode_Int_1_argbuf_r,
          q1a8s_3_1_argbuf_r,
          q2a8t_2_1_argbuf_r,
          q3a8u_1_1_argbuf_r,
          call_main_mask_Int_goMux3_r} = (go_8_goMux_choice_2_r ? mska8r_goMux_mux_onehot :
                                          5'd0);
  
  /* mux (Ty C5,
     Ty Pointer_CTmain_mask_Int) : (go_8_goMux_choice_3,C5) [(call_main_mask_Int_goMux4,Pointer_CTmain_mask_Int),
                                                             (sca2_2_1_argbuf,Pointer_CTmain_mask_Int),
                                                             (sca1_2_1_argbuf,Pointer_CTmain_mask_Int),
                                                             (sca0_2_1_argbuf,Pointer_CTmain_mask_Int),
                                                             (sca3_2_1_argbuf,Pointer_CTmain_mask_Int)] > (sc_0_2_goMux_mux,Pointer_CTmain_mask_Int) */
  logic [16:0] sc_0_2_goMux_mux_mux;
  logic [4:0] sc_0_2_goMux_mux_onehot;
  always_comb
    unique case (go_8_goMux_choice_3_d[3:1])
      3'd0:
        {sc_0_2_goMux_mux_onehot, sc_0_2_goMux_mux_mux} = {5'd1,
                                                           call_main_mask_Int_goMux4_d};
      3'd1:
        {sc_0_2_goMux_mux_onehot, sc_0_2_goMux_mux_mux} = {5'd2,
                                                           sca2_2_1_argbuf_d};
      3'd2:
        {sc_0_2_goMux_mux_onehot, sc_0_2_goMux_mux_mux} = {5'd4,
                                                           sca1_2_1_argbuf_d};
      3'd3:
        {sc_0_2_goMux_mux_onehot, sc_0_2_goMux_mux_mux} = {5'd8,
                                                           sca0_2_1_argbuf_d};
      3'd4:
        {sc_0_2_goMux_mux_onehot, sc_0_2_goMux_mux_mux} = {5'd16,
                                                           sca3_2_1_argbuf_d};
      default:
        {sc_0_2_goMux_mux_onehot, sc_0_2_goMux_mux_mux} = {5'd0,
                                                           {16'd0, 1'd0}};
    endcase
  assign sc_0_2_goMux_mux_d = {sc_0_2_goMux_mux_mux[16:1],
                               (sc_0_2_goMux_mux_mux[0] && go_8_goMux_choice_3_d[0])};
  assign go_8_goMux_choice_3_r = (sc_0_2_goMux_mux_d[0] && sc_0_2_goMux_mux_r);
  assign {sca3_2_1_argbuf_r,
          sca0_2_1_argbuf_r,
          sca1_2_1_argbuf_r,
          sca2_2_1_argbuf_r,
          call_main_mask_Int_goMux4_r} = (go_8_goMux_choice_3_r ? sc_0_2_goMux_mux_onehot :
                                          5'd0);
  
  /* dcon (Ty CTmain_mask_Int,
      Dcon Lmain_mask_Intsbos) : [(go_9_1,Go)] > (go_9_1Lmain_mask_Intsbos,CTmain_mask_Int) */
  assign go_9_1Lmain_mask_Intsbos_d = Lmain_mask_Intsbos_dc((& {go_9_1_d[0]}), go_9_1_d);
  assign {go_9_1_r} = {1 {(go_9_1Lmain_mask_Intsbos_r && go_9_1Lmain_mask_Intsbos_d[0])}};
  
  /* buf (Ty CTmain_mask_Int) : (go_9_1Lmain_mask_Intsbos,CTmain_mask_Int) > (lizzieLet21_1_argbuf,CTmain_mask_Int) */
  CTmain_mask_Int_t go_9_1Lmain_mask_Intsbos_bufchan_d;
  logic go_9_1Lmain_mask_Intsbos_bufchan_r;
  assign go_9_1Lmain_mask_Intsbos_r = ((! go_9_1Lmain_mask_Intsbos_bufchan_d[0]) || go_9_1Lmain_mask_Intsbos_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      go_9_1Lmain_mask_Intsbos_bufchan_d <= {115'd0, 1'd0};
    else
      if (go_9_1Lmain_mask_Intsbos_r)
        go_9_1Lmain_mask_Intsbos_bufchan_d <= go_9_1Lmain_mask_Intsbos_d;
  CTmain_mask_Int_t go_9_1Lmain_mask_Intsbos_bufchan_buf;
  assign go_9_1Lmain_mask_Intsbos_bufchan_r = (! go_9_1Lmain_mask_Intsbos_bufchan_buf[0]);
  assign lizzieLet21_1_argbuf_d = (go_9_1Lmain_mask_Intsbos_bufchan_buf[0] ? go_9_1Lmain_mask_Intsbos_bufchan_buf :
                                   go_9_1Lmain_mask_Intsbos_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      go_9_1Lmain_mask_Intsbos_bufchan_buf <= {115'd0, 1'd0};
    else
      if ((lizzieLet21_1_argbuf_r && go_9_1Lmain_mask_Intsbos_bufchan_buf[0]))
        go_9_1Lmain_mask_Intsbos_bufchan_buf <= {115'd0, 1'd0};
      else if (((! lizzieLet21_1_argbuf_r) && (! go_9_1Lmain_mask_Intsbos_bufchan_buf[0])))
        go_9_1Lmain_mask_Intsbos_bufchan_buf <= go_9_1Lmain_mask_Intsbos_bufchan_d;
  
  /* buf (Ty Go) : (go_9_2,Go) > (go_9_2_argbuf,Go) */
  Go_t go_9_2_bufchan_d;
  logic go_9_2_bufchan_r;
  assign go_9_2_r = ((! go_9_2_bufchan_d[0]) || go_9_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_9_2_bufchan_d <= 1'd0;
    else if (go_9_2_r) go_9_2_bufchan_d <= go_9_2_d;
  Go_t go_9_2_bufchan_buf;
  assign go_9_2_bufchan_r = (! go_9_2_bufchan_buf[0]);
  assign go_9_2_argbuf_d = (go_9_2_bufchan_buf[0] ? go_9_2_bufchan_buf :
                            go_9_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_9_2_bufchan_buf <= 1'd0;
    else
      if ((go_9_2_argbuf_r && go_9_2_bufchan_buf[0]))
        go_9_2_bufchan_buf <= 1'd0;
      else if (((! go_9_2_argbuf_r) && (! go_9_2_bufchan_buf[0])))
        go_9_2_bufchan_buf <= go_9_2_bufchan_d;
  
  /* dcon (Ty TupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Int,
      Dcon TupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Int) : [(go_9_2_argbuf,Go),
                                                                                       (ma8q_1_1_argbuf,Pointer_QTree_Int),
                                                                                       (mska8r_1_1_argbuf,Pointer_MaskQTree),
                                                                                       (lizzieLet4_1_1_argbuf,Pointer_CTmain_mask_Int)] > (call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Int_1,TupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Int) */
  assign call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Int_1_d = TupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Int_dc((& {go_9_2_argbuf_d[0],
                                                                                                                                                                                        ma8q_1_1_argbuf_d[0],
                                                                                                                                                                                        mska8r_1_1_argbuf_d[0],
                                                                                                                                                                                        lizzieLet4_1_1_argbuf_d[0]}), go_9_2_argbuf_d, ma8q_1_1_argbuf_d, mska8r_1_1_argbuf_d, lizzieLet4_1_1_argbuf_d);
  assign {go_9_2_argbuf_r,
          ma8q_1_1_argbuf_r,
          mska8r_1_1_argbuf_r,
          lizzieLet4_1_1_argbuf_r} = {4 {(call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Int_1_r && call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Int_1_d[0])}};
  
  /* destruct (Ty QTree_Int,
          Dcon QNode_Int) : (lizzieLet12_1_1QNode_Int,QTree_Int) > [(q1a8C_destruct,Pointer_QTree_Int),
                                                                    (q2a8D_destruct,Pointer_QTree_Int),
                                                                    (q3a8E_destruct,Pointer_QTree_Int),
                                                                    (q4a8F_destruct,Pointer_QTree_Int)] */
  logic [3:0] lizzieLet12_1_1QNode_Int_emitted;
  logic [3:0] lizzieLet12_1_1QNode_Int_done;
  assign q1a8C_destruct_d = {lizzieLet12_1_1QNode_Int_d[18:3],
                             (lizzieLet12_1_1QNode_Int_d[0] && (! lizzieLet12_1_1QNode_Int_emitted[0]))};
  assign q2a8D_destruct_d = {lizzieLet12_1_1QNode_Int_d[34:19],
                             (lizzieLet12_1_1QNode_Int_d[0] && (! lizzieLet12_1_1QNode_Int_emitted[1]))};
  assign q3a8E_destruct_d = {lizzieLet12_1_1QNode_Int_d[50:35],
                             (lizzieLet12_1_1QNode_Int_d[0] && (! lizzieLet12_1_1QNode_Int_emitted[2]))};
  assign q4a8F_destruct_d = {lizzieLet12_1_1QNode_Int_d[66:51],
                             (lizzieLet12_1_1QNode_Int_d[0] && (! lizzieLet12_1_1QNode_Int_emitted[3]))};
  assign lizzieLet12_1_1QNode_Int_done = (lizzieLet12_1_1QNode_Int_emitted | ({q4a8F_destruct_d[0],
                                                                               q3a8E_destruct_d[0],
                                                                               q2a8D_destruct_d[0],
                                                                               q1a8C_destruct_d[0]} & {q4a8F_destruct_r,
                                                                                                       q3a8E_destruct_r,
                                                                                                       q2a8D_destruct_r,
                                                                                                       q1a8C_destruct_r}));
  assign lizzieLet12_1_1QNode_Int_r = (& lizzieLet12_1_1QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet12_1_1QNode_Int_emitted <= 4'd0;
    else
      lizzieLet12_1_1QNode_Int_emitted <= (lizzieLet12_1_1QNode_Int_r ? 4'd0 :
                                           lizzieLet12_1_1QNode_Int_done);
  
  /* demux (Ty QTree_Int,
       Ty QTree_Int) : (lizzieLet12_1_2,QTree_Int) (lizzieLet12_1_1,QTree_Int) > [(_73,QTree_Int),
                                                                                  (_72,QTree_Int),
                                                                                  (lizzieLet12_1_1QNode_Int,QTree_Int),
                                                                                  (_71,QTree_Int)] */
  logic [3:0] lizzieLet12_1_1_onehotd;
  always_comb
    if ((lizzieLet12_1_2_d[0] && lizzieLet12_1_1_d[0]))
      unique case (lizzieLet12_1_2_d[2:1])
        2'd0: lizzieLet12_1_1_onehotd = 4'd1;
        2'd1: lizzieLet12_1_1_onehotd = 4'd2;
        2'd2: lizzieLet12_1_1_onehotd = 4'd4;
        2'd3: lizzieLet12_1_1_onehotd = 4'd8;
        default: lizzieLet12_1_1_onehotd = 4'd0;
      endcase
    else lizzieLet12_1_1_onehotd = 4'd0;
  assign _73_d = {lizzieLet12_1_1_d[66:1],
                  lizzieLet12_1_1_onehotd[0]};
  assign _72_d = {lizzieLet12_1_1_d[66:1],
                  lizzieLet12_1_1_onehotd[1]};
  assign lizzieLet12_1_1QNode_Int_d = {lizzieLet12_1_1_d[66:1],
                                       lizzieLet12_1_1_onehotd[2]};
  assign _71_d = {lizzieLet12_1_1_d[66:1],
                  lizzieLet12_1_1_onehotd[3]};
  assign lizzieLet12_1_1_r = (| (lizzieLet12_1_1_onehotd & {_71_r,
                                                            lizzieLet12_1_1QNode_Int_r,
                                                            _72_r,
                                                            _73_r}));
  assign lizzieLet12_1_2_r = lizzieLet12_1_1_r;
  
  /* demux (Ty QTree_Int,
       Ty Go) : (lizzieLet12_1_3,QTree_Int) (go_7_goMux_data,Go) > [(lizzieLet12_1_3QNone_Int,Go),
                                                                    (lizzieLet12_1_3QVal_Int,Go),
                                                                    (lizzieLet12_1_3QNode_Int,Go),
                                                                    (lizzieLet12_1_3QError_Int,Go)] */
  logic [3:0] go_7_goMux_data_onehotd;
  always_comb
    if ((lizzieLet12_1_3_d[0] && go_7_goMux_data_d[0]))
      unique case (lizzieLet12_1_3_d[2:1])
        2'd0: go_7_goMux_data_onehotd = 4'd1;
        2'd1: go_7_goMux_data_onehotd = 4'd2;
        2'd2: go_7_goMux_data_onehotd = 4'd4;
        2'd3: go_7_goMux_data_onehotd = 4'd8;
        default: go_7_goMux_data_onehotd = 4'd0;
      endcase
    else go_7_goMux_data_onehotd = 4'd0;
  assign lizzieLet12_1_3QNone_Int_d = go_7_goMux_data_onehotd[0];
  assign lizzieLet12_1_3QVal_Int_d = go_7_goMux_data_onehotd[1];
  assign lizzieLet12_1_3QNode_Int_d = go_7_goMux_data_onehotd[2];
  assign lizzieLet12_1_3QError_Int_d = go_7_goMux_data_onehotd[3];
  assign go_7_goMux_data_r = (| (go_7_goMux_data_onehotd & {lizzieLet12_1_3QError_Int_r,
                                                            lizzieLet12_1_3QNode_Int_r,
                                                            lizzieLet12_1_3QVal_Int_r,
                                                            lizzieLet12_1_3QNone_Int_r}));
  assign lizzieLet12_1_3_r = go_7_goMux_data_r;
  
  /* fork (Ty Go) : (lizzieLet12_1_3QError_Int,Go) > [(lizzieLet12_1_3QError_Int_1,Go),
                                                 (lizzieLet12_1_3QError_Int_2,Go)] */
  logic [1:0] lizzieLet12_1_3QError_Int_emitted;
  logic [1:0] lizzieLet12_1_3QError_Int_done;
  assign lizzieLet12_1_3QError_Int_1_d = (lizzieLet12_1_3QError_Int_d[0] && (! lizzieLet12_1_3QError_Int_emitted[0]));
  assign lizzieLet12_1_3QError_Int_2_d = (lizzieLet12_1_3QError_Int_d[0] && (! lizzieLet12_1_3QError_Int_emitted[1]));
  assign lizzieLet12_1_3QError_Int_done = (lizzieLet12_1_3QError_Int_emitted | ({lizzieLet12_1_3QError_Int_2_d[0],
                                                                                 lizzieLet12_1_3QError_Int_1_d[0]} & {lizzieLet12_1_3QError_Int_2_r,
                                                                                                                      lizzieLet12_1_3QError_Int_1_r}));
  assign lizzieLet12_1_3QError_Int_r = (& lizzieLet12_1_3QError_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet12_1_3QError_Int_emitted <= 2'd0;
    else
      lizzieLet12_1_3QError_Int_emitted <= (lizzieLet12_1_3QError_Int_r ? 2'd0 :
                                            lizzieLet12_1_3QError_Int_done);
  
  /* buf (Ty Go) : (lizzieLet12_1_3QError_Int_1,Go) > (lizzieLet12_1_3QError_Int_1_argbuf,Go) */
  Go_t lizzieLet12_1_3QError_Int_1_bufchan_d;
  logic lizzieLet12_1_3QError_Int_1_bufchan_r;
  assign lizzieLet12_1_3QError_Int_1_r = ((! lizzieLet12_1_3QError_Int_1_bufchan_d[0]) || lizzieLet12_1_3QError_Int_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet12_1_3QError_Int_1_bufchan_d <= 1'd0;
    else
      if (lizzieLet12_1_3QError_Int_1_r)
        lizzieLet12_1_3QError_Int_1_bufchan_d <= lizzieLet12_1_3QError_Int_1_d;
  Go_t lizzieLet12_1_3QError_Int_1_bufchan_buf;
  assign lizzieLet12_1_3QError_Int_1_bufchan_r = (! lizzieLet12_1_3QError_Int_1_bufchan_buf[0]);
  assign lizzieLet12_1_3QError_Int_1_argbuf_d = (lizzieLet12_1_3QError_Int_1_bufchan_buf[0] ? lizzieLet12_1_3QError_Int_1_bufchan_buf :
                                                 lizzieLet12_1_3QError_Int_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_1_3QError_Int_1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet12_1_3QError_Int_1_argbuf_r && lizzieLet12_1_3QError_Int_1_bufchan_buf[0]))
        lizzieLet12_1_3QError_Int_1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet12_1_3QError_Int_1_argbuf_r) && (! lizzieLet12_1_3QError_Int_1_bufchan_buf[0])))
        lizzieLet12_1_3QError_Int_1_bufchan_buf <= lizzieLet12_1_3QError_Int_1_bufchan_d;
  
  /* const (Ty Int#,
       Lit 0) : (lizzieLet12_1_3QError_Int_1_argbuf,Go) > (lizzieLet12_1_3QError_Int_1_argbuf_0,Int#) */
  assign lizzieLet12_1_3QError_Int_1_argbuf_0_d = {32'd0,
                                                   lizzieLet12_1_3QError_Int_1_argbuf_d[0]};
  assign lizzieLet12_1_3QError_Int_1_argbuf_r = lizzieLet12_1_3QError_Int_1_argbuf_0_r;
  
  /* buf (Ty Int#) : (lizzieLet12_1_3QError_Int_1_argbuf_0,Int#) > (lizzieLet5_2_1_argbuf,Int#) */
  \Int#_t  lizzieLet12_1_3QError_Int_1_argbuf_0_bufchan_d;
  logic lizzieLet12_1_3QError_Int_1_argbuf_0_bufchan_r;
  assign lizzieLet12_1_3QError_Int_1_argbuf_0_r = ((! lizzieLet12_1_3QError_Int_1_argbuf_0_bufchan_d[0]) || lizzieLet12_1_3QError_Int_1_argbuf_0_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_1_3QError_Int_1_argbuf_0_bufchan_d <= {32'd0, 1'd0};
    else
      if (lizzieLet12_1_3QError_Int_1_argbuf_0_r)
        lizzieLet12_1_3QError_Int_1_argbuf_0_bufchan_d <= lizzieLet12_1_3QError_Int_1_argbuf_0_d;
  \Int#_t  lizzieLet12_1_3QError_Int_1_argbuf_0_bufchan_buf;
  assign lizzieLet12_1_3QError_Int_1_argbuf_0_bufchan_r = (! lizzieLet12_1_3QError_Int_1_argbuf_0_bufchan_buf[0]);
  assign lizzieLet5_2_1_argbuf_d = (lizzieLet12_1_3QError_Int_1_argbuf_0_bufchan_buf[0] ? lizzieLet12_1_3QError_Int_1_argbuf_0_bufchan_buf :
                                    lizzieLet12_1_3QError_Int_1_argbuf_0_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_1_3QError_Int_1_argbuf_0_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((lizzieLet5_2_1_argbuf_r && lizzieLet12_1_3QError_Int_1_argbuf_0_bufchan_buf[0]))
        lizzieLet12_1_3QError_Int_1_argbuf_0_bufchan_buf <= {32'd0, 1'd0};
      else if (((! lizzieLet5_2_1_argbuf_r) && (! lizzieLet12_1_3QError_Int_1_argbuf_0_bufchan_buf[0])))
        lizzieLet12_1_3QError_Int_1_argbuf_0_bufchan_buf <= lizzieLet12_1_3QError_Int_1_argbuf_0_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet12_1_3QError_Int_2,Go) > (lizzieLet12_1_3QError_Int_2_argbuf,Go) */
  Go_t lizzieLet12_1_3QError_Int_2_bufchan_d;
  logic lizzieLet12_1_3QError_Int_2_bufchan_r;
  assign lizzieLet12_1_3QError_Int_2_r = ((! lizzieLet12_1_3QError_Int_2_bufchan_d[0]) || lizzieLet12_1_3QError_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet12_1_3QError_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet12_1_3QError_Int_2_r)
        lizzieLet12_1_3QError_Int_2_bufchan_d <= lizzieLet12_1_3QError_Int_2_d;
  Go_t lizzieLet12_1_3QError_Int_2_bufchan_buf;
  assign lizzieLet12_1_3QError_Int_2_bufchan_r = (! lizzieLet12_1_3QError_Int_2_bufchan_buf[0]);
  assign lizzieLet12_1_3QError_Int_2_argbuf_d = (lizzieLet12_1_3QError_Int_2_bufchan_buf[0] ? lizzieLet12_1_3QError_Int_2_bufchan_buf :
                                                 lizzieLet12_1_3QError_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_1_3QError_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet12_1_3QError_Int_2_argbuf_r && lizzieLet12_1_3QError_Int_2_bufchan_buf[0]))
        lizzieLet12_1_3QError_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet12_1_3QError_Int_2_argbuf_r) && (! lizzieLet12_1_3QError_Int_2_bufchan_buf[0])))
        lizzieLet12_1_3QError_Int_2_bufchan_buf <= lizzieLet12_1_3QError_Int_2_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet12_1_3QNode_Int,Go) > (lizzieLet12_1_3QNode_Int_1_argbuf,Go) */
  Go_t lizzieLet12_1_3QNode_Int_bufchan_d;
  logic lizzieLet12_1_3QNode_Int_bufchan_r;
  assign lizzieLet12_1_3QNode_Int_r = ((! lizzieLet12_1_3QNode_Int_bufchan_d[0]) || lizzieLet12_1_3QNode_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet12_1_3QNode_Int_bufchan_d <= 1'd0;
    else
      if (lizzieLet12_1_3QNode_Int_r)
        lizzieLet12_1_3QNode_Int_bufchan_d <= lizzieLet12_1_3QNode_Int_d;
  Go_t lizzieLet12_1_3QNode_Int_bufchan_buf;
  assign lizzieLet12_1_3QNode_Int_bufchan_r = (! lizzieLet12_1_3QNode_Int_bufchan_buf[0]);
  assign lizzieLet12_1_3QNode_Int_1_argbuf_d = (lizzieLet12_1_3QNode_Int_bufchan_buf[0] ? lizzieLet12_1_3QNode_Int_bufchan_buf :
                                                lizzieLet12_1_3QNode_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet12_1_3QNode_Int_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet12_1_3QNode_Int_1_argbuf_r && lizzieLet12_1_3QNode_Int_bufchan_buf[0]))
        lizzieLet12_1_3QNode_Int_bufchan_buf <= 1'd0;
      else if (((! lizzieLet12_1_3QNode_Int_1_argbuf_r) && (! lizzieLet12_1_3QNode_Int_bufchan_buf[0])))
        lizzieLet12_1_3QNode_Int_bufchan_buf <= lizzieLet12_1_3QNode_Int_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet12_1_3QNone_Int,Go) > [(lizzieLet12_1_3QNone_Int_1,Go),
                                                (lizzieLet12_1_3QNone_Int_2,Go)] */
  logic [1:0] lizzieLet12_1_3QNone_Int_emitted;
  logic [1:0] lizzieLet12_1_3QNone_Int_done;
  assign lizzieLet12_1_3QNone_Int_1_d = (lizzieLet12_1_3QNone_Int_d[0] && (! lizzieLet12_1_3QNone_Int_emitted[0]));
  assign lizzieLet12_1_3QNone_Int_2_d = (lizzieLet12_1_3QNone_Int_d[0] && (! lizzieLet12_1_3QNone_Int_emitted[1]));
  assign lizzieLet12_1_3QNone_Int_done = (lizzieLet12_1_3QNone_Int_emitted | ({lizzieLet12_1_3QNone_Int_2_d[0],
                                                                               lizzieLet12_1_3QNone_Int_1_d[0]} & {lizzieLet12_1_3QNone_Int_2_r,
                                                                                                                   lizzieLet12_1_3QNone_Int_1_r}));
  assign lizzieLet12_1_3QNone_Int_r = (& lizzieLet12_1_3QNone_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet12_1_3QNone_Int_emitted <= 2'd0;
    else
      lizzieLet12_1_3QNone_Int_emitted <= (lizzieLet12_1_3QNone_Int_r ? 2'd0 :
                                           lizzieLet12_1_3QNone_Int_done);
  
  /* buf (Ty Go) : (lizzieLet12_1_3QNone_Int_1,Go) > (lizzieLet12_1_3QNone_Int_1_argbuf,Go) */
  Go_t lizzieLet12_1_3QNone_Int_1_bufchan_d;
  logic lizzieLet12_1_3QNone_Int_1_bufchan_r;
  assign lizzieLet12_1_3QNone_Int_1_r = ((! lizzieLet12_1_3QNone_Int_1_bufchan_d[0]) || lizzieLet12_1_3QNone_Int_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet12_1_3QNone_Int_1_bufchan_d <= 1'd0;
    else
      if (lizzieLet12_1_3QNone_Int_1_r)
        lizzieLet12_1_3QNone_Int_1_bufchan_d <= lizzieLet12_1_3QNone_Int_1_d;
  Go_t lizzieLet12_1_3QNone_Int_1_bufchan_buf;
  assign lizzieLet12_1_3QNone_Int_1_bufchan_r = (! lizzieLet12_1_3QNone_Int_1_bufchan_buf[0]);
  assign lizzieLet12_1_3QNone_Int_1_argbuf_d = (lizzieLet12_1_3QNone_Int_1_bufchan_buf[0] ? lizzieLet12_1_3QNone_Int_1_bufchan_buf :
                                                lizzieLet12_1_3QNone_Int_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_1_3QNone_Int_1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet12_1_3QNone_Int_1_argbuf_r && lizzieLet12_1_3QNone_Int_1_bufchan_buf[0]))
        lizzieLet12_1_3QNone_Int_1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet12_1_3QNone_Int_1_argbuf_r) && (! lizzieLet12_1_3QNone_Int_1_bufchan_buf[0])))
        lizzieLet12_1_3QNone_Int_1_bufchan_buf <= lizzieLet12_1_3QNone_Int_1_bufchan_d;
  
  /* const (Ty Int#,
       Lit 0) : (lizzieLet12_1_3QNone_Int_1_argbuf,Go) > (lizzieLet12_1_3QNone_Int_1_argbuf_0,Int#) */
  assign lizzieLet12_1_3QNone_Int_1_argbuf_0_d = {32'd0,
                                                  lizzieLet12_1_3QNone_Int_1_argbuf_d[0]};
  assign lizzieLet12_1_3QNone_Int_1_argbuf_r = lizzieLet12_1_3QNone_Int_1_argbuf_0_r;
  
  /* buf (Ty Int#) : (lizzieLet12_1_3QNone_Int_1_argbuf_0,Int#) > (lizzieLet5_1_1_argbuf,Int#) */
  \Int#_t  lizzieLet12_1_3QNone_Int_1_argbuf_0_bufchan_d;
  logic lizzieLet12_1_3QNone_Int_1_argbuf_0_bufchan_r;
  assign lizzieLet12_1_3QNone_Int_1_argbuf_0_r = ((! lizzieLet12_1_3QNone_Int_1_argbuf_0_bufchan_d[0]) || lizzieLet12_1_3QNone_Int_1_argbuf_0_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_1_3QNone_Int_1_argbuf_0_bufchan_d <= {32'd0, 1'd0};
    else
      if (lizzieLet12_1_3QNone_Int_1_argbuf_0_r)
        lizzieLet12_1_3QNone_Int_1_argbuf_0_bufchan_d <= lizzieLet12_1_3QNone_Int_1_argbuf_0_d;
  \Int#_t  lizzieLet12_1_3QNone_Int_1_argbuf_0_bufchan_buf;
  assign lizzieLet12_1_3QNone_Int_1_argbuf_0_bufchan_r = (! lizzieLet12_1_3QNone_Int_1_argbuf_0_bufchan_buf[0]);
  assign lizzieLet5_1_1_argbuf_d = (lizzieLet12_1_3QNone_Int_1_argbuf_0_bufchan_buf[0] ? lizzieLet12_1_3QNone_Int_1_argbuf_0_bufchan_buf :
                                    lizzieLet12_1_3QNone_Int_1_argbuf_0_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_1_3QNone_Int_1_argbuf_0_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((lizzieLet5_1_1_argbuf_r && lizzieLet12_1_3QNone_Int_1_argbuf_0_bufchan_buf[0]))
        lizzieLet12_1_3QNone_Int_1_argbuf_0_bufchan_buf <= {32'd0, 1'd0};
      else if (((! lizzieLet5_1_1_argbuf_r) && (! lizzieLet12_1_3QNone_Int_1_argbuf_0_bufchan_buf[0])))
        lizzieLet12_1_3QNone_Int_1_argbuf_0_bufchan_buf <= lizzieLet12_1_3QNone_Int_1_argbuf_0_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet12_1_3QNone_Int_2,Go) > (lizzieLet12_1_3QNone_Int_2_argbuf,Go) */
  Go_t lizzieLet12_1_3QNone_Int_2_bufchan_d;
  logic lizzieLet12_1_3QNone_Int_2_bufchan_r;
  assign lizzieLet12_1_3QNone_Int_2_r = ((! lizzieLet12_1_3QNone_Int_2_bufchan_d[0]) || lizzieLet12_1_3QNone_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet12_1_3QNone_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet12_1_3QNone_Int_2_r)
        lizzieLet12_1_3QNone_Int_2_bufchan_d <= lizzieLet12_1_3QNone_Int_2_d;
  Go_t lizzieLet12_1_3QNone_Int_2_bufchan_buf;
  assign lizzieLet12_1_3QNone_Int_2_bufchan_r = (! lizzieLet12_1_3QNone_Int_2_bufchan_buf[0]);
  assign lizzieLet12_1_3QNone_Int_2_argbuf_d = (lizzieLet12_1_3QNone_Int_2_bufchan_buf[0] ? lizzieLet12_1_3QNone_Int_2_bufchan_buf :
                                                lizzieLet12_1_3QNone_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_1_3QNone_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet12_1_3QNone_Int_2_argbuf_r && lizzieLet12_1_3QNone_Int_2_bufchan_buf[0]))
        lizzieLet12_1_3QNone_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet12_1_3QNone_Int_2_argbuf_r) && (! lizzieLet12_1_3QNone_Int_2_bufchan_buf[0])))
        lizzieLet12_1_3QNone_Int_2_bufchan_buf <= lizzieLet12_1_3QNone_Int_2_bufchan_d;
  
  /* mergectrl (Ty C4,Ty Go) : [(lizzieLet12_1_3QNone_Int_2_argbuf,Go),
                           (lizzieLet27_3Lcall_$wnnz_Int0_1_argbuf,Go),
                           (lizzieLet12_1_3QVal_Int_2_argbuf,Go),
                           (lizzieLet12_1_3QError_Int_2_argbuf,Go)] > (go_11_goMux_choice,C4) (go_11_goMux_data,Go) */
  logic [3:0] lizzieLet12_1_3QNone_Int_2_argbuf_select_d;
  assign lizzieLet12_1_3QNone_Int_2_argbuf_select_d = ((| lizzieLet12_1_3QNone_Int_2_argbuf_select_q) ? lizzieLet12_1_3QNone_Int_2_argbuf_select_q :
                                                       (lizzieLet12_1_3QNone_Int_2_argbuf_d[0] ? 4'd1 :
                                                        (lizzieLet27_3Lcall_$wnnz_Int0_1_argbuf_d[0] ? 4'd2 :
                                                         (lizzieLet12_1_3QVal_Int_2_argbuf_d[0] ? 4'd4 :
                                                          (lizzieLet12_1_3QError_Int_2_argbuf_d[0] ? 4'd8 :
                                                           4'd0)))));
  logic [3:0] lizzieLet12_1_3QNone_Int_2_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_1_3QNone_Int_2_argbuf_select_q <= 4'd0;
    else
      lizzieLet12_1_3QNone_Int_2_argbuf_select_q <= (lizzieLet12_1_3QNone_Int_2_argbuf_done ? 4'd0 :
                                                     lizzieLet12_1_3QNone_Int_2_argbuf_select_d);
  logic [1:0] lizzieLet12_1_3QNone_Int_2_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_1_3QNone_Int_2_argbuf_emit_q <= 2'd0;
    else
      lizzieLet12_1_3QNone_Int_2_argbuf_emit_q <= (lizzieLet12_1_3QNone_Int_2_argbuf_done ? 2'd0 :
                                                   lizzieLet12_1_3QNone_Int_2_argbuf_emit_d);
  logic [1:0] lizzieLet12_1_3QNone_Int_2_argbuf_emit_d;
  assign lizzieLet12_1_3QNone_Int_2_argbuf_emit_d = (lizzieLet12_1_3QNone_Int_2_argbuf_emit_q | ({go_11_goMux_choice_d[0],
                                                                                                  go_11_goMux_data_d[0]} & {go_11_goMux_choice_r,
                                                                                                                            go_11_goMux_data_r}));
  logic lizzieLet12_1_3QNone_Int_2_argbuf_done;
  assign lizzieLet12_1_3QNone_Int_2_argbuf_done = (& lizzieLet12_1_3QNone_Int_2_argbuf_emit_d);
  assign {lizzieLet12_1_3QError_Int_2_argbuf_r,
          lizzieLet12_1_3QVal_Int_2_argbuf_r,
          lizzieLet27_3Lcall_$wnnz_Int0_1_argbuf_r,
          lizzieLet12_1_3QNone_Int_2_argbuf_r} = (lizzieLet12_1_3QNone_Int_2_argbuf_done ? lizzieLet12_1_3QNone_Int_2_argbuf_select_d :
                                                  4'd0);
  assign go_11_goMux_data_d = ((lizzieLet12_1_3QNone_Int_2_argbuf_select_d[0] && (! lizzieLet12_1_3QNone_Int_2_argbuf_emit_q[0])) ? lizzieLet12_1_3QNone_Int_2_argbuf_d :
                               ((lizzieLet12_1_3QNone_Int_2_argbuf_select_d[1] && (! lizzieLet12_1_3QNone_Int_2_argbuf_emit_q[0])) ? lizzieLet27_3Lcall_$wnnz_Int0_1_argbuf_d :
                                ((lizzieLet12_1_3QNone_Int_2_argbuf_select_d[2] && (! lizzieLet12_1_3QNone_Int_2_argbuf_emit_q[0])) ? lizzieLet12_1_3QVal_Int_2_argbuf_d :
                                 ((lizzieLet12_1_3QNone_Int_2_argbuf_select_d[3] && (! lizzieLet12_1_3QNone_Int_2_argbuf_emit_q[0])) ? lizzieLet12_1_3QError_Int_2_argbuf_d :
                                  1'd0))));
  assign go_11_goMux_choice_d = ((lizzieLet12_1_3QNone_Int_2_argbuf_select_d[0] && (! lizzieLet12_1_3QNone_Int_2_argbuf_emit_q[1])) ? C1_4_dc(1'd1) :
                                 ((lizzieLet12_1_3QNone_Int_2_argbuf_select_d[1] && (! lizzieLet12_1_3QNone_Int_2_argbuf_emit_q[1])) ? C2_4_dc(1'd1) :
                                  ((lizzieLet12_1_3QNone_Int_2_argbuf_select_d[2] && (! lizzieLet12_1_3QNone_Int_2_argbuf_emit_q[1])) ? C3_4_dc(1'd1) :
                                   ((lizzieLet12_1_3QNone_Int_2_argbuf_select_d[3] && (! lizzieLet12_1_3QNone_Int_2_argbuf_emit_q[1])) ? C4_4_dc(1'd1) :
                                    {2'd0, 1'd0}))));
  
  /* fork (Ty Go) : (lizzieLet12_1_3QVal_Int,Go) > [(lizzieLet12_1_3QVal_Int_1,Go),
                                               (lizzieLet12_1_3QVal_Int_2,Go)] */
  logic [1:0] lizzieLet12_1_3QVal_Int_emitted;
  logic [1:0] lizzieLet12_1_3QVal_Int_done;
  assign lizzieLet12_1_3QVal_Int_1_d = (lizzieLet12_1_3QVal_Int_d[0] && (! lizzieLet12_1_3QVal_Int_emitted[0]));
  assign lizzieLet12_1_3QVal_Int_2_d = (lizzieLet12_1_3QVal_Int_d[0] && (! lizzieLet12_1_3QVal_Int_emitted[1]));
  assign lizzieLet12_1_3QVal_Int_done = (lizzieLet12_1_3QVal_Int_emitted | ({lizzieLet12_1_3QVal_Int_2_d[0],
                                                                             lizzieLet12_1_3QVal_Int_1_d[0]} & {lizzieLet12_1_3QVal_Int_2_r,
                                                                                                                lizzieLet12_1_3QVal_Int_1_r}));
  assign lizzieLet12_1_3QVal_Int_r = (& lizzieLet12_1_3QVal_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet12_1_3QVal_Int_emitted <= 2'd0;
    else
      lizzieLet12_1_3QVal_Int_emitted <= (lizzieLet12_1_3QVal_Int_r ? 2'd0 :
                                          lizzieLet12_1_3QVal_Int_done);
  
  /* buf (Ty Go) : (lizzieLet12_1_3QVal_Int_1,Go) > (lizzieLet12_1_3QVal_Int_1_argbuf,Go) */
  Go_t lizzieLet12_1_3QVal_Int_1_bufchan_d;
  logic lizzieLet12_1_3QVal_Int_1_bufchan_r;
  assign lizzieLet12_1_3QVal_Int_1_r = ((! lizzieLet12_1_3QVal_Int_1_bufchan_d[0]) || lizzieLet12_1_3QVal_Int_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet12_1_3QVal_Int_1_bufchan_d <= 1'd0;
    else
      if (lizzieLet12_1_3QVal_Int_1_r)
        lizzieLet12_1_3QVal_Int_1_bufchan_d <= lizzieLet12_1_3QVal_Int_1_d;
  Go_t lizzieLet12_1_3QVal_Int_1_bufchan_buf;
  assign lizzieLet12_1_3QVal_Int_1_bufchan_r = (! lizzieLet12_1_3QVal_Int_1_bufchan_buf[0]);
  assign lizzieLet12_1_3QVal_Int_1_argbuf_d = (lizzieLet12_1_3QVal_Int_1_bufchan_buf[0] ? lizzieLet12_1_3QVal_Int_1_bufchan_buf :
                                               lizzieLet12_1_3QVal_Int_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet12_1_3QVal_Int_1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet12_1_3QVal_Int_1_argbuf_r && lizzieLet12_1_3QVal_Int_1_bufchan_buf[0]))
        lizzieLet12_1_3QVal_Int_1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet12_1_3QVal_Int_1_argbuf_r) && (! lizzieLet12_1_3QVal_Int_1_bufchan_buf[0])))
        lizzieLet12_1_3QVal_Int_1_bufchan_buf <= lizzieLet12_1_3QVal_Int_1_bufchan_d;
  
  /* const (Ty Int#,
       Lit 1) : (lizzieLet12_1_3QVal_Int_1_argbuf,Go) > (lizzieLet12_1_3QVal_Int_1_argbuf_1,Int#) */
  assign lizzieLet12_1_3QVal_Int_1_argbuf_1_d = {32'd1,
                                                 lizzieLet12_1_3QVal_Int_1_argbuf_d[0]};
  assign lizzieLet12_1_3QVal_Int_1_argbuf_r = lizzieLet12_1_3QVal_Int_1_argbuf_1_r;
  
  /* buf (Ty Int#) : (lizzieLet12_1_3QVal_Int_1_argbuf_1,Int#) > (lizzieLet6_1_1_argbuf,Int#) */
  \Int#_t  lizzieLet12_1_3QVal_Int_1_argbuf_1_bufchan_d;
  logic lizzieLet12_1_3QVal_Int_1_argbuf_1_bufchan_r;
  assign lizzieLet12_1_3QVal_Int_1_argbuf_1_r = ((! lizzieLet12_1_3QVal_Int_1_argbuf_1_bufchan_d[0]) || lizzieLet12_1_3QVal_Int_1_argbuf_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_1_3QVal_Int_1_argbuf_1_bufchan_d <= {32'd0, 1'd0};
    else
      if (lizzieLet12_1_3QVal_Int_1_argbuf_1_r)
        lizzieLet12_1_3QVal_Int_1_argbuf_1_bufchan_d <= lizzieLet12_1_3QVal_Int_1_argbuf_1_d;
  \Int#_t  lizzieLet12_1_3QVal_Int_1_argbuf_1_bufchan_buf;
  assign lizzieLet12_1_3QVal_Int_1_argbuf_1_bufchan_r = (! lizzieLet12_1_3QVal_Int_1_argbuf_1_bufchan_buf[0]);
  assign lizzieLet6_1_1_argbuf_d = (lizzieLet12_1_3QVal_Int_1_argbuf_1_bufchan_buf[0] ? lizzieLet12_1_3QVal_Int_1_argbuf_1_bufchan_buf :
                                    lizzieLet12_1_3QVal_Int_1_argbuf_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_1_3QVal_Int_1_argbuf_1_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((lizzieLet6_1_1_argbuf_r && lizzieLet12_1_3QVal_Int_1_argbuf_1_bufchan_buf[0]))
        lizzieLet12_1_3QVal_Int_1_argbuf_1_bufchan_buf <= {32'd0, 1'd0};
      else if (((! lizzieLet6_1_1_argbuf_r) && (! lizzieLet12_1_3QVal_Int_1_argbuf_1_bufchan_buf[0])))
        lizzieLet12_1_3QVal_Int_1_argbuf_1_bufchan_buf <= lizzieLet12_1_3QVal_Int_1_argbuf_1_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet12_1_3QVal_Int_2,Go) > (lizzieLet12_1_3QVal_Int_2_argbuf,Go) */
  Go_t lizzieLet12_1_3QVal_Int_2_bufchan_d;
  logic lizzieLet12_1_3QVal_Int_2_bufchan_r;
  assign lizzieLet12_1_3QVal_Int_2_r = ((! lizzieLet12_1_3QVal_Int_2_bufchan_d[0]) || lizzieLet12_1_3QVal_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet12_1_3QVal_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet12_1_3QVal_Int_2_r)
        lizzieLet12_1_3QVal_Int_2_bufchan_d <= lizzieLet12_1_3QVal_Int_2_d;
  Go_t lizzieLet12_1_3QVal_Int_2_bufchan_buf;
  assign lizzieLet12_1_3QVal_Int_2_bufchan_r = (! lizzieLet12_1_3QVal_Int_2_bufchan_buf[0]);
  assign lizzieLet12_1_3QVal_Int_2_argbuf_d = (lizzieLet12_1_3QVal_Int_2_bufchan_buf[0] ? lizzieLet12_1_3QVal_Int_2_bufchan_buf :
                                               lizzieLet12_1_3QVal_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet12_1_3QVal_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet12_1_3QVal_Int_2_argbuf_r && lizzieLet12_1_3QVal_Int_2_bufchan_buf[0]))
        lizzieLet12_1_3QVal_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet12_1_3QVal_Int_2_argbuf_r) && (! lizzieLet12_1_3QVal_Int_2_bufchan_buf[0])))
        lizzieLet12_1_3QVal_Int_2_bufchan_buf <= lizzieLet12_1_3QVal_Int_2_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_CT$wnnz_Int) : (lizzieLet12_1_4,QTree_Int) (sc_0_1_goMux_mux,Pointer_CT$wnnz_Int) > [(lizzieLet12_1_4QNone_Int,Pointer_CT$wnnz_Int),
                                                                                                       (lizzieLet12_1_4QVal_Int,Pointer_CT$wnnz_Int),
                                                                                                       (lizzieLet12_1_4QNode_Int,Pointer_CT$wnnz_Int),
                                                                                                       (lizzieLet12_1_4QError_Int,Pointer_CT$wnnz_Int)] */
  logic [3:0] sc_0_1_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet12_1_4_d[0] && sc_0_1_goMux_mux_d[0]))
      unique case (lizzieLet12_1_4_d[2:1])
        2'd0: sc_0_1_goMux_mux_onehotd = 4'd1;
        2'd1: sc_0_1_goMux_mux_onehotd = 4'd2;
        2'd2: sc_0_1_goMux_mux_onehotd = 4'd4;
        2'd3: sc_0_1_goMux_mux_onehotd = 4'd8;
        default: sc_0_1_goMux_mux_onehotd = 4'd0;
      endcase
    else sc_0_1_goMux_mux_onehotd = 4'd0;
  assign lizzieLet12_1_4QNone_Int_d = {sc_0_1_goMux_mux_d[16:1],
                                       sc_0_1_goMux_mux_onehotd[0]};
  assign lizzieLet12_1_4QVal_Int_d = {sc_0_1_goMux_mux_d[16:1],
                                      sc_0_1_goMux_mux_onehotd[1]};
  assign lizzieLet12_1_4QNode_Int_d = {sc_0_1_goMux_mux_d[16:1],
                                       sc_0_1_goMux_mux_onehotd[2]};
  assign lizzieLet12_1_4QError_Int_d = {sc_0_1_goMux_mux_d[16:1],
                                        sc_0_1_goMux_mux_onehotd[3]};
  assign sc_0_1_goMux_mux_r = (| (sc_0_1_goMux_mux_onehotd & {lizzieLet12_1_4QError_Int_r,
                                                              lizzieLet12_1_4QNode_Int_r,
                                                              lizzieLet12_1_4QVal_Int_r,
                                                              lizzieLet12_1_4QNone_Int_r}));
  assign lizzieLet12_1_4_r = sc_0_1_goMux_mux_r;
  
  /* buf (Ty Pointer_CT$wnnz_Int) : (lizzieLet12_1_4QError_Int,Pointer_CT$wnnz_Int) > (lizzieLet12_1_4QError_Int_1_argbuf,Pointer_CT$wnnz_Int) */
  Pointer_CT$wnnz_Int_t lizzieLet12_1_4QError_Int_bufchan_d;
  logic lizzieLet12_1_4QError_Int_bufchan_r;
  assign lizzieLet12_1_4QError_Int_r = ((! lizzieLet12_1_4QError_Int_bufchan_d[0]) || lizzieLet12_1_4QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_1_4QError_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet12_1_4QError_Int_r)
        lizzieLet12_1_4QError_Int_bufchan_d <= lizzieLet12_1_4QError_Int_d;
  Pointer_CT$wnnz_Int_t lizzieLet12_1_4QError_Int_bufchan_buf;
  assign lizzieLet12_1_4QError_Int_bufchan_r = (! lizzieLet12_1_4QError_Int_bufchan_buf[0]);
  assign lizzieLet12_1_4QError_Int_1_argbuf_d = (lizzieLet12_1_4QError_Int_bufchan_buf[0] ? lizzieLet12_1_4QError_Int_bufchan_buf :
                                                 lizzieLet12_1_4QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_1_4QError_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet12_1_4QError_Int_1_argbuf_r && lizzieLet12_1_4QError_Int_bufchan_buf[0]))
        lizzieLet12_1_4QError_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet12_1_4QError_Int_1_argbuf_r) && (! lizzieLet12_1_4QError_Int_bufchan_buf[0])))
        lizzieLet12_1_4QError_Int_bufchan_buf <= lizzieLet12_1_4QError_Int_bufchan_d;
  
  /* dcon (Ty CT$wnnz_Int,
      Dcon Lcall_$wnnz_Int3) : [(lizzieLet12_1_4QNode_Int,Pointer_CT$wnnz_Int),
                                (q4a8F_destruct,Pointer_QTree_Int),
                                (q3a8E_destruct,Pointer_QTree_Int),
                                (q2a8D_destruct,Pointer_QTree_Int)] > (lizzieLet12_1_4QNode_Int_1q4a8F_1q3a8E_1q2a8D_1Lcall_$wnnz_Int3,CT$wnnz_Int) */
  assign lizzieLet12_1_4QNode_Int_1q4a8F_1q3a8E_1q2a8D_1Lcall_$wnnz_Int3_d = Lcall_$wnnz_Int3_dc((& {lizzieLet12_1_4QNode_Int_d[0],
                                                                                                     q4a8F_destruct_d[0],
                                                                                                     q3a8E_destruct_d[0],
                                                                                                     q2a8D_destruct_d[0]}), lizzieLet12_1_4QNode_Int_d, q4a8F_destruct_d, q3a8E_destruct_d, q2a8D_destruct_d);
  assign {lizzieLet12_1_4QNode_Int_r,
          q4a8F_destruct_r,
          q3a8E_destruct_r,
          q2a8D_destruct_r} = {4 {(lizzieLet12_1_4QNode_Int_1q4a8F_1q3a8E_1q2a8D_1Lcall_$wnnz_Int3_r && lizzieLet12_1_4QNode_Int_1q4a8F_1q3a8E_1q2a8D_1Lcall_$wnnz_Int3_d[0])}};
  
  /* buf (Ty CT$wnnz_Int) : (lizzieLet12_1_4QNode_Int_1q4a8F_1q3a8E_1q2a8D_1Lcall_$wnnz_Int3,CT$wnnz_Int) > (lizzieLet13_1_1_argbuf,CT$wnnz_Int) */
  CT$wnnz_Int_t lizzieLet12_1_4QNode_Int_1q4a8F_1q3a8E_1q2a8D_1Lcall_$wnnz_Int3_bufchan_d;
  logic lizzieLet12_1_4QNode_Int_1q4a8F_1q3a8E_1q2a8D_1Lcall_$wnnz_Int3_bufchan_r;
  assign lizzieLet12_1_4QNode_Int_1q4a8F_1q3a8E_1q2a8D_1Lcall_$wnnz_Int3_r = ((! lizzieLet12_1_4QNode_Int_1q4a8F_1q3a8E_1q2a8D_1Lcall_$wnnz_Int3_bufchan_d[0]) || lizzieLet12_1_4QNode_Int_1q4a8F_1q3a8E_1q2a8D_1Lcall_$wnnz_Int3_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_1_4QNode_Int_1q4a8F_1q3a8E_1q2a8D_1Lcall_$wnnz_Int3_bufchan_d <= {115'd0,
                                                                                    1'd0};
    else
      if (lizzieLet12_1_4QNode_Int_1q4a8F_1q3a8E_1q2a8D_1Lcall_$wnnz_Int3_r)
        lizzieLet12_1_4QNode_Int_1q4a8F_1q3a8E_1q2a8D_1Lcall_$wnnz_Int3_bufchan_d <= lizzieLet12_1_4QNode_Int_1q4a8F_1q3a8E_1q2a8D_1Lcall_$wnnz_Int3_d;
  CT$wnnz_Int_t lizzieLet12_1_4QNode_Int_1q4a8F_1q3a8E_1q2a8D_1Lcall_$wnnz_Int3_bufchan_buf;
  assign lizzieLet12_1_4QNode_Int_1q4a8F_1q3a8E_1q2a8D_1Lcall_$wnnz_Int3_bufchan_r = (! lizzieLet12_1_4QNode_Int_1q4a8F_1q3a8E_1q2a8D_1Lcall_$wnnz_Int3_bufchan_buf[0]);
  assign lizzieLet13_1_1_argbuf_d = (lizzieLet12_1_4QNode_Int_1q4a8F_1q3a8E_1q2a8D_1Lcall_$wnnz_Int3_bufchan_buf[0] ? lizzieLet12_1_4QNode_Int_1q4a8F_1q3a8E_1q2a8D_1Lcall_$wnnz_Int3_bufchan_buf :
                                     lizzieLet12_1_4QNode_Int_1q4a8F_1q3a8E_1q2a8D_1Lcall_$wnnz_Int3_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_1_4QNode_Int_1q4a8F_1q3a8E_1q2a8D_1Lcall_$wnnz_Int3_bufchan_buf <= {115'd0,
                                                                                      1'd0};
    else
      if ((lizzieLet13_1_1_argbuf_r && lizzieLet12_1_4QNode_Int_1q4a8F_1q3a8E_1q2a8D_1Lcall_$wnnz_Int3_bufchan_buf[0]))
        lizzieLet12_1_4QNode_Int_1q4a8F_1q3a8E_1q2a8D_1Lcall_$wnnz_Int3_bufchan_buf <= {115'd0,
                                                                                        1'd0};
      else if (((! lizzieLet13_1_1_argbuf_r) && (! lizzieLet12_1_4QNode_Int_1q4a8F_1q3a8E_1q2a8D_1Lcall_$wnnz_Int3_bufchan_buf[0])))
        lizzieLet12_1_4QNode_Int_1q4a8F_1q3a8E_1q2a8D_1Lcall_$wnnz_Int3_bufchan_buf <= lizzieLet12_1_4QNode_Int_1q4a8F_1q3a8E_1q2a8D_1Lcall_$wnnz_Int3_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz_Int) : (lizzieLet12_1_4QNone_Int,Pointer_CT$wnnz_Int) > (lizzieLet12_1_4QNone_Int_1_argbuf,Pointer_CT$wnnz_Int) */
  Pointer_CT$wnnz_Int_t lizzieLet12_1_4QNone_Int_bufchan_d;
  logic lizzieLet12_1_4QNone_Int_bufchan_r;
  assign lizzieLet12_1_4QNone_Int_r = ((! lizzieLet12_1_4QNone_Int_bufchan_d[0]) || lizzieLet12_1_4QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_1_4QNone_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet12_1_4QNone_Int_r)
        lizzieLet12_1_4QNone_Int_bufchan_d <= lizzieLet12_1_4QNone_Int_d;
  Pointer_CT$wnnz_Int_t lizzieLet12_1_4QNone_Int_bufchan_buf;
  assign lizzieLet12_1_4QNone_Int_bufchan_r = (! lizzieLet12_1_4QNone_Int_bufchan_buf[0]);
  assign lizzieLet12_1_4QNone_Int_1_argbuf_d = (lizzieLet12_1_4QNone_Int_bufchan_buf[0] ? lizzieLet12_1_4QNone_Int_bufchan_buf :
                                                lizzieLet12_1_4QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_1_4QNone_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet12_1_4QNone_Int_1_argbuf_r && lizzieLet12_1_4QNone_Int_bufchan_buf[0]))
        lizzieLet12_1_4QNone_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet12_1_4QNone_Int_1_argbuf_r) && (! lizzieLet12_1_4QNone_Int_bufchan_buf[0])))
        lizzieLet12_1_4QNone_Int_bufchan_buf <= lizzieLet12_1_4QNone_Int_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz_Int) : (lizzieLet12_1_4QVal_Int,Pointer_CT$wnnz_Int) > (lizzieLet12_1_4QVal_Int_1_argbuf,Pointer_CT$wnnz_Int) */
  Pointer_CT$wnnz_Int_t lizzieLet12_1_4QVal_Int_bufchan_d;
  logic lizzieLet12_1_4QVal_Int_bufchan_r;
  assign lizzieLet12_1_4QVal_Int_r = ((! lizzieLet12_1_4QVal_Int_bufchan_d[0]) || lizzieLet12_1_4QVal_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_1_4QVal_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet12_1_4QVal_Int_r)
        lizzieLet12_1_4QVal_Int_bufchan_d <= lizzieLet12_1_4QVal_Int_d;
  Pointer_CT$wnnz_Int_t lizzieLet12_1_4QVal_Int_bufchan_buf;
  assign lizzieLet12_1_4QVal_Int_bufchan_r = (! lizzieLet12_1_4QVal_Int_bufchan_buf[0]);
  assign lizzieLet12_1_4QVal_Int_1_argbuf_d = (lizzieLet12_1_4QVal_Int_bufchan_buf[0] ? lizzieLet12_1_4QVal_Int_bufchan_buf :
                                               lizzieLet12_1_4QVal_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_1_4QVal_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet12_1_4QVal_Int_1_argbuf_r && lizzieLet12_1_4QVal_Int_bufchan_buf[0]))
        lizzieLet12_1_4QVal_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet12_1_4QVal_Int_1_argbuf_r) && (! lizzieLet12_1_4QVal_Int_bufchan_buf[0])))
        lizzieLet12_1_4QVal_Int_bufchan_buf <= lizzieLet12_1_4QVal_Int_bufchan_d;
  
  /* destruct (Ty MaskQTree,
          Dcon MQNode) : (lizzieLet14_1_1MQNode,MaskQTree) > [(q1a8s_destruct,Pointer_MaskQTree),
                                                              (q2a8t_destruct,Pointer_MaskQTree),
                                                              (q3a8u_destruct,Pointer_MaskQTree),
                                                              (q4a8v_destruct,Pointer_MaskQTree)] */
  logic [3:0] lizzieLet14_1_1MQNode_emitted;
  logic [3:0] lizzieLet14_1_1MQNode_done;
  assign q1a8s_destruct_d = {lizzieLet14_1_1MQNode_d[18:3],
                             (lizzieLet14_1_1MQNode_d[0] && (! lizzieLet14_1_1MQNode_emitted[0]))};
  assign q2a8t_destruct_d = {lizzieLet14_1_1MQNode_d[34:19],
                             (lizzieLet14_1_1MQNode_d[0] && (! lizzieLet14_1_1MQNode_emitted[1]))};
  assign q3a8u_destruct_d = {lizzieLet14_1_1MQNode_d[50:35],
                             (lizzieLet14_1_1MQNode_d[0] && (! lizzieLet14_1_1MQNode_emitted[2]))};
  assign q4a8v_destruct_d = {lizzieLet14_1_1MQNode_d[66:51],
                             (lizzieLet14_1_1MQNode_d[0] && (! lizzieLet14_1_1MQNode_emitted[3]))};
  assign lizzieLet14_1_1MQNode_done = (lizzieLet14_1_1MQNode_emitted | ({q4a8v_destruct_d[0],
                                                                         q3a8u_destruct_d[0],
                                                                         q2a8t_destruct_d[0],
                                                                         q1a8s_destruct_d[0]} & {q4a8v_destruct_r,
                                                                                                 q3a8u_destruct_r,
                                                                                                 q2a8t_destruct_r,
                                                                                                 q1a8s_destruct_r}));
  assign lizzieLet14_1_1MQNode_r = (& lizzieLet14_1_1MQNode_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet14_1_1MQNode_emitted <= 4'd0;
    else
      lizzieLet14_1_1MQNode_emitted <= (lizzieLet14_1_1MQNode_r ? 4'd0 :
                                        lizzieLet14_1_1MQNode_done);
  
  /* demux (Ty MaskQTree,
       Ty MaskQTree) : (lizzieLet14_1_2,MaskQTree) (lizzieLet14_1_1,MaskQTree) > [(_70,MaskQTree),
                                                                                  (_69,MaskQTree),
                                                                                  (lizzieLet14_1_1MQNode,MaskQTree)] */
  logic [2:0] lizzieLet14_1_1_onehotd;
  always_comb
    if ((lizzieLet14_1_2_d[0] && lizzieLet14_1_1_d[0]))
      unique case (lizzieLet14_1_2_d[2:1])
        2'd0: lizzieLet14_1_1_onehotd = 3'd1;
        2'd1: lizzieLet14_1_1_onehotd = 3'd2;
        2'd2: lizzieLet14_1_1_onehotd = 3'd4;
        default: lizzieLet14_1_1_onehotd = 3'd0;
      endcase
    else lizzieLet14_1_1_onehotd = 3'd0;
  assign _70_d = {lizzieLet14_1_1_d[66:1],
                  lizzieLet14_1_1_onehotd[0]};
  assign _69_d = {lizzieLet14_1_1_d[66:1],
                  lizzieLet14_1_1_onehotd[1]};
  assign lizzieLet14_1_1MQNode_d = {lizzieLet14_1_1_d[66:1],
                                    lizzieLet14_1_1_onehotd[2]};
  assign lizzieLet14_1_1_r = (| (lizzieLet14_1_1_onehotd & {lizzieLet14_1_1MQNode_r,
                                                            _69_r,
                                                            _70_r}));
  assign lizzieLet14_1_2_r = lizzieLet14_1_1_r;
  
  /* demux (Ty MaskQTree,
       Ty Go) : (lizzieLet14_1_3,MaskQTree) (go_8_goMux_data,Go) > [(lizzieLet14_1_3MQNone,Go),
                                                                    (lizzieLet14_1_3MQVal,Go),
                                                                    (lizzieLet14_1_3MQNode,Go)] */
  logic [2:0] go_8_goMux_data_onehotd;
  always_comb
    if ((lizzieLet14_1_3_d[0] && go_8_goMux_data_d[0]))
      unique case (lizzieLet14_1_3_d[2:1])
        2'd0: go_8_goMux_data_onehotd = 3'd1;
        2'd1: go_8_goMux_data_onehotd = 3'd2;
        2'd2: go_8_goMux_data_onehotd = 3'd4;
        default: go_8_goMux_data_onehotd = 3'd0;
      endcase
    else go_8_goMux_data_onehotd = 3'd0;
  assign lizzieLet14_1_3MQNone_d = go_8_goMux_data_onehotd[0];
  assign lizzieLet14_1_3MQVal_d = go_8_goMux_data_onehotd[1];
  assign lizzieLet14_1_3MQNode_d = go_8_goMux_data_onehotd[2];
  assign go_8_goMux_data_r = (| (go_8_goMux_data_onehotd & {lizzieLet14_1_3MQNode_r,
                                                            lizzieLet14_1_3MQVal_r,
                                                            lizzieLet14_1_3MQNone_r}));
  assign lizzieLet14_1_3_r = go_8_goMux_data_r;
  
  /* fork (Ty Go) : (lizzieLet14_1_3MQNone,Go) > [(lizzieLet14_1_3MQNone_1,Go),
                                             (lizzieLet14_1_3MQNone_2,Go)] */
  logic [1:0] lizzieLet14_1_3MQNone_emitted;
  logic [1:0] lizzieLet14_1_3MQNone_done;
  assign lizzieLet14_1_3MQNone_1_d = (lizzieLet14_1_3MQNone_d[0] && (! lizzieLet14_1_3MQNone_emitted[0]));
  assign lizzieLet14_1_3MQNone_2_d = (lizzieLet14_1_3MQNone_d[0] && (! lizzieLet14_1_3MQNone_emitted[1]));
  assign lizzieLet14_1_3MQNone_done = (lizzieLet14_1_3MQNone_emitted | ({lizzieLet14_1_3MQNone_2_d[0],
                                                                         lizzieLet14_1_3MQNone_1_d[0]} & {lizzieLet14_1_3MQNone_2_r,
                                                                                                          lizzieLet14_1_3MQNone_1_r}));
  assign lizzieLet14_1_3MQNone_r = (& lizzieLet14_1_3MQNone_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet14_1_3MQNone_emitted <= 2'd0;
    else
      lizzieLet14_1_3MQNone_emitted <= (lizzieLet14_1_3MQNone_r ? 2'd0 :
                                        lizzieLet14_1_3MQNone_done);
  
  /* dcon (Ty QTree_Int,
      Dcon QNone_Int) : [(lizzieLet14_1_3MQNone_1,Go)] > (lizzieLet14_1_3MQNone_1QNone_Int,QTree_Int) */
  assign lizzieLet14_1_3MQNone_1QNone_Int_d = QNone_Int_dc((& {lizzieLet14_1_3MQNone_1_d[0]}), lizzieLet14_1_3MQNone_1_d);
  assign {lizzieLet14_1_3MQNone_1_r} = {1 {(lizzieLet14_1_3MQNone_1QNone_Int_r && lizzieLet14_1_3MQNone_1QNone_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (lizzieLet14_1_3MQNone_1QNone_Int,QTree_Int) > (lizzieLet15_1_argbuf,QTree_Int) */
  QTree_Int_t lizzieLet14_1_3MQNone_1QNone_Int_bufchan_d;
  logic lizzieLet14_1_3MQNone_1QNone_Int_bufchan_r;
  assign lizzieLet14_1_3MQNone_1QNone_Int_r = ((! lizzieLet14_1_3MQNone_1QNone_Int_bufchan_d[0]) || lizzieLet14_1_3MQNone_1QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet14_1_3MQNone_1QNone_Int_bufchan_d <= {66'd0, 1'd0};
    else
      if (lizzieLet14_1_3MQNone_1QNone_Int_r)
        lizzieLet14_1_3MQNone_1QNone_Int_bufchan_d <= lizzieLet14_1_3MQNone_1QNone_Int_d;
  QTree_Int_t lizzieLet14_1_3MQNone_1QNone_Int_bufchan_buf;
  assign lizzieLet14_1_3MQNone_1QNone_Int_bufchan_r = (! lizzieLet14_1_3MQNone_1QNone_Int_bufchan_buf[0]);
  assign lizzieLet15_1_argbuf_d = (lizzieLet14_1_3MQNone_1QNone_Int_bufchan_buf[0] ? lizzieLet14_1_3MQNone_1QNone_Int_bufchan_buf :
                                   lizzieLet14_1_3MQNone_1QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet14_1_3MQNone_1QNone_Int_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((lizzieLet15_1_argbuf_r && lizzieLet14_1_3MQNone_1QNone_Int_bufchan_buf[0]))
        lizzieLet14_1_3MQNone_1QNone_Int_bufchan_buf <= {66'd0, 1'd0};
      else if (((! lizzieLet15_1_argbuf_r) && (! lizzieLet14_1_3MQNone_1QNone_Int_bufchan_buf[0])))
        lizzieLet14_1_3MQNone_1QNone_Int_bufchan_buf <= lizzieLet14_1_3MQNone_1QNone_Int_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet14_1_3MQNone_2,Go) > (lizzieLet14_1_3MQNone_2_argbuf,Go) */
  Go_t lizzieLet14_1_3MQNone_2_bufchan_d;
  logic lizzieLet14_1_3MQNone_2_bufchan_r;
  assign lizzieLet14_1_3MQNone_2_r = ((! lizzieLet14_1_3MQNone_2_bufchan_d[0]) || lizzieLet14_1_3MQNone_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet14_1_3MQNone_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet14_1_3MQNone_2_r)
        lizzieLet14_1_3MQNone_2_bufchan_d <= lizzieLet14_1_3MQNone_2_d;
  Go_t lizzieLet14_1_3MQNone_2_bufchan_buf;
  assign lizzieLet14_1_3MQNone_2_bufchan_r = (! lizzieLet14_1_3MQNone_2_bufchan_buf[0]);
  assign lizzieLet14_1_3MQNone_2_argbuf_d = (lizzieLet14_1_3MQNone_2_bufchan_buf[0] ? lizzieLet14_1_3MQNone_2_bufchan_buf :
                                             lizzieLet14_1_3MQNone_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet14_1_3MQNone_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet14_1_3MQNone_2_argbuf_r && lizzieLet14_1_3MQNone_2_bufchan_buf[0]))
        lizzieLet14_1_3MQNone_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet14_1_3MQNone_2_argbuf_r) && (! lizzieLet14_1_3MQNone_2_bufchan_buf[0])))
        lizzieLet14_1_3MQNone_2_bufchan_buf <= lizzieLet14_1_3MQNone_2_bufchan_d;
  
  /* mergectrl (Ty C6,Ty Go) : [(lizzieLet14_1_3MQNone_2_argbuf,Go),
                           (lizzieLet31_3Lcall_main_mask_Int0_1_argbuf,Go),
                           (lizzieLet14_1_3MQVal_1_argbuf,Go),
                           (lizzieLet14_1_4MQNode_3QNone_Int_2_argbuf,Go),
                           (lizzieLet14_1_4MQNode_3QVal_Int_2_argbuf,Go),
                           (lizzieLet14_1_4MQNode_3QError_Int_2_argbuf,Go)] > (go_12_goMux_choice,C6) (go_12_goMux_data,Go) */
  logic [5:0] lizzieLet14_1_3MQNone_2_argbuf_select_d;
  assign lizzieLet14_1_3MQNone_2_argbuf_select_d = ((| lizzieLet14_1_3MQNone_2_argbuf_select_q) ? lizzieLet14_1_3MQNone_2_argbuf_select_q :
                                                    (lizzieLet14_1_3MQNone_2_argbuf_d[0] ? 6'd1 :
                                                     (lizzieLet31_3Lcall_main_mask_Int0_1_argbuf_d[0] ? 6'd2 :
                                                      (lizzieLet14_1_3MQVal_1_argbuf_d[0] ? 6'd4 :
                                                       (lizzieLet14_1_4MQNode_3QNone_Int_2_argbuf_d[0] ? 6'd8 :
                                                        (lizzieLet14_1_4MQNode_3QVal_Int_2_argbuf_d[0] ? 6'd16 :
                                                         (lizzieLet14_1_4MQNode_3QError_Int_2_argbuf_d[0] ? 6'd32 :
                                                          6'd0)))))));
  logic [5:0] lizzieLet14_1_3MQNone_2_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet14_1_3MQNone_2_argbuf_select_q <= 6'd0;
    else
      lizzieLet14_1_3MQNone_2_argbuf_select_q <= (lizzieLet14_1_3MQNone_2_argbuf_done ? 6'd0 :
                                                  lizzieLet14_1_3MQNone_2_argbuf_select_d);
  logic [1:0] lizzieLet14_1_3MQNone_2_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet14_1_3MQNone_2_argbuf_emit_q <= 2'd0;
    else
      lizzieLet14_1_3MQNone_2_argbuf_emit_q <= (lizzieLet14_1_3MQNone_2_argbuf_done ? 2'd0 :
                                                lizzieLet14_1_3MQNone_2_argbuf_emit_d);
  logic [1:0] lizzieLet14_1_3MQNone_2_argbuf_emit_d;
  assign lizzieLet14_1_3MQNone_2_argbuf_emit_d = (lizzieLet14_1_3MQNone_2_argbuf_emit_q | ({go_12_goMux_choice_d[0],
                                                                                            go_12_goMux_data_d[0]} & {go_12_goMux_choice_r,
                                                                                                                      go_12_goMux_data_r}));
  logic lizzieLet14_1_3MQNone_2_argbuf_done;
  assign lizzieLet14_1_3MQNone_2_argbuf_done = (& lizzieLet14_1_3MQNone_2_argbuf_emit_d);
  assign {lizzieLet14_1_4MQNode_3QError_Int_2_argbuf_r,
          lizzieLet14_1_4MQNode_3QVal_Int_2_argbuf_r,
          lizzieLet14_1_4MQNode_3QNone_Int_2_argbuf_r,
          lizzieLet14_1_3MQVal_1_argbuf_r,
          lizzieLet31_3Lcall_main_mask_Int0_1_argbuf_r,
          lizzieLet14_1_3MQNone_2_argbuf_r} = (lizzieLet14_1_3MQNone_2_argbuf_done ? lizzieLet14_1_3MQNone_2_argbuf_select_d :
                                               6'd0);
  assign go_12_goMux_data_d = ((lizzieLet14_1_3MQNone_2_argbuf_select_d[0] && (! lizzieLet14_1_3MQNone_2_argbuf_emit_q[0])) ? lizzieLet14_1_3MQNone_2_argbuf_d :
                               ((lizzieLet14_1_3MQNone_2_argbuf_select_d[1] && (! lizzieLet14_1_3MQNone_2_argbuf_emit_q[0])) ? lizzieLet31_3Lcall_main_mask_Int0_1_argbuf_d :
                                ((lizzieLet14_1_3MQNone_2_argbuf_select_d[2] && (! lizzieLet14_1_3MQNone_2_argbuf_emit_q[0])) ? lizzieLet14_1_3MQVal_1_argbuf_d :
                                 ((lizzieLet14_1_3MQNone_2_argbuf_select_d[3] && (! lizzieLet14_1_3MQNone_2_argbuf_emit_q[0])) ? lizzieLet14_1_4MQNode_3QNone_Int_2_argbuf_d :
                                  ((lizzieLet14_1_3MQNone_2_argbuf_select_d[4] && (! lizzieLet14_1_3MQNone_2_argbuf_emit_q[0])) ? lizzieLet14_1_4MQNode_3QVal_Int_2_argbuf_d :
                                   ((lizzieLet14_1_3MQNone_2_argbuf_select_d[5] && (! lizzieLet14_1_3MQNone_2_argbuf_emit_q[0])) ? lizzieLet14_1_4MQNode_3QError_Int_2_argbuf_d :
                                    1'd0))))));
  assign go_12_goMux_choice_d = ((lizzieLet14_1_3MQNone_2_argbuf_select_d[0] && (! lizzieLet14_1_3MQNone_2_argbuf_emit_q[1])) ? C1_6_dc(1'd1) :
                                 ((lizzieLet14_1_3MQNone_2_argbuf_select_d[1] && (! lizzieLet14_1_3MQNone_2_argbuf_emit_q[1])) ? C2_6_dc(1'd1) :
                                  ((lizzieLet14_1_3MQNone_2_argbuf_select_d[2] && (! lizzieLet14_1_3MQNone_2_argbuf_emit_q[1])) ? C3_6_dc(1'd1) :
                                   ((lizzieLet14_1_3MQNone_2_argbuf_select_d[3] && (! lizzieLet14_1_3MQNone_2_argbuf_emit_q[1])) ? C4_6_dc(1'd1) :
                                    ((lizzieLet14_1_3MQNone_2_argbuf_select_d[4] && (! lizzieLet14_1_3MQNone_2_argbuf_emit_q[1])) ? C5_6_dc(1'd1) :
                                     ((lizzieLet14_1_3MQNone_2_argbuf_select_d[5] && (! lizzieLet14_1_3MQNone_2_argbuf_emit_q[1])) ? C6_6_dc(1'd1) :
                                      {3'd0, 1'd0}))))));
  
  /* buf (Ty Go) : (lizzieLet14_1_3MQVal,Go) > (lizzieLet14_1_3MQVal_1_argbuf,Go) */
  Go_t lizzieLet14_1_3MQVal_bufchan_d;
  logic lizzieLet14_1_3MQVal_bufchan_r;
  assign lizzieLet14_1_3MQVal_r = ((! lizzieLet14_1_3MQVal_bufchan_d[0]) || lizzieLet14_1_3MQVal_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet14_1_3MQVal_bufchan_d <= 1'd0;
    else
      if (lizzieLet14_1_3MQVal_r)
        lizzieLet14_1_3MQVal_bufchan_d <= lizzieLet14_1_3MQVal_d;
  Go_t lizzieLet14_1_3MQVal_bufchan_buf;
  assign lizzieLet14_1_3MQVal_bufchan_r = (! lizzieLet14_1_3MQVal_bufchan_buf[0]);
  assign lizzieLet14_1_3MQVal_1_argbuf_d = (lizzieLet14_1_3MQVal_bufchan_buf[0] ? lizzieLet14_1_3MQVal_bufchan_buf :
                                            lizzieLet14_1_3MQVal_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet14_1_3MQVal_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet14_1_3MQVal_1_argbuf_r && lizzieLet14_1_3MQVal_bufchan_buf[0]))
        lizzieLet14_1_3MQVal_bufchan_buf <= 1'd0;
      else if (((! lizzieLet14_1_3MQVal_1_argbuf_r) && (! lizzieLet14_1_3MQVal_bufchan_buf[0])))
        lizzieLet14_1_3MQVal_bufchan_buf <= lizzieLet14_1_3MQVal_bufchan_d;
  
  /* demux (Ty MaskQTree,
       Ty QTree_Int) : (lizzieLet14_1_4,MaskQTree) (readPointer_QTree_Intma8q_1_argbuf_rwb,QTree_Int) > [(_68,QTree_Int),
                                                                                                         (_67,QTree_Int),
                                                                                                         (lizzieLet14_1_4MQNode,QTree_Int)] */
  logic [2:0] readPointer_QTree_Intma8q_1_argbuf_rwb_onehotd;
  always_comb
    if ((lizzieLet14_1_4_d[0] && readPointer_QTree_Intma8q_1_argbuf_rwb_d[0]))
      unique case (lizzieLet14_1_4_d[2:1])
        2'd0: readPointer_QTree_Intma8q_1_argbuf_rwb_onehotd = 3'd1;
        2'd1: readPointer_QTree_Intma8q_1_argbuf_rwb_onehotd = 3'd2;
        2'd2: readPointer_QTree_Intma8q_1_argbuf_rwb_onehotd = 3'd4;
        default: readPointer_QTree_Intma8q_1_argbuf_rwb_onehotd = 3'd0;
      endcase
    else readPointer_QTree_Intma8q_1_argbuf_rwb_onehotd = 3'd0;
  assign _68_d = {readPointer_QTree_Intma8q_1_argbuf_rwb_d[66:1],
                  readPointer_QTree_Intma8q_1_argbuf_rwb_onehotd[0]};
  assign _67_d = {readPointer_QTree_Intma8q_1_argbuf_rwb_d[66:1],
                  readPointer_QTree_Intma8q_1_argbuf_rwb_onehotd[1]};
  assign lizzieLet14_1_4MQNode_d = {readPointer_QTree_Intma8q_1_argbuf_rwb_d[66:1],
                                    readPointer_QTree_Intma8q_1_argbuf_rwb_onehotd[2]};
  assign readPointer_QTree_Intma8q_1_argbuf_rwb_r = (| (readPointer_QTree_Intma8q_1_argbuf_rwb_onehotd & {lizzieLet14_1_4MQNode_r,
                                                                                                          _67_r,
                                                                                                          _68_r}));
  assign lizzieLet14_1_4_r = readPointer_QTree_Intma8q_1_argbuf_rwb_r;
  
  /* fork (Ty QTree_Int) : (lizzieLet14_1_4MQNode,QTree_Int) > [(lizzieLet14_1_4MQNode_1,QTree_Int),
                                                           (lizzieLet14_1_4MQNode_2,QTree_Int),
                                                           (lizzieLet14_1_4MQNode_3,QTree_Int),
                                                           (lizzieLet14_1_4MQNode_4,QTree_Int),
                                                           (lizzieLet14_1_4MQNode_5,QTree_Int),
                                                           (lizzieLet14_1_4MQNode_6,QTree_Int),
                                                           (lizzieLet14_1_4MQNode_7,QTree_Int),
                                                           (lizzieLet14_1_4MQNode_8,QTree_Int)] */
  logic [7:0] lizzieLet14_1_4MQNode_emitted;
  logic [7:0] lizzieLet14_1_4MQNode_done;
  assign lizzieLet14_1_4MQNode_1_d = {lizzieLet14_1_4MQNode_d[66:1],
                                      (lizzieLet14_1_4MQNode_d[0] && (! lizzieLet14_1_4MQNode_emitted[0]))};
  assign lizzieLet14_1_4MQNode_2_d = {lizzieLet14_1_4MQNode_d[66:1],
                                      (lizzieLet14_1_4MQNode_d[0] && (! lizzieLet14_1_4MQNode_emitted[1]))};
  assign lizzieLet14_1_4MQNode_3_d = {lizzieLet14_1_4MQNode_d[66:1],
                                      (lizzieLet14_1_4MQNode_d[0] && (! lizzieLet14_1_4MQNode_emitted[2]))};
  assign lizzieLet14_1_4MQNode_4_d = {lizzieLet14_1_4MQNode_d[66:1],
                                      (lizzieLet14_1_4MQNode_d[0] && (! lizzieLet14_1_4MQNode_emitted[3]))};
  assign lizzieLet14_1_4MQNode_5_d = {lizzieLet14_1_4MQNode_d[66:1],
                                      (lizzieLet14_1_4MQNode_d[0] && (! lizzieLet14_1_4MQNode_emitted[4]))};
  assign lizzieLet14_1_4MQNode_6_d = {lizzieLet14_1_4MQNode_d[66:1],
                                      (lizzieLet14_1_4MQNode_d[0] && (! lizzieLet14_1_4MQNode_emitted[5]))};
  assign lizzieLet14_1_4MQNode_7_d = {lizzieLet14_1_4MQNode_d[66:1],
                                      (lizzieLet14_1_4MQNode_d[0] && (! lizzieLet14_1_4MQNode_emitted[6]))};
  assign lizzieLet14_1_4MQNode_8_d = {lizzieLet14_1_4MQNode_d[66:1],
                                      (lizzieLet14_1_4MQNode_d[0] && (! lizzieLet14_1_4MQNode_emitted[7]))};
  assign lizzieLet14_1_4MQNode_done = (lizzieLet14_1_4MQNode_emitted | ({lizzieLet14_1_4MQNode_8_d[0],
                                                                         lizzieLet14_1_4MQNode_7_d[0],
                                                                         lizzieLet14_1_4MQNode_6_d[0],
                                                                         lizzieLet14_1_4MQNode_5_d[0],
                                                                         lizzieLet14_1_4MQNode_4_d[0],
                                                                         lizzieLet14_1_4MQNode_3_d[0],
                                                                         lizzieLet14_1_4MQNode_2_d[0],
                                                                         lizzieLet14_1_4MQNode_1_d[0]} & {lizzieLet14_1_4MQNode_8_r,
                                                                                                          lizzieLet14_1_4MQNode_7_r,
                                                                                                          lizzieLet14_1_4MQNode_6_r,
                                                                                                          lizzieLet14_1_4MQNode_5_r,
                                                                                                          lizzieLet14_1_4MQNode_4_r,
                                                                                                          lizzieLet14_1_4MQNode_3_r,
                                                                                                          lizzieLet14_1_4MQNode_2_r,
                                                                                                          lizzieLet14_1_4MQNode_1_r}));
  assign lizzieLet14_1_4MQNode_r = (& lizzieLet14_1_4MQNode_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet14_1_4MQNode_emitted <= 8'd0;
    else
      lizzieLet14_1_4MQNode_emitted <= (lizzieLet14_1_4MQNode_r ? 8'd0 :
                                        lizzieLet14_1_4MQNode_done);
  
  /* destruct (Ty QTree_Int,
          Dcon QNode_Int) : (lizzieLet14_1_4MQNode_1QNode_Int,QTree_Int) > [(t1a8x_destruct,Pointer_QTree_Int),
                                                                            (t2a8y_destruct,Pointer_QTree_Int),
                                                                            (t3a8z_destruct,Pointer_QTree_Int),
                                                                            (t4a8A_destruct,Pointer_QTree_Int)] */
  logic [3:0] lizzieLet14_1_4MQNode_1QNode_Int_emitted;
  logic [3:0] lizzieLet14_1_4MQNode_1QNode_Int_done;
  assign t1a8x_destruct_d = {lizzieLet14_1_4MQNode_1QNode_Int_d[18:3],
                             (lizzieLet14_1_4MQNode_1QNode_Int_d[0] && (! lizzieLet14_1_4MQNode_1QNode_Int_emitted[0]))};
  assign t2a8y_destruct_d = {lizzieLet14_1_4MQNode_1QNode_Int_d[34:19],
                             (lizzieLet14_1_4MQNode_1QNode_Int_d[0] && (! lizzieLet14_1_4MQNode_1QNode_Int_emitted[1]))};
  assign t3a8z_destruct_d = {lizzieLet14_1_4MQNode_1QNode_Int_d[50:35],
                             (lizzieLet14_1_4MQNode_1QNode_Int_d[0] && (! lizzieLet14_1_4MQNode_1QNode_Int_emitted[2]))};
  assign t4a8A_destruct_d = {lizzieLet14_1_4MQNode_1QNode_Int_d[66:51],
                             (lizzieLet14_1_4MQNode_1QNode_Int_d[0] && (! lizzieLet14_1_4MQNode_1QNode_Int_emitted[3]))};
  assign lizzieLet14_1_4MQNode_1QNode_Int_done = (lizzieLet14_1_4MQNode_1QNode_Int_emitted | ({t4a8A_destruct_d[0],
                                                                                               t3a8z_destruct_d[0],
                                                                                               t2a8y_destruct_d[0],
                                                                                               t1a8x_destruct_d[0]} & {t4a8A_destruct_r,
                                                                                                                       t3a8z_destruct_r,
                                                                                                                       t2a8y_destruct_r,
                                                                                                                       t1a8x_destruct_r}));
  assign lizzieLet14_1_4MQNode_1QNode_Int_r = (& lizzieLet14_1_4MQNode_1QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet14_1_4MQNode_1QNode_Int_emitted <= 4'd0;
    else
      lizzieLet14_1_4MQNode_1QNode_Int_emitted <= (lizzieLet14_1_4MQNode_1QNode_Int_r ? 4'd0 :
                                                   lizzieLet14_1_4MQNode_1QNode_Int_done);
  
  /* demux (Ty QTree_Int,
       Ty QTree_Int) : (lizzieLet14_1_4MQNode_2,QTree_Int) (lizzieLet14_1_4MQNode_1,QTree_Int) > [(_66,QTree_Int),
                                                                                                  (_65,QTree_Int),
                                                                                                  (lizzieLet14_1_4MQNode_1QNode_Int,QTree_Int),
                                                                                                  (_64,QTree_Int)] */
  logic [3:0] lizzieLet14_1_4MQNode_1_onehotd;
  always_comb
    if ((lizzieLet14_1_4MQNode_2_d[0] && lizzieLet14_1_4MQNode_1_d[0]))
      unique case (lizzieLet14_1_4MQNode_2_d[2:1])
        2'd0: lizzieLet14_1_4MQNode_1_onehotd = 4'd1;
        2'd1: lizzieLet14_1_4MQNode_1_onehotd = 4'd2;
        2'd2: lizzieLet14_1_4MQNode_1_onehotd = 4'd4;
        2'd3: lizzieLet14_1_4MQNode_1_onehotd = 4'd8;
        default: lizzieLet14_1_4MQNode_1_onehotd = 4'd0;
      endcase
    else lizzieLet14_1_4MQNode_1_onehotd = 4'd0;
  assign _66_d = {lizzieLet14_1_4MQNode_1_d[66:1],
                  lizzieLet14_1_4MQNode_1_onehotd[0]};
  assign _65_d = {lizzieLet14_1_4MQNode_1_d[66:1],
                  lizzieLet14_1_4MQNode_1_onehotd[1]};
  assign lizzieLet14_1_4MQNode_1QNode_Int_d = {lizzieLet14_1_4MQNode_1_d[66:1],
                                               lizzieLet14_1_4MQNode_1_onehotd[2]};
  assign _64_d = {lizzieLet14_1_4MQNode_1_d[66:1],
                  lizzieLet14_1_4MQNode_1_onehotd[3]};
  assign lizzieLet14_1_4MQNode_1_r = (| (lizzieLet14_1_4MQNode_1_onehotd & {_64_r,
                                                                            lizzieLet14_1_4MQNode_1QNode_Int_r,
                                                                            _65_r,
                                                                            _66_r}));
  assign lizzieLet14_1_4MQNode_2_r = lizzieLet14_1_4MQNode_1_r;
  
  /* demux (Ty QTree_Int,
       Ty Go) : (lizzieLet14_1_4MQNode_3,QTree_Int) (lizzieLet14_1_3MQNode,Go) > [(lizzieLet14_1_4MQNode_3QNone_Int,Go),
                                                                                  (lizzieLet14_1_4MQNode_3QVal_Int,Go),
                                                                                  (lizzieLet14_1_4MQNode_3QNode_Int,Go),
                                                                                  (lizzieLet14_1_4MQNode_3QError_Int,Go)] */
  logic [3:0] lizzieLet14_1_3MQNode_onehotd;
  always_comb
    if ((lizzieLet14_1_4MQNode_3_d[0] && lizzieLet14_1_3MQNode_d[0]))
      unique case (lizzieLet14_1_4MQNode_3_d[2:1])
        2'd0: lizzieLet14_1_3MQNode_onehotd = 4'd1;
        2'd1: lizzieLet14_1_3MQNode_onehotd = 4'd2;
        2'd2: lizzieLet14_1_3MQNode_onehotd = 4'd4;
        2'd3: lizzieLet14_1_3MQNode_onehotd = 4'd8;
        default: lizzieLet14_1_3MQNode_onehotd = 4'd0;
      endcase
    else lizzieLet14_1_3MQNode_onehotd = 4'd0;
  assign lizzieLet14_1_4MQNode_3QNone_Int_d = lizzieLet14_1_3MQNode_onehotd[0];
  assign lizzieLet14_1_4MQNode_3QVal_Int_d = lizzieLet14_1_3MQNode_onehotd[1];
  assign lizzieLet14_1_4MQNode_3QNode_Int_d = lizzieLet14_1_3MQNode_onehotd[2];
  assign lizzieLet14_1_4MQNode_3QError_Int_d = lizzieLet14_1_3MQNode_onehotd[3];
  assign lizzieLet14_1_3MQNode_r = (| (lizzieLet14_1_3MQNode_onehotd & {lizzieLet14_1_4MQNode_3QError_Int_r,
                                                                        lizzieLet14_1_4MQNode_3QNode_Int_r,
                                                                        lizzieLet14_1_4MQNode_3QVal_Int_r,
                                                                        lizzieLet14_1_4MQNode_3QNone_Int_r}));
  assign lizzieLet14_1_4MQNode_3_r = lizzieLet14_1_3MQNode_r;
  
  /* fork (Ty Go) : (lizzieLet14_1_4MQNode_3QError_Int,Go) > [(lizzieLet14_1_4MQNode_3QError_Int_1,Go),
                                                         (lizzieLet14_1_4MQNode_3QError_Int_2,Go)] */
  logic [1:0] lizzieLet14_1_4MQNode_3QError_Int_emitted;
  logic [1:0] lizzieLet14_1_4MQNode_3QError_Int_done;
  assign lizzieLet14_1_4MQNode_3QError_Int_1_d = (lizzieLet14_1_4MQNode_3QError_Int_d[0] && (! lizzieLet14_1_4MQNode_3QError_Int_emitted[0]));
  assign lizzieLet14_1_4MQNode_3QError_Int_2_d = (lizzieLet14_1_4MQNode_3QError_Int_d[0] && (! lizzieLet14_1_4MQNode_3QError_Int_emitted[1]));
  assign lizzieLet14_1_4MQNode_3QError_Int_done = (lizzieLet14_1_4MQNode_3QError_Int_emitted | ({lizzieLet14_1_4MQNode_3QError_Int_2_d[0],
                                                                                                 lizzieLet14_1_4MQNode_3QError_Int_1_d[0]} & {lizzieLet14_1_4MQNode_3QError_Int_2_r,
                                                                                                                                              lizzieLet14_1_4MQNode_3QError_Int_1_r}));
  assign lizzieLet14_1_4MQNode_3QError_Int_r = (& lizzieLet14_1_4MQNode_3QError_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet14_1_4MQNode_3QError_Int_emitted <= 2'd0;
    else
      lizzieLet14_1_4MQNode_3QError_Int_emitted <= (lizzieLet14_1_4MQNode_3QError_Int_r ? 2'd0 :
                                                    lizzieLet14_1_4MQNode_3QError_Int_done);
  
  /* dcon (Ty QTree_Int,
      Dcon QError_Int) : [(lizzieLet14_1_4MQNode_3QError_Int_1,Go)] > (lizzieLet14_1_4MQNode_3QError_Int_1QError_Int,QTree_Int) */
  assign lizzieLet14_1_4MQNode_3QError_Int_1QError_Int_d = QError_Int_dc((& {lizzieLet14_1_4MQNode_3QError_Int_1_d[0]}), lizzieLet14_1_4MQNode_3QError_Int_1_d);
  assign {lizzieLet14_1_4MQNode_3QError_Int_1_r} = {1 {(lizzieLet14_1_4MQNode_3QError_Int_1QError_Int_r && lizzieLet14_1_4MQNode_3QError_Int_1QError_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (lizzieLet14_1_4MQNode_3QError_Int_1QError_Int,QTree_Int) > (lizzieLet20_1_argbuf,QTree_Int) */
  QTree_Int_t lizzieLet14_1_4MQNode_3QError_Int_1QError_Int_bufchan_d;
  logic lizzieLet14_1_4MQNode_3QError_Int_1QError_Int_bufchan_r;
  assign lizzieLet14_1_4MQNode_3QError_Int_1QError_Int_r = ((! lizzieLet14_1_4MQNode_3QError_Int_1QError_Int_bufchan_d[0]) || lizzieLet14_1_4MQNode_3QError_Int_1QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet14_1_4MQNode_3QError_Int_1QError_Int_bufchan_d <= {66'd0,
                                                                  1'd0};
    else
      if (lizzieLet14_1_4MQNode_3QError_Int_1QError_Int_r)
        lizzieLet14_1_4MQNode_3QError_Int_1QError_Int_bufchan_d <= lizzieLet14_1_4MQNode_3QError_Int_1QError_Int_d;
  QTree_Int_t lizzieLet14_1_4MQNode_3QError_Int_1QError_Int_bufchan_buf;
  assign lizzieLet14_1_4MQNode_3QError_Int_1QError_Int_bufchan_r = (! lizzieLet14_1_4MQNode_3QError_Int_1QError_Int_bufchan_buf[0]);
  assign lizzieLet20_1_argbuf_d = (lizzieLet14_1_4MQNode_3QError_Int_1QError_Int_bufchan_buf[0] ? lizzieLet14_1_4MQNode_3QError_Int_1QError_Int_bufchan_buf :
                                   lizzieLet14_1_4MQNode_3QError_Int_1QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet14_1_4MQNode_3QError_Int_1QError_Int_bufchan_buf <= {66'd0,
                                                                    1'd0};
    else
      if ((lizzieLet20_1_argbuf_r && lizzieLet14_1_4MQNode_3QError_Int_1QError_Int_bufchan_buf[0]))
        lizzieLet14_1_4MQNode_3QError_Int_1QError_Int_bufchan_buf <= {66'd0,
                                                                      1'd0};
      else if (((! lizzieLet20_1_argbuf_r) && (! lizzieLet14_1_4MQNode_3QError_Int_1QError_Int_bufchan_buf[0])))
        lizzieLet14_1_4MQNode_3QError_Int_1QError_Int_bufchan_buf <= lizzieLet14_1_4MQNode_3QError_Int_1QError_Int_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet14_1_4MQNode_3QError_Int_2,Go) > (lizzieLet14_1_4MQNode_3QError_Int_2_argbuf,Go) */
  Go_t lizzieLet14_1_4MQNode_3QError_Int_2_bufchan_d;
  logic lizzieLet14_1_4MQNode_3QError_Int_2_bufchan_r;
  assign lizzieLet14_1_4MQNode_3QError_Int_2_r = ((! lizzieLet14_1_4MQNode_3QError_Int_2_bufchan_d[0]) || lizzieLet14_1_4MQNode_3QError_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet14_1_4MQNode_3QError_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet14_1_4MQNode_3QError_Int_2_r)
        lizzieLet14_1_4MQNode_3QError_Int_2_bufchan_d <= lizzieLet14_1_4MQNode_3QError_Int_2_d;
  Go_t lizzieLet14_1_4MQNode_3QError_Int_2_bufchan_buf;
  assign lizzieLet14_1_4MQNode_3QError_Int_2_bufchan_r = (! lizzieLet14_1_4MQNode_3QError_Int_2_bufchan_buf[0]);
  assign lizzieLet14_1_4MQNode_3QError_Int_2_argbuf_d = (lizzieLet14_1_4MQNode_3QError_Int_2_bufchan_buf[0] ? lizzieLet14_1_4MQNode_3QError_Int_2_bufchan_buf :
                                                         lizzieLet14_1_4MQNode_3QError_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet14_1_4MQNode_3QError_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet14_1_4MQNode_3QError_Int_2_argbuf_r && lizzieLet14_1_4MQNode_3QError_Int_2_bufchan_buf[0]))
        lizzieLet14_1_4MQNode_3QError_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet14_1_4MQNode_3QError_Int_2_argbuf_r) && (! lizzieLet14_1_4MQNode_3QError_Int_2_bufchan_buf[0])))
        lizzieLet14_1_4MQNode_3QError_Int_2_bufchan_buf <= lizzieLet14_1_4MQNode_3QError_Int_2_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet14_1_4MQNode_3QNode_Int,Go) > (lizzieLet14_1_4MQNode_3QNode_Int_1_argbuf,Go) */
  Go_t lizzieLet14_1_4MQNode_3QNode_Int_bufchan_d;
  logic lizzieLet14_1_4MQNode_3QNode_Int_bufchan_r;
  assign lizzieLet14_1_4MQNode_3QNode_Int_r = ((! lizzieLet14_1_4MQNode_3QNode_Int_bufchan_d[0]) || lizzieLet14_1_4MQNode_3QNode_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet14_1_4MQNode_3QNode_Int_bufchan_d <= 1'd0;
    else
      if (lizzieLet14_1_4MQNode_3QNode_Int_r)
        lizzieLet14_1_4MQNode_3QNode_Int_bufchan_d <= lizzieLet14_1_4MQNode_3QNode_Int_d;
  Go_t lizzieLet14_1_4MQNode_3QNode_Int_bufchan_buf;
  assign lizzieLet14_1_4MQNode_3QNode_Int_bufchan_r = (! lizzieLet14_1_4MQNode_3QNode_Int_bufchan_buf[0]);
  assign lizzieLet14_1_4MQNode_3QNode_Int_1_argbuf_d = (lizzieLet14_1_4MQNode_3QNode_Int_bufchan_buf[0] ? lizzieLet14_1_4MQNode_3QNode_Int_bufchan_buf :
                                                        lizzieLet14_1_4MQNode_3QNode_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet14_1_4MQNode_3QNode_Int_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet14_1_4MQNode_3QNode_Int_1_argbuf_r && lizzieLet14_1_4MQNode_3QNode_Int_bufchan_buf[0]))
        lizzieLet14_1_4MQNode_3QNode_Int_bufchan_buf <= 1'd0;
      else if (((! lizzieLet14_1_4MQNode_3QNode_Int_1_argbuf_r) && (! lizzieLet14_1_4MQNode_3QNode_Int_bufchan_buf[0])))
        lizzieLet14_1_4MQNode_3QNode_Int_bufchan_buf <= lizzieLet14_1_4MQNode_3QNode_Int_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet14_1_4MQNode_3QNone_Int,Go) > [(lizzieLet14_1_4MQNode_3QNone_Int_1,Go),
                                                        (lizzieLet14_1_4MQNode_3QNone_Int_2,Go)] */
  logic [1:0] lizzieLet14_1_4MQNode_3QNone_Int_emitted;
  logic [1:0] lizzieLet14_1_4MQNode_3QNone_Int_done;
  assign lizzieLet14_1_4MQNode_3QNone_Int_1_d = (lizzieLet14_1_4MQNode_3QNone_Int_d[0] && (! lizzieLet14_1_4MQNode_3QNone_Int_emitted[0]));
  assign lizzieLet14_1_4MQNode_3QNone_Int_2_d = (lizzieLet14_1_4MQNode_3QNone_Int_d[0] && (! lizzieLet14_1_4MQNode_3QNone_Int_emitted[1]));
  assign lizzieLet14_1_4MQNode_3QNone_Int_done = (lizzieLet14_1_4MQNode_3QNone_Int_emitted | ({lizzieLet14_1_4MQNode_3QNone_Int_2_d[0],
                                                                                               lizzieLet14_1_4MQNode_3QNone_Int_1_d[0]} & {lizzieLet14_1_4MQNode_3QNone_Int_2_r,
                                                                                                                                           lizzieLet14_1_4MQNode_3QNone_Int_1_r}));
  assign lizzieLet14_1_4MQNode_3QNone_Int_r = (& lizzieLet14_1_4MQNode_3QNone_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet14_1_4MQNode_3QNone_Int_emitted <= 2'd0;
    else
      lizzieLet14_1_4MQNode_3QNone_Int_emitted <= (lizzieLet14_1_4MQNode_3QNone_Int_r ? 2'd0 :
                                                   lizzieLet14_1_4MQNode_3QNone_Int_done);
  
  /* dcon (Ty QTree_Int,
      Dcon QNone_Int) : [(lizzieLet14_1_4MQNode_3QNone_Int_1,Go)] > (lizzieLet14_1_4MQNode_3QNone_Int_1QNone_Int,QTree_Int) */
  assign lizzieLet14_1_4MQNode_3QNone_Int_1QNone_Int_d = QNone_Int_dc((& {lizzieLet14_1_4MQNode_3QNone_Int_1_d[0]}), lizzieLet14_1_4MQNode_3QNone_Int_1_d);
  assign {lizzieLet14_1_4MQNode_3QNone_Int_1_r} = {1 {(lizzieLet14_1_4MQNode_3QNone_Int_1QNone_Int_r && lizzieLet14_1_4MQNode_3QNone_Int_1QNone_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (lizzieLet14_1_4MQNode_3QNone_Int_1QNone_Int,QTree_Int) > (lizzieLet17_1_argbuf,QTree_Int) */
  QTree_Int_t lizzieLet14_1_4MQNode_3QNone_Int_1QNone_Int_bufchan_d;
  logic lizzieLet14_1_4MQNode_3QNone_Int_1QNone_Int_bufchan_r;
  assign lizzieLet14_1_4MQNode_3QNone_Int_1QNone_Int_r = ((! lizzieLet14_1_4MQNode_3QNone_Int_1QNone_Int_bufchan_d[0]) || lizzieLet14_1_4MQNode_3QNone_Int_1QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet14_1_4MQNode_3QNone_Int_1QNone_Int_bufchan_d <= {66'd0,
                                                                1'd0};
    else
      if (lizzieLet14_1_4MQNode_3QNone_Int_1QNone_Int_r)
        lizzieLet14_1_4MQNode_3QNone_Int_1QNone_Int_bufchan_d <= lizzieLet14_1_4MQNode_3QNone_Int_1QNone_Int_d;
  QTree_Int_t lizzieLet14_1_4MQNode_3QNone_Int_1QNone_Int_bufchan_buf;
  assign lizzieLet14_1_4MQNode_3QNone_Int_1QNone_Int_bufchan_r = (! lizzieLet14_1_4MQNode_3QNone_Int_1QNone_Int_bufchan_buf[0]);
  assign lizzieLet17_1_argbuf_d = (lizzieLet14_1_4MQNode_3QNone_Int_1QNone_Int_bufchan_buf[0] ? lizzieLet14_1_4MQNode_3QNone_Int_1QNone_Int_bufchan_buf :
                                   lizzieLet14_1_4MQNode_3QNone_Int_1QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet14_1_4MQNode_3QNone_Int_1QNone_Int_bufchan_buf <= {66'd0,
                                                                  1'd0};
    else
      if ((lizzieLet17_1_argbuf_r && lizzieLet14_1_4MQNode_3QNone_Int_1QNone_Int_bufchan_buf[0]))
        lizzieLet14_1_4MQNode_3QNone_Int_1QNone_Int_bufchan_buf <= {66'd0,
                                                                    1'd0};
      else if (((! lizzieLet17_1_argbuf_r) && (! lizzieLet14_1_4MQNode_3QNone_Int_1QNone_Int_bufchan_buf[0])))
        lizzieLet14_1_4MQNode_3QNone_Int_1QNone_Int_bufchan_buf <= lizzieLet14_1_4MQNode_3QNone_Int_1QNone_Int_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet14_1_4MQNode_3QNone_Int_2,Go) > (lizzieLet14_1_4MQNode_3QNone_Int_2_argbuf,Go) */
  Go_t lizzieLet14_1_4MQNode_3QNone_Int_2_bufchan_d;
  logic lizzieLet14_1_4MQNode_3QNone_Int_2_bufchan_r;
  assign lizzieLet14_1_4MQNode_3QNone_Int_2_r = ((! lizzieLet14_1_4MQNode_3QNone_Int_2_bufchan_d[0]) || lizzieLet14_1_4MQNode_3QNone_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet14_1_4MQNode_3QNone_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet14_1_4MQNode_3QNone_Int_2_r)
        lizzieLet14_1_4MQNode_3QNone_Int_2_bufchan_d <= lizzieLet14_1_4MQNode_3QNone_Int_2_d;
  Go_t lizzieLet14_1_4MQNode_3QNone_Int_2_bufchan_buf;
  assign lizzieLet14_1_4MQNode_3QNone_Int_2_bufchan_r = (! lizzieLet14_1_4MQNode_3QNone_Int_2_bufchan_buf[0]);
  assign lizzieLet14_1_4MQNode_3QNone_Int_2_argbuf_d = (lizzieLet14_1_4MQNode_3QNone_Int_2_bufchan_buf[0] ? lizzieLet14_1_4MQNode_3QNone_Int_2_bufchan_buf :
                                                        lizzieLet14_1_4MQNode_3QNone_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet14_1_4MQNode_3QNone_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet14_1_4MQNode_3QNone_Int_2_argbuf_r && lizzieLet14_1_4MQNode_3QNone_Int_2_bufchan_buf[0]))
        lizzieLet14_1_4MQNode_3QNone_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet14_1_4MQNode_3QNone_Int_2_argbuf_r) && (! lizzieLet14_1_4MQNode_3QNone_Int_2_bufchan_buf[0])))
        lizzieLet14_1_4MQNode_3QNone_Int_2_bufchan_buf <= lizzieLet14_1_4MQNode_3QNone_Int_2_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet14_1_4MQNode_3QVal_Int,Go) > [(lizzieLet14_1_4MQNode_3QVal_Int_1,Go),
                                                       (lizzieLet14_1_4MQNode_3QVal_Int_2,Go)] */
  logic [1:0] lizzieLet14_1_4MQNode_3QVal_Int_emitted;
  logic [1:0] lizzieLet14_1_4MQNode_3QVal_Int_done;
  assign lizzieLet14_1_4MQNode_3QVal_Int_1_d = (lizzieLet14_1_4MQNode_3QVal_Int_d[0] && (! lizzieLet14_1_4MQNode_3QVal_Int_emitted[0]));
  assign lizzieLet14_1_4MQNode_3QVal_Int_2_d = (lizzieLet14_1_4MQNode_3QVal_Int_d[0] && (! lizzieLet14_1_4MQNode_3QVal_Int_emitted[1]));
  assign lizzieLet14_1_4MQNode_3QVal_Int_done = (lizzieLet14_1_4MQNode_3QVal_Int_emitted | ({lizzieLet14_1_4MQNode_3QVal_Int_2_d[0],
                                                                                             lizzieLet14_1_4MQNode_3QVal_Int_1_d[0]} & {lizzieLet14_1_4MQNode_3QVal_Int_2_r,
                                                                                                                                        lizzieLet14_1_4MQNode_3QVal_Int_1_r}));
  assign lizzieLet14_1_4MQNode_3QVal_Int_r = (& lizzieLet14_1_4MQNode_3QVal_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet14_1_4MQNode_3QVal_Int_emitted <= 2'd0;
    else
      lizzieLet14_1_4MQNode_3QVal_Int_emitted <= (lizzieLet14_1_4MQNode_3QVal_Int_r ? 2'd0 :
                                                  lizzieLet14_1_4MQNode_3QVal_Int_done);
  
  /* dcon (Ty QTree_Int,
      Dcon QError_Int) : [(lizzieLet14_1_4MQNode_3QVal_Int_1,Go)] > (lizzieLet14_1_4MQNode_3QVal_Int_1QError_Int,QTree_Int) */
  assign lizzieLet14_1_4MQNode_3QVal_Int_1QError_Int_d = QError_Int_dc((& {lizzieLet14_1_4MQNode_3QVal_Int_1_d[0]}), lizzieLet14_1_4MQNode_3QVal_Int_1_d);
  assign {lizzieLet14_1_4MQNode_3QVal_Int_1_r} = {1 {(lizzieLet14_1_4MQNode_3QVal_Int_1QError_Int_r && lizzieLet14_1_4MQNode_3QVal_Int_1QError_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (lizzieLet14_1_4MQNode_3QVal_Int_1QError_Int,QTree_Int) > (lizzieLet18_1_argbuf,QTree_Int) */
  QTree_Int_t lizzieLet14_1_4MQNode_3QVal_Int_1QError_Int_bufchan_d;
  logic lizzieLet14_1_4MQNode_3QVal_Int_1QError_Int_bufchan_r;
  assign lizzieLet14_1_4MQNode_3QVal_Int_1QError_Int_r = ((! lizzieLet14_1_4MQNode_3QVal_Int_1QError_Int_bufchan_d[0]) || lizzieLet14_1_4MQNode_3QVal_Int_1QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet14_1_4MQNode_3QVal_Int_1QError_Int_bufchan_d <= {66'd0,
                                                                1'd0};
    else
      if (lizzieLet14_1_4MQNode_3QVal_Int_1QError_Int_r)
        lizzieLet14_1_4MQNode_3QVal_Int_1QError_Int_bufchan_d <= lizzieLet14_1_4MQNode_3QVal_Int_1QError_Int_d;
  QTree_Int_t lizzieLet14_1_4MQNode_3QVal_Int_1QError_Int_bufchan_buf;
  assign lizzieLet14_1_4MQNode_3QVal_Int_1QError_Int_bufchan_r = (! lizzieLet14_1_4MQNode_3QVal_Int_1QError_Int_bufchan_buf[0]);
  assign lizzieLet18_1_argbuf_d = (lizzieLet14_1_4MQNode_3QVal_Int_1QError_Int_bufchan_buf[0] ? lizzieLet14_1_4MQNode_3QVal_Int_1QError_Int_bufchan_buf :
                                   lizzieLet14_1_4MQNode_3QVal_Int_1QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet14_1_4MQNode_3QVal_Int_1QError_Int_bufchan_buf <= {66'd0,
                                                                  1'd0};
    else
      if ((lizzieLet18_1_argbuf_r && lizzieLet14_1_4MQNode_3QVal_Int_1QError_Int_bufchan_buf[0]))
        lizzieLet14_1_4MQNode_3QVal_Int_1QError_Int_bufchan_buf <= {66'd0,
                                                                    1'd0};
      else if (((! lizzieLet18_1_argbuf_r) && (! lizzieLet14_1_4MQNode_3QVal_Int_1QError_Int_bufchan_buf[0])))
        lizzieLet14_1_4MQNode_3QVal_Int_1QError_Int_bufchan_buf <= lizzieLet14_1_4MQNode_3QVal_Int_1QError_Int_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet14_1_4MQNode_3QVal_Int_2,Go) > (lizzieLet14_1_4MQNode_3QVal_Int_2_argbuf,Go) */
  Go_t lizzieLet14_1_4MQNode_3QVal_Int_2_bufchan_d;
  logic lizzieLet14_1_4MQNode_3QVal_Int_2_bufchan_r;
  assign lizzieLet14_1_4MQNode_3QVal_Int_2_r = ((! lizzieLet14_1_4MQNode_3QVal_Int_2_bufchan_d[0]) || lizzieLet14_1_4MQNode_3QVal_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet14_1_4MQNode_3QVal_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet14_1_4MQNode_3QVal_Int_2_r)
        lizzieLet14_1_4MQNode_3QVal_Int_2_bufchan_d <= lizzieLet14_1_4MQNode_3QVal_Int_2_d;
  Go_t lizzieLet14_1_4MQNode_3QVal_Int_2_bufchan_buf;
  assign lizzieLet14_1_4MQNode_3QVal_Int_2_bufchan_r = (! lizzieLet14_1_4MQNode_3QVal_Int_2_bufchan_buf[0]);
  assign lizzieLet14_1_4MQNode_3QVal_Int_2_argbuf_d = (lizzieLet14_1_4MQNode_3QVal_Int_2_bufchan_buf[0] ? lizzieLet14_1_4MQNode_3QVal_Int_2_bufchan_buf :
                                                       lizzieLet14_1_4MQNode_3QVal_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet14_1_4MQNode_3QVal_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet14_1_4MQNode_3QVal_Int_2_argbuf_r && lizzieLet14_1_4MQNode_3QVal_Int_2_bufchan_buf[0]))
        lizzieLet14_1_4MQNode_3QVal_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet14_1_4MQNode_3QVal_Int_2_argbuf_r) && (! lizzieLet14_1_4MQNode_3QVal_Int_2_bufchan_buf[0])))
        lizzieLet14_1_4MQNode_3QVal_Int_2_bufchan_buf <= lizzieLet14_1_4MQNode_3QVal_Int_2_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_CTmain_mask_Int) : (lizzieLet14_1_4MQNode_4,QTree_Int) (lizzieLet14_1_6MQNode,Pointer_CTmain_mask_Int) > [(lizzieLet14_1_4MQNode_4QNone_Int,Pointer_CTmain_mask_Int),
                                                                                                                            (lizzieLet14_1_4MQNode_4QVal_Int,Pointer_CTmain_mask_Int),
                                                                                                                            (lizzieLet14_1_4MQNode_4QNode_Int,Pointer_CTmain_mask_Int),
                                                                                                                            (lizzieLet14_1_4MQNode_4QError_Int,Pointer_CTmain_mask_Int)] */
  logic [3:0] lizzieLet14_1_6MQNode_onehotd;
  always_comb
    if ((lizzieLet14_1_4MQNode_4_d[0] && lizzieLet14_1_6MQNode_d[0]))
      unique case (lizzieLet14_1_4MQNode_4_d[2:1])
        2'd0: lizzieLet14_1_6MQNode_onehotd = 4'd1;
        2'd1: lizzieLet14_1_6MQNode_onehotd = 4'd2;
        2'd2: lizzieLet14_1_6MQNode_onehotd = 4'd4;
        2'd3: lizzieLet14_1_6MQNode_onehotd = 4'd8;
        default: lizzieLet14_1_6MQNode_onehotd = 4'd0;
      endcase
    else lizzieLet14_1_6MQNode_onehotd = 4'd0;
  assign lizzieLet14_1_4MQNode_4QNone_Int_d = {lizzieLet14_1_6MQNode_d[16:1],
                                               lizzieLet14_1_6MQNode_onehotd[0]};
  assign lizzieLet14_1_4MQNode_4QVal_Int_d = {lizzieLet14_1_6MQNode_d[16:1],
                                              lizzieLet14_1_6MQNode_onehotd[1]};
  assign lizzieLet14_1_4MQNode_4QNode_Int_d = {lizzieLet14_1_6MQNode_d[16:1],
                                               lizzieLet14_1_6MQNode_onehotd[2]};
  assign lizzieLet14_1_4MQNode_4QError_Int_d = {lizzieLet14_1_6MQNode_d[16:1],
                                                lizzieLet14_1_6MQNode_onehotd[3]};
  assign lizzieLet14_1_6MQNode_r = (| (lizzieLet14_1_6MQNode_onehotd & {lizzieLet14_1_4MQNode_4QError_Int_r,
                                                                        lizzieLet14_1_4MQNode_4QNode_Int_r,
                                                                        lizzieLet14_1_4MQNode_4QVal_Int_r,
                                                                        lizzieLet14_1_4MQNode_4QNone_Int_r}));
  assign lizzieLet14_1_4MQNode_4_r = lizzieLet14_1_6MQNode_r;
  
  /* buf (Ty Pointer_CTmain_mask_Int) : (lizzieLet14_1_4MQNode_4QError_Int,Pointer_CTmain_mask_Int) > (lizzieLet14_1_4MQNode_4QError_Int_1_argbuf,Pointer_CTmain_mask_Int) */
  Pointer_CTmain_mask_Int_t lizzieLet14_1_4MQNode_4QError_Int_bufchan_d;
  logic lizzieLet14_1_4MQNode_4QError_Int_bufchan_r;
  assign lizzieLet14_1_4MQNode_4QError_Int_r = ((! lizzieLet14_1_4MQNode_4QError_Int_bufchan_d[0]) || lizzieLet14_1_4MQNode_4QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet14_1_4MQNode_4QError_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet14_1_4MQNode_4QError_Int_r)
        lizzieLet14_1_4MQNode_4QError_Int_bufchan_d <= lizzieLet14_1_4MQNode_4QError_Int_d;
  Pointer_CTmain_mask_Int_t lizzieLet14_1_4MQNode_4QError_Int_bufchan_buf;
  assign lizzieLet14_1_4MQNode_4QError_Int_bufchan_r = (! lizzieLet14_1_4MQNode_4QError_Int_bufchan_buf[0]);
  assign lizzieLet14_1_4MQNode_4QError_Int_1_argbuf_d = (lizzieLet14_1_4MQNode_4QError_Int_bufchan_buf[0] ? lizzieLet14_1_4MQNode_4QError_Int_bufchan_buf :
                                                         lizzieLet14_1_4MQNode_4QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet14_1_4MQNode_4QError_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet14_1_4MQNode_4QError_Int_1_argbuf_r && lizzieLet14_1_4MQNode_4QError_Int_bufchan_buf[0]))
        lizzieLet14_1_4MQNode_4QError_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet14_1_4MQNode_4QError_Int_1_argbuf_r) && (! lizzieLet14_1_4MQNode_4QError_Int_bufchan_buf[0])))
        lizzieLet14_1_4MQNode_4QError_Int_bufchan_buf <= lizzieLet14_1_4MQNode_4QError_Int_bufchan_d;
  
  /* dcon (Ty CTmain_mask_Int,
      Dcon Lcall_main_mask_Int3) : [(lizzieLet14_1_4MQNode_4QNode_Int,Pointer_CTmain_mask_Int),
                                    (t1a8x_destruct,Pointer_QTree_Int),
                                    (lizzieLet14_1_4MQNode_5QNode_Int,Pointer_MaskQTree),
                                    (t2a8y_destruct,Pointer_QTree_Int),
                                    (lizzieLet14_1_4MQNode_6QNode_Int,Pointer_MaskQTree),
                                    (t3a8z_destruct,Pointer_QTree_Int),
                                    (lizzieLet14_1_4MQNode_7QNode_Int,Pointer_MaskQTree)] > (lizzieLet14_1_4MQNode_4QNode_Int_1t1a8x_1lizzieLet14_1_4MQNode_5QNode_Int_1t2a8y_1lizzieLet14_1_4MQNode_6QNode_Int_1t3a8z_1lizzieLet14_1_4MQNode_7QNode_Int_1Lcall_main_mask_Int3,CTmain_mask_Int) */
  assign lizzieLet14_1_4MQNode_4QNode_Int_1t1a8x_1lizzieLet14_1_4MQNode_5QNode_Int_1t2a8y_1lizzieLet14_1_4MQNode_6QNode_Int_1t3a8z_1lizzieLet14_1_4MQNode_7QNode_Int_1Lcall_main_mask_Int3_d = Lcall_main_mask_Int3_dc((& {lizzieLet14_1_4MQNode_4QNode_Int_d[0],
                                                                                                                                                                                                                           t1a8x_destruct_d[0],
                                                                                                                                                                                                                           lizzieLet14_1_4MQNode_5QNode_Int_d[0],
                                                                                                                                                                                                                           t2a8y_destruct_d[0],
                                                                                                                                                                                                                           lizzieLet14_1_4MQNode_6QNode_Int_d[0],
                                                                                                                                                                                                                           t3a8z_destruct_d[0],
                                                                                                                                                                                                                           lizzieLet14_1_4MQNode_7QNode_Int_d[0]}), lizzieLet14_1_4MQNode_4QNode_Int_d, t1a8x_destruct_d, lizzieLet14_1_4MQNode_5QNode_Int_d, t2a8y_destruct_d, lizzieLet14_1_4MQNode_6QNode_Int_d, t3a8z_destruct_d, lizzieLet14_1_4MQNode_7QNode_Int_d);
  assign {lizzieLet14_1_4MQNode_4QNode_Int_r,
          t1a8x_destruct_r,
          lizzieLet14_1_4MQNode_5QNode_Int_r,
          t2a8y_destruct_r,
          lizzieLet14_1_4MQNode_6QNode_Int_r,
          t3a8z_destruct_r,
          lizzieLet14_1_4MQNode_7QNode_Int_r} = {7 {(lizzieLet14_1_4MQNode_4QNode_Int_1t1a8x_1lizzieLet14_1_4MQNode_5QNode_Int_1t2a8y_1lizzieLet14_1_4MQNode_6QNode_Int_1t3a8z_1lizzieLet14_1_4MQNode_7QNode_Int_1Lcall_main_mask_Int3_r && lizzieLet14_1_4MQNode_4QNode_Int_1t1a8x_1lizzieLet14_1_4MQNode_5QNode_Int_1t2a8y_1lizzieLet14_1_4MQNode_6QNode_Int_1t3a8z_1lizzieLet14_1_4MQNode_7QNode_Int_1Lcall_main_mask_Int3_d[0])}};
  
  /* buf (Ty CTmain_mask_Int) : (lizzieLet14_1_4MQNode_4QNode_Int_1t1a8x_1lizzieLet14_1_4MQNode_5QNode_Int_1t2a8y_1lizzieLet14_1_4MQNode_6QNode_Int_1t3a8z_1lizzieLet14_1_4MQNode_7QNode_Int_1Lcall_main_mask_Int3,CTmain_mask_Int) > (lizzieLet19_1_argbuf,CTmain_mask_Int) */
  CTmain_mask_Int_t lizzieLet14_1_4MQNode_4QNode_Int_1t1a8x_1lizzieLet14_1_4MQNode_5QNode_Int_1t2a8y_1lizzieLet14_1_4MQNode_6QNode_Int_1t3a8z_1lizzieLet14_1_4MQNode_7QNode_Int_1Lcall_main_mask_Int3_bufchan_d;
  logic lizzieLet14_1_4MQNode_4QNode_Int_1t1a8x_1lizzieLet14_1_4MQNode_5QNode_Int_1t2a8y_1lizzieLet14_1_4MQNode_6QNode_Int_1t3a8z_1lizzieLet14_1_4MQNode_7QNode_Int_1Lcall_main_mask_Int3_bufchan_r;
  assign lizzieLet14_1_4MQNode_4QNode_Int_1t1a8x_1lizzieLet14_1_4MQNode_5QNode_Int_1t2a8y_1lizzieLet14_1_4MQNode_6QNode_Int_1t3a8z_1lizzieLet14_1_4MQNode_7QNode_Int_1Lcall_main_mask_Int3_r = ((! lizzieLet14_1_4MQNode_4QNode_Int_1t1a8x_1lizzieLet14_1_4MQNode_5QNode_Int_1t2a8y_1lizzieLet14_1_4MQNode_6QNode_Int_1t3a8z_1lizzieLet14_1_4MQNode_7QNode_Int_1Lcall_main_mask_Int3_bufchan_d[0]) || lizzieLet14_1_4MQNode_4QNode_Int_1t1a8x_1lizzieLet14_1_4MQNode_5QNode_Int_1t2a8y_1lizzieLet14_1_4MQNode_6QNode_Int_1t3a8z_1lizzieLet14_1_4MQNode_7QNode_Int_1Lcall_main_mask_Int3_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet14_1_4MQNode_4QNode_Int_1t1a8x_1lizzieLet14_1_4MQNode_5QNode_Int_1t2a8y_1lizzieLet14_1_4MQNode_6QNode_Int_1t3a8z_1lizzieLet14_1_4MQNode_7QNode_Int_1Lcall_main_mask_Int3_bufchan_d <= {115'd0,
                                                                                                                                                                                                      1'd0};
    else
      if (lizzieLet14_1_4MQNode_4QNode_Int_1t1a8x_1lizzieLet14_1_4MQNode_5QNode_Int_1t2a8y_1lizzieLet14_1_4MQNode_6QNode_Int_1t3a8z_1lizzieLet14_1_4MQNode_7QNode_Int_1Lcall_main_mask_Int3_r)
        lizzieLet14_1_4MQNode_4QNode_Int_1t1a8x_1lizzieLet14_1_4MQNode_5QNode_Int_1t2a8y_1lizzieLet14_1_4MQNode_6QNode_Int_1t3a8z_1lizzieLet14_1_4MQNode_7QNode_Int_1Lcall_main_mask_Int3_bufchan_d <= lizzieLet14_1_4MQNode_4QNode_Int_1t1a8x_1lizzieLet14_1_4MQNode_5QNode_Int_1t2a8y_1lizzieLet14_1_4MQNode_6QNode_Int_1t3a8z_1lizzieLet14_1_4MQNode_7QNode_Int_1Lcall_main_mask_Int3_d;
  CTmain_mask_Int_t lizzieLet14_1_4MQNode_4QNode_Int_1t1a8x_1lizzieLet14_1_4MQNode_5QNode_Int_1t2a8y_1lizzieLet14_1_4MQNode_6QNode_Int_1t3a8z_1lizzieLet14_1_4MQNode_7QNode_Int_1Lcall_main_mask_Int3_bufchan_buf;
  assign lizzieLet14_1_4MQNode_4QNode_Int_1t1a8x_1lizzieLet14_1_4MQNode_5QNode_Int_1t2a8y_1lizzieLet14_1_4MQNode_6QNode_Int_1t3a8z_1lizzieLet14_1_4MQNode_7QNode_Int_1Lcall_main_mask_Int3_bufchan_r = (! lizzieLet14_1_4MQNode_4QNode_Int_1t1a8x_1lizzieLet14_1_4MQNode_5QNode_Int_1t2a8y_1lizzieLet14_1_4MQNode_6QNode_Int_1t3a8z_1lizzieLet14_1_4MQNode_7QNode_Int_1Lcall_main_mask_Int3_bufchan_buf[0]);
  assign lizzieLet19_1_argbuf_d = (lizzieLet14_1_4MQNode_4QNode_Int_1t1a8x_1lizzieLet14_1_4MQNode_5QNode_Int_1t2a8y_1lizzieLet14_1_4MQNode_6QNode_Int_1t3a8z_1lizzieLet14_1_4MQNode_7QNode_Int_1Lcall_main_mask_Int3_bufchan_buf[0] ? lizzieLet14_1_4MQNode_4QNode_Int_1t1a8x_1lizzieLet14_1_4MQNode_5QNode_Int_1t2a8y_1lizzieLet14_1_4MQNode_6QNode_Int_1t3a8z_1lizzieLet14_1_4MQNode_7QNode_Int_1Lcall_main_mask_Int3_bufchan_buf :
                                   lizzieLet14_1_4MQNode_4QNode_Int_1t1a8x_1lizzieLet14_1_4MQNode_5QNode_Int_1t2a8y_1lizzieLet14_1_4MQNode_6QNode_Int_1t3a8z_1lizzieLet14_1_4MQNode_7QNode_Int_1Lcall_main_mask_Int3_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet14_1_4MQNode_4QNode_Int_1t1a8x_1lizzieLet14_1_4MQNode_5QNode_Int_1t2a8y_1lizzieLet14_1_4MQNode_6QNode_Int_1t3a8z_1lizzieLet14_1_4MQNode_7QNode_Int_1Lcall_main_mask_Int3_bufchan_buf <= {115'd0,
                                                                                                                                                                                                        1'd0};
    else
      if ((lizzieLet19_1_argbuf_r && lizzieLet14_1_4MQNode_4QNode_Int_1t1a8x_1lizzieLet14_1_4MQNode_5QNode_Int_1t2a8y_1lizzieLet14_1_4MQNode_6QNode_Int_1t3a8z_1lizzieLet14_1_4MQNode_7QNode_Int_1Lcall_main_mask_Int3_bufchan_buf[0]))
        lizzieLet14_1_4MQNode_4QNode_Int_1t1a8x_1lizzieLet14_1_4MQNode_5QNode_Int_1t2a8y_1lizzieLet14_1_4MQNode_6QNode_Int_1t3a8z_1lizzieLet14_1_4MQNode_7QNode_Int_1Lcall_main_mask_Int3_bufchan_buf <= {115'd0,
                                                                                                                                                                                                          1'd0};
      else if (((! lizzieLet19_1_argbuf_r) && (! lizzieLet14_1_4MQNode_4QNode_Int_1t1a8x_1lizzieLet14_1_4MQNode_5QNode_Int_1t2a8y_1lizzieLet14_1_4MQNode_6QNode_Int_1t3a8z_1lizzieLet14_1_4MQNode_7QNode_Int_1Lcall_main_mask_Int3_bufchan_buf[0])))
        lizzieLet14_1_4MQNode_4QNode_Int_1t1a8x_1lizzieLet14_1_4MQNode_5QNode_Int_1t2a8y_1lizzieLet14_1_4MQNode_6QNode_Int_1t3a8z_1lizzieLet14_1_4MQNode_7QNode_Int_1Lcall_main_mask_Int3_bufchan_buf <= lizzieLet14_1_4MQNode_4QNode_Int_1t1a8x_1lizzieLet14_1_4MQNode_5QNode_Int_1t2a8y_1lizzieLet14_1_4MQNode_6QNode_Int_1t3a8z_1lizzieLet14_1_4MQNode_7QNode_Int_1Lcall_main_mask_Int3_bufchan_d;
  
  /* buf (Ty Pointer_CTmain_mask_Int) : (lizzieLet14_1_4MQNode_4QNone_Int,Pointer_CTmain_mask_Int) > (lizzieLet14_1_4MQNode_4QNone_Int_1_argbuf,Pointer_CTmain_mask_Int) */
  Pointer_CTmain_mask_Int_t lizzieLet14_1_4MQNode_4QNone_Int_bufchan_d;
  logic lizzieLet14_1_4MQNode_4QNone_Int_bufchan_r;
  assign lizzieLet14_1_4MQNode_4QNone_Int_r = ((! lizzieLet14_1_4MQNode_4QNone_Int_bufchan_d[0]) || lizzieLet14_1_4MQNode_4QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet14_1_4MQNode_4QNone_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet14_1_4MQNode_4QNone_Int_r)
        lizzieLet14_1_4MQNode_4QNone_Int_bufchan_d <= lizzieLet14_1_4MQNode_4QNone_Int_d;
  Pointer_CTmain_mask_Int_t lizzieLet14_1_4MQNode_4QNone_Int_bufchan_buf;
  assign lizzieLet14_1_4MQNode_4QNone_Int_bufchan_r = (! lizzieLet14_1_4MQNode_4QNone_Int_bufchan_buf[0]);
  assign lizzieLet14_1_4MQNode_4QNone_Int_1_argbuf_d = (lizzieLet14_1_4MQNode_4QNone_Int_bufchan_buf[0] ? lizzieLet14_1_4MQNode_4QNone_Int_bufchan_buf :
                                                        lizzieLet14_1_4MQNode_4QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet14_1_4MQNode_4QNone_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet14_1_4MQNode_4QNone_Int_1_argbuf_r && lizzieLet14_1_4MQNode_4QNone_Int_bufchan_buf[0]))
        lizzieLet14_1_4MQNode_4QNone_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet14_1_4MQNode_4QNone_Int_1_argbuf_r) && (! lizzieLet14_1_4MQNode_4QNone_Int_bufchan_buf[0])))
        lizzieLet14_1_4MQNode_4QNone_Int_bufchan_buf <= lizzieLet14_1_4MQNode_4QNone_Int_bufchan_d;
  
  /* buf (Ty Pointer_CTmain_mask_Int) : (lizzieLet14_1_4MQNode_4QVal_Int,Pointer_CTmain_mask_Int) > (lizzieLet14_1_4MQNode_4QVal_Int_1_argbuf,Pointer_CTmain_mask_Int) */
  Pointer_CTmain_mask_Int_t lizzieLet14_1_4MQNode_4QVal_Int_bufchan_d;
  logic lizzieLet14_1_4MQNode_4QVal_Int_bufchan_r;
  assign lizzieLet14_1_4MQNode_4QVal_Int_r = ((! lizzieLet14_1_4MQNode_4QVal_Int_bufchan_d[0]) || lizzieLet14_1_4MQNode_4QVal_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet14_1_4MQNode_4QVal_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet14_1_4MQNode_4QVal_Int_r)
        lizzieLet14_1_4MQNode_4QVal_Int_bufchan_d <= lizzieLet14_1_4MQNode_4QVal_Int_d;
  Pointer_CTmain_mask_Int_t lizzieLet14_1_4MQNode_4QVal_Int_bufchan_buf;
  assign lizzieLet14_1_4MQNode_4QVal_Int_bufchan_r = (! lizzieLet14_1_4MQNode_4QVal_Int_bufchan_buf[0]);
  assign lizzieLet14_1_4MQNode_4QVal_Int_1_argbuf_d = (lizzieLet14_1_4MQNode_4QVal_Int_bufchan_buf[0] ? lizzieLet14_1_4MQNode_4QVal_Int_bufchan_buf :
                                                       lizzieLet14_1_4MQNode_4QVal_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet14_1_4MQNode_4QVal_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet14_1_4MQNode_4QVal_Int_1_argbuf_r && lizzieLet14_1_4MQNode_4QVal_Int_bufchan_buf[0]))
        lizzieLet14_1_4MQNode_4QVal_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet14_1_4MQNode_4QVal_Int_1_argbuf_r) && (! lizzieLet14_1_4MQNode_4QVal_Int_bufchan_buf[0])))
        lizzieLet14_1_4MQNode_4QVal_Int_bufchan_buf <= lizzieLet14_1_4MQNode_4QVal_Int_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_MaskQTree) : (lizzieLet14_1_4MQNode_5,QTree_Int) (q1a8s_destruct,Pointer_MaskQTree) > [(_63,Pointer_MaskQTree),
                                                                                                         (_62,Pointer_MaskQTree),
                                                                                                         (lizzieLet14_1_4MQNode_5QNode_Int,Pointer_MaskQTree),
                                                                                                         (_61,Pointer_MaskQTree)] */
  logic [3:0] q1a8s_destruct_onehotd;
  always_comb
    if ((lizzieLet14_1_4MQNode_5_d[0] && q1a8s_destruct_d[0]))
      unique case (lizzieLet14_1_4MQNode_5_d[2:1])
        2'd0: q1a8s_destruct_onehotd = 4'd1;
        2'd1: q1a8s_destruct_onehotd = 4'd2;
        2'd2: q1a8s_destruct_onehotd = 4'd4;
        2'd3: q1a8s_destruct_onehotd = 4'd8;
        default: q1a8s_destruct_onehotd = 4'd0;
      endcase
    else q1a8s_destruct_onehotd = 4'd0;
  assign _63_d = {q1a8s_destruct_d[16:1], q1a8s_destruct_onehotd[0]};
  assign _62_d = {q1a8s_destruct_d[16:1], q1a8s_destruct_onehotd[1]};
  assign lizzieLet14_1_4MQNode_5QNode_Int_d = {q1a8s_destruct_d[16:1],
                                               q1a8s_destruct_onehotd[2]};
  assign _61_d = {q1a8s_destruct_d[16:1], q1a8s_destruct_onehotd[3]};
  assign q1a8s_destruct_r = (| (q1a8s_destruct_onehotd & {_61_r,
                                                          lizzieLet14_1_4MQNode_5QNode_Int_r,
                                                          _62_r,
                                                          _63_r}));
  assign lizzieLet14_1_4MQNode_5_r = q1a8s_destruct_r;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_MaskQTree) : (lizzieLet14_1_4MQNode_6,QTree_Int) (q2a8t_destruct,Pointer_MaskQTree) > [(_60,Pointer_MaskQTree),
                                                                                                         (_59,Pointer_MaskQTree),
                                                                                                         (lizzieLet14_1_4MQNode_6QNode_Int,Pointer_MaskQTree),
                                                                                                         (_58,Pointer_MaskQTree)] */
  logic [3:0] q2a8t_destruct_onehotd;
  always_comb
    if ((lizzieLet14_1_4MQNode_6_d[0] && q2a8t_destruct_d[0]))
      unique case (lizzieLet14_1_4MQNode_6_d[2:1])
        2'd0: q2a8t_destruct_onehotd = 4'd1;
        2'd1: q2a8t_destruct_onehotd = 4'd2;
        2'd2: q2a8t_destruct_onehotd = 4'd4;
        2'd3: q2a8t_destruct_onehotd = 4'd8;
        default: q2a8t_destruct_onehotd = 4'd0;
      endcase
    else q2a8t_destruct_onehotd = 4'd0;
  assign _60_d = {q2a8t_destruct_d[16:1], q2a8t_destruct_onehotd[0]};
  assign _59_d = {q2a8t_destruct_d[16:1], q2a8t_destruct_onehotd[1]};
  assign lizzieLet14_1_4MQNode_6QNode_Int_d = {q2a8t_destruct_d[16:1],
                                               q2a8t_destruct_onehotd[2]};
  assign _58_d = {q2a8t_destruct_d[16:1], q2a8t_destruct_onehotd[3]};
  assign q2a8t_destruct_r = (| (q2a8t_destruct_onehotd & {_58_r,
                                                          lizzieLet14_1_4MQNode_6QNode_Int_r,
                                                          _59_r,
                                                          _60_r}));
  assign lizzieLet14_1_4MQNode_6_r = q2a8t_destruct_r;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_MaskQTree) : (lizzieLet14_1_4MQNode_7,QTree_Int) (q3a8u_destruct,Pointer_MaskQTree) > [(_57,Pointer_MaskQTree),
                                                                                                         (_56,Pointer_MaskQTree),
                                                                                                         (lizzieLet14_1_4MQNode_7QNode_Int,Pointer_MaskQTree),
                                                                                                         (_55,Pointer_MaskQTree)] */
  logic [3:0] q3a8u_destruct_onehotd;
  always_comb
    if ((lizzieLet14_1_4MQNode_7_d[0] && q3a8u_destruct_d[0]))
      unique case (lizzieLet14_1_4MQNode_7_d[2:1])
        2'd0: q3a8u_destruct_onehotd = 4'd1;
        2'd1: q3a8u_destruct_onehotd = 4'd2;
        2'd2: q3a8u_destruct_onehotd = 4'd4;
        2'd3: q3a8u_destruct_onehotd = 4'd8;
        default: q3a8u_destruct_onehotd = 4'd0;
      endcase
    else q3a8u_destruct_onehotd = 4'd0;
  assign _57_d = {q3a8u_destruct_d[16:1], q3a8u_destruct_onehotd[0]};
  assign _56_d = {q3a8u_destruct_d[16:1], q3a8u_destruct_onehotd[1]};
  assign lizzieLet14_1_4MQNode_7QNode_Int_d = {q3a8u_destruct_d[16:1],
                                               q3a8u_destruct_onehotd[2]};
  assign _55_d = {q3a8u_destruct_d[16:1], q3a8u_destruct_onehotd[3]};
  assign q3a8u_destruct_r = (| (q3a8u_destruct_onehotd & {_55_r,
                                                          lizzieLet14_1_4MQNode_7QNode_Int_r,
                                                          _56_r,
                                                          _57_r}));
  assign lizzieLet14_1_4MQNode_7_r = q3a8u_destruct_r;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_MaskQTree) : (lizzieLet14_1_4MQNode_8,QTree_Int) (q4a8v_destruct,Pointer_MaskQTree) > [(_54,Pointer_MaskQTree),
                                                                                                         (_53,Pointer_MaskQTree),
                                                                                                         (lizzieLet14_1_4MQNode_8QNode_Int,Pointer_MaskQTree),
                                                                                                         (_52,Pointer_MaskQTree)] */
  logic [3:0] q4a8v_destruct_onehotd;
  always_comb
    if ((lizzieLet14_1_4MQNode_8_d[0] && q4a8v_destruct_d[0]))
      unique case (lizzieLet14_1_4MQNode_8_d[2:1])
        2'd0: q4a8v_destruct_onehotd = 4'd1;
        2'd1: q4a8v_destruct_onehotd = 4'd2;
        2'd2: q4a8v_destruct_onehotd = 4'd4;
        2'd3: q4a8v_destruct_onehotd = 4'd8;
        default: q4a8v_destruct_onehotd = 4'd0;
      endcase
    else q4a8v_destruct_onehotd = 4'd0;
  assign _54_d = {q4a8v_destruct_d[16:1], q4a8v_destruct_onehotd[0]};
  assign _53_d = {q4a8v_destruct_d[16:1], q4a8v_destruct_onehotd[1]};
  assign lizzieLet14_1_4MQNode_8QNode_Int_d = {q4a8v_destruct_d[16:1],
                                               q4a8v_destruct_onehotd[2]};
  assign _52_d = {q4a8v_destruct_d[16:1], q4a8v_destruct_onehotd[3]};
  assign q4a8v_destruct_r = (| (q4a8v_destruct_onehotd & {_52_r,
                                                          lizzieLet14_1_4MQNode_8QNode_Int_r,
                                                          _53_r,
                                                          _54_r}));
  assign lizzieLet14_1_4MQNode_8_r = q4a8v_destruct_r;
  
  /* buf (Ty Pointer_MaskQTree) : (lizzieLet14_1_4MQNode_8QNode_Int,Pointer_MaskQTree) > (lizzieLet14_1_4MQNode_8QNode_Int_1_argbuf,Pointer_MaskQTree) */
  Pointer_MaskQTree_t lizzieLet14_1_4MQNode_8QNode_Int_bufchan_d;
  logic lizzieLet14_1_4MQNode_8QNode_Int_bufchan_r;
  assign lizzieLet14_1_4MQNode_8QNode_Int_r = ((! lizzieLet14_1_4MQNode_8QNode_Int_bufchan_d[0]) || lizzieLet14_1_4MQNode_8QNode_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet14_1_4MQNode_8QNode_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet14_1_4MQNode_8QNode_Int_r)
        lizzieLet14_1_4MQNode_8QNode_Int_bufchan_d <= lizzieLet14_1_4MQNode_8QNode_Int_d;
  Pointer_MaskQTree_t lizzieLet14_1_4MQNode_8QNode_Int_bufchan_buf;
  assign lizzieLet14_1_4MQNode_8QNode_Int_bufchan_r = (! lizzieLet14_1_4MQNode_8QNode_Int_bufchan_buf[0]);
  assign lizzieLet14_1_4MQNode_8QNode_Int_1_argbuf_d = (lizzieLet14_1_4MQNode_8QNode_Int_bufchan_buf[0] ? lizzieLet14_1_4MQNode_8QNode_Int_bufchan_buf :
                                                        lizzieLet14_1_4MQNode_8QNode_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet14_1_4MQNode_8QNode_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet14_1_4MQNode_8QNode_Int_1_argbuf_r && lizzieLet14_1_4MQNode_8QNode_Int_bufchan_buf[0]))
        lizzieLet14_1_4MQNode_8QNode_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet14_1_4MQNode_8QNode_Int_1_argbuf_r) && (! lizzieLet14_1_4MQNode_8QNode_Int_bufchan_buf[0])))
        lizzieLet14_1_4MQNode_8QNode_Int_bufchan_buf <= lizzieLet14_1_4MQNode_8QNode_Int_bufchan_d;
  
  /* demux (Ty MaskQTree,
       Ty Pointer_QTree_Int) : (lizzieLet14_1_5,MaskQTree) (ma8q_2,Pointer_QTree_Int) > [(_51,Pointer_QTree_Int),
                                                                                         (lizzieLet14_1_5MQVal,Pointer_QTree_Int),
                                                                                         (_50,Pointer_QTree_Int)] */
  logic [2:0] ma8q_2_onehotd;
  always_comb
    if ((lizzieLet14_1_5_d[0] && ma8q_2_d[0]))
      unique case (lizzieLet14_1_5_d[2:1])
        2'd0: ma8q_2_onehotd = 3'd1;
        2'd1: ma8q_2_onehotd = 3'd2;
        2'd2: ma8q_2_onehotd = 3'd4;
        default: ma8q_2_onehotd = 3'd0;
      endcase
    else ma8q_2_onehotd = 3'd0;
  assign _51_d = {ma8q_2_d[16:1], ma8q_2_onehotd[0]};
  assign lizzieLet14_1_5MQVal_d = {ma8q_2_d[16:1],
                                   ma8q_2_onehotd[1]};
  assign _50_d = {ma8q_2_d[16:1], ma8q_2_onehotd[2]};
  assign ma8q_2_r = (| (ma8q_2_onehotd & {_50_r,
                                          lizzieLet14_1_5MQVal_r,
                                          _51_r}));
  assign lizzieLet14_1_5_r = ma8q_2_r;
  
  /* buf (Ty Pointer_QTree_Int) : (lizzieLet14_1_5MQVal,Pointer_QTree_Int) > (lizzieLet14_1_5MQVal_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t lizzieLet14_1_5MQVal_bufchan_d;
  logic lizzieLet14_1_5MQVal_bufchan_r;
  assign lizzieLet14_1_5MQVal_r = ((! lizzieLet14_1_5MQVal_bufchan_d[0]) || lizzieLet14_1_5MQVal_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet14_1_5MQVal_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet14_1_5MQVal_r)
        lizzieLet14_1_5MQVal_bufchan_d <= lizzieLet14_1_5MQVal_d;
  Pointer_QTree_Int_t lizzieLet14_1_5MQVal_bufchan_buf;
  assign lizzieLet14_1_5MQVal_bufchan_r = (! lizzieLet14_1_5MQVal_bufchan_buf[0]);
  assign lizzieLet14_1_5MQVal_1_argbuf_d = (lizzieLet14_1_5MQVal_bufchan_buf[0] ? lizzieLet14_1_5MQVal_bufchan_buf :
                                            lizzieLet14_1_5MQVal_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet14_1_5MQVal_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet14_1_5MQVal_1_argbuf_r && lizzieLet14_1_5MQVal_bufchan_buf[0]))
        lizzieLet14_1_5MQVal_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet14_1_5MQVal_1_argbuf_r) && (! lizzieLet14_1_5MQVal_bufchan_buf[0])))
        lizzieLet14_1_5MQVal_bufchan_buf <= lizzieLet14_1_5MQVal_bufchan_d;
  
  /* demux (Ty MaskQTree,
       Ty Pointer_CTmain_mask_Int) : (lizzieLet14_1_6,MaskQTree) (sc_0_2_goMux_mux,Pointer_CTmain_mask_Int) > [(lizzieLet14_1_6MQNone,Pointer_CTmain_mask_Int),
                                                                                                               (lizzieLet14_1_6MQVal,Pointer_CTmain_mask_Int),
                                                                                                               (lizzieLet14_1_6MQNode,Pointer_CTmain_mask_Int)] */
  logic [2:0] sc_0_2_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet14_1_6_d[0] && sc_0_2_goMux_mux_d[0]))
      unique case (lizzieLet14_1_6_d[2:1])
        2'd0: sc_0_2_goMux_mux_onehotd = 3'd1;
        2'd1: sc_0_2_goMux_mux_onehotd = 3'd2;
        2'd2: sc_0_2_goMux_mux_onehotd = 3'd4;
        default: sc_0_2_goMux_mux_onehotd = 3'd0;
      endcase
    else sc_0_2_goMux_mux_onehotd = 3'd0;
  assign lizzieLet14_1_6MQNone_d = {sc_0_2_goMux_mux_d[16:1],
                                    sc_0_2_goMux_mux_onehotd[0]};
  assign lizzieLet14_1_6MQVal_d = {sc_0_2_goMux_mux_d[16:1],
                                   sc_0_2_goMux_mux_onehotd[1]};
  assign lizzieLet14_1_6MQNode_d = {sc_0_2_goMux_mux_d[16:1],
                                    sc_0_2_goMux_mux_onehotd[2]};
  assign sc_0_2_goMux_mux_r = (| (sc_0_2_goMux_mux_onehotd & {lizzieLet14_1_6MQNode_r,
                                                              lizzieLet14_1_6MQVal_r,
                                                              lizzieLet14_1_6MQNone_r}));
  assign lizzieLet14_1_6_r = sc_0_2_goMux_mux_r;
  
  /* buf (Ty Pointer_CTmain_mask_Int) : (lizzieLet14_1_6MQNone,Pointer_CTmain_mask_Int) > (lizzieLet14_1_6MQNone_1_argbuf,Pointer_CTmain_mask_Int) */
  Pointer_CTmain_mask_Int_t lizzieLet14_1_6MQNone_bufchan_d;
  logic lizzieLet14_1_6MQNone_bufchan_r;
  assign lizzieLet14_1_6MQNone_r = ((! lizzieLet14_1_6MQNone_bufchan_d[0]) || lizzieLet14_1_6MQNone_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet14_1_6MQNone_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet14_1_6MQNone_r)
        lizzieLet14_1_6MQNone_bufchan_d <= lizzieLet14_1_6MQNone_d;
  Pointer_CTmain_mask_Int_t lizzieLet14_1_6MQNone_bufchan_buf;
  assign lizzieLet14_1_6MQNone_bufchan_r = (! lizzieLet14_1_6MQNone_bufchan_buf[0]);
  assign lizzieLet14_1_6MQNone_1_argbuf_d = (lizzieLet14_1_6MQNone_bufchan_buf[0] ? lizzieLet14_1_6MQNone_bufchan_buf :
                                             lizzieLet14_1_6MQNone_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet14_1_6MQNone_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet14_1_6MQNone_1_argbuf_r && lizzieLet14_1_6MQNone_bufchan_buf[0]))
        lizzieLet14_1_6MQNone_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet14_1_6MQNone_1_argbuf_r) && (! lizzieLet14_1_6MQNone_bufchan_buf[0])))
        lizzieLet14_1_6MQNone_bufchan_buf <= lizzieLet14_1_6MQNone_bufchan_d;
  
  /* buf (Ty Pointer_CTmain_mask_Int) : (lizzieLet14_1_6MQVal,Pointer_CTmain_mask_Int) > (lizzieLet14_1_6MQVal_1_argbuf,Pointer_CTmain_mask_Int) */
  Pointer_CTmain_mask_Int_t lizzieLet14_1_6MQVal_bufchan_d;
  logic lizzieLet14_1_6MQVal_bufchan_r;
  assign lizzieLet14_1_6MQVal_r = ((! lizzieLet14_1_6MQVal_bufchan_d[0]) || lizzieLet14_1_6MQVal_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet14_1_6MQVal_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet14_1_6MQVal_r)
        lizzieLet14_1_6MQVal_bufchan_d <= lizzieLet14_1_6MQVal_d;
  Pointer_CTmain_mask_Int_t lizzieLet14_1_6MQVal_bufchan_buf;
  assign lizzieLet14_1_6MQVal_bufchan_r = (! lizzieLet14_1_6MQVal_bufchan_buf[0]);
  assign lizzieLet14_1_6MQVal_1_argbuf_d = (lizzieLet14_1_6MQVal_bufchan_buf[0] ? lizzieLet14_1_6MQVal_bufchan_buf :
                                            lizzieLet14_1_6MQVal_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet14_1_6MQVal_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet14_1_6MQVal_1_argbuf_r && lizzieLet14_1_6MQVal_bufchan_buf[0]))
        lizzieLet14_1_6MQVal_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet14_1_6MQVal_1_argbuf_r) && (! lizzieLet14_1_6MQVal_bufchan_buf[0])))
        lizzieLet14_1_6MQVal_bufchan_buf <= lizzieLet14_1_6MQVal_bufchan_d;
  
  /* destruct (Ty CT$wmAdd_Int,
          Dcon Lcall_$wmAdd_Int0) : (lizzieLet22_1Lcall_$wmAdd_Int0,CT$wmAdd_Int) > [(es_2_destruct,Pointer_QTree_Int),
                                                                                     (es_3_2_destruct,Pointer_QTree_Int),
                                                                                     (es_4_2_destruct,Pointer_QTree_Int),
                                                                                     (sc_0_6_destruct,Pointer_CT$wmAdd_Int)] */
  logic [3:0] lizzieLet22_1Lcall_$wmAdd_Int0_emitted;
  logic [3:0] lizzieLet22_1Lcall_$wmAdd_Int0_done;
  assign es_2_destruct_d = {lizzieLet22_1Lcall_$wmAdd_Int0_d[19:4],
                            (lizzieLet22_1Lcall_$wmAdd_Int0_d[0] && (! lizzieLet22_1Lcall_$wmAdd_Int0_emitted[0]))};
  assign es_3_2_destruct_d = {lizzieLet22_1Lcall_$wmAdd_Int0_d[35:20],
                              (lizzieLet22_1Lcall_$wmAdd_Int0_d[0] && (! lizzieLet22_1Lcall_$wmAdd_Int0_emitted[1]))};
  assign es_4_2_destruct_d = {lizzieLet22_1Lcall_$wmAdd_Int0_d[51:36],
                              (lizzieLet22_1Lcall_$wmAdd_Int0_d[0] && (! lizzieLet22_1Lcall_$wmAdd_Int0_emitted[2]))};
  assign sc_0_6_destruct_d = {lizzieLet22_1Lcall_$wmAdd_Int0_d[67:52],
                              (lizzieLet22_1Lcall_$wmAdd_Int0_d[0] && (! lizzieLet22_1Lcall_$wmAdd_Int0_emitted[3]))};
  assign lizzieLet22_1Lcall_$wmAdd_Int0_done = (lizzieLet22_1Lcall_$wmAdd_Int0_emitted | ({sc_0_6_destruct_d[0],
                                                                                           es_4_2_destruct_d[0],
                                                                                           es_3_2_destruct_d[0],
                                                                                           es_2_destruct_d[0]} & {sc_0_6_destruct_r,
                                                                                                                  es_4_2_destruct_r,
                                                                                                                  es_3_2_destruct_r,
                                                                                                                  es_2_destruct_r}));
  assign lizzieLet22_1Lcall_$wmAdd_Int0_r = (& lizzieLet22_1Lcall_$wmAdd_Int0_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet22_1Lcall_$wmAdd_Int0_emitted <= 4'd0;
    else
      lizzieLet22_1Lcall_$wmAdd_Int0_emitted <= (lizzieLet22_1Lcall_$wmAdd_Int0_r ? 4'd0 :
                                                 lizzieLet22_1Lcall_$wmAdd_Int0_done);
  
  /* destruct (Ty CT$wmAdd_Int,
          Dcon Lcall_$wmAdd_Int1) : (lizzieLet22_1Lcall_$wmAdd_Int1,CT$wmAdd_Int) > [(es_3_1_destruct,Pointer_QTree_Int),
                                                                                     (es_4_1_destruct,Pointer_QTree_Int),
                                                                                     (sc_0_5_destruct,Pointer_CT$wmAdd_Int),
                                                                                     (wsie_4_destruct,MyDTInt_Int_Int),
                                                                                     (q1a8h_3_destruct,Pointer_QTree_Int),
                                                                                     (t1a8m_3_destruct,Pointer_QTree_Int)] */
  logic [5:0] lizzieLet22_1Lcall_$wmAdd_Int1_emitted;
  logic [5:0] lizzieLet22_1Lcall_$wmAdd_Int1_done;
  assign es_3_1_destruct_d = {lizzieLet22_1Lcall_$wmAdd_Int1_d[19:4],
                              (lizzieLet22_1Lcall_$wmAdd_Int1_d[0] && (! lizzieLet22_1Lcall_$wmAdd_Int1_emitted[0]))};
  assign es_4_1_destruct_d = {lizzieLet22_1Lcall_$wmAdd_Int1_d[35:20],
                              (lizzieLet22_1Lcall_$wmAdd_Int1_d[0] && (! lizzieLet22_1Lcall_$wmAdd_Int1_emitted[1]))};
  assign sc_0_5_destruct_d = {lizzieLet22_1Lcall_$wmAdd_Int1_d[51:36],
                              (lizzieLet22_1Lcall_$wmAdd_Int1_d[0] && (! lizzieLet22_1Lcall_$wmAdd_Int1_emitted[2]))};
  assign wsie_4_destruct_d = (lizzieLet22_1Lcall_$wmAdd_Int1_d[0] && (! lizzieLet22_1Lcall_$wmAdd_Int1_emitted[3]));
  assign q1a8h_3_destruct_d = {lizzieLet22_1Lcall_$wmAdd_Int1_d[67:52],
                               (lizzieLet22_1Lcall_$wmAdd_Int1_d[0] && (! lizzieLet22_1Lcall_$wmAdd_Int1_emitted[4]))};
  assign t1a8m_3_destruct_d = {lizzieLet22_1Lcall_$wmAdd_Int1_d[83:68],
                               (lizzieLet22_1Lcall_$wmAdd_Int1_d[0] && (! lizzieLet22_1Lcall_$wmAdd_Int1_emitted[5]))};
  assign lizzieLet22_1Lcall_$wmAdd_Int1_done = (lizzieLet22_1Lcall_$wmAdd_Int1_emitted | ({t1a8m_3_destruct_d[0],
                                                                                           q1a8h_3_destruct_d[0],
                                                                                           wsie_4_destruct_d[0],
                                                                                           sc_0_5_destruct_d[0],
                                                                                           es_4_1_destruct_d[0],
                                                                                           es_3_1_destruct_d[0]} & {t1a8m_3_destruct_r,
                                                                                                                    q1a8h_3_destruct_r,
                                                                                                                    wsie_4_destruct_r,
                                                                                                                    sc_0_5_destruct_r,
                                                                                                                    es_4_1_destruct_r,
                                                                                                                    es_3_1_destruct_r}));
  assign lizzieLet22_1Lcall_$wmAdd_Int1_r = (& lizzieLet22_1Lcall_$wmAdd_Int1_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet22_1Lcall_$wmAdd_Int1_emitted <= 6'd0;
    else
      lizzieLet22_1Lcall_$wmAdd_Int1_emitted <= (lizzieLet22_1Lcall_$wmAdd_Int1_r ? 6'd0 :
                                                 lizzieLet22_1Lcall_$wmAdd_Int1_done);
  
  /* destruct (Ty CT$wmAdd_Int,
          Dcon Lcall_$wmAdd_Int2) : (lizzieLet22_1Lcall_$wmAdd_Int2,CT$wmAdd_Int) > [(es_4_destruct,Pointer_QTree_Int),
                                                                                     (sc_0_4_destruct,Pointer_CT$wmAdd_Int),
                                                                                     (wsie_3_destruct,MyDTInt_Int_Int),
                                                                                     (q1a8h_2_destruct,Pointer_QTree_Int),
                                                                                     (t1a8m_2_destruct,Pointer_QTree_Int),
                                                                                     (q2a8i_2_destruct,Pointer_QTree_Int),
                                                                                     (t2a8n_2_destruct,Pointer_QTree_Int)] */
  logic [6:0] lizzieLet22_1Lcall_$wmAdd_Int2_emitted;
  logic [6:0] lizzieLet22_1Lcall_$wmAdd_Int2_done;
  assign es_4_destruct_d = {lizzieLet22_1Lcall_$wmAdd_Int2_d[19:4],
                            (lizzieLet22_1Lcall_$wmAdd_Int2_d[0] && (! lizzieLet22_1Lcall_$wmAdd_Int2_emitted[0]))};
  assign sc_0_4_destruct_d = {lizzieLet22_1Lcall_$wmAdd_Int2_d[35:20],
                              (lizzieLet22_1Lcall_$wmAdd_Int2_d[0] && (! lizzieLet22_1Lcall_$wmAdd_Int2_emitted[1]))};
  assign wsie_3_destruct_d = (lizzieLet22_1Lcall_$wmAdd_Int2_d[0] && (! lizzieLet22_1Lcall_$wmAdd_Int2_emitted[2]));
  assign q1a8h_2_destruct_d = {lizzieLet22_1Lcall_$wmAdd_Int2_d[51:36],
                               (lizzieLet22_1Lcall_$wmAdd_Int2_d[0] && (! lizzieLet22_1Lcall_$wmAdd_Int2_emitted[3]))};
  assign t1a8m_2_destruct_d = {lizzieLet22_1Lcall_$wmAdd_Int2_d[67:52],
                               (lizzieLet22_1Lcall_$wmAdd_Int2_d[0] && (! lizzieLet22_1Lcall_$wmAdd_Int2_emitted[4]))};
  assign q2a8i_2_destruct_d = {lizzieLet22_1Lcall_$wmAdd_Int2_d[83:68],
                               (lizzieLet22_1Lcall_$wmAdd_Int2_d[0] && (! lizzieLet22_1Lcall_$wmAdd_Int2_emitted[5]))};
  assign t2a8n_2_destruct_d = {lizzieLet22_1Lcall_$wmAdd_Int2_d[99:84],
                               (lizzieLet22_1Lcall_$wmAdd_Int2_d[0] && (! lizzieLet22_1Lcall_$wmAdd_Int2_emitted[6]))};
  assign lizzieLet22_1Lcall_$wmAdd_Int2_done = (lizzieLet22_1Lcall_$wmAdd_Int2_emitted | ({t2a8n_2_destruct_d[0],
                                                                                           q2a8i_2_destruct_d[0],
                                                                                           t1a8m_2_destruct_d[0],
                                                                                           q1a8h_2_destruct_d[0],
                                                                                           wsie_3_destruct_d[0],
                                                                                           sc_0_4_destruct_d[0],
                                                                                           es_4_destruct_d[0]} & {t2a8n_2_destruct_r,
                                                                                                                  q2a8i_2_destruct_r,
                                                                                                                  t1a8m_2_destruct_r,
                                                                                                                  q1a8h_2_destruct_r,
                                                                                                                  wsie_3_destruct_r,
                                                                                                                  sc_0_4_destruct_r,
                                                                                                                  es_4_destruct_r}));
  assign lizzieLet22_1Lcall_$wmAdd_Int2_r = (& lizzieLet22_1Lcall_$wmAdd_Int2_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet22_1Lcall_$wmAdd_Int2_emitted <= 7'd0;
    else
      lizzieLet22_1Lcall_$wmAdd_Int2_emitted <= (lizzieLet22_1Lcall_$wmAdd_Int2_r ? 7'd0 :
                                                 lizzieLet22_1Lcall_$wmAdd_Int2_done);
  
  /* destruct (Ty CT$wmAdd_Int,
          Dcon Lcall_$wmAdd_Int3) : (lizzieLet22_1Lcall_$wmAdd_Int3,CT$wmAdd_Int) > [(sc_0_3_destruct,Pointer_CT$wmAdd_Int),
                                                                                     (wsie_2_destruct,MyDTInt_Int_Int),
                                                                                     (q1a8h_1_destruct,Pointer_QTree_Int),
                                                                                     (t1a8m_1_destruct,Pointer_QTree_Int),
                                                                                     (q2a8i_1_destruct,Pointer_QTree_Int),
                                                                                     (t2a8n_1_destruct,Pointer_QTree_Int),
                                                                                     (q3a8j_1_destruct,Pointer_QTree_Int),
                                                                                     (t3a8o_1_destruct,Pointer_QTree_Int)] */
  logic [7:0] lizzieLet22_1Lcall_$wmAdd_Int3_emitted;
  logic [7:0] lizzieLet22_1Lcall_$wmAdd_Int3_done;
  assign sc_0_3_destruct_d = {lizzieLet22_1Lcall_$wmAdd_Int3_d[19:4],
                              (lizzieLet22_1Lcall_$wmAdd_Int3_d[0] && (! lizzieLet22_1Lcall_$wmAdd_Int3_emitted[0]))};
  assign wsie_2_destruct_d = (lizzieLet22_1Lcall_$wmAdd_Int3_d[0] && (! lizzieLet22_1Lcall_$wmAdd_Int3_emitted[1]));
  assign q1a8h_1_destruct_d = {lizzieLet22_1Lcall_$wmAdd_Int3_d[35:20],
                               (lizzieLet22_1Lcall_$wmAdd_Int3_d[0] && (! lizzieLet22_1Lcall_$wmAdd_Int3_emitted[2]))};
  assign t1a8m_1_destruct_d = {lizzieLet22_1Lcall_$wmAdd_Int3_d[51:36],
                               (lizzieLet22_1Lcall_$wmAdd_Int3_d[0] && (! lizzieLet22_1Lcall_$wmAdd_Int3_emitted[3]))};
  assign q2a8i_1_destruct_d = {lizzieLet22_1Lcall_$wmAdd_Int3_d[67:52],
                               (lizzieLet22_1Lcall_$wmAdd_Int3_d[0] && (! lizzieLet22_1Lcall_$wmAdd_Int3_emitted[4]))};
  assign t2a8n_1_destruct_d = {lizzieLet22_1Lcall_$wmAdd_Int3_d[83:68],
                               (lizzieLet22_1Lcall_$wmAdd_Int3_d[0] && (! lizzieLet22_1Lcall_$wmAdd_Int3_emitted[5]))};
  assign q3a8j_1_destruct_d = {lizzieLet22_1Lcall_$wmAdd_Int3_d[99:84],
                               (lizzieLet22_1Lcall_$wmAdd_Int3_d[0] && (! lizzieLet22_1Lcall_$wmAdd_Int3_emitted[6]))};
  assign t3a8o_1_destruct_d = {lizzieLet22_1Lcall_$wmAdd_Int3_d[115:100],
                               (lizzieLet22_1Lcall_$wmAdd_Int3_d[0] && (! lizzieLet22_1Lcall_$wmAdd_Int3_emitted[7]))};
  assign lizzieLet22_1Lcall_$wmAdd_Int3_done = (lizzieLet22_1Lcall_$wmAdd_Int3_emitted | ({t3a8o_1_destruct_d[0],
                                                                                           q3a8j_1_destruct_d[0],
                                                                                           t2a8n_1_destruct_d[0],
                                                                                           q2a8i_1_destruct_d[0],
                                                                                           t1a8m_1_destruct_d[0],
                                                                                           q1a8h_1_destruct_d[0],
                                                                                           wsie_2_destruct_d[0],
                                                                                           sc_0_3_destruct_d[0]} & {t3a8o_1_destruct_r,
                                                                                                                    q3a8j_1_destruct_r,
                                                                                                                    t2a8n_1_destruct_r,
                                                                                                                    q2a8i_1_destruct_r,
                                                                                                                    t1a8m_1_destruct_r,
                                                                                                                    q1a8h_1_destruct_r,
                                                                                                                    wsie_2_destruct_r,
                                                                                                                    sc_0_3_destruct_r}));
  assign lizzieLet22_1Lcall_$wmAdd_Int3_r = (& lizzieLet22_1Lcall_$wmAdd_Int3_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet22_1Lcall_$wmAdd_Int3_emitted <= 8'd0;
    else
      lizzieLet22_1Lcall_$wmAdd_Int3_emitted <= (lizzieLet22_1Lcall_$wmAdd_Int3_r ? 8'd0 :
                                                 lizzieLet22_1Lcall_$wmAdd_Int3_done);
  
  /* demux (Ty CT$wmAdd_Int,
       Ty CT$wmAdd_Int) : (lizzieLet22_2,CT$wmAdd_Int) (lizzieLet22_1,CT$wmAdd_Int) > [(_49,CT$wmAdd_Int),
                                                                                       (lizzieLet22_1Lcall_$wmAdd_Int3,CT$wmAdd_Int),
                                                                                       (lizzieLet22_1Lcall_$wmAdd_Int2,CT$wmAdd_Int),
                                                                                       (lizzieLet22_1Lcall_$wmAdd_Int1,CT$wmAdd_Int),
                                                                                       (lizzieLet22_1Lcall_$wmAdd_Int0,CT$wmAdd_Int)] */
  logic [4:0] lizzieLet22_1_onehotd;
  always_comb
    if ((lizzieLet22_2_d[0] && lizzieLet22_1_d[0]))
      unique case (lizzieLet22_2_d[3:1])
        3'd0: lizzieLet22_1_onehotd = 5'd1;
        3'd1: lizzieLet22_1_onehotd = 5'd2;
        3'd2: lizzieLet22_1_onehotd = 5'd4;
        3'd3: lizzieLet22_1_onehotd = 5'd8;
        3'd4: lizzieLet22_1_onehotd = 5'd16;
        default: lizzieLet22_1_onehotd = 5'd0;
      endcase
    else lizzieLet22_1_onehotd = 5'd0;
  assign _49_d = {lizzieLet22_1_d[115:1], lizzieLet22_1_onehotd[0]};
  assign lizzieLet22_1Lcall_$wmAdd_Int3_d = {lizzieLet22_1_d[115:1],
                                             lizzieLet22_1_onehotd[1]};
  assign lizzieLet22_1Lcall_$wmAdd_Int2_d = {lizzieLet22_1_d[115:1],
                                             lizzieLet22_1_onehotd[2]};
  assign lizzieLet22_1Lcall_$wmAdd_Int1_d = {lizzieLet22_1_d[115:1],
                                             lizzieLet22_1_onehotd[3]};
  assign lizzieLet22_1Lcall_$wmAdd_Int0_d = {lizzieLet22_1_d[115:1],
                                             lizzieLet22_1_onehotd[4]};
  assign lizzieLet22_1_r = (| (lizzieLet22_1_onehotd & {lizzieLet22_1Lcall_$wmAdd_Int0_r,
                                                        lizzieLet22_1Lcall_$wmAdd_Int1_r,
                                                        lizzieLet22_1Lcall_$wmAdd_Int2_r,
                                                        lizzieLet22_1Lcall_$wmAdd_Int3_r,
                                                        _49_r}));
  assign lizzieLet22_2_r = lizzieLet22_1_r;
  
  /* demux (Ty CT$wmAdd_Int,
       Ty Go) : (lizzieLet22_3,CT$wmAdd_Int) (go_10_goMux_data,Go) > [(_48,Go),
                                                                      (lizzieLet22_3Lcall_$wmAdd_Int3,Go),
                                                                      (lizzieLet22_3Lcall_$wmAdd_Int2,Go),
                                                                      (lizzieLet22_3Lcall_$wmAdd_Int1,Go),
                                                                      (lizzieLet22_3Lcall_$wmAdd_Int0,Go)] */
  logic [4:0] go_10_goMux_data_onehotd;
  always_comb
    if ((lizzieLet22_3_d[0] && go_10_goMux_data_d[0]))
      unique case (lizzieLet22_3_d[3:1])
        3'd0: go_10_goMux_data_onehotd = 5'd1;
        3'd1: go_10_goMux_data_onehotd = 5'd2;
        3'd2: go_10_goMux_data_onehotd = 5'd4;
        3'd3: go_10_goMux_data_onehotd = 5'd8;
        3'd4: go_10_goMux_data_onehotd = 5'd16;
        default: go_10_goMux_data_onehotd = 5'd0;
      endcase
    else go_10_goMux_data_onehotd = 5'd0;
  assign _48_d = go_10_goMux_data_onehotd[0];
  assign lizzieLet22_3Lcall_$wmAdd_Int3_d = go_10_goMux_data_onehotd[1];
  assign lizzieLet22_3Lcall_$wmAdd_Int2_d = go_10_goMux_data_onehotd[2];
  assign lizzieLet22_3Lcall_$wmAdd_Int1_d = go_10_goMux_data_onehotd[3];
  assign lizzieLet22_3Lcall_$wmAdd_Int0_d = go_10_goMux_data_onehotd[4];
  assign go_10_goMux_data_r = (| (go_10_goMux_data_onehotd & {lizzieLet22_3Lcall_$wmAdd_Int0_r,
                                                              lizzieLet22_3Lcall_$wmAdd_Int1_r,
                                                              lizzieLet22_3Lcall_$wmAdd_Int2_r,
                                                              lizzieLet22_3Lcall_$wmAdd_Int3_r,
                                                              _48_r}));
  assign lizzieLet22_3_r = go_10_goMux_data_r;
  
  /* buf (Ty Go) : (lizzieLet22_3Lcall_$wmAdd_Int0,Go) > (lizzieLet22_3Lcall_$wmAdd_Int0_1_argbuf,Go) */
  Go_t lizzieLet22_3Lcall_$wmAdd_Int0_bufchan_d;
  logic lizzieLet22_3Lcall_$wmAdd_Int0_bufchan_r;
  assign lizzieLet22_3Lcall_$wmAdd_Int0_r = ((! lizzieLet22_3Lcall_$wmAdd_Int0_bufchan_d[0]) || lizzieLet22_3Lcall_$wmAdd_Int0_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet22_3Lcall_$wmAdd_Int0_bufchan_d <= 1'd0;
    else
      if (lizzieLet22_3Lcall_$wmAdd_Int0_r)
        lizzieLet22_3Lcall_$wmAdd_Int0_bufchan_d <= lizzieLet22_3Lcall_$wmAdd_Int0_d;
  Go_t lizzieLet22_3Lcall_$wmAdd_Int0_bufchan_buf;
  assign lizzieLet22_3Lcall_$wmAdd_Int0_bufchan_r = (! lizzieLet22_3Lcall_$wmAdd_Int0_bufchan_buf[0]);
  assign lizzieLet22_3Lcall_$wmAdd_Int0_1_argbuf_d = (lizzieLet22_3Lcall_$wmAdd_Int0_bufchan_buf[0] ? lizzieLet22_3Lcall_$wmAdd_Int0_bufchan_buf :
                                                      lizzieLet22_3Lcall_$wmAdd_Int0_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet22_3Lcall_$wmAdd_Int0_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet22_3Lcall_$wmAdd_Int0_1_argbuf_r && lizzieLet22_3Lcall_$wmAdd_Int0_bufchan_buf[0]))
        lizzieLet22_3Lcall_$wmAdd_Int0_bufchan_buf <= 1'd0;
      else if (((! lizzieLet22_3Lcall_$wmAdd_Int0_1_argbuf_r) && (! lizzieLet22_3Lcall_$wmAdd_Int0_bufchan_buf[0])))
        lizzieLet22_3Lcall_$wmAdd_Int0_bufchan_buf <= lizzieLet22_3Lcall_$wmAdd_Int0_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet22_3Lcall_$wmAdd_Int1,Go) > (lizzieLet22_3Lcall_$wmAdd_Int1_1_argbuf,Go) */
  Go_t lizzieLet22_3Lcall_$wmAdd_Int1_bufchan_d;
  logic lizzieLet22_3Lcall_$wmAdd_Int1_bufchan_r;
  assign lizzieLet22_3Lcall_$wmAdd_Int1_r = ((! lizzieLet22_3Lcall_$wmAdd_Int1_bufchan_d[0]) || lizzieLet22_3Lcall_$wmAdd_Int1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet22_3Lcall_$wmAdd_Int1_bufchan_d <= 1'd0;
    else
      if (lizzieLet22_3Lcall_$wmAdd_Int1_r)
        lizzieLet22_3Lcall_$wmAdd_Int1_bufchan_d <= lizzieLet22_3Lcall_$wmAdd_Int1_d;
  Go_t lizzieLet22_3Lcall_$wmAdd_Int1_bufchan_buf;
  assign lizzieLet22_3Lcall_$wmAdd_Int1_bufchan_r = (! lizzieLet22_3Lcall_$wmAdd_Int1_bufchan_buf[0]);
  assign lizzieLet22_3Lcall_$wmAdd_Int1_1_argbuf_d = (lizzieLet22_3Lcall_$wmAdd_Int1_bufchan_buf[0] ? lizzieLet22_3Lcall_$wmAdd_Int1_bufchan_buf :
                                                      lizzieLet22_3Lcall_$wmAdd_Int1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet22_3Lcall_$wmAdd_Int1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet22_3Lcall_$wmAdd_Int1_1_argbuf_r && lizzieLet22_3Lcall_$wmAdd_Int1_bufchan_buf[0]))
        lizzieLet22_3Lcall_$wmAdd_Int1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet22_3Lcall_$wmAdd_Int1_1_argbuf_r) && (! lizzieLet22_3Lcall_$wmAdd_Int1_bufchan_buf[0])))
        lizzieLet22_3Lcall_$wmAdd_Int1_bufchan_buf <= lizzieLet22_3Lcall_$wmAdd_Int1_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet22_3Lcall_$wmAdd_Int2,Go) > (lizzieLet22_3Lcall_$wmAdd_Int2_1_argbuf,Go) */
  Go_t lizzieLet22_3Lcall_$wmAdd_Int2_bufchan_d;
  logic lizzieLet22_3Lcall_$wmAdd_Int2_bufchan_r;
  assign lizzieLet22_3Lcall_$wmAdd_Int2_r = ((! lizzieLet22_3Lcall_$wmAdd_Int2_bufchan_d[0]) || lizzieLet22_3Lcall_$wmAdd_Int2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet22_3Lcall_$wmAdd_Int2_bufchan_d <= 1'd0;
    else
      if (lizzieLet22_3Lcall_$wmAdd_Int2_r)
        lizzieLet22_3Lcall_$wmAdd_Int2_bufchan_d <= lizzieLet22_3Lcall_$wmAdd_Int2_d;
  Go_t lizzieLet22_3Lcall_$wmAdd_Int2_bufchan_buf;
  assign lizzieLet22_3Lcall_$wmAdd_Int2_bufchan_r = (! lizzieLet22_3Lcall_$wmAdd_Int2_bufchan_buf[0]);
  assign lizzieLet22_3Lcall_$wmAdd_Int2_1_argbuf_d = (lizzieLet22_3Lcall_$wmAdd_Int2_bufchan_buf[0] ? lizzieLet22_3Lcall_$wmAdd_Int2_bufchan_buf :
                                                      lizzieLet22_3Lcall_$wmAdd_Int2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet22_3Lcall_$wmAdd_Int2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet22_3Lcall_$wmAdd_Int2_1_argbuf_r && lizzieLet22_3Lcall_$wmAdd_Int2_bufchan_buf[0]))
        lizzieLet22_3Lcall_$wmAdd_Int2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet22_3Lcall_$wmAdd_Int2_1_argbuf_r) && (! lizzieLet22_3Lcall_$wmAdd_Int2_bufchan_buf[0])))
        lizzieLet22_3Lcall_$wmAdd_Int2_bufchan_buf <= lizzieLet22_3Lcall_$wmAdd_Int2_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet22_3Lcall_$wmAdd_Int3,Go) > (lizzieLet22_3Lcall_$wmAdd_Int3_1_argbuf,Go) */
  Go_t lizzieLet22_3Lcall_$wmAdd_Int3_bufchan_d;
  logic lizzieLet22_3Lcall_$wmAdd_Int3_bufchan_r;
  assign lizzieLet22_3Lcall_$wmAdd_Int3_r = ((! lizzieLet22_3Lcall_$wmAdd_Int3_bufchan_d[0]) || lizzieLet22_3Lcall_$wmAdd_Int3_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet22_3Lcall_$wmAdd_Int3_bufchan_d <= 1'd0;
    else
      if (lizzieLet22_3Lcall_$wmAdd_Int3_r)
        lizzieLet22_3Lcall_$wmAdd_Int3_bufchan_d <= lizzieLet22_3Lcall_$wmAdd_Int3_d;
  Go_t lizzieLet22_3Lcall_$wmAdd_Int3_bufchan_buf;
  assign lizzieLet22_3Lcall_$wmAdd_Int3_bufchan_r = (! lizzieLet22_3Lcall_$wmAdd_Int3_bufchan_buf[0]);
  assign lizzieLet22_3Lcall_$wmAdd_Int3_1_argbuf_d = (lizzieLet22_3Lcall_$wmAdd_Int3_bufchan_buf[0] ? lizzieLet22_3Lcall_$wmAdd_Int3_bufchan_buf :
                                                      lizzieLet22_3Lcall_$wmAdd_Int3_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet22_3Lcall_$wmAdd_Int3_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet22_3Lcall_$wmAdd_Int3_1_argbuf_r && lizzieLet22_3Lcall_$wmAdd_Int3_bufchan_buf[0]))
        lizzieLet22_3Lcall_$wmAdd_Int3_bufchan_buf <= 1'd0;
      else if (((! lizzieLet22_3Lcall_$wmAdd_Int3_1_argbuf_r) && (! lizzieLet22_3Lcall_$wmAdd_Int3_bufchan_buf[0])))
        lizzieLet22_3Lcall_$wmAdd_Int3_bufchan_buf <= lizzieLet22_3Lcall_$wmAdd_Int3_bufchan_d;
  
  /* demux (Ty CT$wmAdd_Int,
       Ty Pointer_QTree_Int) : (lizzieLet22_4,CT$wmAdd_Int) (srtarg_0_goMux_mux,Pointer_QTree_Int) > [(lizzieLet22_4L$wmAdd_Intsbos,Pointer_QTree_Int),
                                                                                                      (lizzieLet22_4Lcall_$wmAdd_Int3,Pointer_QTree_Int),
                                                                                                      (lizzieLet22_4Lcall_$wmAdd_Int2,Pointer_QTree_Int),
                                                                                                      (lizzieLet22_4Lcall_$wmAdd_Int1,Pointer_QTree_Int),
                                                                                                      (lizzieLet22_4Lcall_$wmAdd_Int0,Pointer_QTree_Int)] */
  logic [4:0] srtarg_0_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet22_4_d[0] && srtarg_0_goMux_mux_d[0]))
      unique case (lizzieLet22_4_d[3:1])
        3'd0: srtarg_0_goMux_mux_onehotd = 5'd1;
        3'd1: srtarg_0_goMux_mux_onehotd = 5'd2;
        3'd2: srtarg_0_goMux_mux_onehotd = 5'd4;
        3'd3: srtarg_0_goMux_mux_onehotd = 5'd8;
        3'd4: srtarg_0_goMux_mux_onehotd = 5'd16;
        default: srtarg_0_goMux_mux_onehotd = 5'd0;
      endcase
    else srtarg_0_goMux_mux_onehotd = 5'd0;
  assign lizzieLet22_4L$wmAdd_Intsbos_d = {srtarg_0_goMux_mux_d[16:1],
                                           srtarg_0_goMux_mux_onehotd[0]};
  assign lizzieLet22_4Lcall_$wmAdd_Int3_d = {srtarg_0_goMux_mux_d[16:1],
                                             srtarg_0_goMux_mux_onehotd[1]};
  assign lizzieLet22_4Lcall_$wmAdd_Int2_d = {srtarg_0_goMux_mux_d[16:1],
                                             srtarg_0_goMux_mux_onehotd[2]};
  assign lizzieLet22_4Lcall_$wmAdd_Int1_d = {srtarg_0_goMux_mux_d[16:1],
                                             srtarg_0_goMux_mux_onehotd[3]};
  assign lizzieLet22_4Lcall_$wmAdd_Int0_d = {srtarg_0_goMux_mux_d[16:1],
                                             srtarg_0_goMux_mux_onehotd[4]};
  assign srtarg_0_goMux_mux_r = (| (srtarg_0_goMux_mux_onehotd & {lizzieLet22_4Lcall_$wmAdd_Int0_r,
                                                                  lizzieLet22_4Lcall_$wmAdd_Int1_r,
                                                                  lizzieLet22_4Lcall_$wmAdd_Int2_r,
                                                                  lizzieLet22_4Lcall_$wmAdd_Int3_r,
                                                                  lizzieLet22_4L$wmAdd_Intsbos_r}));
  assign lizzieLet22_4_r = srtarg_0_goMux_mux_r;
  
  /* fork (Ty Pointer_QTree_Int) : (lizzieLet22_4L$wmAdd_Intsbos,Pointer_QTree_Int) > [(lizzieLet22_4L$wmAdd_Intsbos_1_merge_merge_fork_1,Pointer_QTree_Int),
                                                                                  (lizzieLet22_4L$wmAdd_Intsbos_1_merge_merge_fork_2,Pointer_QTree_Int)] */
  logic [1:0] lizzieLet22_4L$wmAdd_Intsbos_emitted;
  logic [1:0] lizzieLet22_4L$wmAdd_Intsbos_done;
  assign lizzieLet22_4L$wmAdd_Intsbos_1_merge_merge_fork_1_d = {lizzieLet22_4L$wmAdd_Intsbos_d[16:1],
                                                                (lizzieLet22_4L$wmAdd_Intsbos_d[0] && (! lizzieLet22_4L$wmAdd_Intsbos_emitted[0]))};
  assign lizzieLet22_4L$wmAdd_Intsbos_1_merge_merge_fork_2_d = {lizzieLet22_4L$wmAdd_Intsbos_d[16:1],
                                                                (lizzieLet22_4L$wmAdd_Intsbos_d[0] && (! lizzieLet22_4L$wmAdd_Intsbos_emitted[1]))};
  assign lizzieLet22_4L$wmAdd_Intsbos_done = (lizzieLet22_4L$wmAdd_Intsbos_emitted | ({lizzieLet22_4L$wmAdd_Intsbos_1_merge_merge_fork_2_d[0],
                                                                                       lizzieLet22_4L$wmAdd_Intsbos_1_merge_merge_fork_1_d[0]} & {lizzieLet22_4L$wmAdd_Intsbos_1_merge_merge_fork_2_r,
                                                                                                                                                  lizzieLet22_4L$wmAdd_Intsbos_1_merge_merge_fork_1_r}));
  assign lizzieLet22_4L$wmAdd_Intsbos_r = (& lizzieLet22_4L$wmAdd_Intsbos_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet22_4L$wmAdd_Intsbos_emitted <= 2'd0;
    else
      lizzieLet22_4L$wmAdd_Intsbos_emitted <= (lizzieLet22_4L$wmAdd_Intsbos_r ? 2'd0 :
                                               lizzieLet22_4L$wmAdd_Intsbos_done);
  
  /* togo (Ty Pointer_QTree_Int) : (lizzieLet22_4L$wmAdd_Intsbos_1_merge_merge_fork_1,Pointer_QTree_Int) > (call_$wmAdd_Int_goConst,Go) */
  assign call_$wmAdd_Int_goConst_d = lizzieLet22_4L$wmAdd_Intsbos_1_merge_merge_fork_1_d[0];
  assign lizzieLet22_4L$wmAdd_Intsbos_1_merge_merge_fork_1_r = call_$wmAdd_Int_goConst_r;
  
  /* buf (Ty Pointer_QTree_Int) : (lizzieLet22_4L$wmAdd_Intsbos_1_merge_merge_fork_2,Pointer_QTree_Int) > ($wmAdd_Int_resbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t lizzieLet22_4L$wmAdd_Intsbos_1_merge_merge_fork_2_bufchan_d;
  logic lizzieLet22_4L$wmAdd_Intsbos_1_merge_merge_fork_2_bufchan_r;
  assign lizzieLet22_4L$wmAdd_Intsbos_1_merge_merge_fork_2_r = ((! lizzieLet22_4L$wmAdd_Intsbos_1_merge_merge_fork_2_bufchan_d[0]) || lizzieLet22_4L$wmAdd_Intsbos_1_merge_merge_fork_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet22_4L$wmAdd_Intsbos_1_merge_merge_fork_2_bufchan_d <= {16'd0,
                                                                      1'd0};
    else
      if (lizzieLet22_4L$wmAdd_Intsbos_1_merge_merge_fork_2_r)
        lizzieLet22_4L$wmAdd_Intsbos_1_merge_merge_fork_2_bufchan_d <= lizzieLet22_4L$wmAdd_Intsbos_1_merge_merge_fork_2_d;
  Pointer_QTree_Int_t lizzieLet22_4L$wmAdd_Intsbos_1_merge_merge_fork_2_bufchan_buf;
  assign lizzieLet22_4L$wmAdd_Intsbos_1_merge_merge_fork_2_bufchan_r = (! lizzieLet22_4L$wmAdd_Intsbos_1_merge_merge_fork_2_bufchan_buf[0]);
  assign \$wmAdd_Int_resbuf_d  = (lizzieLet22_4L$wmAdd_Intsbos_1_merge_merge_fork_2_bufchan_buf[0] ? lizzieLet22_4L$wmAdd_Intsbos_1_merge_merge_fork_2_bufchan_buf :
                                  lizzieLet22_4L$wmAdd_Intsbos_1_merge_merge_fork_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet22_4L$wmAdd_Intsbos_1_merge_merge_fork_2_bufchan_buf <= {16'd0,
                                                                        1'd0};
    else
      if ((\$wmAdd_Int_resbuf_r  && lizzieLet22_4L$wmAdd_Intsbos_1_merge_merge_fork_2_bufchan_buf[0]))
        lizzieLet22_4L$wmAdd_Intsbos_1_merge_merge_fork_2_bufchan_buf <= {16'd0,
                                                                          1'd0};
      else if (((! \$wmAdd_Int_resbuf_r ) && (! lizzieLet22_4L$wmAdd_Intsbos_1_merge_merge_fork_2_bufchan_buf[0])))
        lizzieLet22_4L$wmAdd_Intsbos_1_merge_merge_fork_2_bufchan_buf <= lizzieLet22_4L$wmAdd_Intsbos_1_merge_merge_fork_2_bufchan_d;
  
  /* dcon (Ty QTree_Int,
      Dcon QNode_Int) : [(lizzieLet22_4Lcall_$wmAdd_Int0,Pointer_QTree_Int),
                         (es_2_destruct,Pointer_QTree_Int),
                         (es_3_2_destruct,Pointer_QTree_Int),
                         (es_4_2_destruct,Pointer_QTree_Int)] > (lizzieLet22_4Lcall_$wmAdd_Int0_1es_2_1es_3_2_1es_4_2_1QNode_Int,QTree_Int) */
  assign lizzieLet22_4Lcall_$wmAdd_Int0_1es_2_1es_3_2_1es_4_2_1QNode_Int_d = QNode_Int_dc((& {lizzieLet22_4Lcall_$wmAdd_Int0_d[0],
                                                                                              es_2_destruct_d[0],
                                                                                              es_3_2_destruct_d[0],
                                                                                              es_4_2_destruct_d[0]}), lizzieLet22_4Lcall_$wmAdd_Int0_d, es_2_destruct_d, es_3_2_destruct_d, es_4_2_destruct_d);
  assign {lizzieLet22_4Lcall_$wmAdd_Int0_r,
          es_2_destruct_r,
          es_3_2_destruct_r,
          es_4_2_destruct_r} = {4 {(lizzieLet22_4Lcall_$wmAdd_Int0_1es_2_1es_3_2_1es_4_2_1QNode_Int_r && lizzieLet22_4Lcall_$wmAdd_Int0_1es_2_1es_3_2_1es_4_2_1QNode_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (lizzieLet22_4Lcall_$wmAdd_Int0_1es_2_1es_3_2_1es_4_2_1QNode_Int,QTree_Int) > (lizzieLet26_1_argbuf,QTree_Int) */
  QTree_Int_t lizzieLet22_4Lcall_$wmAdd_Int0_1es_2_1es_3_2_1es_4_2_1QNode_Int_bufchan_d;
  logic lizzieLet22_4Lcall_$wmAdd_Int0_1es_2_1es_3_2_1es_4_2_1QNode_Int_bufchan_r;
  assign lizzieLet22_4Lcall_$wmAdd_Int0_1es_2_1es_3_2_1es_4_2_1QNode_Int_r = ((! lizzieLet22_4Lcall_$wmAdd_Int0_1es_2_1es_3_2_1es_4_2_1QNode_Int_bufchan_d[0]) || lizzieLet22_4Lcall_$wmAdd_Int0_1es_2_1es_3_2_1es_4_2_1QNode_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet22_4Lcall_$wmAdd_Int0_1es_2_1es_3_2_1es_4_2_1QNode_Int_bufchan_d <= {66'd0,
                                                                                    1'd0};
    else
      if (lizzieLet22_4Lcall_$wmAdd_Int0_1es_2_1es_3_2_1es_4_2_1QNode_Int_r)
        lizzieLet22_4Lcall_$wmAdd_Int0_1es_2_1es_3_2_1es_4_2_1QNode_Int_bufchan_d <= lizzieLet22_4Lcall_$wmAdd_Int0_1es_2_1es_3_2_1es_4_2_1QNode_Int_d;
  QTree_Int_t lizzieLet22_4Lcall_$wmAdd_Int0_1es_2_1es_3_2_1es_4_2_1QNode_Int_bufchan_buf;
  assign lizzieLet22_4Lcall_$wmAdd_Int0_1es_2_1es_3_2_1es_4_2_1QNode_Int_bufchan_r = (! lizzieLet22_4Lcall_$wmAdd_Int0_1es_2_1es_3_2_1es_4_2_1QNode_Int_bufchan_buf[0]);
  assign lizzieLet26_1_argbuf_d = (lizzieLet22_4Lcall_$wmAdd_Int0_1es_2_1es_3_2_1es_4_2_1QNode_Int_bufchan_buf[0] ? lizzieLet22_4Lcall_$wmAdd_Int0_1es_2_1es_3_2_1es_4_2_1QNode_Int_bufchan_buf :
                                   lizzieLet22_4Lcall_$wmAdd_Int0_1es_2_1es_3_2_1es_4_2_1QNode_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet22_4Lcall_$wmAdd_Int0_1es_2_1es_3_2_1es_4_2_1QNode_Int_bufchan_buf <= {66'd0,
                                                                                      1'd0};
    else
      if ((lizzieLet26_1_argbuf_r && lizzieLet22_4Lcall_$wmAdd_Int0_1es_2_1es_3_2_1es_4_2_1QNode_Int_bufchan_buf[0]))
        lizzieLet22_4Lcall_$wmAdd_Int0_1es_2_1es_3_2_1es_4_2_1QNode_Int_bufchan_buf <= {66'd0,
                                                                                        1'd0};
      else if (((! lizzieLet26_1_argbuf_r) && (! lizzieLet22_4Lcall_$wmAdd_Int0_1es_2_1es_3_2_1es_4_2_1QNode_Int_bufchan_buf[0])))
        lizzieLet22_4Lcall_$wmAdd_Int0_1es_2_1es_3_2_1es_4_2_1QNode_Int_bufchan_buf <= lizzieLet22_4Lcall_$wmAdd_Int0_1es_2_1es_3_2_1es_4_2_1QNode_Int_bufchan_d;
  
  /* dcon (Ty CT$wmAdd_Int,
      Dcon Lcall_$wmAdd_Int0) : [(lizzieLet22_4Lcall_$wmAdd_Int1,Pointer_QTree_Int),
                                 (es_3_1_destruct,Pointer_QTree_Int),
                                 (es_4_1_destruct,Pointer_QTree_Int),
                                 (sc_0_5_destruct,Pointer_CT$wmAdd_Int)] > (lizzieLet22_4Lcall_$wmAdd_Int1_1es_3_1_1es_4_1_1sc_0_5_1Lcall_$wmAdd_Int0,CT$wmAdd_Int) */
  assign lizzieLet22_4Lcall_$wmAdd_Int1_1es_3_1_1es_4_1_1sc_0_5_1Lcall_$wmAdd_Int0_d = Lcall_$wmAdd_Int0_dc((& {lizzieLet22_4Lcall_$wmAdd_Int1_d[0],
                                                                                                                es_3_1_destruct_d[0],
                                                                                                                es_4_1_destruct_d[0],
                                                                                                                sc_0_5_destruct_d[0]}), lizzieLet22_4Lcall_$wmAdd_Int1_d, es_3_1_destruct_d, es_4_1_destruct_d, sc_0_5_destruct_d);
  assign {lizzieLet22_4Lcall_$wmAdd_Int1_r,
          es_3_1_destruct_r,
          es_4_1_destruct_r,
          sc_0_5_destruct_r} = {4 {(lizzieLet22_4Lcall_$wmAdd_Int1_1es_3_1_1es_4_1_1sc_0_5_1Lcall_$wmAdd_Int0_r && lizzieLet22_4Lcall_$wmAdd_Int1_1es_3_1_1es_4_1_1sc_0_5_1Lcall_$wmAdd_Int0_d[0])}};
  
  /* buf (Ty CT$wmAdd_Int) : (lizzieLet22_4Lcall_$wmAdd_Int1_1es_3_1_1es_4_1_1sc_0_5_1Lcall_$wmAdd_Int0,CT$wmAdd_Int) > (lizzieLet25_1_argbuf,CT$wmAdd_Int) */
  CT$wmAdd_Int_t lizzieLet22_4Lcall_$wmAdd_Int1_1es_3_1_1es_4_1_1sc_0_5_1Lcall_$wmAdd_Int0_bufchan_d;
  logic lizzieLet22_4Lcall_$wmAdd_Int1_1es_3_1_1es_4_1_1sc_0_5_1Lcall_$wmAdd_Int0_bufchan_r;
  assign lizzieLet22_4Lcall_$wmAdd_Int1_1es_3_1_1es_4_1_1sc_0_5_1Lcall_$wmAdd_Int0_r = ((! lizzieLet22_4Lcall_$wmAdd_Int1_1es_3_1_1es_4_1_1sc_0_5_1Lcall_$wmAdd_Int0_bufchan_d[0]) || lizzieLet22_4Lcall_$wmAdd_Int1_1es_3_1_1es_4_1_1sc_0_5_1Lcall_$wmAdd_Int0_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet22_4Lcall_$wmAdd_Int1_1es_3_1_1es_4_1_1sc_0_5_1Lcall_$wmAdd_Int0_bufchan_d <= {115'd0,
                                                                                              1'd0};
    else
      if (lizzieLet22_4Lcall_$wmAdd_Int1_1es_3_1_1es_4_1_1sc_0_5_1Lcall_$wmAdd_Int0_r)
        lizzieLet22_4Lcall_$wmAdd_Int1_1es_3_1_1es_4_1_1sc_0_5_1Lcall_$wmAdd_Int0_bufchan_d <= lizzieLet22_4Lcall_$wmAdd_Int1_1es_3_1_1es_4_1_1sc_0_5_1Lcall_$wmAdd_Int0_d;
  CT$wmAdd_Int_t lizzieLet22_4Lcall_$wmAdd_Int1_1es_3_1_1es_4_1_1sc_0_5_1Lcall_$wmAdd_Int0_bufchan_buf;
  assign lizzieLet22_4Lcall_$wmAdd_Int1_1es_3_1_1es_4_1_1sc_0_5_1Lcall_$wmAdd_Int0_bufchan_r = (! lizzieLet22_4Lcall_$wmAdd_Int1_1es_3_1_1es_4_1_1sc_0_5_1Lcall_$wmAdd_Int0_bufchan_buf[0]);
  assign lizzieLet25_1_argbuf_d = (lizzieLet22_4Lcall_$wmAdd_Int1_1es_3_1_1es_4_1_1sc_0_5_1Lcall_$wmAdd_Int0_bufchan_buf[0] ? lizzieLet22_4Lcall_$wmAdd_Int1_1es_3_1_1es_4_1_1sc_0_5_1Lcall_$wmAdd_Int0_bufchan_buf :
                                   lizzieLet22_4Lcall_$wmAdd_Int1_1es_3_1_1es_4_1_1sc_0_5_1Lcall_$wmAdd_Int0_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet22_4Lcall_$wmAdd_Int1_1es_3_1_1es_4_1_1sc_0_5_1Lcall_$wmAdd_Int0_bufchan_buf <= {115'd0,
                                                                                                1'd0};
    else
      if ((lizzieLet25_1_argbuf_r && lizzieLet22_4Lcall_$wmAdd_Int1_1es_3_1_1es_4_1_1sc_0_5_1Lcall_$wmAdd_Int0_bufchan_buf[0]))
        lizzieLet22_4Lcall_$wmAdd_Int1_1es_3_1_1es_4_1_1sc_0_5_1Lcall_$wmAdd_Int0_bufchan_buf <= {115'd0,
                                                                                                  1'd0};
      else if (((! lizzieLet25_1_argbuf_r) && (! lizzieLet22_4Lcall_$wmAdd_Int1_1es_3_1_1es_4_1_1sc_0_5_1Lcall_$wmAdd_Int0_bufchan_buf[0])))
        lizzieLet22_4Lcall_$wmAdd_Int1_1es_3_1_1es_4_1_1sc_0_5_1Lcall_$wmAdd_Int0_bufchan_buf <= lizzieLet22_4Lcall_$wmAdd_Int1_1es_3_1_1es_4_1_1sc_0_5_1Lcall_$wmAdd_Int0_bufchan_d;
  
  /* dcon (Ty CT$wmAdd_Int,
      Dcon Lcall_$wmAdd_Int1) : [(lizzieLet22_4Lcall_$wmAdd_Int2,Pointer_QTree_Int),
                                 (es_4_destruct,Pointer_QTree_Int),
                                 (sc_0_4_destruct,Pointer_CT$wmAdd_Int),
                                 (wsie_3_1,MyDTInt_Int_Int),
                                 (q1a8h_2_destruct,Pointer_QTree_Int),
                                 (t1a8m_2_destruct,Pointer_QTree_Int)] > (lizzieLet22_4Lcall_$wmAdd_Int2_1es_4_1sc_0_4_1wsie_3_1q1a8h_2_1t1a8m_2_1Lcall_$wmAdd_Int1,CT$wmAdd_Int) */
  assign lizzieLet22_4Lcall_$wmAdd_Int2_1es_4_1sc_0_4_1wsie_3_1q1a8h_2_1t1a8m_2_1Lcall_$wmAdd_Int1_d = Lcall_$wmAdd_Int1_dc((& {lizzieLet22_4Lcall_$wmAdd_Int2_d[0],
                                                                                                                                es_4_destruct_d[0],
                                                                                                                                sc_0_4_destruct_d[0],
                                                                                                                                wsie_3_1_d[0],
                                                                                                                                q1a8h_2_destruct_d[0],
                                                                                                                                t1a8m_2_destruct_d[0]}), lizzieLet22_4Lcall_$wmAdd_Int2_d, es_4_destruct_d, sc_0_4_destruct_d, wsie_3_1_d, q1a8h_2_destruct_d, t1a8m_2_destruct_d);
  assign {lizzieLet22_4Lcall_$wmAdd_Int2_r,
          es_4_destruct_r,
          sc_0_4_destruct_r,
          wsie_3_1_r,
          q1a8h_2_destruct_r,
          t1a8m_2_destruct_r} = {6 {(lizzieLet22_4Lcall_$wmAdd_Int2_1es_4_1sc_0_4_1wsie_3_1q1a8h_2_1t1a8m_2_1Lcall_$wmAdd_Int1_r && lizzieLet22_4Lcall_$wmAdd_Int2_1es_4_1sc_0_4_1wsie_3_1q1a8h_2_1t1a8m_2_1Lcall_$wmAdd_Int1_d[0])}};
  
  /* buf (Ty CT$wmAdd_Int) : (lizzieLet22_4Lcall_$wmAdd_Int2_1es_4_1sc_0_4_1wsie_3_1q1a8h_2_1t1a8m_2_1Lcall_$wmAdd_Int1,CT$wmAdd_Int) > (lizzieLet24_1_argbuf,CT$wmAdd_Int) */
  CT$wmAdd_Int_t lizzieLet22_4Lcall_$wmAdd_Int2_1es_4_1sc_0_4_1wsie_3_1q1a8h_2_1t1a8m_2_1Lcall_$wmAdd_Int1_bufchan_d;
  logic lizzieLet22_4Lcall_$wmAdd_Int2_1es_4_1sc_0_4_1wsie_3_1q1a8h_2_1t1a8m_2_1Lcall_$wmAdd_Int1_bufchan_r;
  assign lizzieLet22_4Lcall_$wmAdd_Int2_1es_4_1sc_0_4_1wsie_3_1q1a8h_2_1t1a8m_2_1Lcall_$wmAdd_Int1_r = ((! lizzieLet22_4Lcall_$wmAdd_Int2_1es_4_1sc_0_4_1wsie_3_1q1a8h_2_1t1a8m_2_1Lcall_$wmAdd_Int1_bufchan_d[0]) || lizzieLet22_4Lcall_$wmAdd_Int2_1es_4_1sc_0_4_1wsie_3_1q1a8h_2_1t1a8m_2_1Lcall_$wmAdd_Int1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet22_4Lcall_$wmAdd_Int2_1es_4_1sc_0_4_1wsie_3_1q1a8h_2_1t1a8m_2_1Lcall_$wmAdd_Int1_bufchan_d <= {115'd0,
                                                                                                              1'd0};
    else
      if (lizzieLet22_4Lcall_$wmAdd_Int2_1es_4_1sc_0_4_1wsie_3_1q1a8h_2_1t1a8m_2_1Lcall_$wmAdd_Int1_r)
        lizzieLet22_4Lcall_$wmAdd_Int2_1es_4_1sc_0_4_1wsie_3_1q1a8h_2_1t1a8m_2_1Lcall_$wmAdd_Int1_bufchan_d <= lizzieLet22_4Lcall_$wmAdd_Int2_1es_4_1sc_0_4_1wsie_3_1q1a8h_2_1t1a8m_2_1Lcall_$wmAdd_Int1_d;
  CT$wmAdd_Int_t lizzieLet22_4Lcall_$wmAdd_Int2_1es_4_1sc_0_4_1wsie_3_1q1a8h_2_1t1a8m_2_1Lcall_$wmAdd_Int1_bufchan_buf;
  assign lizzieLet22_4Lcall_$wmAdd_Int2_1es_4_1sc_0_4_1wsie_3_1q1a8h_2_1t1a8m_2_1Lcall_$wmAdd_Int1_bufchan_r = (! lizzieLet22_4Lcall_$wmAdd_Int2_1es_4_1sc_0_4_1wsie_3_1q1a8h_2_1t1a8m_2_1Lcall_$wmAdd_Int1_bufchan_buf[0]);
  assign lizzieLet24_1_argbuf_d = (lizzieLet22_4Lcall_$wmAdd_Int2_1es_4_1sc_0_4_1wsie_3_1q1a8h_2_1t1a8m_2_1Lcall_$wmAdd_Int1_bufchan_buf[0] ? lizzieLet22_4Lcall_$wmAdd_Int2_1es_4_1sc_0_4_1wsie_3_1q1a8h_2_1t1a8m_2_1Lcall_$wmAdd_Int1_bufchan_buf :
                                   lizzieLet22_4Lcall_$wmAdd_Int2_1es_4_1sc_0_4_1wsie_3_1q1a8h_2_1t1a8m_2_1Lcall_$wmAdd_Int1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet22_4Lcall_$wmAdd_Int2_1es_4_1sc_0_4_1wsie_3_1q1a8h_2_1t1a8m_2_1Lcall_$wmAdd_Int1_bufchan_buf <= {115'd0,
                                                                                                                1'd0};
    else
      if ((lizzieLet24_1_argbuf_r && lizzieLet22_4Lcall_$wmAdd_Int2_1es_4_1sc_0_4_1wsie_3_1q1a8h_2_1t1a8m_2_1Lcall_$wmAdd_Int1_bufchan_buf[0]))
        lizzieLet22_4Lcall_$wmAdd_Int2_1es_4_1sc_0_4_1wsie_3_1q1a8h_2_1t1a8m_2_1Lcall_$wmAdd_Int1_bufchan_buf <= {115'd0,
                                                                                                                  1'd0};
      else if (((! lizzieLet24_1_argbuf_r) && (! lizzieLet22_4Lcall_$wmAdd_Int2_1es_4_1sc_0_4_1wsie_3_1q1a8h_2_1t1a8m_2_1Lcall_$wmAdd_Int1_bufchan_buf[0])))
        lizzieLet22_4Lcall_$wmAdd_Int2_1es_4_1sc_0_4_1wsie_3_1q1a8h_2_1t1a8m_2_1Lcall_$wmAdd_Int1_bufchan_buf <= lizzieLet22_4Lcall_$wmAdd_Int2_1es_4_1sc_0_4_1wsie_3_1q1a8h_2_1t1a8m_2_1Lcall_$wmAdd_Int1_bufchan_d;
  
  /* dcon (Ty CT$wmAdd_Int,
      Dcon Lcall_$wmAdd_Int2) : [(lizzieLet22_4Lcall_$wmAdd_Int3,Pointer_QTree_Int),
                                 (sc_0_3_destruct,Pointer_CT$wmAdd_Int),
                                 (wsie_2_1,MyDTInt_Int_Int),
                                 (q1a8h_1_destruct,Pointer_QTree_Int),
                                 (t1a8m_1_destruct,Pointer_QTree_Int),
                                 (q2a8i_1_destruct,Pointer_QTree_Int),
                                 (t2a8n_1_destruct,Pointer_QTree_Int)] > (lizzieLet22_4Lcall_$wmAdd_Int3_1sc_0_3_1wsie_2_1q1a8h_1_1t1a8m_1_1q2a8i_1_1t2a8n_1_1Lcall_$wmAdd_Int2,CT$wmAdd_Int) */
  assign lizzieLet22_4Lcall_$wmAdd_Int3_1sc_0_3_1wsie_2_1q1a8h_1_1t1a8m_1_1q2a8i_1_1t2a8n_1_1Lcall_$wmAdd_Int2_d = Lcall_$wmAdd_Int2_dc((& {lizzieLet22_4Lcall_$wmAdd_Int3_d[0],
                                                                                                                                            sc_0_3_destruct_d[0],
                                                                                                                                            wsie_2_1_d[0],
                                                                                                                                            q1a8h_1_destruct_d[0],
                                                                                                                                            t1a8m_1_destruct_d[0],
                                                                                                                                            q2a8i_1_destruct_d[0],
                                                                                                                                            t2a8n_1_destruct_d[0]}), lizzieLet22_4Lcall_$wmAdd_Int3_d, sc_0_3_destruct_d, wsie_2_1_d, q1a8h_1_destruct_d, t1a8m_1_destruct_d, q2a8i_1_destruct_d, t2a8n_1_destruct_d);
  assign {lizzieLet22_4Lcall_$wmAdd_Int3_r,
          sc_0_3_destruct_r,
          wsie_2_1_r,
          q1a8h_1_destruct_r,
          t1a8m_1_destruct_r,
          q2a8i_1_destruct_r,
          t2a8n_1_destruct_r} = {7 {(lizzieLet22_4Lcall_$wmAdd_Int3_1sc_0_3_1wsie_2_1q1a8h_1_1t1a8m_1_1q2a8i_1_1t2a8n_1_1Lcall_$wmAdd_Int2_r && lizzieLet22_4Lcall_$wmAdd_Int3_1sc_0_3_1wsie_2_1q1a8h_1_1t1a8m_1_1q2a8i_1_1t2a8n_1_1Lcall_$wmAdd_Int2_d[0])}};
  
  /* buf (Ty CT$wmAdd_Int) : (lizzieLet22_4Lcall_$wmAdd_Int3_1sc_0_3_1wsie_2_1q1a8h_1_1t1a8m_1_1q2a8i_1_1t2a8n_1_1Lcall_$wmAdd_Int2,CT$wmAdd_Int) > (lizzieLet23_1_argbuf,CT$wmAdd_Int) */
  CT$wmAdd_Int_t lizzieLet22_4Lcall_$wmAdd_Int3_1sc_0_3_1wsie_2_1q1a8h_1_1t1a8m_1_1q2a8i_1_1t2a8n_1_1Lcall_$wmAdd_Int2_bufchan_d;
  logic lizzieLet22_4Lcall_$wmAdd_Int3_1sc_0_3_1wsie_2_1q1a8h_1_1t1a8m_1_1q2a8i_1_1t2a8n_1_1Lcall_$wmAdd_Int2_bufchan_r;
  assign lizzieLet22_4Lcall_$wmAdd_Int3_1sc_0_3_1wsie_2_1q1a8h_1_1t1a8m_1_1q2a8i_1_1t2a8n_1_1Lcall_$wmAdd_Int2_r = ((! lizzieLet22_4Lcall_$wmAdd_Int3_1sc_0_3_1wsie_2_1q1a8h_1_1t1a8m_1_1q2a8i_1_1t2a8n_1_1Lcall_$wmAdd_Int2_bufchan_d[0]) || lizzieLet22_4Lcall_$wmAdd_Int3_1sc_0_3_1wsie_2_1q1a8h_1_1t1a8m_1_1q2a8i_1_1t2a8n_1_1Lcall_$wmAdd_Int2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet22_4Lcall_$wmAdd_Int3_1sc_0_3_1wsie_2_1q1a8h_1_1t1a8m_1_1q2a8i_1_1t2a8n_1_1Lcall_$wmAdd_Int2_bufchan_d <= {115'd0,
                                                                                                                          1'd0};
    else
      if (lizzieLet22_4Lcall_$wmAdd_Int3_1sc_0_3_1wsie_2_1q1a8h_1_1t1a8m_1_1q2a8i_1_1t2a8n_1_1Lcall_$wmAdd_Int2_r)
        lizzieLet22_4Lcall_$wmAdd_Int3_1sc_0_3_1wsie_2_1q1a8h_1_1t1a8m_1_1q2a8i_1_1t2a8n_1_1Lcall_$wmAdd_Int2_bufchan_d <= lizzieLet22_4Lcall_$wmAdd_Int3_1sc_0_3_1wsie_2_1q1a8h_1_1t1a8m_1_1q2a8i_1_1t2a8n_1_1Lcall_$wmAdd_Int2_d;
  CT$wmAdd_Int_t lizzieLet22_4Lcall_$wmAdd_Int3_1sc_0_3_1wsie_2_1q1a8h_1_1t1a8m_1_1q2a8i_1_1t2a8n_1_1Lcall_$wmAdd_Int2_bufchan_buf;
  assign lizzieLet22_4Lcall_$wmAdd_Int3_1sc_0_3_1wsie_2_1q1a8h_1_1t1a8m_1_1q2a8i_1_1t2a8n_1_1Lcall_$wmAdd_Int2_bufchan_r = (! lizzieLet22_4Lcall_$wmAdd_Int3_1sc_0_3_1wsie_2_1q1a8h_1_1t1a8m_1_1q2a8i_1_1t2a8n_1_1Lcall_$wmAdd_Int2_bufchan_buf[0]);
  assign lizzieLet23_1_argbuf_d = (lizzieLet22_4Lcall_$wmAdd_Int3_1sc_0_3_1wsie_2_1q1a8h_1_1t1a8m_1_1q2a8i_1_1t2a8n_1_1Lcall_$wmAdd_Int2_bufchan_buf[0] ? lizzieLet22_4Lcall_$wmAdd_Int3_1sc_0_3_1wsie_2_1q1a8h_1_1t1a8m_1_1q2a8i_1_1t2a8n_1_1Lcall_$wmAdd_Int2_bufchan_buf :
                                   lizzieLet22_4Lcall_$wmAdd_Int3_1sc_0_3_1wsie_2_1q1a8h_1_1t1a8m_1_1q2a8i_1_1t2a8n_1_1Lcall_$wmAdd_Int2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet22_4Lcall_$wmAdd_Int3_1sc_0_3_1wsie_2_1q1a8h_1_1t1a8m_1_1q2a8i_1_1t2a8n_1_1Lcall_$wmAdd_Int2_bufchan_buf <= {115'd0,
                                                                                                                            1'd0};
    else
      if ((lizzieLet23_1_argbuf_r && lizzieLet22_4Lcall_$wmAdd_Int3_1sc_0_3_1wsie_2_1q1a8h_1_1t1a8m_1_1q2a8i_1_1t2a8n_1_1Lcall_$wmAdd_Int2_bufchan_buf[0]))
        lizzieLet22_4Lcall_$wmAdd_Int3_1sc_0_3_1wsie_2_1q1a8h_1_1t1a8m_1_1q2a8i_1_1t2a8n_1_1Lcall_$wmAdd_Int2_bufchan_buf <= {115'd0,
                                                                                                                              1'd0};
      else if (((! lizzieLet23_1_argbuf_r) && (! lizzieLet22_4Lcall_$wmAdd_Int3_1sc_0_3_1wsie_2_1q1a8h_1_1t1a8m_1_1q2a8i_1_1t2a8n_1_1Lcall_$wmAdd_Int2_bufchan_buf[0])))
        lizzieLet22_4Lcall_$wmAdd_Int3_1sc_0_3_1wsie_2_1q1a8h_1_1t1a8m_1_1q2a8i_1_1t2a8n_1_1Lcall_$wmAdd_Int2_bufchan_buf <= lizzieLet22_4Lcall_$wmAdd_Int3_1sc_0_3_1wsie_2_1q1a8h_1_1t1a8m_1_1q2a8i_1_1t2a8n_1_1Lcall_$wmAdd_Int2_bufchan_d;
  
  /* destruct (Ty CT$wnnz_Int,
          Dcon Lcall_$wnnz_Int0) : (lizzieLet27_1Lcall_$wnnz_Int0,CT$wnnz_Int) > [(wwsim_4_destruct,Int#),
                                                                                  (ww1XiS_2_destruct,Int#),
                                                                                  (ww2XiV_1_destruct,Int#),
                                                                                  (sc_0_10_destruct,Pointer_CT$wnnz_Int)] */
  logic [3:0] lizzieLet27_1Lcall_$wnnz_Int0_emitted;
  logic [3:0] lizzieLet27_1Lcall_$wnnz_Int0_done;
  assign wwsim_4_destruct_d = {lizzieLet27_1Lcall_$wnnz_Int0_d[35:4],
                               (lizzieLet27_1Lcall_$wnnz_Int0_d[0] && (! lizzieLet27_1Lcall_$wnnz_Int0_emitted[0]))};
  assign ww1XiS_2_destruct_d = {lizzieLet27_1Lcall_$wnnz_Int0_d[67:36],
                                (lizzieLet27_1Lcall_$wnnz_Int0_d[0] && (! lizzieLet27_1Lcall_$wnnz_Int0_emitted[1]))};
  assign ww2XiV_1_destruct_d = {lizzieLet27_1Lcall_$wnnz_Int0_d[99:68],
                                (lizzieLet27_1Lcall_$wnnz_Int0_d[0] && (! lizzieLet27_1Lcall_$wnnz_Int0_emitted[2]))};
  assign sc_0_10_destruct_d = {lizzieLet27_1Lcall_$wnnz_Int0_d[115:100],
                               (lizzieLet27_1Lcall_$wnnz_Int0_d[0] && (! lizzieLet27_1Lcall_$wnnz_Int0_emitted[3]))};
  assign lizzieLet27_1Lcall_$wnnz_Int0_done = (lizzieLet27_1Lcall_$wnnz_Int0_emitted | ({sc_0_10_destruct_d[0],
                                                                                         ww2XiV_1_destruct_d[0],
                                                                                         ww1XiS_2_destruct_d[0],
                                                                                         wwsim_4_destruct_d[0]} & {sc_0_10_destruct_r,
                                                                                                                   ww2XiV_1_destruct_r,
                                                                                                                   ww1XiS_2_destruct_r,
                                                                                                                   wwsim_4_destruct_r}));
  assign lizzieLet27_1Lcall_$wnnz_Int0_r = (& lizzieLet27_1Lcall_$wnnz_Int0_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet27_1Lcall_$wnnz_Int0_emitted <= 4'd0;
    else
      lizzieLet27_1Lcall_$wnnz_Int0_emitted <= (lizzieLet27_1Lcall_$wnnz_Int0_r ? 4'd0 :
                                                lizzieLet27_1Lcall_$wnnz_Int0_done);
  
  /* destruct (Ty CT$wnnz_Int,
          Dcon Lcall_$wnnz_Int1) : (lizzieLet27_1Lcall_$wnnz_Int1,CT$wnnz_Int) > [(wwsim_3_destruct,Int#),
                                                                                  (ww1XiS_1_destruct,Int#),
                                                                                  (sc_0_9_destruct,Pointer_CT$wnnz_Int),
                                                                                  (q4a8F_3_destruct,Pointer_QTree_Int)] */
  logic [3:0] lizzieLet27_1Lcall_$wnnz_Int1_emitted;
  logic [3:0] lizzieLet27_1Lcall_$wnnz_Int1_done;
  assign wwsim_3_destruct_d = {lizzieLet27_1Lcall_$wnnz_Int1_d[35:4],
                               (lizzieLet27_1Lcall_$wnnz_Int1_d[0] && (! lizzieLet27_1Lcall_$wnnz_Int1_emitted[0]))};
  assign ww1XiS_1_destruct_d = {lizzieLet27_1Lcall_$wnnz_Int1_d[67:36],
                                (lizzieLet27_1Lcall_$wnnz_Int1_d[0] && (! lizzieLet27_1Lcall_$wnnz_Int1_emitted[1]))};
  assign sc_0_9_destruct_d = {lizzieLet27_1Lcall_$wnnz_Int1_d[83:68],
                              (lizzieLet27_1Lcall_$wnnz_Int1_d[0] && (! lizzieLet27_1Lcall_$wnnz_Int1_emitted[2]))};
  assign q4a8F_3_destruct_d = {lizzieLet27_1Lcall_$wnnz_Int1_d[99:84],
                               (lizzieLet27_1Lcall_$wnnz_Int1_d[0] && (! lizzieLet27_1Lcall_$wnnz_Int1_emitted[3]))};
  assign lizzieLet27_1Lcall_$wnnz_Int1_done = (lizzieLet27_1Lcall_$wnnz_Int1_emitted | ({q4a8F_3_destruct_d[0],
                                                                                         sc_0_9_destruct_d[0],
                                                                                         ww1XiS_1_destruct_d[0],
                                                                                         wwsim_3_destruct_d[0]} & {q4a8F_3_destruct_r,
                                                                                                                   sc_0_9_destruct_r,
                                                                                                                   ww1XiS_1_destruct_r,
                                                                                                                   wwsim_3_destruct_r}));
  assign lizzieLet27_1Lcall_$wnnz_Int1_r = (& lizzieLet27_1Lcall_$wnnz_Int1_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet27_1Lcall_$wnnz_Int1_emitted <= 4'd0;
    else
      lizzieLet27_1Lcall_$wnnz_Int1_emitted <= (lizzieLet27_1Lcall_$wnnz_Int1_r ? 4'd0 :
                                                lizzieLet27_1Lcall_$wnnz_Int1_done);
  
  /* destruct (Ty CT$wnnz_Int,
          Dcon Lcall_$wnnz_Int2) : (lizzieLet27_1Lcall_$wnnz_Int2,CT$wnnz_Int) > [(wwsim_2_destruct,Int#),
                                                                                  (sc_0_8_destruct,Pointer_CT$wnnz_Int),
                                                                                  (q4a8F_2_destruct,Pointer_QTree_Int),
                                                                                  (q3a8E_2_destruct,Pointer_QTree_Int)] */
  logic [3:0] lizzieLet27_1Lcall_$wnnz_Int2_emitted;
  logic [3:0] lizzieLet27_1Lcall_$wnnz_Int2_done;
  assign wwsim_2_destruct_d = {lizzieLet27_1Lcall_$wnnz_Int2_d[35:4],
                               (lizzieLet27_1Lcall_$wnnz_Int2_d[0] && (! lizzieLet27_1Lcall_$wnnz_Int2_emitted[0]))};
  assign sc_0_8_destruct_d = {lizzieLet27_1Lcall_$wnnz_Int2_d[51:36],
                              (lizzieLet27_1Lcall_$wnnz_Int2_d[0] && (! lizzieLet27_1Lcall_$wnnz_Int2_emitted[1]))};
  assign q4a8F_2_destruct_d = {lizzieLet27_1Lcall_$wnnz_Int2_d[67:52],
                               (lizzieLet27_1Lcall_$wnnz_Int2_d[0] && (! lizzieLet27_1Lcall_$wnnz_Int2_emitted[2]))};
  assign q3a8E_2_destruct_d = {lizzieLet27_1Lcall_$wnnz_Int2_d[83:68],
                               (lizzieLet27_1Lcall_$wnnz_Int2_d[0] && (! lizzieLet27_1Lcall_$wnnz_Int2_emitted[3]))};
  assign lizzieLet27_1Lcall_$wnnz_Int2_done = (lizzieLet27_1Lcall_$wnnz_Int2_emitted | ({q3a8E_2_destruct_d[0],
                                                                                         q4a8F_2_destruct_d[0],
                                                                                         sc_0_8_destruct_d[0],
                                                                                         wwsim_2_destruct_d[0]} & {q3a8E_2_destruct_r,
                                                                                                                   q4a8F_2_destruct_r,
                                                                                                                   sc_0_8_destruct_r,
                                                                                                                   wwsim_2_destruct_r}));
  assign lizzieLet27_1Lcall_$wnnz_Int2_r = (& lizzieLet27_1Lcall_$wnnz_Int2_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet27_1Lcall_$wnnz_Int2_emitted <= 4'd0;
    else
      lizzieLet27_1Lcall_$wnnz_Int2_emitted <= (lizzieLet27_1Lcall_$wnnz_Int2_r ? 4'd0 :
                                                lizzieLet27_1Lcall_$wnnz_Int2_done);
  
  /* destruct (Ty CT$wnnz_Int,
          Dcon Lcall_$wnnz_Int3) : (lizzieLet27_1Lcall_$wnnz_Int3,CT$wnnz_Int) > [(sc_0_7_destruct,Pointer_CT$wnnz_Int),
                                                                                  (q4a8F_1_destruct,Pointer_QTree_Int),
                                                                                  (q3a8E_1_destruct,Pointer_QTree_Int),
                                                                                  (q2a8D_1_destruct,Pointer_QTree_Int)] */
  logic [3:0] lizzieLet27_1Lcall_$wnnz_Int3_emitted;
  logic [3:0] lizzieLet27_1Lcall_$wnnz_Int3_done;
  assign sc_0_7_destruct_d = {lizzieLet27_1Lcall_$wnnz_Int3_d[19:4],
                              (lizzieLet27_1Lcall_$wnnz_Int3_d[0] && (! lizzieLet27_1Lcall_$wnnz_Int3_emitted[0]))};
  assign q4a8F_1_destruct_d = {lizzieLet27_1Lcall_$wnnz_Int3_d[35:20],
                               (lizzieLet27_1Lcall_$wnnz_Int3_d[0] && (! lizzieLet27_1Lcall_$wnnz_Int3_emitted[1]))};
  assign q3a8E_1_destruct_d = {lizzieLet27_1Lcall_$wnnz_Int3_d[51:36],
                               (lizzieLet27_1Lcall_$wnnz_Int3_d[0] && (! lizzieLet27_1Lcall_$wnnz_Int3_emitted[2]))};
  assign q2a8D_1_destruct_d = {lizzieLet27_1Lcall_$wnnz_Int3_d[67:52],
                               (lizzieLet27_1Lcall_$wnnz_Int3_d[0] && (! lizzieLet27_1Lcall_$wnnz_Int3_emitted[3]))};
  assign lizzieLet27_1Lcall_$wnnz_Int3_done = (lizzieLet27_1Lcall_$wnnz_Int3_emitted | ({q2a8D_1_destruct_d[0],
                                                                                         q3a8E_1_destruct_d[0],
                                                                                         q4a8F_1_destruct_d[0],
                                                                                         sc_0_7_destruct_d[0]} & {q2a8D_1_destruct_r,
                                                                                                                  q3a8E_1_destruct_r,
                                                                                                                  q4a8F_1_destruct_r,
                                                                                                                  sc_0_7_destruct_r}));
  assign lizzieLet27_1Lcall_$wnnz_Int3_r = (& lizzieLet27_1Lcall_$wnnz_Int3_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet27_1Lcall_$wnnz_Int3_emitted <= 4'd0;
    else
      lizzieLet27_1Lcall_$wnnz_Int3_emitted <= (lizzieLet27_1Lcall_$wnnz_Int3_r ? 4'd0 :
                                                lizzieLet27_1Lcall_$wnnz_Int3_done);
  
  /* demux (Ty CT$wnnz_Int,
       Ty CT$wnnz_Int) : (lizzieLet27_2,CT$wnnz_Int) (lizzieLet27_1,CT$wnnz_Int) > [(_47,CT$wnnz_Int),
                                                                                    (lizzieLet27_1Lcall_$wnnz_Int3,CT$wnnz_Int),
                                                                                    (lizzieLet27_1Lcall_$wnnz_Int2,CT$wnnz_Int),
                                                                                    (lizzieLet27_1Lcall_$wnnz_Int1,CT$wnnz_Int),
                                                                                    (lizzieLet27_1Lcall_$wnnz_Int0,CT$wnnz_Int)] */
  logic [4:0] lizzieLet27_1_onehotd;
  always_comb
    if ((lizzieLet27_2_d[0] && lizzieLet27_1_d[0]))
      unique case (lizzieLet27_2_d[3:1])
        3'd0: lizzieLet27_1_onehotd = 5'd1;
        3'd1: lizzieLet27_1_onehotd = 5'd2;
        3'd2: lizzieLet27_1_onehotd = 5'd4;
        3'd3: lizzieLet27_1_onehotd = 5'd8;
        3'd4: lizzieLet27_1_onehotd = 5'd16;
        default: lizzieLet27_1_onehotd = 5'd0;
      endcase
    else lizzieLet27_1_onehotd = 5'd0;
  assign _47_d = {lizzieLet27_1_d[115:1], lizzieLet27_1_onehotd[0]};
  assign lizzieLet27_1Lcall_$wnnz_Int3_d = {lizzieLet27_1_d[115:1],
                                            lizzieLet27_1_onehotd[1]};
  assign lizzieLet27_1Lcall_$wnnz_Int2_d = {lizzieLet27_1_d[115:1],
                                            lizzieLet27_1_onehotd[2]};
  assign lizzieLet27_1Lcall_$wnnz_Int1_d = {lizzieLet27_1_d[115:1],
                                            lizzieLet27_1_onehotd[3]};
  assign lizzieLet27_1Lcall_$wnnz_Int0_d = {lizzieLet27_1_d[115:1],
                                            lizzieLet27_1_onehotd[4]};
  assign lizzieLet27_1_r = (| (lizzieLet27_1_onehotd & {lizzieLet27_1Lcall_$wnnz_Int0_r,
                                                        lizzieLet27_1Lcall_$wnnz_Int1_r,
                                                        lizzieLet27_1Lcall_$wnnz_Int2_r,
                                                        lizzieLet27_1Lcall_$wnnz_Int3_r,
                                                        _47_r}));
  assign lizzieLet27_2_r = lizzieLet27_1_r;
  
  /* demux (Ty CT$wnnz_Int,
       Ty Go) : (lizzieLet27_3,CT$wnnz_Int) (go_11_goMux_data,Go) > [(_46,Go),
                                                                     (lizzieLet27_3Lcall_$wnnz_Int3,Go),
                                                                     (lizzieLet27_3Lcall_$wnnz_Int2,Go),
                                                                     (lizzieLet27_3Lcall_$wnnz_Int1,Go),
                                                                     (lizzieLet27_3Lcall_$wnnz_Int0,Go)] */
  logic [4:0] go_11_goMux_data_onehotd;
  always_comb
    if ((lizzieLet27_3_d[0] && go_11_goMux_data_d[0]))
      unique case (lizzieLet27_3_d[3:1])
        3'd0: go_11_goMux_data_onehotd = 5'd1;
        3'd1: go_11_goMux_data_onehotd = 5'd2;
        3'd2: go_11_goMux_data_onehotd = 5'd4;
        3'd3: go_11_goMux_data_onehotd = 5'd8;
        3'd4: go_11_goMux_data_onehotd = 5'd16;
        default: go_11_goMux_data_onehotd = 5'd0;
      endcase
    else go_11_goMux_data_onehotd = 5'd0;
  assign _46_d = go_11_goMux_data_onehotd[0];
  assign lizzieLet27_3Lcall_$wnnz_Int3_d = go_11_goMux_data_onehotd[1];
  assign lizzieLet27_3Lcall_$wnnz_Int2_d = go_11_goMux_data_onehotd[2];
  assign lizzieLet27_3Lcall_$wnnz_Int1_d = go_11_goMux_data_onehotd[3];
  assign lizzieLet27_3Lcall_$wnnz_Int0_d = go_11_goMux_data_onehotd[4];
  assign go_11_goMux_data_r = (| (go_11_goMux_data_onehotd & {lizzieLet27_3Lcall_$wnnz_Int0_r,
                                                              lizzieLet27_3Lcall_$wnnz_Int1_r,
                                                              lizzieLet27_3Lcall_$wnnz_Int2_r,
                                                              lizzieLet27_3Lcall_$wnnz_Int3_r,
                                                              _46_r}));
  assign lizzieLet27_3_r = go_11_goMux_data_r;
  
  /* buf (Ty Go) : (lizzieLet27_3Lcall_$wnnz_Int0,Go) > (lizzieLet27_3Lcall_$wnnz_Int0_1_argbuf,Go) */
  Go_t lizzieLet27_3Lcall_$wnnz_Int0_bufchan_d;
  logic lizzieLet27_3Lcall_$wnnz_Int0_bufchan_r;
  assign lizzieLet27_3Lcall_$wnnz_Int0_r = ((! lizzieLet27_3Lcall_$wnnz_Int0_bufchan_d[0]) || lizzieLet27_3Lcall_$wnnz_Int0_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet27_3Lcall_$wnnz_Int0_bufchan_d <= 1'd0;
    else
      if (lizzieLet27_3Lcall_$wnnz_Int0_r)
        lizzieLet27_3Lcall_$wnnz_Int0_bufchan_d <= lizzieLet27_3Lcall_$wnnz_Int0_d;
  Go_t lizzieLet27_3Lcall_$wnnz_Int0_bufchan_buf;
  assign lizzieLet27_3Lcall_$wnnz_Int0_bufchan_r = (! lizzieLet27_3Lcall_$wnnz_Int0_bufchan_buf[0]);
  assign lizzieLet27_3Lcall_$wnnz_Int0_1_argbuf_d = (lizzieLet27_3Lcall_$wnnz_Int0_bufchan_buf[0] ? lizzieLet27_3Lcall_$wnnz_Int0_bufchan_buf :
                                                     lizzieLet27_3Lcall_$wnnz_Int0_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet27_3Lcall_$wnnz_Int0_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet27_3Lcall_$wnnz_Int0_1_argbuf_r && lizzieLet27_3Lcall_$wnnz_Int0_bufchan_buf[0]))
        lizzieLet27_3Lcall_$wnnz_Int0_bufchan_buf <= 1'd0;
      else if (((! lizzieLet27_3Lcall_$wnnz_Int0_1_argbuf_r) && (! lizzieLet27_3Lcall_$wnnz_Int0_bufchan_buf[0])))
        lizzieLet27_3Lcall_$wnnz_Int0_bufchan_buf <= lizzieLet27_3Lcall_$wnnz_Int0_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet27_3Lcall_$wnnz_Int1,Go) > (lizzieLet27_3Lcall_$wnnz_Int1_1_argbuf,Go) */
  Go_t lizzieLet27_3Lcall_$wnnz_Int1_bufchan_d;
  logic lizzieLet27_3Lcall_$wnnz_Int1_bufchan_r;
  assign lizzieLet27_3Lcall_$wnnz_Int1_r = ((! lizzieLet27_3Lcall_$wnnz_Int1_bufchan_d[0]) || lizzieLet27_3Lcall_$wnnz_Int1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet27_3Lcall_$wnnz_Int1_bufchan_d <= 1'd0;
    else
      if (lizzieLet27_3Lcall_$wnnz_Int1_r)
        lizzieLet27_3Lcall_$wnnz_Int1_bufchan_d <= lizzieLet27_3Lcall_$wnnz_Int1_d;
  Go_t lizzieLet27_3Lcall_$wnnz_Int1_bufchan_buf;
  assign lizzieLet27_3Lcall_$wnnz_Int1_bufchan_r = (! lizzieLet27_3Lcall_$wnnz_Int1_bufchan_buf[0]);
  assign lizzieLet27_3Lcall_$wnnz_Int1_1_argbuf_d = (lizzieLet27_3Lcall_$wnnz_Int1_bufchan_buf[0] ? lizzieLet27_3Lcall_$wnnz_Int1_bufchan_buf :
                                                     lizzieLet27_3Lcall_$wnnz_Int1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet27_3Lcall_$wnnz_Int1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet27_3Lcall_$wnnz_Int1_1_argbuf_r && lizzieLet27_3Lcall_$wnnz_Int1_bufchan_buf[0]))
        lizzieLet27_3Lcall_$wnnz_Int1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet27_3Lcall_$wnnz_Int1_1_argbuf_r) && (! lizzieLet27_3Lcall_$wnnz_Int1_bufchan_buf[0])))
        lizzieLet27_3Lcall_$wnnz_Int1_bufchan_buf <= lizzieLet27_3Lcall_$wnnz_Int1_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet27_3Lcall_$wnnz_Int2,Go) > (lizzieLet27_3Lcall_$wnnz_Int2_1_argbuf,Go) */
  Go_t lizzieLet27_3Lcall_$wnnz_Int2_bufchan_d;
  logic lizzieLet27_3Lcall_$wnnz_Int2_bufchan_r;
  assign lizzieLet27_3Lcall_$wnnz_Int2_r = ((! lizzieLet27_3Lcall_$wnnz_Int2_bufchan_d[0]) || lizzieLet27_3Lcall_$wnnz_Int2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet27_3Lcall_$wnnz_Int2_bufchan_d <= 1'd0;
    else
      if (lizzieLet27_3Lcall_$wnnz_Int2_r)
        lizzieLet27_3Lcall_$wnnz_Int2_bufchan_d <= lizzieLet27_3Lcall_$wnnz_Int2_d;
  Go_t lizzieLet27_3Lcall_$wnnz_Int2_bufchan_buf;
  assign lizzieLet27_3Lcall_$wnnz_Int2_bufchan_r = (! lizzieLet27_3Lcall_$wnnz_Int2_bufchan_buf[0]);
  assign lizzieLet27_3Lcall_$wnnz_Int2_1_argbuf_d = (lizzieLet27_3Lcall_$wnnz_Int2_bufchan_buf[0] ? lizzieLet27_3Lcall_$wnnz_Int2_bufchan_buf :
                                                     lizzieLet27_3Lcall_$wnnz_Int2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet27_3Lcall_$wnnz_Int2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet27_3Lcall_$wnnz_Int2_1_argbuf_r && lizzieLet27_3Lcall_$wnnz_Int2_bufchan_buf[0]))
        lizzieLet27_3Lcall_$wnnz_Int2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet27_3Lcall_$wnnz_Int2_1_argbuf_r) && (! lizzieLet27_3Lcall_$wnnz_Int2_bufchan_buf[0])))
        lizzieLet27_3Lcall_$wnnz_Int2_bufchan_buf <= lizzieLet27_3Lcall_$wnnz_Int2_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet27_3Lcall_$wnnz_Int3,Go) > (lizzieLet27_3Lcall_$wnnz_Int3_1_argbuf,Go) */
  Go_t lizzieLet27_3Lcall_$wnnz_Int3_bufchan_d;
  logic lizzieLet27_3Lcall_$wnnz_Int3_bufchan_r;
  assign lizzieLet27_3Lcall_$wnnz_Int3_r = ((! lizzieLet27_3Lcall_$wnnz_Int3_bufchan_d[0]) || lizzieLet27_3Lcall_$wnnz_Int3_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet27_3Lcall_$wnnz_Int3_bufchan_d <= 1'd0;
    else
      if (lizzieLet27_3Lcall_$wnnz_Int3_r)
        lizzieLet27_3Lcall_$wnnz_Int3_bufchan_d <= lizzieLet27_3Lcall_$wnnz_Int3_d;
  Go_t lizzieLet27_3Lcall_$wnnz_Int3_bufchan_buf;
  assign lizzieLet27_3Lcall_$wnnz_Int3_bufchan_r = (! lizzieLet27_3Lcall_$wnnz_Int3_bufchan_buf[0]);
  assign lizzieLet27_3Lcall_$wnnz_Int3_1_argbuf_d = (lizzieLet27_3Lcall_$wnnz_Int3_bufchan_buf[0] ? lizzieLet27_3Lcall_$wnnz_Int3_bufchan_buf :
                                                     lizzieLet27_3Lcall_$wnnz_Int3_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet27_3Lcall_$wnnz_Int3_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet27_3Lcall_$wnnz_Int3_1_argbuf_r && lizzieLet27_3Lcall_$wnnz_Int3_bufchan_buf[0]))
        lizzieLet27_3Lcall_$wnnz_Int3_bufchan_buf <= 1'd0;
      else if (((! lizzieLet27_3Lcall_$wnnz_Int3_1_argbuf_r) && (! lizzieLet27_3Lcall_$wnnz_Int3_bufchan_buf[0])))
        lizzieLet27_3Lcall_$wnnz_Int3_bufchan_buf <= lizzieLet27_3Lcall_$wnnz_Int3_bufchan_d;
  
  /* demux (Ty CT$wnnz_Int,
       Ty Int#) : (lizzieLet27_4,CT$wnnz_Int) (srtarg_0_1_goMux_mux,Int#) > [(lizzieLet27_4L$wnnz_Intsbos,Int#),
                                                                             (lizzieLet27_4Lcall_$wnnz_Int3,Int#),
                                                                             (lizzieLet27_4Lcall_$wnnz_Int2,Int#),
                                                                             (lizzieLet27_4Lcall_$wnnz_Int1,Int#),
                                                                             (lizzieLet27_4Lcall_$wnnz_Int0,Int#)] */
  logic [4:0] srtarg_0_1_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet27_4_d[0] && srtarg_0_1_goMux_mux_d[0]))
      unique case (lizzieLet27_4_d[3:1])
        3'd0: srtarg_0_1_goMux_mux_onehotd = 5'd1;
        3'd1: srtarg_0_1_goMux_mux_onehotd = 5'd2;
        3'd2: srtarg_0_1_goMux_mux_onehotd = 5'd4;
        3'd3: srtarg_0_1_goMux_mux_onehotd = 5'd8;
        3'd4: srtarg_0_1_goMux_mux_onehotd = 5'd16;
        default: srtarg_0_1_goMux_mux_onehotd = 5'd0;
      endcase
    else srtarg_0_1_goMux_mux_onehotd = 5'd0;
  assign lizzieLet27_4L$wnnz_Intsbos_d = {srtarg_0_1_goMux_mux_d[32:1],
                                          srtarg_0_1_goMux_mux_onehotd[0]};
  assign lizzieLet27_4Lcall_$wnnz_Int3_d = {srtarg_0_1_goMux_mux_d[32:1],
                                            srtarg_0_1_goMux_mux_onehotd[1]};
  assign lizzieLet27_4Lcall_$wnnz_Int2_d = {srtarg_0_1_goMux_mux_d[32:1],
                                            srtarg_0_1_goMux_mux_onehotd[2]};
  assign lizzieLet27_4Lcall_$wnnz_Int1_d = {srtarg_0_1_goMux_mux_d[32:1],
                                            srtarg_0_1_goMux_mux_onehotd[3]};
  assign lizzieLet27_4Lcall_$wnnz_Int0_d = {srtarg_0_1_goMux_mux_d[32:1],
                                            srtarg_0_1_goMux_mux_onehotd[4]};
  assign srtarg_0_1_goMux_mux_r = (| (srtarg_0_1_goMux_mux_onehotd & {lizzieLet27_4Lcall_$wnnz_Int0_r,
                                                                      lizzieLet27_4Lcall_$wnnz_Int1_r,
                                                                      lizzieLet27_4Lcall_$wnnz_Int2_r,
                                                                      lizzieLet27_4Lcall_$wnnz_Int3_r,
                                                                      lizzieLet27_4L$wnnz_Intsbos_r}));
  assign lizzieLet27_4_r = srtarg_0_1_goMux_mux_r;
  
  /* fork (Ty Int#) : (lizzieLet27_4L$wnnz_Intsbos,Int#) > [(lizzieLet27_4L$wnnz_Intsbos_1_merge_merge_fork_1,Int#),
                                                       (lizzieLet27_4L$wnnz_Intsbos_1_merge_merge_fork_2,Int#)] */
  logic [1:0] lizzieLet27_4L$wnnz_Intsbos_emitted;
  logic [1:0] lizzieLet27_4L$wnnz_Intsbos_done;
  assign lizzieLet27_4L$wnnz_Intsbos_1_merge_merge_fork_1_d = {lizzieLet27_4L$wnnz_Intsbos_d[32:1],
                                                               (lizzieLet27_4L$wnnz_Intsbos_d[0] && (! lizzieLet27_4L$wnnz_Intsbos_emitted[0]))};
  assign lizzieLet27_4L$wnnz_Intsbos_1_merge_merge_fork_2_d = {lizzieLet27_4L$wnnz_Intsbos_d[32:1],
                                                               (lizzieLet27_4L$wnnz_Intsbos_d[0] && (! lizzieLet27_4L$wnnz_Intsbos_emitted[1]))};
  assign lizzieLet27_4L$wnnz_Intsbos_done = (lizzieLet27_4L$wnnz_Intsbos_emitted | ({lizzieLet27_4L$wnnz_Intsbos_1_merge_merge_fork_2_d[0],
                                                                                     lizzieLet27_4L$wnnz_Intsbos_1_merge_merge_fork_1_d[0]} & {lizzieLet27_4L$wnnz_Intsbos_1_merge_merge_fork_2_r,
                                                                                                                                               lizzieLet27_4L$wnnz_Intsbos_1_merge_merge_fork_1_r}));
  assign lizzieLet27_4L$wnnz_Intsbos_r = (& lizzieLet27_4L$wnnz_Intsbos_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet27_4L$wnnz_Intsbos_emitted <= 2'd0;
    else
      lizzieLet27_4L$wnnz_Intsbos_emitted <= (lizzieLet27_4L$wnnz_Intsbos_r ? 2'd0 :
                                              lizzieLet27_4L$wnnz_Intsbos_done);
  
  /* togo (Ty Int#) : (lizzieLet27_4L$wnnz_Intsbos_1_merge_merge_fork_1,Int#) > (call_$wnnz_Int_goConst,Go) */
  assign call_$wnnz_Int_goConst_d = lizzieLet27_4L$wnnz_Intsbos_1_merge_merge_fork_1_d[0];
  assign lizzieLet27_4L$wnnz_Intsbos_1_merge_merge_fork_1_r = call_$wnnz_Int_goConst_r;
  
  /* buf (Ty Int#) : (lizzieLet27_4L$wnnz_Intsbos_1_merge_merge_fork_2,Int#) > ($wnnz_Int_resbuf,Int#) */
  \Int#_t  lizzieLet27_4L$wnnz_Intsbos_1_merge_merge_fork_2_bufchan_d;
  logic lizzieLet27_4L$wnnz_Intsbos_1_merge_merge_fork_2_bufchan_r;
  assign lizzieLet27_4L$wnnz_Intsbos_1_merge_merge_fork_2_r = ((! lizzieLet27_4L$wnnz_Intsbos_1_merge_merge_fork_2_bufchan_d[0]) || lizzieLet27_4L$wnnz_Intsbos_1_merge_merge_fork_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet27_4L$wnnz_Intsbos_1_merge_merge_fork_2_bufchan_d <= {32'd0,
                                                                     1'd0};
    else
      if (lizzieLet27_4L$wnnz_Intsbos_1_merge_merge_fork_2_r)
        lizzieLet27_4L$wnnz_Intsbos_1_merge_merge_fork_2_bufchan_d <= lizzieLet27_4L$wnnz_Intsbos_1_merge_merge_fork_2_d;
  \Int#_t  lizzieLet27_4L$wnnz_Intsbos_1_merge_merge_fork_2_bufchan_buf;
  assign lizzieLet27_4L$wnnz_Intsbos_1_merge_merge_fork_2_bufchan_r = (! lizzieLet27_4L$wnnz_Intsbos_1_merge_merge_fork_2_bufchan_buf[0]);
  assign \$wnnz_Int_resbuf_d  = (lizzieLet27_4L$wnnz_Intsbos_1_merge_merge_fork_2_bufchan_buf[0] ? lizzieLet27_4L$wnnz_Intsbos_1_merge_merge_fork_2_bufchan_buf :
                                 lizzieLet27_4L$wnnz_Intsbos_1_merge_merge_fork_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet27_4L$wnnz_Intsbos_1_merge_merge_fork_2_bufchan_buf <= {32'd0,
                                                                       1'd0};
    else
      if ((\$wnnz_Int_resbuf_r  && lizzieLet27_4L$wnnz_Intsbos_1_merge_merge_fork_2_bufchan_buf[0]))
        lizzieLet27_4L$wnnz_Intsbos_1_merge_merge_fork_2_bufchan_buf <= {32'd0,
                                                                         1'd0};
      else if (((! \$wnnz_Int_resbuf_r ) && (! lizzieLet27_4L$wnnz_Intsbos_1_merge_merge_fork_2_bufchan_buf[0])))
        lizzieLet27_4L$wnnz_Intsbos_1_merge_merge_fork_2_bufchan_buf <= lizzieLet27_4L$wnnz_Intsbos_1_merge_merge_fork_2_bufchan_d;
  
  /* dcon (Ty CT$wnnz_Int,
      Dcon Lcall_$wnnz_Int2) : [(lizzieLet27_4Lcall_$wnnz_Int3,Int#),
                                (sc_0_7_destruct,Pointer_CT$wnnz_Int),
                                (q4a8F_1_destruct,Pointer_QTree_Int),
                                (q3a8E_1_destruct,Pointer_QTree_Int)] > (lizzieLet27_4Lcall_$wnnz_Int3_1sc_0_7_1q4a8F_1_1q3a8E_1_1Lcall_$wnnz_Int2,CT$wnnz_Int) */
  assign lizzieLet27_4Lcall_$wnnz_Int3_1sc_0_7_1q4a8F_1_1q3a8E_1_1Lcall_$wnnz_Int2_d = Lcall_$wnnz_Int2_dc((& {lizzieLet27_4Lcall_$wnnz_Int3_d[0],
                                                                                                               sc_0_7_destruct_d[0],
                                                                                                               q4a8F_1_destruct_d[0],
                                                                                                               q3a8E_1_destruct_d[0]}), lizzieLet27_4Lcall_$wnnz_Int3_d, sc_0_7_destruct_d, q4a8F_1_destruct_d, q3a8E_1_destruct_d);
  assign {lizzieLet27_4Lcall_$wnnz_Int3_r,
          sc_0_7_destruct_r,
          q4a8F_1_destruct_r,
          q3a8E_1_destruct_r} = {4 {(lizzieLet27_4Lcall_$wnnz_Int3_1sc_0_7_1q4a8F_1_1q3a8E_1_1Lcall_$wnnz_Int2_r && lizzieLet27_4Lcall_$wnnz_Int3_1sc_0_7_1q4a8F_1_1q3a8E_1_1Lcall_$wnnz_Int2_d[0])}};
  
  /* buf (Ty CT$wnnz_Int) : (lizzieLet27_4Lcall_$wnnz_Int3_1sc_0_7_1q4a8F_1_1q3a8E_1_1Lcall_$wnnz_Int2,CT$wnnz_Int) > (lizzieLet28_1_argbuf,CT$wnnz_Int) */
  CT$wnnz_Int_t lizzieLet27_4Lcall_$wnnz_Int3_1sc_0_7_1q4a8F_1_1q3a8E_1_1Lcall_$wnnz_Int2_bufchan_d;
  logic lizzieLet27_4Lcall_$wnnz_Int3_1sc_0_7_1q4a8F_1_1q3a8E_1_1Lcall_$wnnz_Int2_bufchan_r;
  assign lizzieLet27_4Lcall_$wnnz_Int3_1sc_0_7_1q4a8F_1_1q3a8E_1_1Lcall_$wnnz_Int2_r = ((! lizzieLet27_4Lcall_$wnnz_Int3_1sc_0_7_1q4a8F_1_1q3a8E_1_1Lcall_$wnnz_Int2_bufchan_d[0]) || lizzieLet27_4Lcall_$wnnz_Int3_1sc_0_7_1q4a8F_1_1q3a8E_1_1Lcall_$wnnz_Int2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet27_4Lcall_$wnnz_Int3_1sc_0_7_1q4a8F_1_1q3a8E_1_1Lcall_$wnnz_Int2_bufchan_d <= {115'd0,
                                                                                              1'd0};
    else
      if (lizzieLet27_4Lcall_$wnnz_Int3_1sc_0_7_1q4a8F_1_1q3a8E_1_1Lcall_$wnnz_Int2_r)
        lizzieLet27_4Lcall_$wnnz_Int3_1sc_0_7_1q4a8F_1_1q3a8E_1_1Lcall_$wnnz_Int2_bufchan_d <= lizzieLet27_4Lcall_$wnnz_Int3_1sc_0_7_1q4a8F_1_1q3a8E_1_1Lcall_$wnnz_Int2_d;
  CT$wnnz_Int_t lizzieLet27_4Lcall_$wnnz_Int3_1sc_0_7_1q4a8F_1_1q3a8E_1_1Lcall_$wnnz_Int2_bufchan_buf;
  assign lizzieLet27_4Lcall_$wnnz_Int3_1sc_0_7_1q4a8F_1_1q3a8E_1_1Lcall_$wnnz_Int2_bufchan_r = (! lizzieLet27_4Lcall_$wnnz_Int3_1sc_0_7_1q4a8F_1_1q3a8E_1_1Lcall_$wnnz_Int2_bufchan_buf[0]);
  assign lizzieLet28_1_argbuf_d = (lizzieLet27_4Lcall_$wnnz_Int3_1sc_0_7_1q4a8F_1_1q3a8E_1_1Lcall_$wnnz_Int2_bufchan_buf[0] ? lizzieLet27_4Lcall_$wnnz_Int3_1sc_0_7_1q4a8F_1_1q3a8E_1_1Lcall_$wnnz_Int2_bufchan_buf :
                                   lizzieLet27_4Lcall_$wnnz_Int3_1sc_0_7_1q4a8F_1_1q3a8E_1_1Lcall_$wnnz_Int2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet27_4Lcall_$wnnz_Int3_1sc_0_7_1q4a8F_1_1q3a8E_1_1Lcall_$wnnz_Int2_bufchan_buf <= {115'd0,
                                                                                                1'd0};
    else
      if ((lizzieLet28_1_argbuf_r && lizzieLet27_4Lcall_$wnnz_Int3_1sc_0_7_1q4a8F_1_1q3a8E_1_1Lcall_$wnnz_Int2_bufchan_buf[0]))
        lizzieLet27_4Lcall_$wnnz_Int3_1sc_0_7_1q4a8F_1_1q3a8E_1_1Lcall_$wnnz_Int2_bufchan_buf <= {115'd0,
                                                                                                  1'd0};
      else if (((! lizzieLet28_1_argbuf_r) && (! lizzieLet27_4Lcall_$wnnz_Int3_1sc_0_7_1q4a8F_1_1q3a8E_1_1Lcall_$wnnz_Int2_bufchan_buf[0])))
        lizzieLet27_4Lcall_$wnnz_Int3_1sc_0_7_1q4a8F_1_1q3a8E_1_1Lcall_$wnnz_Int2_bufchan_buf <= lizzieLet27_4Lcall_$wnnz_Int3_1sc_0_7_1q4a8F_1_1q3a8E_1_1Lcall_$wnnz_Int2_bufchan_d;
  
  /* destruct (Ty QTree_Int,
          Dcon QNode_Int) : (lizzieLet2_1QNode_Int,QTree_Int) > [(q1a8h_destruct,Pointer_QTree_Int),
                                                                 (q2a8i_destruct,Pointer_QTree_Int),
                                                                 (q3a8j_destruct,Pointer_QTree_Int),
                                                                 (q4a8k_destruct,Pointer_QTree_Int)] */
  logic [3:0] lizzieLet2_1QNode_Int_emitted;
  logic [3:0] lizzieLet2_1QNode_Int_done;
  assign q1a8h_destruct_d = {lizzieLet2_1QNode_Int_d[18:3],
                             (lizzieLet2_1QNode_Int_d[0] && (! lizzieLet2_1QNode_Int_emitted[0]))};
  assign q2a8i_destruct_d = {lizzieLet2_1QNode_Int_d[34:19],
                             (lizzieLet2_1QNode_Int_d[0] && (! lizzieLet2_1QNode_Int_emitted[1]))};
  assign q3a8j_destruct_d = {lizzieLet2_1QNode_Int_d[50:35],
                             (lizzieLet2_1QNode_Int_d[0] && (! lizzieLet2_1QNode_Int_emitted[2]))};
  assign q4a8k_destruct_d = {lizzieLet2_1QNode_Int_d[66:51],
                             (lizzieLet2_1QNode_Int_d[0] && (! lizzieLet2_1QNode_Int_emitted[3]))};
  assign lizzieLet2_1QNode_Int_done = (lizzieLet2_1QNode_Int_emitted | ({q4a8k_destruct_d[0],
                                                                         q3a8j_destruct_d[0],
                                                                         q2a8i_destruct_d[0],
                                                                         q1a8h_destruct_d[0]} & {q4a8k_destruct_r,
                                                                                                 q3a8j_destruct_r,
                                                                                                 q2a8i_destruct_r,
                                                                                                 q1a8h_destruct_r}));
  assign lizzieLet2_1QNode_Int_r = (& lizzieLet2_1QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet2_1QNode_Int_emitted <= 4'd0;
    else
      lizzieLet2_1QNode_Int_emitted <= (lizzieLet2_1QNode_Int_r ? 4'd0 :
                                        lizzieLet2_1QNode_Int_done);
  
  /* destruct (Ty QTree_Int,
          Dcon QVal_Int) : (lizzieLet2_1QVal_Int,QTree_Int) > [(v1a8b_destruct,Int)] */
  assign v1a8b_destruct_d = {lizzieLet2_1QVal_Int_d[34:3],
                             lizzieLet2_1QVal_Int_d[0]};
  assign lizzieLet2_1QVal_Int_r = v1a8b_destruct_r;
  
  /* demux (Ty QTree_Int,
       Ty QTree_Int) : (lizzieLet2_2,QTree_Int) (lizzieLet2_1,QTree_Int) > [(_45,QTree_Int),
                                                                            (lizzieLet2_1QVal_Int,QTree_Int),
                                                                            (lizzieLet2_1QNode_Int,QTree_Int),
                                                                            (_44,QTree_Int)] */
  logic [3:0] lizzieLet2_1_onehotd;
  always_comb
    if ((lizzieLet2_2_d[0] && lizzieLet2_1_d[0]))
      unique case (lizzieLet2_2_d[2:1])
        2'd0: lizzieLet2_1_onehotd = 4'd1;
        2'd1: lizzieLet2_1_onehotd = 4'd2;
        2'd2: lizzieLet2_1_onehotd = 4'd4;
        2'd3: lizzieLet2_1_onehotd = 4'd8;
        default: lizzieLet2_1_onehotd = 4'd0;
      endcase
    else lizzieLet2_1_onehotd = 4'd0;
  assign _45_d = {lizzieLet2_1_d[66:1], lizzieLet2_1_onehotd[0]};
  assign lizzieLet2_1QVal_Int_d = {lizzieLet2_1_d[66:1],
                                   lizzieLet2_1_onehotd[1]};
  assign lizzieLet2_1QNode_Int_d = {lizzieLet2_1_d[66:1],
                                    lizzieLet2_1_onehotd[2]};
  assign _44_d = {lizzieLet2_1_d[66:1], lizzieLet2_1_onehotd[3]};
  assign lizzieLet2_1_r = (| (lizzieLet2_1_onehotd & {_44_r,
                                                      lizzieLet2_1QNode_Int_r,
                                                      lizzieLet2_1QVal_Int_r,
                                                      _45_r}));
  assign lizzieLet2_2_r = lizzieLet2_1_r;
  
  /* demux (Ty QTree_Int,
       Ty Go) : (lizzieLet2_3,QTree_Int) (go_6_goMux_data,Go) > [(lizzieLet2_3QNone_Int,Go),
                                                                 (lizzieLet2_3QVal_Int,Go),
                                                                 (lizzieLet2_3QNode_Int,Go),
                                                                 (lizzieLet2_3QError_Int,Go)] */
  logic [3:0] go_6_goMux_data_onehotd;
  always_comb
    if ((lizzieLet2_3_d[0] && go_6_goMux_data_d[0]))
      unique case (lizzieLet2_3_d[2:1])
        2'd0: go_6_goMux_data_onehotd = 4'd1;
        2'd1: go_6_goMux_data_onehotd = 4'd2;
        2'd2: go_6_goMux_data_onehotd = 4'd4;
        2'd3: go_6_goMux_data_onehotd = 4'd8;
        default: go_6_goMux_data_onehotd = 4'd0;
      endcase
    else go_6_goMux_data_onehotd = 4'd0;
  assign lizzieLet2_3QNone_Int_d = go_6_goMux_data_onehotd[0];
  assign lizzieLet2_3QVal_Int_d = go_6_goMux_data_onehotd[1];
  assign lizzieLet2_3QNode_Int_d = go_6_goMux_data_onehotd[2];
  assign lizzieLet2_3QError_Int_d = go_6_goMux_data_onehotd[3];
  assign go_6_goMux_data_r = (| (go_6_goMux_data_onehotd & {lizzieLet2_3QError_Int_r,
                                                            lizzieLet2_3QNode_Int_r,
                                                            lizzieLet2_3QVal_Int_r,
                                                            lizzieLet2_3QNone_Int_r}));
  assign lizzieLet2_3_r = go_6_goMux_data_r;
  
  /* fork (Ty Go) : (lizzieLet2_3QError_Int,Go) > [(lizzieLet2_3QError_Int_1,Go),
                                              (lizzieLet2_3QError_Int_2,Go)] */
  logic [1:0] lizzieLet2_3QError_Int_emitted;
  logic [1:0] lizzieLet2_3QError_Int_done;
  assign lizzieLet2_3QError_Int_1_d = (lizzieLet2_3QError_Int_d[0] && (! lizzieLet2_3QError_Int_emitted[0]));
  assign lizzieLet2_3QError_Int_2_d = (lizzieLet2_3QError_Int_d[0] && (! lizzieLet2_3QError_Int_emitted[1]));
  assign lizzieLet2_3QError_Int_done = (lizzieLet2_3QError_Int_emitted | ({lizzieLet2_3QError_Int_2_d[0],
                                                                           lizzieLet2_3QError_Int_1_d[0]} & {lizzieLet2_3QError_Int_2_r,
                                                                                                             lizzieLet2_3QError_Int_1_r}));
  assign lizzieLet2_3QError_Int_r = (& lizzieLet2_3QError_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet2_3QError_Int_emitted <= 2'd0;
    else
      lizzieLet2_3QError_Int_emitted <= (lizzieLet2_3QError_Int_r ? 2'd0 :
                                         lizzieLet2_3QError_Int_done);
  
  /* dcon (Ty QTree_Int,
      Dcon QError_Int) : [(lizzieLet2_3QError_Int_1,Go)] > (lizzieLet2_3QError_Int_1QError_Int,QTree_Int) */
  assign lizzieLet2_3QError_Int_1QError_Int_d = QError_Int_dc((& {lizzieLet2_3QError_Int_1_d[0]}), lizzieLet2_3QError_Int_1_d);
  assign {lizzieLet2_3QError_Int_1_r} = {1 {(lizzieLet2_3QError_Int_1QError_Int_r && lizzieLet2_3QError_Int_1QError_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (lizzieLet2_3QError_Int_1QError_Int,QTree_Int) > (lizzieLet11_1_1_argbuf,QTree_Int) */
  QTree_Int_t lizzieLet2_3QError_Int_1QError_Int_bufchan_d;
  logic lizzieLet2_3QError_Int_1QError_Int_bufchan_r;
  assign lizzieLet2_3QError_Int_1QError_Int_r = ((! lizzieLet2_3QError_Int_1QError_Int_bufchan_d[0]) || lizzieLet2_3QError_Int_1QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet2_3QError_Int_1QError_Int_bufchan_d <= {66'd0, 1'd0};
    else
      if (lizzieLet2_3QError_Int_1QError_Int_r)
        lizzieLet2_3QError_Int_1QError_Int_bufchan_d <= lizzieLet2_3QError_Int_1QError_Int_d;
  QTree_Int_t lizzieLet2_3QError_Int_1QError_Int_bufchan_buf;
  assign lizzieLet2_3QError_Int_1QError_Int_bufchan_r = (! lizzieLet2_3QError_Int_1QError_Int_bufchan_buf[0]);
  assign lizzieLet11_1_1_argbuf_d = (lizzieLet2_3QError_Int_1QError_Int_bufchan_buf[0] ? lizzieLet2_3QError_Int_1QError_Int_bufchan_buf :
                                     lizzieLet2_3QError_Int_1QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet2_3QError_Int_1QError_Int_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((lizzieLet11_1_1_argbuf_r && lizzieLet2_3QError_Int_1QError_Int_bufchan_buf[0]))
        lizzieLet2_3QError_Int_1QError_Int_bufchan_buf <= {66'd0, 1'd0};
      else if (((! lizzieLet11_1_1_argbuf_r) && (! lizzieLet2_3QError_Int_1QError_Int_bufchan_buf[0])))
        lizzieLet2_3QError_Int_1QError_Int_bufchan_buf <= lizzieLet2_3QError_Int_1QError_Int_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet2_3QError_Int_2,Go) > (lizzieLet2_3QError_Int_2_argbuf,Go) */
  Go_t lizzieLet2_3QError_Int_2_bufchan_d;
  logic lizzieLet2_3QError_Int_2_bufchan_r;
  assign lizzieLet2_3QError_Int_2_r = ((! lizzieLet2_3QError_Int_2_bufchan_d[0]) || lizzieLet2_3QError_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet2_3QError_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet2_3QError_Int_2_r)
        lizzieLet2_3QError_Int_2_bufchan_d <= lizzieLet2_3QError_Int_2_d;
  Go_t lizzieLet2_3QError_Int_2_bufchan_buf;
  assign lizzieLet2_3QError_Int_2_bufchan_r = (! lizzieLet2_3QError_Int_2_bufchan_buf[0]);
  assign lizzieLet2_3QError_Int_2_argbuf_d = (lizzieLet2_3QError_Int_2_bufchan_buf[0] ? lizzieLet2_3QError_Int_2_bufchan_buf :
                                              lizzieLet2_3QError_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet2_3QError_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet2_3QError_Int_2_argbuf_r && lizzieLet2_3QError_Int_2_bufchan_buf[0]))
        lizzieLet2_3QError_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet2_3QError_Int_2_argbuf_r) && (! lizzieLet2_3QError_Int_2_bufchan_buf[0])))
        lizzieLet2_3QError_Int_2_bufchan_buf <= lizzieLet2_3QError_Int_2_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet2_3QNone_Int,Go) > (lizzieLet2_3QNone_Int_1_argbuf,Go) */
  Go_t lizzieLet2_3QNone_Int_bufchan_d;
  logic lizzieLet2_3QNone_Int_bufchan_r;
  assign lizzieLet2_3QNone_Int_r = ((! lizzieLet2_3QNone_Int_bufchan_d[0]) || lizzieLet2_3QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet2_3QNone_Int_bufchan_d <= 1'd0;
    else
      if (lizzieLet2_3QNone_Int_r)
        lizzieLet2_3QNone_Int_bufchan_d <= lizzieLet2_3QNone_Int_d;
  Go_t lizzieLet2_3QNone_Int_bufchan_buf;
  assign lizzieLet2_3QNone_Int_bufchan_r = (! lizzieLet2_3QNone_Int_bufchan_buf[0]);
  assign lizzieLet2_3QNone_Int_1_argbuf_d = (lizzieLet2_3QNone_Int_bufchan_buf[0] ? lizzieLet2_3QNone_Int_bufchan_buf :
                                             lizzieLet2_3QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet2_3QNone_Int_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet2_3QNone_Int_1_argbuf_r && lizzieLet2_3QNone_Int_bufchan_buf[0]))
        lizzieLet2_3QNone_Int_bufchan_buf <= 1'd0;
      else if (((! lizzieLet2_3QNone_Int_1_argbuf_r) && (! lizzieLet2_3QNone_Int_bufchan_buf[0])))
        lizzieLet2_3QNone_Int_bufchan_buf <= lizzieLet2_3QNone_Int_bufchan_d;
  
  /* mergectrl (Ty C10,Ty Go) : [(lizzieLet2_3QNone_Int_1_argbuf,Go),
                            (lizzieLet22_3Lcall_$wmAdd_Int0_1_argbuf,Go),
                            (lizzieLet2_4QVal_Int_3QNone_Int_1_argbuf,Go),
                            (lizzieLet2_4QVal_Int_3QVal_Int_1_argbuf,Go),
                            (lizzieLet2_4QVal_Int_3QNode_Int_2_argbuf,Go),
                            (lizzieLet2_4QVal_Int_3QError_Int_2_argbuf,Go),
                            (lizzieLet2_4QNode_Int_3QNone_Int_1_argbuf,Go),
                            (lizzieLet2_4QNode_Int_3QVal_Int_2_argbuf,Go),
                            (lizzieLet2_4QNode_Int_3QError_Int_2_argbuf,Go),
                            (lizzieLet2_3QError_Int_2_argbuf,Go)] > (go_10_goMux_choice,C10) (go_10_goMux_data,Go) */
  logic [9:0] lizzieLet2_3QNone_Int_1_argbuf_select_d;
  assign lizzieLet2_3QNone_Int_1_argbuf_select_d = ((| lizzieLet2_3QNone_Int_1_argbuf_select_q) ? lizzieLet2_3QNone_Int_1_argbuf_select_q :
                                                    (lizzieLet2_3QNone_Int_1_argbuf_d[0] ? 10'd1 :
                                                     (lizzieLet22_3Lcall_$wmAdd_Int0_1_argbuf_d[0] ? 10'd2 :
                                                      (lizzieLet2_4QVal_Int_3QNone_Int_1_argbuf_d[0] ? 10'd4 :
                                                       (lizzieLet2_4QVal_Int_3QVal_Int_1_argbuf_d[0] ? 10'd8 :
                                                        (lizzieLet2_4QVal_Int_3QNode_Int_2_argbuf_d[0] ? 10'd16 :
                                                         (lizzieLet2_4QVal_Int_3QError_Int_2_argbuf_d[0] ? 10'd32 :
                                                          (lizzieLet2_4QNode_Int_3QNone_Int_1_argbuf_d[0] ? 10'd64 :
                                                           (lizzieLet2_4QNode_Int_3QVal_Int_2_argbuf_d[0] ? 10'd128 :
                                                            (lizzieLet2_4QNode_Int_3QError_Int_2_argbuf_d[0] ? 10'd256 :
                                                             (lizzieLet2_3QError_Int_2_argbuf_d[0] ? 10'd512 :
                                                              10'd0)))))))))));
  logic [9:0] lizzieLet2_3QNone_Int_1_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet2_3QNone_Int_1_argbuf_select_q <= 10'd0;
    else
      lizzieLet2_3QNone_Int_1_argbuf_select_q <= (lizzieLet2_3QNone_Int_1_argbuf_done ? 10'd0 :
                                                  lizzieLet2_3QNone_Int_1_argbuf_select_d);
  logic [1:0] lizzieLet2_3QNone_Int_1_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet2_3QNone_Int_1_argbuf_emit_q <= 2'd0;
    else
      lizzieLet2_3QNone_Int_1_argbuf_emit_q <= (lizzieLet2_3QNone_Int_1_argbuf_done ? 2'd0 :
                                                lizzieLet2_3QNone_Int_1_argbuf_emit_d);
  logic [1:0] lizzieLet2_3QNone_Int_1_argbuf_emit_d;
  assign lizzieLet2_3QNone_Int_1_argbuf_emit_d = (lizzieLet2_3QNone_Int_1_argbuf_emit_q | ({go_10_goMux_choice_d[0],
                                                                                            go_10_goMux_data_d[0]} & {go_10_goMux_choice_r,
                                                                                                                      go_10_goMux_data_r}));
  logic lizzieLet2_3QNone_Int_1_argbuf_done;
  assign lizzieLet2_3QNone_Int_1_argbuf_done = (& lizzieLet2_3QNone_Int_1_argbuf_emit_d);
  assign {lizzieLet2_3QError_Int_2_argbuf_r,
          lizzieLet2_4QNode_Int_3QError_Int_2_argbuf_r,
          lizzieLet2_4QNode_Int_3QVal_Int_2_argbuf_r,
          lizzieLet2_4QNode_Int_3QNone_Int_1_argbuf_r,
          lizzieLet2_4QVal_Int_3QError_Int_2_argbuf_r,
          lizzieLet2_4QVal_Int_3QNode_Int_2_argbuf_r,
          lizzieLet2_4QVal_Int_3QVal_Int_1_argbuf_r,
          lizzieLet2_4QVal_Int_3QNone_Int_1_argbuf_r,
          lizzieLet22_3Lcall_$wmAdd_Int0_1_argbuf_r,
          lizzieLet2_3QNone_Int_1_argbuf_r} = (lizzieLet2_3QNone_Int_1_argbuf_done ? lizzieLet2_3QNone_Int_1_argbuf_select_d :
                                               10'd0);
  assign go_10_goMux_data_d = ((lizzieLet2_3QNone_Int_1_argbuf_select_d[0] && (! lizzieLet2_3QNone_Int_1_argbuf_emit_q[0])) ? lizzieLet2_3QNone_Int_1_argbuf_d :
                               ((lizzieLet2_3QNone_Int_1_argbuf_select_d[1] && (! lizzieLet2_3QNone_Int_1_argbuf_emit_q[0])) ? lizzieLet22_3Lcall_$wmAdd_Int0_1_argbuf_d :
                                ((lizzieLet2_3QNone_Int_1_argbuf_select_d[2] && (! lizzieLet2_3QNone_Int_1_argbuf_emit_q[0])) ? lizzieLet2_4QVal_Int_3QNone_Int_1_argbuf_d :
                                 ((lizzieLet2_3QNone_Int_1_argbuf_select_d[3] && (! lizzieLet2_3QNone_Int_1_argbuf_emit_q[0])) ? lizzieLet2_4QVal_Int_3QVal_Int_1_argbuf_d :
                                  ((lizzieLet2_3QNone_Int_1_argbuf_select_d[4] && (! lizzieLet2_3QNone_Int_1_argbuf_emit_q[0])) ? lizzieLet2_4QVal_Int_3QNode_Int_2_argbuf_d :
                                   ((lizzieLet2_3QNone_Int_1_argbuf_select_d[5] && (! lizzieLet2_3QNone_Int_1_argbuf_emit_q[0])) ? lizzieLet2_4QVal_Int_3QError_Int_2_argbuf_d :
                                    ((lizzieLet2_3QNone_Int_1_argbuf_select_d[6] && (! lizzieLet2_3QNone_Int_1_argbuf_emit_q[0])) ? lizzieLet2_4QNode_Int_3QNone_Int_1_argbuf_d :
                                     ((lizzieLet2_3QNone_Int_1_argbuf_select_d[7] && (! lizzieLet2_3QNone_Int_1_argbuf_emit_q[0])) ? lizzieLet2_4QNode_Int_3QVal_Int_2_argbuf_d :
                                      ((lizzieLet2_3QNone_Int_1_argbuf_select_d[8] && (! lizzieLet2_3QNone_Int_1_argbuf_emit_q[0])) ? lizzieLet2_4QNode_Int_3QError_Int_2_argbuf_d :
                                       ((lizzieLet2_3QNone_Int_1_argbuf_select_d[9] && (! lizzieLet2_3QNone_Int_1_argbuf_emit_q[0])) ? lizzieLet2_3QError_Int_2_argbuf_d :
                                        1'd0))))))))));
  assign go_10_goMux_choice_d = ((lizzieLet2_3QNone_Int_1_argbuf_select_d[0] && (! lizzieLet2_3QNone_Int_1_argbuf_emit_q[1])) ? C1_10_dc(1'd1) :
                                 ((lizzieLet2_3QNone_Int_1_argbuf_select_d[1] && (! lizzieLet2_3QNone_Int_1_argbuf_emit_q[1])) ? C2_10_dc(1'd1) :
                                  ((lizzieLet2_3QNone_Int_1_argbuf_select_d[2] && (! lizzieLet2_3QNone_Int_1_argbuf_emit_q[1])) ? C3_10_dc(1'd1) :
                                   ((lizzieLet2_3QNone_Int_1_argbuf_select_d[3] && (! lizzieLet2_3QNone_Int_1_argbuf_emit_q[1])) ? C4_10_dc(1'd1) :
                                    ((lizzieLet2_3QNone_Int_1_argbuf_select_d[4] && (! lizzieLet2_3QNone_Int_1_argbuf_emit_q[1])) ? C5_10_dc(1'd1) :
                                     ((lizzieLet2_3QNone_Int_1_argbuf_select_d[5] && (! lizzieLet2_3QNone_Int_1_argbuf_emit_q[1])) ? C6_10_dc(1'd1) :
                                      ((lizzieLet2_3QNone_Int_1_argbuf_select_d[6] && (! lizzieLet2_3QNone_Int_1_argbuf_emit_q[1])) ? C7_10_dc(1'd1) :
                                       ((lizzieLet2_3QNone_Int_1_argbuf_select_d[7] && (! lizzieLet2_3QNone_Int_1_argbuf_emit_q[1])) ? C8_10_dc(1'd1) :
                                        ((lizzieLet2_3QNone_Int_1_argbuf_select_d[8] && (! lizzieLet2_3QNone_Int_1_argbuf_emit_q[1])) ? C9_10_dc(1'd1) :
                                         ((lizzieLet2_3QNone_Int_1_argbuf_select_d[9] && (! lizzieLet2_3QNone_Int_1_argbuf_emit_q[1])) ? C10_10_dc(1'd1) :
                                          {4'd0, 1'd0}))))))))));
  
  /* demux (Ty QTree_Int,
       Ty QTree_Int) : (lizzieLet2_4,QTree_Int) (readPointer_QTree_Intw2sig_1_1_argbuf_rwb,QTree_Int) > [(_43,QTree_Int),
                                                                                                         (lizzieLet2_4QVal_Int,QTree_Int),
                                                                                                         (lizzieLet2_4QNode_Int,QTree_Int),
                                                                                                         (_42,QTree_Int)] */
  logic [3:0] readPointer_QTree_Intw2sig_1_1_argbuf_rwb_onehotd;
  always_comb
    if ((lizzieLet2_4_d[0] && readPointer_QTree_Intw2sig_1_1_argbuf_rwb_d[0]))
      unique case (lizzieLet2_4_d[2:1])
        2'd0: readPointer_QTree_Intw2sig_1_1_argbuf_rwb_onehotd = 4'd1;
        2'd1: readPointer_QTree_Intw2sig_1_1_argbuf_rwb_onehotd = 4'd2;
        2'd2: readPointer_QTree_Intw2sig_1_1_argbuf_rwb_onehotd = 4'd4;
        2'd3: readPointer_QTree_Intw2sig_1_1_argbuf_rwb_onehotd = 4'd8;
        default: readPointer_QTree_Intw2sig_1_1_argbuf_rwb_onehotd = 4'd0;
      endcase
    else readPointer_QTree_Intw2sig_1_1_argbuf_rwb_onehotd = 4'd0;
  assign _43_d = {readPointer_QTree_Intw2sig_1_1_argbuf_rwb_d[66:1],
                  readPointer_QTree_Intw2sig_1_1_argbuf_rwb_onehotd[0]};
  assign lizzieLet2_4QVal_Int_d = {readPointer_QTree_Intw2sig_1_1_argbuf_rwb_d[66:1],
                                   readPointer_QTree_Intw2sig_1_1_argbuf_rwb_onehotd[1]};
  assign lizzieLet2_4QNode_Int_d = {readPointer_QTree_Intw2sig_1_1_argbuf_rwb_d[66:1],
                                    readPointer_QTree_Intw2sig_1_1_argbuf_rwb_onehotd[2]};
  assign _42_d = {readPointer_QTree_Intw2sig_1_1_argbuf_rwb_d[66:1],
                  readPointer_QTree_Intw2sig_1_1_argbuf_rwb_onehotd[3]};
  assign readPointer_QTree_Intw2sig_1_1_argbuf_rwb_r = (| (readPointer_QTree_Intw2sig_1_1_argbuf_rwb_onehotd & {_42_r,
                                                                                                                lizzieLet2_4QNode_Int_r,
                                                                                                                lizzieLet2_4QVal_Int_r,
                                                                                                                _43_r}));
  assign lizzieLet2_4_r = readPointer_QTree_Intw2sig_1_1_argbuf_rwb_r;
  
  /* fork (Ty QTree_Int) : (lizzieLet2_4QNode_Int,QTree_Int) > [(lizzieLet2_4QNode_Int_1,QTree_Int),
                                                           (lizzieLet2_4QNode_Int_2,QTree_Int),
                                                           (lizzieLet2_4QNode_Int_3,QTree_Int),
                                                           (lizzieLet2_4QNode_Int_4,QTree_Int),
                                                           (lizzieLet2_4QNode_Int_5,QTree_Int),
                                                           (lizzieLet2_4QNode_Int_6,QTree_Int),
                                                           (lizzieLet2_4QNode_Int_7,QTree_Int),
                                                           (lizzieLet2_4QNode_Int_8,QTree_Int),
                                                           (lizzieLet2_4QNode_Int_9,QTree_Int),
                                                           (lizzieLet2_4QNode_Int_10,QTree_Int)] */
  logic [9:0] lizzieLet2_4QNode_Int_emitted;
  logic [9:0] lizzieLet2_4QNode_Int_done;
  assign lizzieLet2_4QNode_Int_1_d = {lizzieLet2_4QNode_Int_d[66:1],
                                      (lizzieLet2_4QNode_Int_d[0] && (! lizzieLet2_4QNode_Int_emitted[0]))};
  assign lizzieLet2_4QNode_Int_2_d = {lizzieLet2_4QNode_Int_d[66:1],
                                      (lizzieLet2_4QNode_Int_d[0] && (! lizzieLet2_4QNode_Int_emitted[1]))};
  assign lizzieLet2_4QNode_Int_3_d = {lizzieLet2_4QNode_Int_d[66:1],
                                      (lizzieLet2_4QNode_Int_d[0] && (! lizzieLet2_4QNode_Int_emitted[2]))};
  assign lizzieLet2_4QNode_Int_4_d = {lizzieLet2_4QNode_Int_d[66:1],
                                      (lizzieLet2_4QNode_Int_d[0] && (! lizzieLet2_4QNode_Int_emitted[3]))};
  assign lizzieLet2_4QNode_Int_5_d = {lizzieLet2_4QNode_Int_d[66:1],
                                      (lizzieLet2_4QNode_Int_d[0] && (! lizzieLet2_4QNode_Int_emitted[4]))};
  assign lizzieLet2_4QNode_Int_6_d = {lizzieLet2_4QNode_Int_d[66:1],
                                      (lizzieLet2_4QNode_Int_d[0] && (! lizzieLet2_4QNode_Int_emitted[5]))};
  assign lizzieLet2_4QNode_Int_7_d = {lizzieLet2_4QNode_Int_d[66:1],
                                      (lizzieLet2_4QNode_Int_d[0] && (! lizzieLet2_4QNode_Int_emitted[6]))};
  assign lizzieLet2_4QNode_Int_8_d = {lizzieLet2_4QNode_Int_d[66:1],
                                      (lizzieLet2_4QNode_Int_d[0] && (! lizzieLet2_4QNode_Int_emitted[7]))};
  assign lizzieLet2_4QNode_Int_9_d = {lizzieLet2_4QNode_Int_d[66:1],
                                      (lizzieLet2_4QNode_Int_d[0] && (! lizzieLet2_4QNode_Int_emitted[8]))};
  assign lizzieLet2_4QNode_Int_10_d = {lizzieLet2_4QNode_Int_d[66:1],
                                       (lizzieLet2_4QNode_Int_d[0] && (! lizzieLet2_4QNode_Int_emitted[9]))};
  assign lizzieLet2_4QNode_Int_done = (lizzieLet2_4QNode_Int_emitted | ({lizzieLet2_4QNode_Int_10_d[0],
                                                                         lizzieLet2_4QNode_Int_9_d[0],
                                                                         lizzieLet2_4QNode_Int_8_d[0],
                                                                         lizzieLet2_4QNode_Int_7_d[0],
                                                                         lizzieLet2_4QNode_Int_6_d[0],
                                                                         lizzieLet2_4QNode_Int_5_d[0],
                                                                         lizzieLet2_4QNode_Int_4_d[0],
                                                                         lizzieLet2_4QNode_Int_3_d[0],
                                                                         lizzieLet2_4QNode_Int_2_d[0],
                                                                         lizzieLet2_4QNode_Int_1_d[0]} & {lizzieLet2_4QNode_Int_10_r,
                                                                                                          lizzieLet2_4QNode_Int_9_r,
                                                                                                          lizzieLet2_4QNode_Int_8_r,
                                                                                                          lizzieLet2_4QNode_Int_7_r,
                                                                                                          lizzieLet2_4QNode_Int_6_r,
                                                                                                          lizzieLet2_4QNode_Int_5_r,
                                                                                                          lizzieLet2_4QNode_Int_4_r,
                                                                                                          lizzieLet2_4QNode_Int_3_r,
                                                                                                          lizzieLet2_4QNode_Int_2_r,
                                                                                                          lizzieLet2_4QNode_Int_1_r}));
  assign lizzieLet2_4QNode_Int_r = (& lizzieLet2_4QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet2_4QNode_Int_emitted <= 10'd0;
    else
      lizzieLet2_4QNode_Int_emitted <= (lizzieLet2_4QNode_Int_r ? 10'd0 :
                                        lizzieLet2_4QNode_Int_done);
  
  /* demux (Ty QTree_Int,
       Ty Pointer_QTree_Int) : (lizzieLet2_4QNode_Int_10,QTree_Int) (q4a8k_destruct,Pointer_QTree_Int) > [(_41,Pointer_QTree_Int),
                                                                                                          (_40,Pointer_QTree_Int),
                                                                                                          (lizzieLet2_4QNode_Int_10QNode_Int,Pointer_QTree_Int),
                                                                                                          (_39,Pointer_QTree_Int)] */
  logic [3:0] q4a8k_destruct_onehotd;
  always_comb
    if ((lizzieLet2_4QNode_Int_10_d[0] && q4a8k_destruct_d[0]))
      unique case (lizzieLet2_4QNode_Int_10_d[2:1])
        2'd0: q4a8k_destruct_onehotd = 4'd1;
        2'd1: q4a8k_destruct_onehotd = 4'd2;
        2'd2: q4a8k_destruct_onehotd = 4'd4;
        2'd3: q4a8k_destruct_onehotd = 4'd8;
        default: q4a8k_destruct_onehotd = 4'd0;
      endcase
    else q4a8k_destruct_onehotd = 4'd0;
  assign _41_d = {q4a8k_destruct_d[16:1], q4a8k_destruct_onehotd[0]};
  assign _40_d = {q4a8k_destruct_d[16:1], q4a8k_destruct_onehotd[1]};
  assign lizzieLet2_4QNode_Int_10QNode_Int_d = {q4a8k_destruct_d[16:1],
                                                q4a8k_destruct_onehotd[2]};
  assign _39_d = {q4a8k_destruct_d[16:1], q4a8k_destruct_onehotd[3]};
  assign q4a8k_destruct_r = (| (q4a8k_destruct_onehotd & {_39_r,
                                                          lizzieLet2_4QNode_Int_10QNode_Int_r,
                                                          _40_r,
                                                          _41_r}));
  assign lizzieLet2_4QNode_Int_10_r = q4a8k_destruct_r;
  
  /* buf (Ty Pointer_QTree_Int) : (lizzieLet2_4QNode_Int_10QNode_Int,Pointer_QTree_Int) > (lizzieLet2_4QNode_Int_10QNode_Int_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t lizzieLet2_4QNode_Int_10QNode_Int_bufchan_d;
  logic lizzieLet2_4QNode_Int_10QNode_Int_bufchan_r;
  assign lizzieLet2_4QNode_Int_10QNode_Int_r = ((! lizzieLet2_4QNode_Int_10QNode_Int_bufchan_d[0]) || lizzieLet2_4QNode_Int_10QNode_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet2_4QNode_Int_10QNode_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet2_4QNode_Int_10QNode_Int_r)
        lizzieLet2_4QNode_Int_10QNode_Int_bufchan_d <= lizzieLet2_4QNode_Int_10QNode_Int_d;
  Pointer_QTree_Int_t lizzieLet2_4QNode_Int_10QNode_Int_bufchan_buf;
  assign lizzieLet2_4QNode_Int_10QNode_Int_bufchan_r = (! lizzieLet2_4QNode_Int_10QNode_Int_bufchan_buf[0]);
  assign lizzieLet2_4QNode_Int_10QNode_Int_1_argbuf_d = (lizzieLet2_4QNode_Int_10QNode_Int_bufchan_buf[0] ? lizzieLet2_4QNode_Int_10QNode_Int_bufchan_buf :
                                                         lizzieLet2_4QNode_Int_10QNode_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet2_4QNode_Int_10QNode_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet2_4QNode_Int_10QNode_Int_1_argbuf_r && lizzieLet2_4QNode_Int_10QNode_Int_bufchan_buf[0]))
        lizzieLet2_4QNode_Int_10QNode_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet2_4QNode_Int_10QNode_Int_1_argbuf_r) && (! lizzieLet2_4QNode_Int_10QNode_Int_bufchan_buf[0])))
        lizzieLet2_4QNode_Int_10QNode_Int_bufchan_buf <= lizzieLet2_4QNode_Int_10QNode_Int_bufchan_d;
  
  /* destruct (Ty QTree_Int,
          Dcon QNode_Int) : (lizzieLet2_4QNode_Int_1QNode_Int,QTree_Int) > [(t1a8m_destruct,Pointer_QTree_Int),
                                                                            (t2a8n_destruct,Pointer_QTree_Int),
                                                                            (t3a8o_destruct,Pointer_QTree_Int),
                                                                            (t4a8p_destruct,Pointer_QTree_Int)] */
  logic [3:0] lizzieLet2_4QNode_Int_1QNode_Int_emitted;
  logic [3:0] lizzieLet2_4QNode_Int_1QNode_Int_done;
  assign t1a8m_destruct_d = {lizzieLet2_4QNode_Int_1QNode_Int_d[18:3],
                             (lizzieLet2_4QNode_Int_1QNode_Int_d[0] && (! lizzieLet2_4QNode_Int_1QNode_Int_emitted[0]))};
  assign t2a8n_destruct_d = {lizzieLet2_4QNode_Int_1QNode_Int_d[34:19],
                             (lizzieLet2_4QNode_Int_1QNode_Int_d[0] && (! lizzieLet2_4QNode_Int_1QNode_Int_emitted[1]))};
  assign t3a8o_destruct_d = {lizzieLet2_4QNode_Int_1QNode_Int_d[50:35],
                             (lizzieLet2_4QNode_Int_1QNode_Int_d[0] && (! lizzieLet2_4QNode_Int_1QNode_Int_emitted[2]))};
  assign t4a8p_destruct_d = {lizzieLet2_4QNode_Int_1QNode_Int_d[66:51],
                             (lizzieLet2_4QNode_Int_1QNode_Int_d[0] && (! lizzieLet2_4QNode_Int_1QNode_Int_emitted[3]))};
  assign lizzieLet2_4QNode_Int_1QNode_Int_done = (lizzieLet2_4QNode_Int_1QNode_Int_emitted | ({t4a8p_destruct_d[0],
                                                                                               t3a8o_destruct_d[0],
                                                                                               t2a8n_destruct_d[0],
                                                                                               t1a8m_destruct_d[0]} & {t4a8p_destruct_r,
                                                                                                                       t3a8o_destruct_r,
                                                                                                                       t2a8n_destruct_r,
                                                                                                                       t1a8m_destruct_r}));
  assign lizzieLet2_4QNode_Int_1QNode_Int_r = (& lizzieLet2_4QNode_Int_1QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet2_4QNode_Int_1QNode_Int_emitted <= 4'd0;
    else
      lizzieLet2_4QNode_Int_1QNode_Int_emitted <= (lizzieLet2_4QNode_Int_1QNode_Int_r ? 4'd0 :
                                                   lizzieLet2_4QNode_Int_1QNode_Int_done);
  
  /* demux (Ty QTree_Int,
       Ty QTree_Int) : (lizzieLet2_4QNode_Int_2,QTree_Int) (lizzieLet2_4QNode_Int_1,QTree_Int) > [(_38,QTree_Int),
                                                                                                  (_37,QTree_Int),
                                                                                                  (lizzieLet2_4QNode_Int_1QNode_Int,QTree_Int),
                                                                                                  (_36,QTree_Int)] */
  logic [3:0] lizzieLet2_4QNode_Int_1_onehotd;
  always_comb
    if ((lizzieLet2_4QNode_Int_2_d[0] && lizzieLet2_4QNode_Int_1_d[0]))
      unique case (lizzieLet2_4QNode_Int_2_d[2:1])
        2'd0: lizzieLet2_4QNode_Int_1_onehotd = 4'd1;
        2'd1: lizzieLet2_4QNode_Int_1_onehotd = 4'd2;
        2'd2: lizzieLet2_4QNode_Int_1_onehotd = 4'd4;
        2'd3: lizzieLet2_4QNode_Int_1_onehotd = 4'd8;
        default: lizzieLet2_4QNode_Int_1_onehotd = 4'd0;
      endcase
    else lizzieLet2_4QNode_Int_1_onehotd = 4'd0;
  assign _38_d = {lizzieLet2_4QNode_Int_1_d[66:1],
                  lizzieLet2_4QNode_Int_1_onehotd[0]};
  assign _37_d = {lizzieLet2_4QNode_Int_1_d[66:1],
                  lizzieLet2_4QNode_Int_1_onehotd[1]};
  assign lizzieLet2_4QNode_Int_1QNode_Int_d = {lizzieLet2_4QNode_Int_1_d[66:1],
                                               lizzieLet2_4QNode_Int_1_onehotd[2]};
  assign _36_d = {lizzieLet2_4QNode_Int_1_d[66:1],
                  lizzieLet2_4QNode_Int_1_onehotd[3]};
  assign lizzieLet2_4QNode_Int_1_r = (| (lizzieLet2_4QNode_Int_1_onehotd & {_36_r,
                                                                            lizzieLet2_4QNode_Int_1QNode_Int_r,
                                                                            _37_r,
                                                                            _38_r}));
  assign lizzieLet2_4QNode_Int_2_r = lizzieLet2_4QNode_Int_1_r;
  
  /* demux (Ty QTree_Int,
       Ty Go) : (lizzieLet2_4QNode_Int_3,QTree_Int) (lizzieLet2_3QNode_Int,Go) > [(lizzieLet2_4QNode_Int_3QNone_Int,Go),
                                                                                  (lizzieLet2_4QNode_Int_3QVal_Int,Go),
                                                                                  (lizzieLet2_4QNode_Int_3QNode_Int,Go),
                                                                                  (lizzieLet2_4QNode_Int_3QError_Int,Go)] */
  logic [3:0] lizzieLet2_3QNode_Int_onehotd;
  always_comb
    if ((lizzieLet2_4QNode_Int_3_d[0] && lizzieLet2_3QNode_Int_d[0]))
      unique case (lizzieLet2_4QNode_Int_3_d[2:1])
        2'd0: lizzieLet2_3QNode_Int_onehotd = 4'd1;
        2'd1: lizzieLet2_3QNode_Int_onehotd = 4'd2;
        2'd2: lizzieLet2_3QNode_Int_onehotd = 4'd4;
        2'd3: lizzieLet2_3QNode_Int_onehotd = 4'd8;
        default: lizzieLet2_3QNode_Int_onehotd = 4'd0;
      endcase
    else lizzieLet2_3QNode_Int_onehotd = 4'd0;
  assign lizzieLet2_4QNode_Int_3QNone_Int_d = lizzieLet2_3QNode_Int_onehotd[0];
  assign lizzieLet2_4QNode_Int_3QVal_Int_d = lizzieLet2_3QNode_Int_onehotd[1];
  assign lizzieLet2_4QNode_Int_3QNode_Int_d = lizzieLet2_3QNode_Int_onehotd[2];
  assign lizzieLet2_4QNode_Int_3QError_Int_d = lizzieLet2_3QNode_Int_onehotd[3];
  assign lizzieLet2_3QNode_Int_r = (| (lizzieLet2_3QNode_Int_onehotd & {lizzieLet2_4QNode_Int_3QError_Int_r,
                                                                        lizzieLet2_4QNode_Int_3QNode_Int_r,
                                                                        lizzieLet2_4QNode_Int_3QVal_Int_r,
                                                                        lizzieLet2_4QNode_Int_3QNone_Int_r}));
  assign lizzieLet2_4QNode_Int_3_r = lizzieLet2_3QNode_Int_r;
  
  /* fork (Ty Go) : (lizzieLet2_4QNode_Int_3QError_Int,Go) > [(lizzieLet2_4QNode_Int_3QError_Int_1,Go),
                                                         (lizzieLet2_4QNode_Int_3QError_Int_2,Go)] */
  logic [1:0] lizzieLet2_4QNode_Int_3QError_Int_emitted;
  logic [1:0] lizzieLet2_4QNode_Int_3QError_Int_done;
  assign lizzieLet2_4QNode_Int_3QError_Int_1_d = (lizzieLet2_4QNode_Int_3QError_Int_d[0] && (! lizzieLet2_4QNode_Int_3QError_Int_emitted[0]));
  assign lizzieLet2_4QNode_Int_3QError_Int_2_d = (lizzieLet2_4QNode_Int_3QError_Int_d[0] && (! lizzieLet2_4QNode_Int_3QError_Int_emitted[1]));
  assign lizzieLet2_4QNode_Int_3QError_Int_done = (lizzieLet2_4QNode_Int_3QError_Int_emitted | ({lizzieLet2_4QNode_Int_3QError_Int_2_d[0],
                                                                                                 lizzieLet2_4QNode_Int_3QError_Int_1_d[0]} & {lizzieLet2_4QNode_Int_3QError_Int_2_r,
                                                                                                                                              lizzieLet2_4QNode_Int_3QError_Int_1_r}));
  assign lizzieLet2_4QNode_Int_3QError_Int_r = (& lizzieLet2_4QNode_Int_3QError_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet2_4QNode_Int_3QError_Int_emitted <= 2'd0;
    else
      lizzieLet2_4QNode_Int_3QError_Int_emitted <= (lizzieLet2_4QNode_Int_3QError_Int_r ? 2'd0 :
                                                    lizzieLet2_4QNode_Int_3QError_Int_done);
  
  /* dcon (Ty QTree_Int,
      Dcon QError_Int) : [(lizzieLet2_4QNode_Int_3QError_Int_1,Go)] > (lizzieLet2_4QNode_Int_3QError_Int_1QError_Int,QTree_Int) */
  assign lizzieLet2_4QNode_Int_3QError_Int_1QError_Int_d = QError_Int_dc((& {lizzieLet2_4QNode_Int_3QError_Int_1_d[0]}), lizzieLet2_4QNode_Int_3QError_Int_1_d);
  assign {lizzieLet2_4QNode_Int_3QError_Int_1_r} = {1 {(lizzieLet2_4QNode_Int_3QError_Int_1QError_Int_r && lizzieLet2_4QNode_Int_3QError_Int_1QError_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (lizzieLet2_4QNode_Int_3QError_Int_1QError_Int,QTree_Int) > (lizzieLet10_1_1_argbuf,QTree_Int) */
  QTree_Int_t lizzieLet2_4QNode_Int_3QError_Int_1QError_Int_bufchan_d;
  logic lizzieLet2_4QNode_Int_3QError_Int_1QError_Int_bufchan_r;
  assign lizzieLet2_4QNode_Int_3QError_Int_1QError_Int_r = ((! lizzieLet2_4QNode_Int_3QError_Int_1QError_Int_bufchan_d[0]) || lizzieLet2_4QNode_Int_3QError_Int_1QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet2_4QNode_Int_3QError_Int_1QError_Int_bufchan_d <= {66'd0,
                                                                  1'd0};
    else
      if (lizzieLet2_4QNode_Int_3QError_Int_1QError_Int_r)
        lizzieLet2_4QNode_Int_3QError_Int_1QError_Int_bufchan_d <= lizzieLet2_4QNode_Int_3QError_Int_1QError_Int_d;
  QTree_Int_t lizzieLet2_4QNode_Int_3QError_Int_1QError_Int_bufchan_buf;
  assign lizzieLet2_4QNode_Int_3QError_Int_1QError_Int_bufchan_r = (! lizzieLet2_4QNode_Int_3QError_Int_1QError_Int_bufchan_buf[0]);
  assign lizzieLet10_1_1_argbuf_d = (lizzieLet2_4QNode_Int_3QError_Int_1QError_Int_bufchan_buf[0] ? lizzieLet2_4QNode_Int_3QError_Int_1QError_Int_bufchan_buf :
                                     lizzieLet2_4QNode_Int_3QError_Int_1QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet2_4QNode_Int_3QError_Int_1QError_Int_bufchan_buf <= {66'd0,
                                                                    1'd0};
    else
      if ((lizzieLet10_1_1_argbuf_r && lizzieLet2_4QNode_Int_3QError_Int_1QError_Int_bufchan_buf[0]))
        lizzieLet2_4QNode_Int_3QError_Int_1QError_Int_bufchan_buf <= {66'd0,
                                                                      1'd0};
      else if (((! lizzieLet10_1_1_argbuf_r) && (! lizzieLet2_4QNode_Int_3QError_Int_1QError_Int_bufchan_buf[0])))
        lizzieLet2_4QNode_Int_3QError_Int_1QError_Int_bufchan_buf <= lizzieLet2_4QNode_Int_3QError_Int_1QError_Int_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet2_4QNode_Int_3QError_Int_2,Go) > (lizzieLet2_4QNode_Int_3QError_Int_2_argbuf,Go) */
  Go_t lizzieLet2_4QNode_Int_3QError_Int_2_bufchan_d;
  logic lizzieLet2_4QNode_Int_3QError_Int_2_bufchan_r;
  assign lizzieLet2_4QNode_Int_3QError_Int_2_r = ((! lizzieLet2_4QNode_Int_3QError_Int_2_bufchan_d[0]) || lizzieLet2_4QNode_Int_3QError_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet2_4QNode_Int_3QError_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet2_4QNode_Int_3QError_Int_2_r)
        lizzieLet2_4QNode_Int_3QError_Int_2_bufchan_d <= lizzieLet2_4QNode_Int_3QError_Int_2_d;
  Go_t lizzieLet2_4QNode_Int_3QError_Int_2_bufchan_buf;
  assign lizzieLet2_4QNode_Int_3QError_Int_2_bufchan_r = (! lizzieLet2_4QNode_Int_3QError_Int_2_bufchan_buf[0]);
  assign lizzieLet2_4QNode_Int_3QError_Int_2_argbuf_d = (lizzieLet2_4QNode_Int_3QError_Int_2_bufchan_buf[0] ? lizzieLet2_4QNode_Int_3QError_Int_2_bufchan_buf :
                                                         lizzieLet2_4QNode_Int_3QError_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet2_4QNode_Int_3QError_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet2_4QNode_Int_3QError_Int_2_argbuf_r && lizzieLet2_4QNode_Int_3QError_Int_2_bufchan_buf[0]))
        lizzieLet2_4QNode_Int_3QError_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet2_4QNode_Int_3QError_Int_2_argbuf_r) && (! lizzieLet2_4QNode_Int_3QError_Int_2_bufchan_buf[0])))
        lizzieLet2_4QNode_Int_3QError_Int_2_bufchan_buf <= lizzieLet2_4QNode_Int_3QError_Int_2_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet2_4QNode_Int_3QNode_Int,Go) > (lizzieLet2_4QNode_Int_3QNode_Int_1_argbuf,Go) */
  Go_t lizzieLet2_4QNode_Int_3QNode_Int_bufchan_d;
  logic lizzieLet2_4QNode_Int_3QNode_Int_bufchan_r;
  assign lizzieLet2_4QNode_Int_3QNode_Int_r = ((! lizzieLet2_4QNode_Int_3QNode_Int_bufchan_d[0]) || lizzieLet2_4QNode_Int_3QNode_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet2_4QNode_Int_3QNode_Int_bufchan_d <= 1'd0;
    else
      if (lizzieLet2_4QNode_Int_3QNode_Int_r)
        lizzieLet2_4QNode_Int_3QNode_Int_bufchan_d <= lizzieLet2_4QNode_Int_3QNode_Int_d;
  Go_t lizzieLet2_4QNode_Int_3QNode_Int_bufchan_buf;
  assign lizzieLet2_4QNode_Int_3QNode_Int_bufchan_r = (! lizzieLet2_4QNode_Int_3QNode_Int_bufchan_buf[0]);
  assign lizzieLet2_4QNode_Int_3QNode_Int_1_argbuf_d = (lizzieLet2_4QNode_Int_3QNode_Int_bufchan_buf[0] ? lizzieLet2_4QNode_Int_3QNode_Int_bufchan_buf :
                                                        lizzieLet2_4QNode_Int_3QNode_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet2_4QNode_Int_3QNode_Int_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet2_4QNode_Int_3QNode_Int_1_argbuf_r && lizzieLet2_4QNode_Int_3QNode_Int_bufchan_buf[0]))
        lizzieLet2_4QNode_Int_3QNode_Int_bufchan_buf <= 1'd0;
      else if (((! lizzieLet2_4QNode_Int_3QNode_Int_1_argbuf_r) && (! lizzieLet2_4QNode_Int_3QNode_Int_bufchan_buf[0])))
        lizzieLet2_4QNode_Int_3QNode_Int_bufchan_buf <= lizzieLet2_4QNode_Int_3QNode_Int_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet2_4QNode_Int_3QNone_Int,Go) > (lizzieLet2_4QNode_Int_3QNone_Int_1_argbuf,Go) */
  Go_t lizzieLet2_4QNode_Int_3QNone_Int_bufchan_d;
  logic lizzieLet2_4QNode_Int_3QNone_Int_bufchan_r;
  assign lizzieLet2_4QNode_Int_3QNone_Int_r = ((! lizzieLet2_4QNode_Int_3QNone_Int_bufchan_d[0]) || lizzieLet2_4QNode_Int_3QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet2_4QNode_Int_3QNone_Int_bufchan_d <= 1'd0;
    else
      if (lizzieLet2_4QNode_Int_3QNone_Int_r)
        lizzieLet2_4QNode_Int_3QNone_Int_bufchan_d <= lizzieLet2_4QNode_Int_3QNone_Int_d;
  Go_t lizzieLet2_4QNode_Int_3QNone_Int_bufchan_buf;
  assign lizzieLet2_4QNode_Int_3QNone_Int_bufchan_r = (! lizzieLet2_4QNode_Int_3QNone_Int_bufchan_buf[0]);
  assign lizzieLet2_4QNode_Int_3QNone_Int_1_argbuf_d = (lizzieLet2_4QNode_Int_3QNone_Int_bufchan_buf[0] ? lizzieLet2_4QNode_Int_3QNone_Int_bufchan_buf :
                                                        lizzieLet2_4QNode_Int_3QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet2_4QNode_Int_3QNone_Int_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet2_4QNode_Int_3QNone_Int_1_argbuf_r && lizzieLet2_4QNode_Int_3QNone_Int_bufchan_buf[0]))
        lizzieLet2_4QNode_Int_3QNone_Int_bufchan_buf <= 1'd0;
      else if (((! lizzieLet2_4QNode_Int_3QNone_Int_1_argbuf_r) && (! lizzieLet2_4QNode_Int_3QNone_Int_bufchan_buf[0])))
        lizzieLet2_4QNode_Int_3QNone_Int_bufchan_buf <= lizzieLet2_4QNode_Int_3QNone_Int_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet2_4QNode_Int_3QVal_Int,Go) > [(lizzieLet2_4QNode_Int_3QVal_Int_1,Go),
                                                       (lizzieLet2_4QNode_Int_3QVal_Int_2,Go)] */
  logic [1:0] lizzieLet2_4QNode_Int_3QVal_Int_emitted;
  logic [1:0] lizzieLet2_4QNode_Int_3QVal_Int_done;
  assign lizzieLet2_4QNode_Int_3QVal_Int_1_d = (lizzieLet2_4QNode_Int_3QVal_Int_d[0] && (! lizzieLet2_4QNode_Int_3QVal_Int_emitted[0]));
  assign lizzieLet2_4QNode_Int_3QVal_Int_2_d = (lizzieLet2_4QNode_Int_3QVal_Int_d[0] && (! lizzieLet2_4QNode_Int_3QVal_Int_emitted[1]));
  assign lizzieLet2_4QNode_Int_3QVal_Int_done = (lizzieLet2_4QNode_Int_3QVal_Int_emitted | ({lizzieLet2_4QNode_Int_3QVal_Int_2_d[0],
                                                                                             lizzieLet2_4QNode_Int_3QVal_Int_1_d[0]} & {lizzieLet2_4QNode_Int_3QVal_Int_2_r,
                                                                                                                                        lizzieLet2_4QNode_Int_3QVal_Int_1_r}));
  assign lizzieLet2_4QNode_Int_3QVal_Int_r = (& lizzieLet2_4QNode_Int_3QVal_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet2_4QNode_Int_3QVal_Int_emitted <= 2'd0;
    else
      lizzieLet2_4QNode_Int_3QVal_Int_emitted <= (lizzieLet2_4QNode_Int_3QVal_Int_r ? 2'd0 :
                                                  lizzieLet2_4QNode_Int_3QVal_Int_done);
  
  /* dcon (Ty QTree_Int,
      Dcon QError_Int) : [(lizzieLet2_4QNode_Int_3QVal_Int_1,Go)] > (lizzieLet2_4QNode_Int_3QVal_Int_1QError_Int,QTree_Int) */
  assign lizzieLet2_4QNode_Int_3QVal_Int_1QError_Int_d = QError_Int_dc((& {lizzieLet2_4QNode_Int_3QVal_Int_1_d[0]}), lizzieLet2_4QNode_Int_3QVal_Int_1_d);
  assign {lizzieLet2_4QNode_Int_3QVal_Int_1_r} = {1 {(lizzieLet2_4QNode_Int_3QVal_Int_1QError_Int_r && lizzieLet2_4QNode_Int_3QVal_Int_1QError_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (lizzieLet2_4QNode_Int_3QVal_Int_1QError_Int,QTree_Int) > (lizzieLet8_1_1_argbuf,QTree_Int) */
  QTree_Int_t lizzieLet2_4QNode_Int_3QVal_Int_1QError_Int_bufchan_d;
  logic lizzieLet2_4QNode_Int_3QVal_Int_1QError_Int_bufchan_r;
  assign lizzieLet2_4QNode_Int_3QVal_Int_1QError_Int_r = ((! lizzieLet2_4QNode_Int_3QVal_Int_1QError_Int_bufchan_d[0]) || lizzieLet2_4QNode_Int_3QVal_Int_1QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet2_4QNode_Int_3QVal_Int_1QError_Int_bufchan_d <= {66'd0,
                                                                1'd0};
    else
      if (lizzieLet2_4QNode_Int_3QVal_Int_1QError_Int_r)
        lizzieLet2_4QNode_Int_3QVal_Int_1QError_Int_bufchan_d <= lizzieLet2_4QNode_Int_3QVal_Int_1QError_Int_d;
  QTree_Int_t lizzieLet2_4QNode_Int_3QVal_Int_1QError_Int_bufchan_buf;
  assign lizzieLet2_4QNode_Int_3QVal_Int_1QError_Int_bufchan_r = (! lizzieLet2_4QNode_Int_3QVal_Int_1QError_Int_bufchan_buf[0]);
  assign lizzieLet8_1_1_argbuf_d = (lizzieLet2_4QNode_Int_3QVal_Int_1QError_Int_bufchan_buf[0] ? lizzieLet2_4QNode_Int_3QVal_Int_1QError_Int_bufchan_buf :
                                    lizzieLet2_4QNode_Int_3QVal_Int_1QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet2_4QNode_Int_3QVal_Int_1QError_Int_bufchan_buf <= {66'd0,
                                                                  1'd0};
    else
      if ((lizzieLet8_1_1_argbuf_r && lizzieLet2_4QNode_Int_3QVal_Int_1QError_Int_bufchan_buf[0]))
        lizzieLet2_4QNode_Int_3QVal_Int_1QError_Int_bufchan_buf <= {66'd0,
                                                                    1'd0};
      else if (((! lizzieLet8_1_1_argbuf_r) && (! lizzieLet2_4QNode_Int_3QVal_Int_1QError_Int_bufchan_buf[0])))
        lizzieLet2_4QNode_Int_3QVal_Int_1QError_Int_bufchan_buf <= lizzieLet2_4QNode_Int_3QVal_Int_1QError_Int_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet2_4QNode_Int_3QVal_Int_2,Go) > (lizzieLet2_4QNode_Int_3QVal_Int_2_argbuf,Go) */
  Go_t lizzieLet2_4QNode_Int_3QVal_Int_2_bufchan_d;
  logic lizzieLet2_4QNode_Int_3QVal_Int_2_bufchan_r;
  assign lizzieLet2_4QNode_Int_3QVal_Int_2_r = ((! lizzieLet2_4QNode_Int_3QVal_Int_2_bufchan_d[0]) || lizzieLet2_4QNode_Int_3QVal_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet2_4QNode_Int_3QVal_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet2_4QNode_Int_3QVal_Int_2_r)
        lizzieLet2_4QNode_Int_3QVal_Int_2_bufchan_d <= lizzieLet2_4QNode_Int_3QVal_Int_2_d;
  Go_t lizzieLet2_4QNode_Int_3QVal_Int_2_bufchan_buf;
  assign lizzieLet2_4QNode_Int_3QVal_Int_2_bufchan_r = (! lizzieLet2_4QNode_Int_3QVal_Int_2_bufchan_buf[0]);
  assign lizzieLet2_4QNode_Int_3QVal_Int_2_argbuf_d = (lizzieLet2_4QNode_Int_3QVal_Int_2_bufchan_buf[0] ? lizzieLet2_4QNode_Int_3QVal_Int_2_bufchan_buf :
                                                       lizzieLet2_4QNode_Int_3QVal_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet2_4QNode_Int_3QVal_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet2_4QNode_Int_3QVal_Int_2_argbuf_r && lizzieLet2_4QNode_Int_3QVal_Int_2_bufchan_buf[0]))
        lizzieLet2_4QNode_Int_3QVal_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet2_4QNode_Int_3QVal_Int_2_argbuf_r) && (! lizzieLet2_4QNode_Int_3QVal_Int_2_bufchan_buf[0])))
        lizzieLet2_4QNode_Int_3QVal_Int_2_bufchan_buf <= lizzieLet2_4QNode_Int_3QVal_Int_2_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_CT$wmAdd_Int) : (lizzieLet2_4QNode_Int_4,QTree_Int) (lizzieLet2_5QNode_Int,Pointer_CT$wmAdd_Int) > [(lizzieLet2_4QNode_Int_4QNone_Int,Pointer_CT$wmAdd_Int),
                                                                                                                      (lizzieLet2_4QNode_Int_4QVal_Int,Pointer_CT$wmAdd_Int),
                                                                                                                      (lizzieLet2_4QNode_Int_4QNode_Int,Pointer_CT$wmAdd_Int),
                                                                                                                      (lizzieLet2_4QNode_Int_4QError_Int,Pointer_CT$wmAdd_Int)] */
  logic [3:0] lizzieLet2_5QNode_Int_onehotd;
  always_comb
    if ((lizzieLet2_4QNode_Int_4_d[0] && lizzieLet2_5QNode_Int_d[0]))
      unique case (lizzieLet2_4QNode_Int_4_d[2:1])
        2'd0: lizzieLet2_5QNode_Int_onehotd = 4'd1;
        2'd1: lizzieLet2_5QNode_Int_onehotd = 4'd2;
        2'd2: lizzieLet2_5QNode_Int_onehotd = 4'd4;
        2'd3: lizzieLet2_5QNode_Int_onehotd = 4'd8;
        default: lizzieLet2_5QNode_Int_onehotd = 4'd0;
      endcase
    else lizzieLet2_5QNode_Int_onehotd = 4'd0;
  assign lizzieLet2_4QNode_Int_4QNone_Int_d = {lizzieLet2_5QNode_Int_d[16:1],
                                               lizzieLet2_5QNode_Int_onehotd[0]};
  assign lizzieLet2_4QNode_Int_4QVal_Int_d = {lizzieLet2_5QNode_Int_d[16:1],
                                              lizzieLet2_5QNode_Int_onehotd[1]};
  assign lizzieLet2_4QNode_Int_4QNode_Int_d = {lizzieLet2_5QNode_Int_d[16:1],
                                               lizzieLet2_5QNode_Int_onehotd[2]};
  assign lizzieLet2_4QNode_Int_4QError_Int_d = {lizzieLet2_5QNode_Int_d[16:1],
                                                lizzieLet2_5QNode_Int_onehotd[3]};
  assign lizzieLet2_5QNode_Int_r = (| (lizzieLet2_5QNode_Int_onehotd & {lizzieLet2_4QNode_Int_4QError_Int_r,
                                                                        lizzieLet2_4QNode_Int_4QNode_Int_r,
                                                                        lizzieLet2_4QNode_Int_4QVal_Int_r,
                                                                        lizzieLet2_4QNode_Int_4QNone_Int_r}));
  assign lizzieLet2_4QNode_Int_4_r = lizzieLet2_5QNode_Int_r;
  
  /* buf (Ty Pointer_CT$wmAdd_Int) : (lizzieLet2_4QNode_Int_4QError_Int,Pointer_CT$wmAdd_Int) > (lizzieLet2_4QNode_Int_4QError_Int_1_argbuf,Pointer_CT$wmAdd_Int) */
  Pointer_CT$wmAdd_Int_t lizzieLet2_4QNode_Int_4QError_Int_bufchan_d;
  logic lizzieLet2_4QNode_Int_4QError_Int_bufchan_r;
  assign lizzieLet2_4QNode_Int_4QError_Int_r = ((! lizzieLet2_4QNode_Int_4QError_Int_bufchan_d[0]) || lizzieLet2_4QNode_Int_4QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet2_4QNode_Int_4QError_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet2_4QNode_Int_4QError_Int_r)
        lizzieLet2_4QNode_Int_4QError_Int_bufchan_d <= lizzieLet2_4QNode_Int_4QError_Int_d;
  Pointer_CT$wmAdd_Int_t lizzieLet2_4QNode_Int_4QError_Int_bufchan_buf;
  assign lizzieLet2_4QNode_Int_4QError_Int_bufchan_r = (! lizzieLet2_4QNode_Int_4QError_Int_bufchan_buf[0]);
  assign lizzieLet2_4QNode_Int_4QError_Int_1_argbuf_d = (lizzieLet2_4QNode_Int_4QError_Int_bufchan_buf[0] ? lizzieLet2_4QNode_Int_4QError_Int_bufchan_buf :
                                                         lizzieLet2_4QNode_Int_4QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet2_4QNode_Int_4QError_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet2_4QNode_Int_4QError_Int_1_argbuf_r && lizzieLet2_4QNode_Int_4QError_Int_bufchan_buf[0]))
        lizzieLet2_4QNode_Int_4QError_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet2_4QNode_Int_4QError_Int_1_argbuf_r) && (! lizzieLet2_4QNode_Int_4QError_Int_bufchan_buf[0])))
        lizzieLet2_4QNode_Int_4QError_Int_bufchan_buf <= lizzieLet2_4QNode_Int_4QError_Int_bufchan_d;
  
  /* dcon (Ty CT$wmAdd_Int,
      Dcon Lcall_$wmAdd_Int3) : [(lizzieLet2_4QNode_Int_4QNode_Int,Pointer_CT$wmAdd_Int),
                                 (lizzieLet2_4QNode_Int_6QNode_Int_1,MyDTInt_Int_Int),
                                 (lizzieLet2_4QNode_Int_7QNode_Int,Pointer_QTree_Int),
                                 (t1a8m_destruct,Pointer_QTree_Int),
                                 (lizzieLet2_4QNode_Int_8QNode_Int,Pointer_QTree_Int),
                                 (t2a8n_destruct,Pointer_QTree_Int),
                                 (lizzieLet2_4QNode_Int_9QNode_Int,Pointer_QTree_Int),
                                 (t3a8o_destruct,Pointer_QTree_Int)] > (lizzieLet2_4QNode_Int_4QNode_Int_1lizzieLet2_4QNode_Int_6QNode_Int_1lizzieLet2_4QNode_Int_7QNode_Int_1t1a8m_1lizzieLet2_4QNode_Int_8QNode_Int_1t2a8n_1lizzieLet2_4QNode_Int_9QNode_Int_1t3a8o_1Lcall_$wmAdd_Int3,CT$wmAdd_Int) */
  assign lizzieLet2_4QNode_Int_4QNode_Int_1lizzieLet2_4QNode_Int_6QNode_Int_1lizzieLet2_4QNode_Int_7QNode_Int_1t1a8m_1lizzieLet2_4QNode_Int_8QNode_Int_1t2a8n_1lizzieLet2_4QNode_Int_9QNode_Int_1t3a8o_1Lcall_$wmAdd_Int3_d = Lcall_$wmAdd_Int3_dc((& {lizzieLet2_4QNode_Int_4QNode_Int_d[0],
                                                                                                                                                                                                                                                       lizzieLet2_4QNode_Int_6QNode_Int_1_d[0],
                                                                                                                                                                                                                                                       lizzieLet2_4QNode_Int_7QNode_Int_d[0],
                                                                                                                                                                                                                                                       t1a8m_destruct_d[0],
                                                                                                                                                                                                                                                       lizzieLet2_4QNode_Int_8QNode_Int_d[0],
                                                                                                                                                                                                                                                       t2a8n_destruct_d[0],
                                                                                                                                                                                                                                                       lizzieLet2_4QNode_Int_9QNode_Int_d[0],
                                                                                                                                                                                                                                                       t3a8o_destruct_d[0]}), lizzieLet2_4QNode_Int_4QNode_Int_d, lizzieLet2_4QNode_Int_6QNode_Int_1_d, lizzieLet2_4QNode_Int_7QNode_Int_d, t1a8m_destruct_d, lizzieLet2_4QNode_Int_8QNode_Int_d, t2a8n_destruct_d, lizzieLet2_4QNode_Int_9QNode_Int_d, t3a8o_destruct_d);
  assign {lizzieLet2_4QNode_Int_4QNode_Int_r,
          lizzieLet2_4QNode_Int_6QNode_Int_1_r,
          lizzieLet2_4QNode_Int_7QNode_Int_r,
          t1a8m_destruct_r,
          lizzieLet2_4QNode_Int_8QNode_Int_r,
          t2a8n_destruct_r,
          lizzieLet2_4QNode_Int_9QNode_Int_r,
          t3a8o_destruct_r} = {8 {(lizzieLet2_4QNode_Int_4QNode_Int_1lizzieLet2_4QNode_Int_6QNode_Int_1lizzieLet2_4QNode_Int_7QNode_Int_1t1a8m_1lizzieLet2_4QNode_Int_8QNode_Int_1t2a8n_1lizzieLet2_4QNode_Int_9QNode_Int_1t3a8o_1Lcall_$wmAdd_Int3_r && lizzieLet2_4QNode_Int_4QNode_Int_1lizzieLet2_4QNode_Int_6QNode_Int_1lizzieLet2_4QNode_Int_7QNode_Int_1t1a8m_1lizzieLet2_4QNode_Int_8QNode_Int_1t2a8n_1lizzieLet2_4QNode_Int_9QNode_Int_1t3a8o_1Lcall_$wmAdd_Int3_d[0])}};
  
  /* buf (Ty CT$wmAdd_Int) : (lizzieLet2_4QNode_Int_4QNode_Int_1lizzieLet2_4QNode_Int_6QNode_Int_1lizzieLet2_4QNode_Int_7QNode_Int_1t1a8m_1lizzieLet2_4QNode_Int_8QNode_Int_1t2a8n_1lizzieLet2_4QNode_Int_9QNode_Int_1t3a8o_1Lcall_$wmAdd_Int3,CT$wmAdd_Int) > (lizzieLet9_1_1_argbuf,CT$wmAdd_Int) */
  CT$wmAdd_Int_t lizzieLet2_4QNode_Int_4QNode_Int_1lizzieLet2_4QNode_Int_6QNode_Int_1lizzieLet2_4QNode_Int_7QNode_Int_1t1a8m_1lizzieLet2_4QNode_Int_8QNode_Int_1t2a8n_1lizzieLet2_4QNode_Int_9QNode_Int_1t3a8o_1Lcall_$wmAdd_Int3_bufchan_d;
  logic lizzieLet2_4QNode_Int_4QNode_Int_1lizzieLet2_4QNode_Int_6QNode_Int_1lizzieLet2_4QNode_Int_7QNode_Int_1t1a8m_1lizzieLet2_4QNode_Int_8QNode_Int_1t2a8n_1lizzieLet2_4QNode_Int_9QNode_Int_1t3a8o_1Lcall_$wmAdd_Int3_bufchan_r;
  assign lizzieLet2_4QNode_Int_4QNode_Int_1lizzieLet2_4QNode_Int_6QNode_Int_1lizzieLet2_4QNode_Int_7QNode_Int_1t1a8m_1lizzieLet2_4QNode_Int_8QNode_Int_1t2a8n_1lizzieLet2_4QNode_Int_9QNode_Int_1t3a8o_1Lcall_$wmAdd_Int3_r = ((! lizzieLet2_4QNode_Int_4QNode_Int_1lizzieLet2_4QNode_Int_6QNode_Int_1lizzieLet2_4QNode_Int_7QNode_Int_1t1a8m_1lizzieLet2_4QNode_Int_8QNode_Int_1t2a8n_1lizzieLet2_4QNode_Int_9QNode_Int_1t3a8o_1Lcall_$wmAdd_Int3_bufchan_d[0]) || lizzieLet2_4QNode_Int_4QNode_Int_1lizzieLet2_4QNode_Int_6QNode_Int_1lizzieLet2_4QNode_Int_7QNode_Int_1t1a8m_1lizzieLet2_4QNode_Int_8QNode_Int_1t2a8n_1lizzieLet2_4QNode_Int_9QNode_Int_1t3a8o_1Lcall_$wmAdd_Int3_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet2_4QNode_Int_4QNode_Int_1lizzieLet2_4QNode_Int_6QNode_Int_1lizzieLet2_4QNode_Int_7QNode_Int_1t1a8m_1lizzieLet2_4QNode_Int_8QNode_Int_1t2a8n_1lizzieLet2_4QNode_Int_9QNode_Int_1t3a8o_1Lcall_$wmAdd_Int3_bufchan_d <= {115'd0,
                                                                                                                                                                                                                                     1'd0};
    else
      if (lizzieLet2_4QNode_Int_4QNode_Int_1lizzieLet2_4QNode_Int_6QNode_Int_1lizzieLet2_4QNode_Int_7QNode_Int_1t1a8m_1lizzieLet2_4QNode_Int_8QNode_Int_1t2a8n_1lizzieLet2_4QNode_Int_9QNode_Int_1t3a8o_1Lcall_$wmAdd_Int3_r)
        lizzieLet2_4QNode_Int_4QNode_Int_1lizzieLet2_4QNode_Int_6QNode_Int_1lizzieLet2_4QNode_Int_7QNode_Int_1t1a8m_1lizzieLet2_4QNode_Int_8QNode_Int_1t2a8n_1lizzieLet2_4QNode_Int_9QNode_Int_1t3a8o_1Lcall_$wmAdd_Int3_bufchan_d <= lizzieLet2_4QNode_Int_4QNode_Int_1lizzieLet2_4QNode_Int_6QNode_Int_1lizzieLet2_4QNode_Int_7QNode_Int_1t1a8m_1lizzieLet2_4QNode_Int_8QNode_Int_1t2a8n_1lizzieLet2_4QNode_Int_9QNode_Int_1t3a8o_1Lcall_$wmAdd_Int3_d;
  CT$wmAdd_Int_t lizzieLet2_4QNode_Int_4QNode_Int_1lizzieLet2_4QNode_Int_6QNode_Int_1lizzieLet2_4QNode_Int_7QNode_Int_1t1a8m_1lizzieLet2_4QNode_Int_8QNode_Int_1t2a8n_1lizzieLet2_4QNode_Int_9QNode_Int_1t3a8o_1Lcall_$wmAdd_Int3_bufchan_buf;
  assign lizzieLet2_4QNode_Int_4QNode_Int_1lizzieLet2_4QNode_Int_6QNode_Int_1lizzieLet2_4QNode_Int_7QNode_Int_1t1a8m_1lizzieLet2_4QNode_Int_8QNode_Int_1t2a8n_1lizzieLet2_4QNode_Int_9QNode_Int_1t3a8o_1Lcall_$wmAdd_Int3_bufchan_r = (! lizzieLet2_4QNode_Int_4QNode_Int_1lizzieLet2_4QNode_Int_6QNode_Int_1lizzieLet2_4QNode_Int_7QNode_Int_1t1a8m_1lizzieLet2_4QNode_Int_8QNode_Int_1t2a8n_1lizzieLet2_4QNode_Int_9QNode_Int_1t3a8o_1Lcall_$wmAdd_Int3_bufchan_buf[0]);
  assign lizzieLet9_1_1_argbuf_d = (lizzieLet2_4QNode_Int_4QNode_Int_1lizzieLet2_4QNode_Int_6QNode_Int_1lizzieLet2_4QNode_Int_7QNode_Int_1t1a8m_1lizzieLet2_4QNode_Int_8QNode_Int_1t2a8n_1lizzieLet2_4QNode_Int_9QNode_Int_1t3a8o_1Lcall_$wmAdd_Int3_bufchan_buf[0] ? lizzieLet2_4QNode_Int_4QNode_Int_1lizzieLet2_4QNode_Int_6QNode_Int_1lizzieLet2_4QNode_Int_7QNode_Int_1t1a8m_1lizzieLet2_4QNode_Int_8QNode_Int_1t2a8n_1lizzieLet2_4QNode_Int_9QNode_Int_1t3a8o_1Lcall_$wmAdd_Int3_bufchan_buf :
                                    lizzieLet2_4QNode_Int_4QNode_Int_1lizzieLet2_4QNode_Int_6QNode_Int_1lizzieLet2_4QNode_Int_7QNode_Int_1t1a8m_1lizzieLet2_4QNode_Int_8QNode_Int_1t2a8n_1lizzieLet2_4QNode_Int_9QNode_Int_1t3a8o_1Lcall_$wmAdd_Int3_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet2_4QNode_Int_4QNode_Int_1lizzieLet2_4QNode_Int_6QNode_Int_1lizzieLet2_4QNode_Int_7QNode_Int_1t1a8m_1lizzieLet2_4QNode_Int_8QNode_Int_1t2a8n_1lizzieLet2_4QNode_Int_9QNode_Int_1t3a8o_1Lcall_$wmAdd_Int3_bufchan_buf <= {115'd0,
                                                                                                                                                                                                                                       1'd0};
    else
      if ((lizzieLet9_1_1_argbuf_r && lizzieLet2_4QNode_Int_4QNode_Int_1lizzieLet2_4QNode_Int_6QNode_Int_1lizzieLet2_4QNode_Int_7QNode_Int_1t1a8m_1lizzieLet2_4QNode_Int_8QNode_Int_1t2a8n_1lizzieLet2_4QNode_Int_9QNode_Int_1t3a8o_1Lcall_$wmAdd_Int3_bufchan_buf[0]))
        lizzieLet2_4QNode_Int_4QNode_Int_1lizzieLet2_4QNode_Int_6QNode_Int_1lizzieLet2_4QNode_Int_7QNode_Int_1t1a8m_1lizzieLet2_4QNode_Int_8QNode_Int_1t2a8n_1lizzieLet2_4QNode_Int_9QNode_Int_1t3a8o_1Lcall_$wmAdd_Int3_bufchan_buf <= {115'd0,
                                                                                                                                                                                                                                         1'd0};
      else if (((! lizzieLet9_1_1_argbuf_r) && (! lizzieLet2_4QNode_Int_4QNode_Int_1lizzieLet2_4QNode_Int_6QNode_Int_1lizzieLet2_4QNode_Int_7QNode_Int_1t1a8m_1lizzieLet2_4QNode_Int_8QNode_Int_1t2a8n_1lizzieLet2_4QNode_Int_9QNode_Int_1t3a8o_1Lcall_$wmAdd_Int3_bufchan_buf[0])))
        lizzieLet2_4QNode_Int_4QNode_Int_1lizzieLet2_4QNode_Int_6QNode_Int_1lizzieLet2_4QNode_Int_7QNode_Int_1t1a8m_1lizzieLet2_4QNode_Int_8QNode_Int_1t2a8n_1lizzieLet2_4QNode_Int_9QNode_Int_1t3a8o_1Lcall_$wmAdd_Int3_bufchan_buf <= lizzieLet2_4QNode_Int_4QNode_Int_1lizzieLet2_4QNode_Int_6QNode_Int_1lizzieLet2_4QNode_Int_7QNode_Int_1t1a8m_1lizzieLet2_4QNode_Int_8QNode_Int_1t2a8n_1lizzieLet2_4QNode_Int_9QNode_Int_1t3a8o_1Lcall_$wmAdd_Int3_bufchan_d;
  
  /* buf (Ty Pointer_CT$wmAdd_Int) : (lizzieLet2_4QNode_Int_4QNone_Int,Pointer_CT$wmAdd_Int) > (lizzieLet2_4QNode_Int_4QNone_Int_1_argbuf,Pointer_CT$wmAdd_Int) */
  Pointer_CT$wmAdd_Int_t lizzieLet2_4QNode_Int_4QNone_Int_bufchan_d;
  logic lizzieLet2_4QNode_Int_4QNone_Int_bufchan_r;
  assign lizzieLet2_4QNode_Int_4QNone_Int_r = ((! lizzieLet2_4QNode_Int_4QNone_Int_bufchan_d[0]) || lizzieLet2_4QNode_Int_4QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet2_4QNode_Int_4QNone_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet2_4QNode_Int_4QNone_Int_r)
        lizzieLet2_4QNode_Int_4QNone_Int_bufchan_d <= lizzieLet2_4QNode_Int_4QNone_Int_d;
  Pointer_CT$wmAdd_Int_t lizzieLet2_4QNode_Int_4QNone_Int_bufchan_buf;
  assign lizzieLet2_4QNode_Int_4QNone_Int_bufchan_r = (! lizzieLet2_4QNode_Int_4QNone_Int_bufchan_buf[0]);
  assign lizzieLet2_4QNode_Int_4QNone_Int_1_argbuf_d = (lizzieLet2_4QNode_Int_4QNone_Int_bufchan_buf[0] ? lizzieLet2_4QNode_Int_4QNone_Int_bufchan_buf :
                                                        lizzieLet2_4QNode_Int_4QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet2_4QNode_Int_4QNone_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet2_4QNode_Int_4QNone_Int_1_argbuf_r && lizzieLet2_4QNode_Int_4QNone_Int_bufchan_buf[0]))
        lizzieLet2_4QNode_Int_4QNone_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet2_4QNode_Int_4QNone_Int_1_argbuf_r) && (! lizzieLet2_4QNode_Int_4QNone_Int_bufchan_buf[0])))
        lizzieLet2_4QNode_Int_4QNone_Int_bufchan_buf <= lizzieLet2_4QNode_Int_4QNone_Int_bufchan_d;
  
  /* buf (Ty Pointer_CT$wmAdd_Int) : (lizzieLet2_4QNode_Int_4QVal_Int,Pointer_CT$wmAdd_Int) > (lizzieLet2_4QNode_Int_4QVal_Int_1_argbuf,Pointer_CT$wmAdd_Int) */
  Pointer_CT$wmAdd_Int_t lizzieLet2_4QNode_Int_4QVal_Int_bufchan_d;
  logic lizzieLet2_4QNode_Int_4QVal_Int_bufchan_r;
  assign lizzieLet2_4QNode_Int_4QVal_Int_r = ((! lizzieLet2_4QNode_Int_4QVal_Int_bufchan_d[0]) || lizzieLet2_4QNode_Int_4QVal_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet2_4QNode_Int_4QVal_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet2_4QNode_Int_4QVal_Int_r)
        lizzieLet2_4QNode_Int_4QVal_Int_bufchan_d <= lizzieLet2_4QNode_Int_4QVal_Int_d;
  Pointer_CT$wmAdd_Int_t lizzieLet2_4QNode_Int_4QVal_Int_bufchan_buf;
  assign lizzieLet2_4QNode_Int_4QVal_Int_bufchan_r = (! lizzieLet2_4QNode_Int_4QVal_Int_bufchan_buf[0]);
  assign lizzieLet2_4QNode_Int_4QVal_Int_1_argbuf_d = (lizzieLet2_4QNode_Int_4QVal_Int_bufchan_buf[0] ? lizzieLet2_4QNode_Int_4QVal_Int_bufchan_buf :
                                                       lizzieLet2_4QNode_Int_4QVal_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet2_4QNode_Int_4QVal_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet2_4QNode_Int_4QVal_Int_1_argbuf_r && lizzieLet2_4QNode_Int_4QVal_Int_bufchan_buf[0]))
        lizzieLet2_4QNode_Int_4QVal_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet2_4QNode_Int_4QVal_Int_1_argbuf_r) && (! lizzieLet2_4QNode_Int_4QVal_Int_bufchan_buf[0])))
        lizzieLet2_4QNode_Int_4QVal_Int_bufchan_buf <= lizzieLet2_4QNode_Int_4QVal_Int_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_QTree_Int) : (lizzieLet2_4QNode_Int_5,QTree_Int) (lizzieLet2_6QNode_Int,Pointer_QTree_Int) > [(lizzieLet2_4QNode_Int_5QNone_Int,Pointer_QTree_Int),
                                                                                                                (_35,Pointer_QTree_Int),
                                                                                                                (_34,Pointer_QTree_Int),
                                                                                                                (_33,Pointer_QTree_Int)] */
  logic [3:0] lizzieLet2_6QNode_Int_onehotd;
  always_comb
    if ((lizzieLet2_4QNode_Int_5_d[0] && lizzieLet2_6QNode_Int_d[0]))
      unique case (lizzieLet2_4QNode_Int_5_d[2:1])
        2'd0: lizzieLet2_6QNode_Int_onehotd = 4'd1;
        2'd1: lizzieLet2_6QNode_Int_onehotd = 4'd2;
        2'd2: lizzieLet2_6QNode_Int_onehotd = 4'd4;
        2'd3: lizzieLet2_6QNode_Int_onehotd = 4'd8;
        default: lizzieLet2_6QNode_Int_onehotd = 4'd0;
      endcase
    else lizzieLet2_6QNode_Int_onehotd = 4'd0;
  assign lizzieLet2_4QNode_Int_5QNone_Int_d = {lizzieLet2_6QNode_Int_d[16:1],
                                               lizzieLet2_6QNode_Int_onehotd[0]};
  assign _35_d = {lizzieLet2_6QNode_Int_d[16:1],
                  lizzieLet2_6QNode_Int_onehotd[1]};
  assign _34_d = {lizzieLet2_6QNode_Int_d[16:1],
                  lizzieLet2_6QNode_Int_onehotd[2]};
  assign _33_d = {lizzieLet2_6QNode_Int_d[16:1],
                  lizzieLet2_6QNode_Int_onehotd[3]};
  assign lizzieLet2_6QNode_Int_r = (| (lizzieLet2_6QNode_Int_onehotd & {_33_r,
                                                                        _34_r,
                                                                        _35_r,
                                                                        lizzieLet2_4QNode_Int_5QNone_Int_r}));
  assign lizzieLet2_4QNode_Int_5_r = lizzieLet2_6QNode_Int_r;
  
  /* buf (Ty Pointer_QTree_Int) : (lizzieLet2_4QNode_Int_5QNone_Int,Pointer_QTree_Int) > (lizzieLet2_4QNode_Int_5QNone_Int_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t lizzieLet2_4QNode_Int_5QNone_Int_bufchan_d;
  logic lizzieLet2_4QNode_Int_5QNone_Int_bufchan_r;
  assign lizzieLet2_4QNode_Int_5QNone_Int_r = ((! lizzieLet2_4QNode_Int_5QNone_Int_bufchan_d[0]) || lizzieLet2_4QNode_Int_5QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet2_4QNode_Int_5QNone_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet2_4QNode_Int_5QNone_Int_r)
        lizzieLet2_4QNode_Int_5QNone_Int_bufchan_d <= lizzieLet2_4QNode_Int_5QNone_Int_d;
  Pointer_QTree_Int_t lizzieLet2_4QNode_Int_5QNone_Int_bufchan_buf;
  assign lizzieLet2_4QNode_Int_5QNone_Int_bufchan_r = (! lizzieLet2_4QNode_Int_5QNone_Int_bufchan_buf[0]);
  assign lizzieLet2_4QNode_Int_5QNone_Int_1_argbuf_d = (lizzieLet2_4QNode_Int_5QNone_Int_bufchan_buf[0] ? lizzieLet2_4QNode_Int_5QNone_Int_bufchan_buf :
                                                        lizzieLet2_4QNode_Int_5QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet2_4QNode_Int_5QNone_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet2_4QNode_Int_5QNone_Int_1_argbuf_r && lizzieLet2_4QNode_Int_5QNone_Int_bufchan_buf[0]))
        lizzieLet2_4QNode_Int_5QNone_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet2_4QNode_Int_5QNone_Int_1_argbuf_r) && (! lizzieLet2_4QNode_Int_5QNone_Int_bufchan_buf[0])))
        lizzieLet2_4QNode_Int_5QNone_Int_bufchan_buf <= lizzieLet2_4QNode_Int_5QNone_Int_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty MyDTInt_Int_Int) : (lizzieLet2_4QNode_Int_6,QTree_Int) (lizzieLet2_8QNode_Int,MyDTInt_Int_Int) > [(_32,MyDTInt_Int_Int),
                                                                                                            (_31,MyDTInt_Int_Int),
                                                                                                            (lizzieLet2_4QNode_Int_6QNode_Int,MyDTInt_Int_Int),
                                                                                                            (_30,MyDTInt_Int_Int)] */
  logic [3:0] lizzieLet2_8QNode_Int_onehotd;
  always_comb
    if ((lizzieLet2_4QNode_Int_6_d[0] && lizzieLet2_8QNode_Int_d[0]))
      unique case (lizzieLet2_4QNode_Int_6_d[2:1])
        2'd0: lizzieLet2_8QNode_Int_onehotd = 4'd1;
        2'd1: lizzieLet2_8QNode_Int_onehotd = 4'd2;
        2'd2: lizzieLet2_8QNode_Int_onehotd = 4'd4;
        2'd3: lizzieLet2_8QNode_Int_onehotd = 4'd8;
        default: lizzieLet2_8QNode_Int_onehotd = 4'd0;
      endcase
    else lizzieLet2_8QNode_Int_onehotd = 4'd0;
  assign _32_d = lizzieLet2_8QNode_Int_onehotd[0];
  assign _31_d = lizzieLet2_8QNode_Int_onehotd[1];
  assign lizzieLet2_4QNode_Int_6QNode_Int_d = lizzieLet2_8QNode_Int_onehotd[2];
  assign _30_d = lizzieLet2_8QNode_Int_onehotd[3];
  assign lizzieLet2_8QNode_Int_r = (| (lizzieLet2_8QNode_Int_onehotd & {_30_r,
                                                                        lizzieLet2_4QNode_Int_6QNode_Int_r,
                                                                        _31_r,
                                                                        _32_r}));
  assign lizzieLet2_4QNode_Int_6_r = lizzieLet2_8QNode_Int_r;
  
  /* fork (Ty MyDTInt_Int_Int) : (lizzieLet2_4QNode_Int_6QNode_Int,MyDTInt_Int_Int) > [(lizzieLet2_4QNode_Int_6QNode_Int_1,MyDTInt_Int_Int),
                                                                                  (lizzieLet2_4QNode_Int_6QNode_Int_2,MyDTInt_Int_Int)] */
  logic [1:0] lizzieLet2_4QNode_Int_6QNode_Int_emitted;
  logic [1:0] lizzieLet2_4QNode_Int_6QNode_Int_done;
  assign lizzieLet2_4QNode_Int_6QNode_Int_1_d = (lizzieLet2_4QNode_Int_6QNode_Int_d[0] && (! lizzieLet2_4QNode_Int_6QNode_Int_emitted[0]));
  assign lizzieLet2_4QNode_Int_6QNode_Int_2_d = (lizzieLet2_4QNode_Int_6QNode_Int_d[0] && (! lizzieLet2_4QNode_Int_6QNode_Int_emitted[1]));
  assign lizzieLet2_4QNode_Int_6QNode_Int_done = (lizzieLet2_4QNode_Int_6QNode_Int_emitted | ({lizzieLet2_4QNode_Int_6QNode_Int_2_d[0],
                                                                                               lizzieLet2_4QNode_Int_6QNode_Int_1_d[0]} & {lizzieLet2_4QNode_Int_6QNode_Int_2_r,
                                                                                                                                           lizzieLet2_4QNode_Int_6QNode_Int_1_r}));
  assign lizzieLet2_4QNode_Int_6QNode_Int_r = (& lizzieLet2_4QNode_Int_6QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet2_4QNode_Int_6QNode_Int_emitted <= 2'd0;
    else
      lizzieLet2_4QNode_Int_6QNode_Int_emitted <= (lizzieLet2_4QNode_Int_6QNode_Int_r ? 2'd0 :
                                                   lizzieLet2_4QNode_Int_6QNode_Int_done);
  
  /* buf (Ty MyDTInt_Int_Int) : (lizzieLet2_4QNode_Int_6QNode_Int_2,MyDTInt_Int_Int) > (lizzieLet2_4QNode_Int_6QNode_Int_2_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t lizzieLet2_4QNode_Int_6QNode_Int_2_bufchan_d;
  logic lizzieLet2_4QNode_Int_6QNode_Int_2_bufchan_r;
  assign lizzieLet2_4QNode_Int_6QNode_Int_2_r = ((! lizzieLet2_4QNode_Int_6QNode_Int_2_bufchan_d[0]) || lizzieLet2_4QNode_Int_6QNode_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet2_4QNode_Int_6QNode_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet2_4QNode_Int_6QNode_Int_2_r)
        lizzieLet2_4QNode_Int_6QNode_Int_2_bufchan_d <= lizzieLet2_4QNode_Int_6QNode_Int_2_d;
  MyDTInt_Int_Int_t lizzieLet2_4QNode_Int_6QNode_Int_2_bufchan_buf;
  assign lizzieLet2_4QNode_Int_6QNode_Int_2_bufchan_r = (! lizzieLet2_4QNode_Int_6QNode_Int_2_bufchan_buf[0]);
  assign lizzieLet2_4QNode_Int_6QNode_Int_2_argbuf_d = (lizzieLet2_4QNode_Int_6QNode_Int_2_bufchan_buf[0] ? lizzieLet2_4QNode_Int_6QNode_Int_2_bufchan_buf :
                                                        lizzieLet2_4QNode_Int_6QNode_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet2_4QNode_Int_6QNode_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet2_4QNode_Int_6QNode_Int_2_argbuf_r && lizzieLet2_4QNode_Int_6QNode_Int_2_bufchan_buf[0]))
        lizzieLet2_4QNode_Int_6QNode_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet2_4QNode_Int_6QNode_Int_2_argbuf_r) && (! lizzieLet2_4QNode_Int_6QNode_Int_2_bufchan_buf[0])))
        lizzieLet2_4QNode_Int_6QNode_Int_2_bufchan_buf <= lizzieLet2_4QNode_Int_6QNode_Int_2_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_QTree_Int) : (lizzieLet2_4QNode_Int_7,QTree_Int) (q1a8h_destruct,Pointer_QTree_Int) > [(_29,Pointer_QTree_Int),
                                                                                                         (_28,Pointer_QTree_Int),
                                                                                                         (lizzieLet2_4QNode_Int_7QNode_Int,Pointer_QTree_Int),
                                                                                                         (_27,Pointer_QTree_Int)] */
  logic [3:0] q1a8h_destruct_onehotd;
  always_comb
    if ((lizzieLet2_4QNode_Int_7_d[0] && q1a8h_destruct_d[0]))
      unique case (lizzieLet2_4QNode_Int_7_d[2:1])
        2'd0: q1a8h_destruct_onehotd = 4'd1;
        2'd1: q1a8h_destruct_onehotd = 4'd2;
        2'd2: q1a8h_destruct_onehotd = 4'd4;
        2'd3: q1a8h_destruct_onehotd = 4'd8;
        default: q1a8h_destruct_onehotd = 4'd0;
      endcase
    else q1a8h_destruct_onehotd = 4'd0;
  assign _29_d = {q1a8h_destruct_d[16:1], q1a8h_destruct_onehotd[0]};
  assign _28_d = {q1a8h_destruct_d[16:1], q1a8h_destruct_onehotd[1]};
  assign lizzieLet2_4QNode_Int_7QNode_Int_d = {q1a8h_destruct_d[16:1],
                                               q1a8h_destruct_onehotd[2]};
  assign _27_d = {q1a8h_destruct_d[16:1], q1a8h_destruct_onehotd[3]};
  assign q1a8h_destruct_r = (| (q1a8h_destruct_onehotd & {_27_r,
                                                          lizzieLet2_4QNode_Int_7QNode_Int_r,
                                                          _28_r,
                                                          _29_r}));
  assign lizzieLet2_4QNode_Int_7_r = q1a8h_destruct_r;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_QTree_Int) : (lizzieLet2_4QNode_Int_8,QTree_Int) (q2a8i_destruct,Pointer_QTree_Int) > [(_26,Pointer_QTree_Int),
                                                                                                         (_25,Pointer_QTree_Int),
                                                                                                         (lizzieLet2_4QNode_Int_8QNode_Int,Pointer_QTree_Int),
                                                                                                         (_24,Pointer_QTree_Int)] */
  logic [3:0] q2a8i_destruct_onehotd;
  always_comb
    if ((lizzieLet2_4QNode_Int_8_d[0] && q2a8i_destruct_d[0]))
      unique case (lizzieLet2_4QNode_Int_8_d[2:1])
        2'd0: q2a8i_destruct_onehotd = 4'd1;
        2'd1: q2a8i_destruct_onehotd = 4'd2;
        2'd2: q2a8i_destruct_onehotd = 4'd4;
        2'd3: q2a8i_destruct_onehotd = 4'd8;
        default: q2a8i_destruct_onehotd = 4'd0;
      endcase
    else q2a8i_destruct_onehotd = 4'd0;
  assign _26_d = {q2a8i_destruct_d[16:1], q2a8i_destruct_onehotd[0]};
  assign _25_d = {q2a8i_destruct_d[16:1], q2a8i_destruct_onehotd[1]};
  assign lizzieLet2_4QNode_Int_8QNode_Int_d = {q2a8i_destruct_d[16:1],
                                               q2a8i_destruct_onehotd[2]};
  assign _24_d = {q2a8i_destruct_d[16:1], q2a8i_destruct_onehotd[3]};
  assign q2a8i_destruct_r = (| (q2a8i_destruct_onehotd & {_24_r,
                                                          lizzieLet2_4QNode_Int_8QNode_Int_r,
                                                          _25_r,
                                                          _26_r}));
  assign lizzieLet2_4QNode_Int_8_r = q2a8i_destruct_r;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_QTree_Int) : (lizzieLet2_4QNode_Int_9,QTree_Int) (q3a8j_destruct,Pointer_QTree_Int) > [(_23,Pointer_QTree_Int),
                                                                                                         (_22,Pointer_QTree_Int),
                                                                                                         (lizzieLet2_4QNode_Int_9QNode_Int,Pointer_QTree_Int),
                                                                                                         (_21,Pointer_QTree_Int)] */
  logic [3:0] q3a8j_destruct_onehotd;
  always_comb
    if ((lizzieLet2_4QNode_Int_9_d[0] && q3a8j_destruct_d[0]))
      unique case (lizzieLet2_4QNode_Int_9_d[2:1])
        2'd0: q3a8j_destruct_onehotd = 4'd1;
        2'd1: q3a8j_destruct_onehotd = 4'd2;
        2'd2: q3a8j_destruct_onehotd = 4'd4;
        2'd3: q3a8j_destruct_onehotd = 4'd8;
        default: q3a8j_destruct_onehotd = 4'd0;
      endcase
    else q3a8j_destruct_onehotd = 4'd0;
  assign _23_d = {q3a8j_destruct_d[16:1], q3a8j_destruct_onehotd[0]};
  assign _22_d = {q3a8j_destruct_d[16:1], q3a8j_destruct_onehotd[1]};
  assign lizzieLet2_4QNode_Int_9QNode_Int_d = {q3a8j_destruct_d[16:1],
                                               q3a8j_destruct_onehotd[2]};
  assign _21_d = {q3a8j_destruct_d[16:1], q3a8j_destruct_onehotd[3]};
  assign q3a8j_destruct_r = (| (q3a8j_destruct_onehotd & {_21_r,
                                                          lizzieLet2_4QNode_Int_9QNode_Int_r,
                                                          _22_r,
                                                          _23_r}));
  assign lizzieLet2_4QNode_Int_9_r = q3a8j_destruct_r;
  
  /* fork (Ty QTree_Int) : (lizzieLet2_4QVal_Int,QTree_Int) > [(lizzieLet2_4QVal_Int_1,QTree_Int),
                                                          (lizzieLet2_4QVal_Int_2,QTree_Int),
                                                          (lizzieLet2_4QVal_Int_3,QTree_Int),
                                                          (lizzieLet2_4QVal_Int_4,QTree_Int),
                                                          (lizzieLet2_4QVal_Int_5,QTree_Int),
                                                          (lizzieLet2_4QVal_Int_6,QTree_Int),
                                                          (lizzieLet2_4QVal_Int_7,QTree_Int)] */
  logic [6:0] lizzieLet2_4QVal_Int_emitted;
  logic [6:0] lizzieLet2_4QVal_Int_done;
  assign lizzieLet2_4QVal_Int_1_d = {lizzieLet2_4QVal_Int_d[66:1],
                                     (lizzieLet2_4QVal_Int_d[0] && (! lizzieLet2_4QVal_Int_emitted[0]))};
  assign lizzieLet2_4QVal_Int_2_d = {lizzieLet2_4QVal_Int_d[66:1],
                                     (lizzieLet2_4QVal_Int_d[0] && (! lizzieLet2_4QVal_Int_emitted[1]))};
  assign lizzieLet2_4QVal_Int_3_d = {lizzieLet2_4QVal_Int_d[66:1],
                                     (lizzieLet2_4QVal_Int_d[0] && (! lizzieLet2_4QVal_Int_emitted[2]))};
  assign lizzieLet2_4QVal_Int_4_d = {lizzieLet2_4QVal_Int_d[66:1],
                                     (lizzieLet2_4QVal_Int_d[0] && (! lizzieLet2_4QVal_Int_emitted[3]))};
  assign lizzieLet2_4QVal_Int_5_d = {lizzieLet2_4QVal_Int_d[66:1],
                                     (lizzieLet2_4QVal_Int_d[0] && (! lizzieLet2_4QVal_Int_emitted[4]))};
  assign lizzieLet2_4QVal_Int_6_d = {lizzieLet2_4QVal_Int_d[66:1],
                                     (lizzieLet2_4QVal_Int_d[0] && (! lizzieLet2_4QVal_Int_emitted[5]))};
  assign lizzieLet2_4QVal_Int_7_d = {lizzieLet2_4QVal_Int_d[66:1],
                                     (lizzieLet2_4QVal_Int_d[0] && (! lizzieLet2_4QVal_Int_emitted[6]))};
  assign lizzieLet2_4QVal_Int_done = (lizzieLet2_4QVal_Int_emitted | ({lizzieLet2_4QVal_Int_7_d[0],
                                                                       lizzieLet2_4QVal_Int_6_d[0],
                                                                       lizzieLet2_4QVal_Int_5_d[0],
                                                                       lizzieLet2_4QVal_Int_4_d[0],
                                                                       lizzieLet2_4QVal_Int_3_d[0],
                                                                       lizzieLet2_4QVal_Int_2_d[0],
                                                                       lizzieLet2_4QVal_Int_1_d[0]} & {lizzieLet2_4QVal_Int_7_r,
                                                                                                       lizzieLet2_4QVal_Int_6_r,
                                                                                                       lizzieLet2_4QVal_Int_5_r,
                                                                                                       lizzieLet2_4QVal_Int_4_r,
                                                                                                       lizzieLet2_4QVal_Int_3_r,
                                                                                                       lizzieLet2_4QVal_Int_2_r,
                                                                                                       lizzieLet2_4QVal_Int_1_r}));
  assign lizzieLet2_4QVal_Int_r = (& lizzieLet2_4QVal_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet2_4QVal_Int_emitted <= 7'd0;
    else
      lizzieLet2_4QVal_Int_emitted <= (lizzieLet2_4QVal_Int_r ? 7'd0 :
                                       lizzieLet2_4QVal_Int_done);
  
  /* destruct (Ty QTree_Int,
          Dcon QVal_Int) : (lizzieLet2_4QVal_Int_1QVal_Int,QTree_Int) > [(va8c_destruct,Int)] */
  assign va8c_destruct_d = {lizzieLet2_4QVal_Int_1QVal_Int_d[34:3],
                            lizzieLet2_4QVal_Int_1QVal_Int_d[0]};
  assign lizzieLet2_4QVal_Int_1QVal_Int_r = va8c_destruct_r;
  
  /* demux (Ty QTree_Int,
       Ty QTree_Int) : (lizzieLet2_4QVal_Int_2,QTree_Int) (lizzieLet2_4QVal_Int_1,QTree_Int) > [(_20,QTree_Int),
                                                                                                (lizzieLet2_4QVal_Int_1QVal_Int,QTree_Int),
                                                                                                (_19,QTree_Int),
                                                                                                (_18,QTree_Int)] */
  logic [3:0] lizzieLet2_4QVal_Int_1_onehotd;
  always_comb
    if ((lizzieLet2_4QVal_Int_2_d[0] && lizzieLet2_4QVal_Int_1_d[0]))
      unique case (lizzieLet2_4QVal_Int_2_d[2:1])
        2'd0: lizzieLet2_4QVal_Int_1_onehotd = 4'd1;
        2'd1: lizzieLet2_4QVal_Int_1_onehotd = 4'd2;
        2'd2: lizzieLet2_4QVal_Int_1_onehotd = 4'd4;
        2'd3: lizzieLet2_4QVal_Int_1_onehotd = 4'd8;
        default: lizzieLet2_4QVal_Int_1_onehotd = 4'd0;
      endcase
    else lizzieLet2_4QVal_Int_1_onehotd = 4'd0;
  assign _20_d = {lizzieLet2_4QVal_Int_1_d[66:1],
                  lizzieLet2_4QVal_Int_1_onehotd[0]};
  assign lizzieLet2_4QVal_Int_1QVal_Int_d = {lizzieLet2_4QVal_Int_1_d[66:1],
                                             lizzieLet2_4QVal_Int_1_onehotd[1]};
  assign _19_d = {lizzieLet2_4QVal_Int_1_d[66:1],
                  lizzieLet2_4QVal_Int_1_onehotd[2]};
  assign _18_d = {lizzieLet2_4QVal_Int_1_d[66:1],
                  lizzieLet2_4QVal_Int_1_onehotd[3]};
  assign lizzieLet2_4QVal_Int_1_r = (| (lizzieLet2_4QVal_Int_1_onehotd & {_18_r,
                                                                          _19_r,
                                                                          lizzieLet2_4QVal_Int_1QVal_Int_r,
                                                                          _20_r}));
  assign lizzieLet2_4QVal_Int_2_r = lizzieLet2_4QVal_Int_1_r;
  
  /* demux (Ty QTree_Int,
       Ty Go) : (lizzieLet2_4QVal_Int_3,QTree_Int) (lizzieLet2_3QVal_Int,Go) > [(lizzieLet2_4QVal_Int_3QNone_Int,Go),
                                                                                (lizzieLet2_4QVal_Int_3QVal_Int,Go),
                                                                                (lizzieLet2_4QVal_Int_3QNode_Int,Go),
                                                                                (lizzieLet2_4QVal_Int_3QError_Int,Go)] */
  logic [3:0] lizzieLet2_3QVal_Int_onehotd;
  always_comb
    if ((lizzieLet2_4QVal_Int_3_d[0] && lizzieLet2_3QVal_Int_d[0]))
      unique case (lizzieLet2_4QVal_Int_3_d[2:1])
        2'd0: lizzieLet2_3QVal_Int_onehotd = 4'd1;
        2'd1: lizzieLet2_3QVal_Int_onehotd = 4'd2;
        2'd2: lizzieLet2_3QVal_Int_onehotd = 4'd4;
        2'd3: lizzieLet2_3QVal_Int_onehotd = 4'd8;
        default: lizzieLet2_3QVal_Int_onehotd = 4'd0;
      endcase
    else lizzieLet2_3QVal_Int_onehotd = 4'd0;
  assign lizzieLet2_4QVal_Int_3QNone_Int_d = lizzieLet2_3QVal_Int_onehotd[0];
  assign lizzieLet2_4QVal_Int_3QVal_Int_d = lizzieLet2_3QVal_Int_onehotd[1];
  assign lizzieLet2_4QVal_Int_3QNode_Int_d = lizzieLet2_3QVal_Int_onehotd[2];
  assign lizzieLet2_4QVal_Int_3QError_Int_d = lizzieLet2_3QVal_Int_onehotd[3];
  assign lizzieLet2_3QVal_Int_r = (| (lizzieLet2_3QVal_Int_onehotd & {lizzieLet2_4QVal_Int_3QError_Int_r,
                                                                      lizzieLet2_4QVal_Int_3QNode_Int_r,
                                                                      lizzieLet2_4QVal_Int_3QVal_Int_r,
                                                                      lizzieLet2_4QVal_Int_3QNone_Int_r}));
  assign lizzieLet2_4QVal_Int_3_r = lizzieLet2_3QVal_Int_r;
  
  /* fork (Ty Go) : (lizzieLet2_4QVal_Int_3QError_Int,Go) > [(lizzieLet2_4QVal_Int_3QError_Int_1,Go),
                                                        (lizzieLet2_4QVal_Int_3QError_Int_2,Go)] */
  logic [1:0] lizzieLet2_4QVal_Int_3QError_Int_emitted;
  logic [1:0] lizzieLet2_4QVal_Int_3QError_Int_done;
  assign lizzieLet2_4QVal_Int_3QError_Int_1_d = (lizzieLet2_4QVal_Int_3QError_Int_d[0] && (! lizzieLet2_4QVal_Int_3QError_Int_emitted[0]));
  assign lizzieLet2_4QVal_Int_3QError_Int_2_d = (lizzieLet2_4QVal_Int_3QError_Int_d[0] && (! lizzieLet2_4QVal_Int_3QError_Int_emitted[1]));
  assign lizzieLet2_4QVal_Int_3QError_Int_done = (lizzieLet2_4QVal_Int_3QError_Int_emitted | ({lizzieLet2_4QVal_Int_3QError_Int_2_d[0],
                                                                                               lizzieLet2_4QVal_Int_3QError_Int_1_d[0]} & {lizzieLet2_4QVal_Int_3QError_Int_2_r,
                                                                                                                                           lizzieLet2_4QVal_Int_3QError_Int_1_r}));
  assign lizzieLet2_4QVal_Int_3QError_Int_r = (& lizzieLet2_4QVal_Int_3QError_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet2_4QVal_Int_3QError_Int_emitted <= 2'd0;
    else
      lizzieLet2_4QVal_Int_3QError_Int_emitted <= (lizzieLet2_4QVal_Int_3QError_Int_r ? 2'd0 :
                                                   lizzieLet2_4QVal_Int_3QError_Int_done);
  
  /* dcon (Ty QTree_Int,
      Dcon QError_Int) : [(lizzieLet2_4QVal_Int_3QError_Int_1,Go)] > (lizzieLet2_4QVal_Int_3QError_Int_1QError_Int,QTree_Int) */
  assign lizzieLet2_4QVal_Int_3QError_Int_1QError_Int_d = QError_Int_dc((& {lizzieLet2_4QVal_Int_3QError_Int_1_d[0]}), lizzieLet2_4QVal_Int_3QError_Int_1_d);
  assign {lizzieLet2_4QVal_Int_3QError_Int_1_r} = {1 {(lizzieLet2_4QVal_Int_3QError_Int_1QError_Int_r && lizzieLet2_4QVal_Int_3QError_Int_1QError_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (lizzieLet2_4QVal_Int_3QError_Int_1QError_Int,QTree_Int) > (lizzieLet6_1_argbuf,QTree_Int) */
  QTree_Int_t lizzieLet2_4QVal_Int_3QError_Int_1QError_Int_bufchan_d;
  logic lizzieLet2_4QVal_Int_3QError_Int_1QError_Int_bufchan_r;
  assign lizzieLet2_4QVal_Int_3QError_Int_1QError_Int_r = ((! lizzieLet2_4QVal_Int_3QError_Int_1QError_Int_bufchan_d[0]) || lizzieLet2_4QVal_Int_3QError_Int_1QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet2_4QVal_Int_3QError_Int_1QError_Int_bufchan_d <= {66'd0,
                                                                 1'd0};
    else
      if (lizzieLet2_4QVal_Int_3QError_Int_1QError_Int_r)
        lizzieLet2_4QVal_Int_3QError_Int_1QError_Int_bufchan_d <= lizzieLet2_4QVal_Int_3QError_Int_1QError_Int_d;
  QTree_Int_t lizzieLet2_4QVal_Int_3QError_Int_1QError_Int_bufchan_buf;
  assign lizzieLet2_4QVal_Int_3QError_Int_1QError_Int_bufchan_r = (! lizzieLet2_4QVal_Int_3QError_Int_1QError_Int_bufchan_buf[0]);
  assign lizzieLet6_1_argbuf_d = (lizzieLet2_4QVal_Int_3QError_Int_1QError_Int_bufchan_buf[0] ? lizzieLet2_4QVal_Int_3QError_Int_1QError_Int_bufchan_buf :
                                  lizzieLet2_4QVal_Int_3QError_Int_1QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet2_4QVal_Int_3QError_Int_1QError_Int_bufchan_buf <= {66'd0,
                                                                   1'd0};
    else
      if ((lizzieLet6_1_argbuf_r && lizzieLet2_4QVal_Int_3QError_Int_1QError_Int_bufchan_buf[0]))
        lizzieLet2_4QVal_Int_3QError_Int_1QError_Int_bufchan_buf <= {66'd0,
                                                                     1'd0};
      else if (((! lizzieLet6_1_argbuf_r) && (! lizzieLet2_4QVal_Int_3QError_Int_1QError_Int_bufchan_buf[0])))
        lizzieLet2_4QVal_Int_3QError_Int_1QError_Int_bufchan_buf <= lizzieLet2_4QVal_Int_3QError_Int_1QError_Int_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet2_4QVal_Int_3QError_Int_2,Go) > (lizzieLet2_4QVal_Int_3QError_Int_2_argbuf,Go) */
  Go_t lizzieLet2_4QVal_Int_3QError_Int_2_bufchan_d;
  logic lizzieLet2_4QVal_Int_3QError_Int_2_bufchan_r;
  assign lizzieLet2_4QVal_Int_3QError_Int_2_r = ((! lizzieLet2_4QVal_Int_3QError_Int_2_bufchan_d[0]) || lizzieLet2_4QVal_Int_3QError_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet2_4QVal_Int_3QError_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet2_4QVal_Int_3QError_Int_2_r)
        lizzieLet2_4QVal_Int_3QError_Int_2_bufchan_d <= lizzieLet2_4QVal_Int_3QError_Int_2_d;
  Go_t lizzieLet2_4QVal_Int_3QError_Int_2_bufchan_buf;
  assign lizzieLet2_4QVal_Int_3QError_Int_2_bufchan_r = (! lizzieLet2_4QVal_Int_3QError_Int_2_bufchan_buf[0]);
  assign lizzieLet2_4QVal_Int_3QError_Int_2_argbuf_d = (lizzieLet2_4QVal_Int_3QError_Int_2_bufchan_buf[0] ? lizzieLet2_4QVal_Int_3QError_Int_2_bufchan_buf :
                                                        lizzieLet2_4QVal_Int_3QError_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet2_4QVal_Int_3QError_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet2_4QVal_Int_3QError_Int_2_argbuf_r && lizzieLet2_4QVal_Int_3QError_Int_2_bufchan_buf[0]))
        lizzieLet2_4QVal_Int_3QError_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet2_4QVal_Int_3QError_Int_2_argbuf_r) && (! lizzieLet2_4QVal_Int_3QError_Int_2_bufchan_buf[0])))
        lizzieLet2_4QVal_Int_3QError_Int_2_bufchan_buf <= lizzieLet2_4QVal_Int_3QError_Int_2_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet2_4QVal_Int_3QNode_Int,Go) > [(lizzieLet2_4QVal_Int_3QNode_Int_1,Go),
                                                       (lizzieLet2_4QVal_Int_3QNode_Int_2,Go)] */
  logic [1:0] lizzieLet2_4QVal_Int_3QNode_Int_emitted;
  logic [1:0] lizzieLet2_4QVal_Int_3QNode_Int_done;
  assign lizzieLet2_4QVal_Int_3QNode_Int_1_d = (lizzieLet2_4QVal_Int_3QNode_Int_d[0] && (! lizzieLet2_4QVal_Int_3QNode_Int_emitted[0]));
  assign lizzieLet2_4QVal_Int_3QNode_Int_2_d = (lizzieLet2_4QVal_Int_3QNode_Int_d[0] && (! lizzieLet2_4QVal_Int_3QNode_Int_emitted[1]));
  assign lizzieLet2_4QVal_Int_3QNode_Int_done = (lizzieLet2_4QVal_Int_3QNode_Int_emitted | ({lizzieLet2_4QVal_Int_3QNode_Int_2_d[0],
                                                                                             lizzieLet2_4QVal_Int_3QNode_Int_1_d[0]} & {lizzieLet2_4QVal_Int_3QNode_Int_2_r,
                                                                                                                                        lizzieLet2_4QVal_Int_3QNode_Int_1_r}));
  assign lizzieLet2_4QVal_Int_3QNode_Int_r = (& lizzieLet2_4QVal_Int_3QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet2_4QVal_Int_3QNode_Int_emitted <= 2'd0;
    else
      lizzieLet2_4QVal_Int_3QNode_Int_emitted <= (lizzieLet2_4QVal_Int_3QNode_Int_r ? 2'd0 :
                                                  lizzieLet2_4QVal_Int_3QNode_Int_done);
  
  /* dcon (Ty QTree_Int,
      Dcon QError_Int) : [(lizzieLet2_4QVal_Int_3QNode_Int_1,Go)] > (lizzieLet2_4QVal_Int_3QNode_Int_1QError_Int,QTree_Int) */
  assign lizzieLet2_4QVal_Int_3QNode_Int_1QError_Int_d = QError_Int_dc((& {lizzieLet2_4QVal_Int_3QNode_Int_1_d[0]}), lizzieLet2_4QVal_Int_3QNode_Int_1_d);
  assign {lizzieLet2_4QVal_Int_3QNode_Int_1_r} = {1 {(lizzieLet2_4QVal_Int_3QNode_Int_1QError_Int_r && lizzieLet2_4QVal_Int_3QNode_Int_1QError_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (lizzieLet2_4QVal_Int_3QNode_Int_1QError_Int,QTree_Int) > (lizzieLet5_1_argbuf,QTree_Int) */
  QTree_Int_t lizzieLet2_4QVal_Int_3QNode_Int_1QError_Int_bufchan_d;
  logic lizzieLet2_4QVal_Int_3QNode_Int_1QError_Int_bufchan_r;
  assign lizzieLet2_4QVal_Int_3QNode_Int_1QError_Int_r = ((! lizzieLet2_4QVal_Int_3QNode_Int_1QError_Int_bufchan_d[0]) || lizzieLet2_4QVal_Int_3QNode_Int_1QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet2_4QVal_Int_3QNode_Int_1QError_Int_bufchan_d <= {66'd0,
                                                                1'd0};
    else
      if (lizzieLet2_4QVal_Int_3QNode_Int_1QError_Int_r)
        lizzieLet2_4QVal_Int_3QNode_Int_1QError_Int_bufchan_d <= lizzieLet2_4QVal_Int_3QNode_Int_1QError_Int_d;
  QTree_Int_t lizzieLet2_4QVal_Int_3QNode_Int_1QError_Int_bufchan_buf;
  assign lizzieLet2_4QVal_Int_3QNode_Int_1QError_Int_bufchan_r = (! lizzieLet2_4QVal_Int_3QNode_Int_1QError_Int_bufchan_buf[0]);
  assign lizzieLet5_1_argbuf_d = (lizzieLet2_4QVal_Int_3QNode_Int_1QError_Int_bufchan_buf[0] ? lizzieLet2_4QVal_Int_3QNode_Int_1QError_Int_bufchan_buf :
                                  lizzieLet2_4QVal_Int_3QNode_Int_1QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet2_4QVal_Int_3QNode_Int_1QError_Int_bufchan_buf <= {66'd0,
                                                                  1'd0};
    else
      if ((lizzieLet5_1_argbuf_r && lizzieLet2_4QVal_Int_3QNode_Int_1QError_Int_bufchan_buf[0]))
        lizzieLet2_4QVal_Int_3QNode_Int_1QError_Int_bufchan_buf <= {66'd0,
                                                                    1'd0};
      else if (((! lizzieLet5_1_argbuf_r) && (! lizzieLet2_4QVal_Int_3QNode_Int_1QError_Int_bufchan_buf[0])))
        lizzieLet2_4QVal_Int_3QNode_Int_1QError_Int_bufchan_buf <= lizzieLet2_4QVal_Int_3QNode_Int_1QError_Int_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet2_4QVal_Int_3QNode_Int_2,Go) > (lizzieLet2_4QVal_Int_3QNode_Int_2_argbuf,Go) */
  Go_t lizzieLet2_4QVal_Int_3QNode_Int_2_bufchan_d;
  logic lizzieLet2_4QVal_Int_3QNode_Int_2_bufchan_r;
  assign lizzieLet2_4QVal_Int_3QNode_Int_2_r = ((! lizzieLet2_4QVal_Int_3QNode_Int_2_bufchan_d[0]) || lizzieLet2_4QVal_Int_3QNode_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet2_4QVal_Int_3QNode_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet2_4QVal_Int_3QNode_Int_2_r)
        lizzieLet2_4QVal_Int_3QNode_Int_2_bufchan_d <= lizzieLet2_4QVal_Int_3QNode_Int_2_d;
  Go_t lizzieLet2_4QVal_Int_3QNode_Int_2_bufchan_buf;
  assign lizzieLet2_4QVal_Int_3QNode_Int_2_bufchan_r = (! lizzieLet2_4QVal_Int_3QNode_Int_2_bufchan_buf[0]);
  assign lizzieLet2_4QVal_Int_3QNode_Int_2_argbuf_d = (lizzieLet2_4QVal_Int_3QNode_Int_2_bufchan_buf[0] ? lizzieLet2_4QVal_Int_3QNode_Int_2_bufchan_buf :
                                                       lizzieLet2_4QVal_Int_3QNode_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet2_4QVal_Int_3QNode_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet2_4QVal_Int_3QNode_Int_2_argbuf_r && lizzieLet2_4QVal_Int_3QNode_Int_2_bufchan_buf[0]))
        lizzieLet2_4QVal_Int_3QNode_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet2_4QVal_Int_3QNode_Int_2_argbuf_r) && (! lizzieLet2_4QVal_Int_3QNode_Int_2_bufchan_buf[0])))
        lizzieLet2_4QVal_Int_3QNode_Int_2_bufchan_buf <= lizzieLet2_4QVal_Int_3QNode_Int_2_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet2_4QVal_Int_3QNone_Int,Go) > (lizzieLet2_4QVal_Int_3QNone_Int_1_argbuf,Go) */
  Go_t lizzieLet2_4QVal_Int_3QNone_Int_bufchan_d;
  logic lizzieLet2_4QVal_Int_3QNone_Int_bufchan_r;
  assign lizzieLet2_4QVal_Int_3QNone_Int_r = ((! lizzieLet2_4QVal_Int_3QNone_Int_bufchan_d[0]) || lizzieLet2_4QVal_Int_3QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet2_4QVal_Int_3QNone_Int_bufchan_d <= 1'd0;
    else
      if (lizzieLet2_4QVal_Int_3QNone_Int_r)
        lizzieLet2_4QVal_Int_3QNone_Int_bufchan_d <= lizzieLet2_4QVal_Int_3QNone_Int_d;
  Go_t lizzieLet2_4QVal_Int_3QNone_Int_bufchan_buf;
  assign lizzieLet2_4QVal_Int_3QNone_Int_bufchan_r = (! lizzieLet2_4QVal_Int_3QNone_Int_bufchan_buf[0]);
  assign lizzieLet2_4QVal_Int_3QNone_Int_1_argbuf_d = (lizzieLet2_4QVal_Int_3QNone_Int_bufchan_buf[0] ? lizzieLet2_4QVal_Int_3QNone_Int_bufchan_buf :
                                                       lizzieLet2_4QVal_Int_3QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet2_4QVal_Int_3QNone_Int_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet2_4QVal_Int_3QNone_Int_1_argbuf_r && lizzieLet2_4QVal_Int_3QNone_Int_bufchan_buf[0]))
        lizzieLet2_4QVal_Int_3QNone_Int_bufchan_buf <= 1'd0;
      else if (((! lizzieLet2_4QVal_Int_3QNone_Int_1_argbuf_r) && (! lizzieLet2_4QVal_Int_3QNone_Int_bufchan_buf[0])))
        lizzieLet2_4QVal_Int_3QNone_Int_bufchan_buf <= lizzieLet2_4QVal_Int_3QNone_Int_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet2_4QVal_Int_3QVal_Int,Go) > (lizzieLet2_4QVal_Int_3QVal_Int_1_argbuf,Go) */
  Go_t lizzieLet2_4QVal_Int_3QVal_Int_bufchan_d;
  logic lizzieLet2_4QVal_Int_3QVal_Int_bufchan_r;
  assign lizzieLet2_4QVal_Int_3QVal_Int_r = ((! lizzieLet2_4QVal_Int_3QVal_Int_bufchan_d[0]) || lizzieLet2_4QVal_Int_3QVal_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet2_4QVal_Int_3QVal_Int_bufchan_d <= 1'd0;
    else
      if (lizzieLet2_4QVal_Int_3QVal_Int_r)
        lizzieLet2_4QVal_Int_3QVal_Int_bufchan_d <= lizzieLet2_4QVal_Int_3QVal_Int_d;
  Go_t lizzieLet2_4QVal_Int_3QVal_Int_bufchan_buf;
  assign lizzieLet2_4QVal_Int_3QVal_Int_bufchan_r = (! lizzieLet2_4QVal_Int_3QVal_Int_bufchan_buf[0]);
  assign lizzieLet2_4QVal_Int_3QVal_Int_1_argbuf_d = (lizzieLet2_4QVal_Int_3QVal_Int_bufchan_buf[0] ? lizzieLet2_4QVal_Int_3QVal_Int_bufchan_buf :
                                                      lizzieLet2_4QVal_Int_3QVal_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet2_4QVal_Int_3QVal_Int_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet2_4QVal_Int_3QVal_Int_1_argbuf_r && lizzieLet2_4QVal_Int_3QVal_Int_bufchan_buf[0]))
        lizzieLet2_4QVal_Int_3QVal_Int_bufchan_buf <= 1'd0;
      else if (((! lizzieLet2_4QVal_Int_3QVal_Int_1_argbuf_r) && (! lizzieLet2_4QVal_Int_3QVal_Int_bufchan_buf[0])))
        lizzieLet2_4QVal_Int_3QVal_Int_bufchan_buf <= lizzieLet2_4QVal_Int_3QVal_Int_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_CT$wmAdd_Int) : (lizzieLet2_4QVal_Int_4,QTree_Int) (lizzieLet2_5QVal_Int,Pointer_CT$wmAdd_Int) > [(lizzieLet2_4QVal_Int_4QNone_Int,Pointer_CT$wmAdd_Int),
                                                                                                                    (lizzieLet2_4QVal_Int_4QVal_Int,Pointer_CT$wmAdd_Int),
                                                                                                                    (lizzieLet2_4QVal_Int_4QNode_Int,Pointer_CT$wmAdd_Int),
                                                                                                                    (lizzieLet2_4QVal_Int_4QError_Int,Pointer_CT$wmAdd_Int)] */
  logic [3:0] lizzieLet2_5QVal_Int_onehotd;
  always_comb
    if ((lizzieLet2_4QVal_Int_4_d[0] && lizzieLet2_5QVal_Int_d[0]))
      unique case (lizzieLet2_4QVal_Int_4_d[2:1])
        2'd0: lizzieLet2_5QVal_Int_onehotd = 4'd1;
        2'd1: lizzieLet2_5QVal_Int_onehotd = 4'd2;
        2'd2: lizzieLet2_5QVal_Int_onehotd = 4'd4;
        2'd3: lizzieLet2_5QVal_Int_onehotd = 4'd8;
        default: lizzieLet2_5QVal_Int_onehotd = 4'd0;
      endcase
    else lizzieLet2_5QVal_Int_onehotd = 4'd0;
  assign lizzieLet2_4QVal_Int_4QNone_Int_d = {lizzieLet2_5QVal_Int_d[16:1],
                                              lizzieLet2_5QVal_Int_onehotd[0]};
  assign lizzieLet2_4QVal_Int_4QVal_Int_d = {lizzieLet2_5QVal_Int_d[16:1],
                                             lizzieLet2_5QVal_Int_onehotd[1]};
  assign lizzieLet2_4QVal_Int_4QNode_Int_d = {lizzieLet2_5QVal_Int_d[16:1],
                                              lizzieLet2_5QVal_Int_onehotd[2]};
  assign lizzieLet2_4QVal_Int_4QError_Int_d = {lizzieLet2_5QVal_Int_d[16:1],
                                               lizzieLet2_5QVal_Int_onehotd[3]};
  assign lizzieLet2_5QVal_Int_r = (| (lizzieLet2_5QVal_Int_onehotd & {lizzieLet2_4QVal_Int_4QError_Int_r,
                                                                      lizzieLet2_4QVal_Int_4QNode_Int_r,
                                                                      lizzieLet2_4QVal_Int_4QVal_Int_r,
                                                                      lizzieLet2_4QVal_Int_4QNone_Int_r}));
  assign lizzieLet2_4QVal_Int_4_r = lizzieLet2_5QVal_Int_r;
  
  /* buf (Ty Pointer_CT$wmAdd_Int) : (lizzieLet2_4QVal_Int_4QError_Int,Pointer_CT$wmAdd_Int) > (lizzieLet2_4QVal_Int_4QError_Int_1_argbuf,Pointer_CT$wmAdd_Int) */
  Pointer_CT$wmAdd_Int_t lizzieLet2_4QVal_Int_4QError_Int_bufchan_d;
  logic lizzieLet2_4QVal_Int_4QError_Int_bufchan_r;
  assign lizzieLet2_4QVal_Int_4QError_Int_r = ((! lizzieLet2_4QVal_Int_4QError_Int_bufchan_d[0]) || lizzieLet2_4QVal_Int_4QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet2_4QVal_Int_4QError_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet2_4QVal_Int_4QError_Int_r)
        lizzieLet2_4QVal_Int_4QError_Int_bufchan_d <= lizzieLet2_4QVal_Int_4QError_Int_d;
  Pointer_CT$wmAdd_Int_t lizzieLet2_4QVal_Int_4QError_Int_bufchan_buf;
  assign lizzieLet2_4QVal_Int_4QError_Int_bufchan_r = (! lizzieLet2_4QVal_Int_4QError_Int_bufchan_buf[0]);
  assign lizzieLet2_4QVal_Int_4QError_Int_1_argbuf_d = (lizzieLet2_4QVal_Int_4QError_Int_bufchan_buf[0] ? lizzieLet2_4QVal_Int_4QError_Int_bufchan_buf :
                                                        lizzieLet2_4QVal_Int_4QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet2_4QVal_Int_4QError_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet2_4QVal_Int_4QError_Int_1_argbuf_r && lizzieLet2_4QVal_Int_4QError_Int_bufchan_buf[0]))
        lizzieLet2_4QVal_Int_4QError_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet2_4QVal_Int_4QError_Int_1_argbuf_r) && (! lizzieLet2_4QVal_Int_4QError_Int_bufchan_buf[0])))
        lizzieLet2_4QVal_Int_4QError_Int_bufchan_buf <= lizzieLet2_4QVal_Int_4QError_Int_bufchan_d;
  
  /* buf (Ty Pointer_CT$wmAdd_Int) : (lizzieLet2_4QVal_Int_4QNode_Int,Pointer_CT$wmAdd_Int) > (lizzieLet2_4QVal_Int_4QNode_Int_1_argbuf,Pointer_CT$wmAdd_Int) */
  Pointer_CT$wmAdd_Int_t lizzieLet2_4QVal_Int_4QNode_Int_bufchan_d;
  logic lizzieLet2_4QVal_Int_4QNode_Int_bufchan_r;
  assign lizzieLet2_4QVal_Int_4QNode_Int_r = ((! lizzieLet2_4QVal_Int_4QNode_Int_bufchan_d[0]) || lizzieLet2_4QVal_Int_4QNode_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet2_4QVal_Int_4QNode_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet2_4QVal_Int_4QNode_Int_r)
        lizzieLet2_4QVal_Int_4QNode_Int_bufchan_d <= lizzieLet2_4QVal_Int_4QNode_Int_d;
  Pointer_CT$wmAdd_Int_t lizzieLet2_4QVal_Int_4QNode_Int_bufchan_buf;
  assign lizzieLet2_4QVal_Int_4QNode_Int_bufchan_r = (! lizzieLet2_4QVal_Int_4QNode_Int_bufchan_buf[0]);
  assign lizzieLet2_4QVal_Int_4QNode_Int_1_argbuf_d = (lizzieLet2_4QVal_Int_4QNode_Int_bufchan_buf[0] ? lizzieLet2_4QVal_Int_4QNode_Int_bufchan_buf :
                                                       lizzieLet2_4QVal_Int_4QNode_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet2_4QVal_Int_4QNode_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet2_4QVal_Int_4QNode_Int_1_argbuf_r && lizzieLet2_4QVal_Int_4QNode_Int_bufchan_buf[0]))
        lizzieLet2_4QVal_Int_4QNode_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet2_4QVal_Int_4QNode_Int_1_argbuf_r) && (! lizzieLet2_4QVal_Int_4QNode_Int_bufchan_buf[0])))
        lizzieLet2_4QVal_Int_4QNode_Int_bufchan_buf <= lizzieLet2_4QVal_Int_4QNode_Int_bufchan_d;
  
  /* buf (Ty Pointer_CT$wmAdd_Int) : (lizzieLet2_4QVal_Int_4QNone_Int,Pointer_CT$wmAdd_Int) > (lizzieLet2_4QVal_Int_4QNone_Int_1_argbuf,Pointer_CT$wmAdd_Int) */
  Pointer_CT$wmAdd_Int_t lizzieLet2_4QVal_Int_4QNone_Int_bufchan_d;
  logic lizzieLet2_4QVal_Int_4QNone_Int_bufchan_r;
  assign lizzieLet2_4QVal_Int_4QNone_Int_r = ((! lizzieLet2_4QVal_Int_4QNone_Int_bufchan_d[0]) || lizzieLet2_4QVal_Int_4QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet2_4QVal_Int_4QNone_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet2_4QVal_Int_4QNone_Int_r)
        lizzieLet2_4QVal_Int_4QNone_Int_bufchan_d <= lizzieLet2_4QVal_Int_4QNone_Int_d;
  Pointer_CT$wmAdd_Int_t lizzieLet2_4QVal_Int_4QNone_Int_bufchan_buf;
  assign lizzieLet2_4QVal_Int_4QNone_Int_bufchan_r = (! lizzieLet2_4QVal_Int_4QNone_Int_bufchan_buf[0]);
  assign lizzieLet2_4QVal_Int_4QNone_Int_1_argbuf_d = (lizzieLet2_4QVal_Int_4QNone_Int_bufchan_buf[0] ? lizzieLet2_4QVal_Int_4QNone_Int_bufchan_buf :
                                                       lizzieLet2_4QVal_Int_4QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet2_4QVal_Int_4QNone_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet2_4QVal_Int_4QNone_Int_1_argbuf_r && lizzieLet2_4QVal_Int_4QNone_Int_bufchan_buf[0]))
        lizzieLet2_4QVal_Int_4QNone_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet2_4QVal_Int_4QNone_Int_1_argbuf_r) && (! lizzieLet2_4QVal_Int_4QNone_Int_bufchan_buf[0])))
        lizzieLet2_4QVal_Int_4QNone_Int_bufchan_buf <= lizzieLet2_4QVal_Int_4QNone_Int_bufchan_d;
  
  /* buf (Ty Pointer_CT$wmAdd_Int) : (lizzieLet2_4QVal_Int_4QVal_Int,Pointer_CT$wmAdd_Int) > (lizzieLet2_4QVal_Int_4QVal_Int_1_argbuf,Pointer_CT$wmAdd_Int) */
  Pointer_CT$wmAdd_Int_t lizzieLet2_4QVal_Int_4QVal_Int_bufchan_d;
  logic lizzieLet2_4QVal_Int_4QVal_Int_bufchan_r;
  assign lizzieLet2_4QVal_Int_4QVal_Int_r = ((! lizzieLet2_4QVal_Int_4QVal_Int_bufchan_d[0]) || lizzieLet2_4QVal_Int_4QVal_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet2_4QVal_Int_4QVal_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet2_4QVal_Int_4QVal_Int_r)
        lizzieLet2_4QVal_Int_4QVal_Int_bufchan_d <= lizzieLet2_4QVal_Int_4QVal_Int_d;
  Pointer_CT$wmAdd_Int_t lizzieLet2_4QVal_Int_4QVal_Int_bufchan_buf;
  assign lizzieLet2_4QVal_Int_4QVal_Int_bufchan_r = (! lizzieLet2_4QVal_Int_4QVal_Int_bufchan_buf[0]);
  assign lizzieLet2_4QVal_Int_4QVal_Int_1_argbuf_d = (lizzieLet2_4QVal_Int_4QVal_Int_bufchan_buf[0] ? lizzieLet2_4QVal_Int_4QVal_Int_bufchan_buf :
                                                      lizzieLet2_4QVal_Int_4QVal_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet2_4QVal_Int_4QVal_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet2_4QVal_Int_4QVal_Int_1_argbuf_r && lizzieLet2_4QVal_Int_4QVal_Int_bufchan_buf[0]))
        lizzieLet2_4QVal_Int_4QVal_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet2_4QVal_Int_4QVal_Int_1_argbuf_r) && (! lizzieLet2_4QVal_Int_4QVal_Int_bufchan_buf[0])))
        lizzieLet2_4QVal_Int_4QVal_Int_bufchan_buf <= lizzieLet2_4QVal_Int_4QVal_Int_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_QTree_Int) : (lizzieLet2_4QVal_Int_5,QTree_Int) (lizzieLet2_6QVal_Int,Pointer_QTree_Int) > [(lizzieLet2_4QVal_Int_5QNone_Int,Pointer_QTree_Int),
                                                                                                              (_17,Pointer_QTree_Int),
                                                                                                              (_16,Pointer_QTree_Int),
                                                                                                              (_15,Pointer_QTree_Int)] */
  logic [3:0] lizzieLet2_6QVal_Int_onehotd;
  always_comb
    if ((lizzieLet2_4QVal_Int_5_d[0] && lizzieLet2_6QVal_Int_d[0]))
      unique case (lizzieLet2_4QVal_Int_5_d[2:1])
        2'd0: lizzieLet2_6QVal_Int_onehotd = 4'd1;
        2'd1: lizzieLet2_6QVal_Int_onehotd = 4'd2;
        2'd2: lizzieLet2_6QVal_Int_onehotd = 4'd4;
        2'd3: lizzieLet2_6QVal_Int_onehotd = 4'd8;
        default: lizzieLet2_6QVal_Int_onehotd = 4'd0;
      endcase
    else lizzieLet2_6QVal_Int_onehotd = 4'd0;
  assign lizzieLet2_4QVal_Int_5QNone_Int_d = {lizzieLet2_6QVal_Int_d[16:1],
                                              lizzieLet2_6QVal_Int_onehotd[0]};
  assign _17_d = {lizzieLet2_6QVal_Int_d[16:1],
                  lizzieLet2_6QVal_Int_onehotd[1]};
  assign _16_d = {lizzieLet2_6QVal_Int_d[16:1],
                  lizzieLet2_6QVal_Int_onehotd[2]};
  assign _15_d = {lizzieLet2_6QVal_Int_d[16:1],
                  lizzieLet2_6QVal_Int_onehotd[3]};
  assign lizzieLet2_6QVal_Int_r = (| (lizzieLet2_6QVal_Int_onehotd & {_15_r,
                                                                      _16_r,
                                                                      _17_r,
                                                                      lizzieLet2_4QVal_Int_5QNone_Int_r}));
  assign lizzieLet2_4QVal_Int_5_r = lizzieLet2_6QVal_Int_r;
  
  /* buf (Ty Pointer_QTree_Int) : (lizzieLet2_4QVal_Int_5QNone_Int,Pointer_QTree_Int) > (lizzieLet2_4QVal_Int_5QNone_Int_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t lizzieLet2_4QVal_Int_5QNone_Int_bufchan_d;
  logic lizzieLet2_4QVal_Int_5QNone_Int_bufchan_r;
  assign lizzieLet2_4QVal_Int_5QNone_Int_r = ((! lizzieLet2_4QVal_Int_5QNone_Int_bufchan_d[0]) || lizzieLet2_4QVal_Int_5QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet2_4QVal_Int_5QNone_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet2_4QVal_Int_5QNone_Int_r)
        lizzieLet2_4QVal_Int_5QNone_Int_bufchan_d <= lizzieLet2_4QVal_Int_5QNone_Int_d;
  Pointer_QTree_Int_t lizzieLet2_4QVal_Int_5QNone_Int_bufchan_buf;
  assign lizzieLet2_4QVal_Int_5QNone_Int_bufchan_r = (! lizzieLet2_4QVal_Int_5QNone_Int_bufchan_buf[0]);
  assign lizzieLet2_4QVal_Int_5QNone_Int_1_argbuf_d = (lizzieLet2_4QVal_Int_5QNone_Int_bufchan_buf[0] ? lizzieLet2_4QVal_Int_5QNone_Int_bufchan_buf :
                                                       lizzieLet2_4QVal_Int_5QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet2_4QVal_Int_5QNone_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet2_4QVal_Int_5QNone_Int_1_argbuf_r && lizzieLet2_4QVal_Int_5QNone_Int_bufchan_buf[0]))
        lizzieLet2_4QVal_Int_5QNone_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet2_4QVal_Int_5QNone_Int_1_argbuf_r) && (! lizzieLet2_4QVal_Int_5QNone_Int_bufchan_buf[0])))
        lizzieLet2_4QVal_Int_5QNone_Int_bufchan_buf <= lizzieLet2_4QVal_Int_5QNone_Int_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty MyDTInt_Int_Int) : (lizzieLet2_4QVal_Int_6,QTree_Int) (lizzieLet2_8QVal_Int,MyDTInt_Int_Int) > [(_14,MyDTInt_Int_Int),
                                                                                                          (lizzieLet2_4QVal_Int_6QVal_Int,MyDTInt_Int_Int),
                                                                                                          (_13,MyDTInt_Int_Int),
                                                                                                          (_12,MyDTInt_Int_Int)] */
  logic [3:0] lizzieLet2_8QVal_Int_onehotd;
  always_comb
    if ((lizzieLet2_4QVal_Int_6_d[0] && lizzieLet2_8QVal_Int_d[0]))
      unique case (lizzieLet2_4QVal_Int_6_d[2:1])
        2'd0: lizzieLet2_8QVal_Int_onehotd = 4'd1;
        2'd1: lizzieLet2_8QVal_Int_onehotd = 4'd2;
        2'd2: lizzieLet2_8QVal_Int_onehotd = 4'd4;
        2'd3: lizzieLet2_8QVal_Int_onehotd = 4'd8;
        default: lizzieLet2_8QVal_Int_onehotd = 4'd0;
      endcase
    else lizzieLet2_8QVal_Int_onehotd = 4'd0;
  assign _14_d = lizzieLet2_8QVal_Int_onehotd[0];
  assign lizzieLet2_4QVal_Int_6QVal_Int_d = lizzieLet2_8QVal_Int_onehotd[1];
  assign _13_d = lizzieLet2_8QVal_Int_onehotd[2];
  assign _12_d = lizzieLet2_8QVal_Int_onehotd[3];
  assign lizzieLet2_8QVal_Int_r = (| (lizzieLet2_8QVal_Int_onehotd & {_12_r,
                                                                      _13_r,
                                                                      lizzieLet2_4QVal_Int_6QVal_Int_r,
                                                                      _14_r}));
  assign lizzieLet2_4QVal_Int_6_r = lizzieLet2_8QVal_Int_r;
  
  /* buf (Ty MyDTInt_Int_Int) : (lizzieLet2_4QVal_Int_6QVal_Int,MyDTInt_Int_Int) > (lizzieLet2_4QVal_Int_6QVal_Int_1_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t lizzieLet2_4QVal_Int_6QVal_Int_bufchan_d;
  logic lizzieLet2_4QVal_Int_6QVal_Int_bufchan_r;
  assign lizzieLet2_4QVal_Int_6QVal_Int_r = ((! lizzieLet2_4QVal_Int_6QVal_Int_bufchan_d[0]) || lizzieLet2_4QVal_Int_6QVal_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet2_4QVal_Int_6QVal_Int_bufchan_d <= 1'd0;
    else
      if (lizzieLet2_4QVal_Int_6QVal_Int_r)
        lizzieLet2_4QVal_Int_6QVal_Int_bufchan_d <= lizzieLet2_4QVal_Int_6QVal_Int_d;
  MyDTInt_Int_Int_t lizzieLet2_4QVal_Int_6QVal_Int_bufchan_buf;
  assign lizzieLet2_4QVal_Int_6QVal_Int_bufchan_r = (! lizzieLet2_4QVal_Int_6QVal_Int_bufchan_buf[0]);
  assign lizzieLet2_4QVal_Int_6QVal_Int_1_argbuf_d = (lizzieLet2_4QVal_Int_6QVal_Int_bufchan_buf[0] ? lizzieLet2_4QVal_Int_6QVal_Int_bufchan_buf :
                                                      lizzieLet2_4QVal_Int_6QVal_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet2_4QVal_Int_6QVal_Int_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet2_4QVal_Int_6QVal_Int_1_argbuf_r && lizzieLet2_4QVal_Int_6QVal_Int_bufchan_buf[0]))
        lizzieLet2_4QVal_Int_6QVal_Int_bufchan_buf <= 1'd0;
      else if (((! lizzieLet2_4QVal_Int_6QVal_Int_1_argbuf_r) && (! lizzieLet2_4QVal_Int_6QVal_Int_bufchan_buf[0])))
        lizzieLet2_4QVal_Int_6QVal_Int_bufchan_buf <= lizzieLet2_4QVal_Int_6QVal_Int_bufchan_d;
  
  /* dcon (Ty TupMyDTInt_Int_Int___Int___Int,
      Dcon TupMyDTInt_Int_Int___Int___Int) : [(lizzieLet2_4QVal_Int_6QVal_Int_1_argbuf,MyDTInt_Int_Int),
                                              (lizzieLet2_4QVal_Int_7QVal_Int_1_argbuf,Int),
                                              (va8c_1_argbuf,Int)] > (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1,TupMyDTInt_Int_Int___Int___Int) */
  assign applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_d = TupMyDTInt_Int_Int___Int___Int_dc((& {lizzieLet2_4QVal_Int_6QVal_Int_1_argbuf_d[0],
                                                                                                        lizzieLet2_4QVal_Int_7QVal_Int_1_argbuf_d[0],
                                                                                                        va8c_1_argbuf_d[0]}), lizzieLet2_4QVal_Int_6QVal_Int_1_argbuf_d, lizzieLet2_4QVal_Int_7QVal_Int_1_argbuf_d, va8c_1_argbuf_d);
  assign {lizzieLet2_4QVal_Int_6QVal_Int_1_argbuf_r,
          lizzieLet2_4QVal_Int_7QVal_Int_1_argbuf_r,
          va8c_1_argbuf_r} = {3 {(applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_r && applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_d[0])}};
  
  /* demux (Ty QTree_Int,
       Ty Int) : (lizzieLet2_4QVal_Int_7,QTree_Int) (v1a8b_destruct,Int) > [(_11,Int),
                                                                            (lizzieLet2_4QVal_Int_7QVal_Int,Int),
                                                                            (_10,Int),
                                                                            (_9,Int)] */
  logic [3:0] v1a8b_destruct_onehotd;
  always_comb
    if ((lizzieLet2_4QVal_Int_7_d[0] && v1a8b_destruct_d[0]))
      unique case (lizzieLet2_4QVal_Int_7_d[2:1])
        2'd0: v1a8b_destruct_onehotd = 4'd1;
        2'd1: v1a8b_destruct_onehotd = 4'd2;
        2'd2: v1a8b_destruct_onehotd = 4'd4;
        2'd3: v1a8b_destruct_onehotd = 4'd8;
        default: v1a8b_destruct_onehotd = 4'd0;
      endcase
    else v1a8b_destruct_onehotd = 4'd0;
  assign _11_d = {v1a8b_destruct_d[32:1], v1a8b_destruct_onehotd[0]};
  assign lizzieLet2_4QVal_Int_7QVal_Int_d = {v1a8b_destruct_d[32:1],
                                             v1a8b_destruct_onehotd[1]};
  assign _10_d = {v1a8b_destruct_d[32:1], v1a8b_destruct_onehotd[2]};
  assign _9_d = {v1a8b_destruct_d[32:1], v1a8b_destruct_onehotd[3]};
  assign v1a8b_destruct_r = (| (v1a8b_destruct_onehotd & {_9_r,
                                                          _10_r,
                                                          lizzieLet2_4QVal_Int_7QVal_Int_r,
                                                          _11_r}));
  assign lizzieLet2_4QVal_Int_7_r = v1a8b_destruct_r;
  
  /* buf (Ty Int) : (lizzieLet2_4QVal_Int_7QVal_Int,Int) > (lizzieLet2_4QVal_Int_7QVal_Int_1_argbuf,Int) */
  Int_t lizzieLet2_4QVal_Int_7QVal_Int_bufchan_d;
  logic lizzieLet2_4QVal_Int_7QVal_Int_bufchan_r;
  assign lizzieLet2_4QVal_Int_7QVal_Int_r = ((! lizzieLet2_4QVal_Int_7QVal_Int_bufchan_d[0]) || lizzieLet2_4QVal_Int_7QVal_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet2_4QVal_Int_7QVal_Int_bufchan_d <= {32'd0, 1'd0};
    else
      if (lizzieLet2_4QVal_Int_7QVal_Int_r)
        lizzieLet2_4QVal_Int_7QVal_Int_bufchan_d <= lizzieLet2_4QVal_Int_7QVal_Int_d;
  Int_t lizzieLet2_4QVal_Int_7QVal_Int_bufchan_buf;
  assign lizzieLet2_4QVal_Int_7QVal_Int_bufchan_r = (! lizzieLet2_4QVal_Int_7QVal_Int_bufchan_buf[0]);
  assign lizzieLet2_4QVal_Int_7QVal_Int_1_argbuf_d = (lizzieLet2_4QVal_Int_7QVal_Int_bufchan_buf[0] ? lizzieLet2_4QVal_Int_7QVal_Int_bufchan_buf :
                                                      lizzieLet2_4QVal_Int_7QVal_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet2_4QVal_Int_7QVal_Int_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((lizzieLet2_4QVal_Int_7QVal_Int_1_argbuf_r && lizzieLet2_4QVal_Int_7QVal_Int_bufchan_buf[0]))
        lizzieLet2_4QVal_Int_7QVal_Int_bufchan_buf <= {32'd0, 1'd0};
      else if (((! lizzieLet2_4QVal_Int_7QVal_Int_1_argbuf_r) && (! lizzieLet2_4QVal_Int_7QVal_Int_bufchan_buf[0])))
        lizzieLet2_4QVal_Int_7QVal_Int_bufchan_buf <= lizzieLet2_4QVal_Int_7QVal_Int_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_CT$wmAdd_Int) : (lizzieLet2_5,QTree_Int) (sc_0_goMux_mux,Pointer_CT$wmAdd_Int) > [(lizzieLet2_5QNone_Int,Pointer_CT$wmAdd_Int),
                                                                                                    (lizzieLet2_5QVal_Int,Pointer_CT$wmAdd_Int),
                                                                                                    (lizzieLet2_5QNode_Int,Pointer_CT$wmAdd_Int),
                                                                                                    (lizzieLet2_5QError_Int,Pointer_CT$wmAdd_Int)] */
  logic [3:0] sc_0_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet2_5_d[0] && sc_0_goMux_mux_d[0]))
      unique case (lizzieLet2_5_d[2:1])
        2'd0: sc_0_goMux_mux_onehotd = 4'd1;
        2'd1: sc_0_goMux_mux_onehotd = 4'd2;
        2'd2: sc_0_goMux_mux_onehotd = 4'd4;
        2'd3: sc_0_goMux_mux_onehotd = 4'd8;
        default: sc_0_goMux_mux_onehotd = 4'd0;
      endcase
    else sc_0_goMux_mux_onehotd = 4'd0;
  assign lizzieLet2_5QNone_Int_d = {sc_0_goMux_mux_d[16:1],
                                    sc_0_goMux_mux_onehotd[0]};
  assign lizzieLet2_5QVal_Int_d = {sc_0_goMux_mux_d[16:1],
                                   sc_0_goMux_mux_onehotd[1]};
  assign lizzieLet2_5QNode_Int_d = {sc_0_goMux_mux_d[16:1],
                                    sc_0_goMux_mux_onehotd[2]};
  assign lizzieLet2_5QError_Int_d = {sc_0_goMux_mux_d[16:1],
                                     sc_0_goMux_mux_onehotd[3]};
  assign sc_0_goMux_mux_r = (| (sc_0_goMux_mux_onehotd & {lizzieLet2_5QError_Int_r,
                                                          lizzieLet2_5QNode_Int_r,
                                                          lizzieLet2_5QVal_Int_r,
                                                          lizzieLet2_5QNone_Int_r}));
  assign lizzieLet2_5_r = sc_0_goMux_mux_r;
  
  /* buf (Ty Pointer_CT$wmAdd_Int) : (lizzieLet2_5QError_Int,Pointer_CT$wmAdd_Int) > (lizzieLet2_5QError_Int_1_argbuf,Pointer_CT$wmAdd_Int) */
  Pointer_CT$wmAdd_Int_t lizzieLet2_5QError_Int_bufchan_d;
  logic lizzieLet2_5QError_Int_bufchan_r;
  assign lizzieLet2_5QError_Int_r = ((! lizzieLet2_5QError_Int_bufchan_d[0]) || lizzieLet2_5QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet2_5QError_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet2_5QError_Int_r)
        lizzieLet2_5QError_Int_bufchan_d <= lizzieLet2_5QError_Int_d;
  Pointer_CT$wmAdd_Int_t lizzieLet2_5QError_Int_bufchan_buf;
  assign lizzieLet2_5QError_Int_bufchan_r = (! lizzieLet2_5QError_Int_bufchan_buf[0]);
  assign lizzieLet2_5QError_Int_1_argbuf_d = (lizzieLet2_5QError_Int_bufchan_buf[0] ? lizzieLet2_5QError_Int_bufchan_buf :
                                              lizzieLet2_5QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet2_5QError_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet2_5QError_Int_1_argbuf_r && lizzieLet2_5QError_Int_bufchan_buf[0]))
        lizzieLet2_5QError_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet2_5QError_Int_1_argbuf_r) && (! lizzieLet2_5QError_Int_bufchan_buf[0])))
        lizzieLet2_5QError_Int_bufchan_buf <= lizzieLet2_5QError_Int_bufchan_d;
  
  /* buf (Ty Pointer_CT$wmAdd_Int) : (lizzieLet2_5QNone_Int,Pointer_CT$wmAdd_Int) > (lizzieLet2_5QNone_Int_1_argbuf,Pointer_CT$wmAdd_Int) */
  Pointer_CT$wmAdd_Int_t lizzieLet2_5QNone_Int_bufchan_d;
  logic lizzieLet2_5QNone_Int_bufchan_r;
  assign lizzieLet2_5QNone_Int_r = ((! lizzieLet2_5QNone_Int_bufchan_d[0]) || lizzieLet2_5QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet2_5QNone_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet2_5QNone_Int_r)
        lizzieLet2_5QNone_Int_bufchan_d <= lizzieLet2_5QNone_Int_d;
  Pointer_CT$wmAdd_Int_t lizzieLet2_5QNone_Int_bufchan_buf;
  assign lizzieLet2_5QNone_Int_bufchan_r = (! lizzieLet2_5QNone_Int_bufchan_buf[0]);
  assign lizzieLet2_5QNone_Int_1_argbuf_d = (lizzieLet2_5QNone_Int_bufchan_buf[0] ? lizzieLet2_5QNone_Int_bufchan_buf :
                                             lizzieLet2_5QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet2_5QNone_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet2_5QNone_Int_1_argbuf_r && lizzieLet2_5QNone_Int_bufchan_buf[0]))
        lizzieLet2_5QNone_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet2_5QNone_Int_1_argbuf_r) && (! lizzieLet2_5QNone_Int_bufchan_buf[0])))
        lizzieLet2_5QNone_Int_bufchan_buf <= lizzieLet2_5QNone_Int_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_QTree_Int) : (lizzieLet2_6,QTree_Int) (w1sif_1_2,Pointer_QTree_Int) > [(_8,Pointer_QTree_Int),
                                                                                         (lizzieLet2_6QVal_Int,Pointer_QTree_Int),
                                                                                         (lizzieLet2_6QNode_Int,Pointer_QTree_Int),
                                                                                         (_7,Pointer_QTree_Int)] */
  logic [3:0] w1sif_1_2_onehotd;
  always_comb
    if ((lizzieLet2_6_d[0] && w1sif_1_2_d[0]))
      unique case (lizzieLet2_6_d[2:1])
        2'd0: w1sif_1_2_onehotd = 4'd1;
        2'd1: w1sif_1_2_onehotd = 4'd2;
        2'd2: w1sif_1_2_onehotd = 4'd4;
        2'd3: w1sif_1_2_onehotd = 4'd8;
        default: w1sif_1_2_onehotd = 4'd0;
      endcase
    else w1sif_1_2_onehotd = 4'd0;
  assign _8_d = {w1sif_1_2_d[16:1], w1sif_1_2_onehotd[0]};
  assign lizzieLet2_6QVal_Int_d = {w1sif_1_2_d[16:1],
                                   w1sif_1_2_onehotd[1]};
  assign lizzieLet2_6QNode_Int_d = {w1sif_1_2_d[16:1],
                                    w1sif_1_2_onehotd[2]};
  assign _7_d = {w1sif_1_2_d[16:1], w1sif_1_2_onehotd[3]};
  assign w1sif_1_2_r = (| (w1sif_1_2_onehotd & {_7_r,
                                                lizzieLet2_6QNode_Int_r,
                                                lizzieLet2_6QVal_Int_r,
                                                _8_r}));
  assign lizzieLet2_6_r = w1sif_1_2_r;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_QTree_Int) : (lizzieLet2_7,QTree_Int) (w2sig_1_2,Pointer_QTree_Int) > [(lizzieLet2_7QNone_Int,Pointer_QTree_Int),
                                                                                         (_6,Pointer_QTree_Int),
                                                                                         (_5,Pointer_QTree_Int),
                                                                                         (_4,Pointer_QTree_Int)] */
  logic [3:0] w2sig_1_2_onehotd;
  always_comb
    if ((lizzieLet2_7_d[0] && w2sig_1_2_d[0]))
      unique case (lizzieLet2_7_d[2:1])
        2'd0: w2sig_1_2_onehotd = 4'd1;
        2'd1: w2sig_1_2_onehotd = 4'd2;
        2'd2: w2sig_1_2_onehotd = 4'd4;
        2'd3: w2sig_1_2_onehotd = 4'd8;
        default: w2sig_1_2_onehotd = 4'd0;
      endcase
    else w2sig_1_2_onehotd = 4'd0;
  assign lizzieLet2_7QNone_Int_d = {w2sig_1_2_d[16:1],
                                    w2sig_1_2_onehotd[0]};
  assign _6_d = {w2sig_1_2_d[16:1], w2sig_1_2_onehotd[1]};
  assign _5_d = {w2sig_1_2_d[16:1], w2sig_1_2_onehotd[2]};
  assign _4_d = {w2sig_1_2_d[16:1], w2sig_1_2_onehotd[3]};
  assign w2sig_1_2_r = (| (w2sig_1_2_onehotd & {_4_r,
                                                _5_r,
                                                _6_r,
                                                lizzieLet2_7QNone_Int_r}));
  assign lizzieLet2_7_r = w2sig_1_2_r;
  
  /* buf (Ty Pointer_QTree_Int) : (lizzieLet2_7QNone_Int,Pointer_QTree_Int) > (lizzieLet2_7QNone_Int_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t lizzieLet2_7QNone_Int_bufchan_d;
  logic lizzieLet2_7QNone_Int_bufchan_r;
  assign lizzieLet2_7QNone_Int_r = ((! lizzieLet2_7QNone_Int_bufchan_d[0]) || lizzieLet2_7QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet2_7QNone_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet2_7QNone_Int_r)
        lizzieLet2_7QNone_Int_bufchan_d <= lizzieLet2_7QNone_Int_d;
  Pointer_QTree_Int_t lizzieLet2_7QNone_Int_bufchan_buf;
  assign lizzieLet2_7QNone_Int_bufchan_r = (! lizzieLet2_7QNone_Int_bufchan_buf[0]);
  assign lizzieLet2_7QNone_Int_1_argbuf_d = (lizzieLet2_7QNone_Int_bufchan_buf[0] ? lizzieLet2_7QNone_Int_bufchan_buf :
                                             lizzieLet2_7QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet2_7QNone_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet2_7QNone_Int_1_argbuf_r && lizzieLet2_7QNone_Int_bufchan_buf[0]))
        lizzieLet2_7QNone_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet2_7QNone_Int_1_argbuf_r) && (! lizzieLet2_7QNone_Int_bufchan_buf[0])))
        lizzieLet2_7QNone_Int_bufchan_buf <= lizzieLet2_7QNone_Int_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty MyDTInt_Int_Int) : (lizzieLet2_8,QTree_Int) (wsie_1_goMux_mux,MyDTInt_Int_Int) > [(_3,MyDTInt_Int_Int),
                                                                                            (lizzieLet2_8QVal_Int,MyDTInt_Int_Int),
                                                                                            (lizzieLet2_8QNode_Int,MyDTInt_Int_Int),
                                                                                            (_2,MyDTInt_Int_Int)] */
  logic [3:0] wsie_1_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet2_8_d[0] && wsie_1_goMux_mux_d[0]))
      unique case (lizzieLet2_8_d[2:1])
        2'd0: wsie_1_goMux_mux_onehotd = 4'd1;
        2'd1: wsie_1_goMux_mux_onehotd = 4'd2;
        2'd2: wsie_1_goMux_mux_onehotd = 4'd4;
        2'd3: wsie_1_goMux_mux_onehotd = 4'd8;
        default: wsie_1_goMux_mux_onehotd = 4'd0;
      endcase
    else wsie_1_goMux_mux_onehotd = 4'd0;
  assign _3_d = wsie_1_goMux_mux_onehotd[0];
  assign lizzieLet2_8QVal_Int_d = wsie_1_goMux_mux_onehotd[1];
  assign lizzieLet2_8QNode_Int_d = wsie_1_goMux_mux_onehotd[2];
  assign _2_d = wsie_1_goMux_mux_onehotd[3];
  assign wsie_1_goMux_mux_r = (| (wsie_1_goMux_mux_onehotd & {_2_r,
                                                              lizzieLet2_8QNode_Int_r,
                                                              lizzieLet2_8QVal_Int_r,
                                                              _3_r}));
  assign lizzieLet2_8_r = wsie_1_goMux_mux_r;
  
  /* destruct (Ty CTmain_mask_Int,
          Dcon Lcall_main_mask_Int0) : (lizzieLet31_1Lcall_main_mask_Int0,CTmain_mask_Int) > [(es_1_1_destruct,Pointer_QTree_Int),
                                                                                              (es_2_2_destruct,Pointer_QTree_Int),
                                                                                              (es_3_5_destruct,Pointer_QTree_Int),
                                                                                              (sc_0_14_destruct,Pointer_CTmain_mask_Int)] */
  logic [3:0] lizzieLet31_1Lcall_main_mask_Int0_emitted;
  logic [3:0] lizzieLet31_1Lcall_main_mask_Int0_done;
  assign es_1_1_destruct_d = {lizzieLet31_1Lcall_main_mask_Int0_d[19:4],
                              (lizzieLet31_1Lcall_main_mask_Int0_d[0] && (! lizzieLet31_1Lcall_main_mask_Int0_emitted[0]))};
  assign es_2_2_destruct_d = {lizzieLet31_1Lcall_main_mask_Int0_d[35:20],
                              (lizzieLet31_1Lcall_main_mask_Int0_d[0] && (! lizzieLet31_1Lcall_main_mask_Int0_emitted[1]))};
  assign es_3_5_destruct_d = {lizzieLet31_1Lcall_main_mask_Int0_d[51:36],
                              (lizzieLet31_1Lcall_main_mask_Int0_d[0] && (! lizzieLet31_1Lcall_main_mask_Int0_emitted[2]))};
  assign sc_0_14_destruct_d = {lizzieLet31_1Lcall_main_mask_Int0_d[67:52],
                               (lizzieLet31_1Lcall_main_mask_Int0_d[0] && (! lizzieLet31_1Lcall_main_mask_Int0_emitted[3]))};
  assign lizzieLet31_1Lcall_main_mask_Int0_done = (lizzieLet31_1Lcall_main_mask_Int0_emitted | ({sc_0_14_destruct_d[0],
                                                                                                 es_3_5_destruct_d[0],
                                                                                                 es_2_2_destruct_d[0],
                                                                                                 es_1_1_destruct_d[0]} & {sc_0_14_destruct_r,
                                                                                                                          es_3_5_destruct_r,
                                                                                                                          es_2_2_destruct_r,
                                                                                                                          es_1_1_destruct_r}));
  assign lizzieLet31_1Lcall_main_mask_Int0_r = (& lizzieLet31_1Lcall_main_mask_Int0_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet31_1Lcall_main_mask_Int0_emitted <= 4'd0;
    else
      lizzieLet31_1Lcall_main_mask_Int0_emitted <= (lizzieLet31_1Lcall_main_mask_Int0_r ? 4'd0 :
                                                    lizzieLet31_1Lcall_main_mask_Int0_done);
  
  /* destruct (Ty CTmain_mask_Int,
          Dcon Lcall_main_mask_Int1) : (lizzieLet31_1Lcall_main_mask_Int1,CTmain_mask_Int) > [(es_2_1_destruct,Pointer_QTree_Int),
                                                                                              (es_3_4_destruct,Pointer_QTree_Int),
                                                                                              (sc_0_13_destruct,Pointer_CTmain_mask_Int),
                                                                                              (t1a8x_3_destruct,Pointer_QTree_Int),
                                                                                              (q1a8s_3_destruct,Pointer_MaskQTree)] */
  logic [4:0] lizzieLet31_1Lcall_main_mask_Int1_emitted;
  logic [4:0] lizzieLet31_1Lcall_main_mask_Int1_done;
  assign es_2_1_destruct_d = {lizzieLet31_1Lcall_main_mask_Int1_d[19:4],
                              (lizzieLet31_1Lcall_main_mask_Int1_d[0] && (! lizzieLet31_1Lcall_main_mask_Int1_emitted[0]))};
  assign es_3_4_destruct_d = {lizzieLet31_1Lcall_main_mask_Int1_d[35:20],
                              (lizzieLet31_1Lcall_main_mask_Int1_d[0] && (! lizzieLet31_1Lcall_main_mask_Int1_emitted[1]))};
  assign sc_0_13_destruct_d = {lizzieLet31_1Lcall_main_mask_Int1_d[51:36],
                               (lizzieLet31_1Lcall_main_mask_Int1_d[0] && (! lizzieLet31_1Lcall_main_mask_Int1_emitted[2]))};
  assign t1a8x_3_destruct_d = {lizzieLet31_1Lcall_main_mask_Int1_d[67:52],
                               (lizzieLet31_1Lcall_main_mask_Int1_d[0] && (! lizzieLet31_1Lcall_main_mask_Int1_emitted[3]))};
  assign q1a8s_3_destruct_d = {lizzieLet31_1Lcall_main_mask_Int1_d[83:68],
                               (lizzieLet31_1Lcall_main_mask_Int1_d[0] && (! lizzieLet31_1Lcall_main_mask_Int1_emitted[4]))};
  assign lizzieLet31_1Lcall_main_mask_Int1_done = (lizzieLet31_1Lcall_main_mask_Int1_emitted | ({q1a8s_3_destruct_d[0],
                                                                                                 t1a8x_3_destruct_d[0],
                                                                                                 sc_0_13_destruct_d[0],
                                                                                                 es_3_4_destruct_d[0],
                                                                                                 es_2_1_destruct_d[0]} & {q1a8s_3_destruct_r,
                                                                                                                          t1a8x_3_destruct_r,
                                                                                                                          sc_0_13_destruct_r,
                                                                                                                          es_3_4_destruct_r,
                                                                                                                          es_2_1_destruct_r}));
  assign lizzieLet31_1Lcall_main_mask_Int1_r = (& lizzieLet31_1Lcall_main_mask_Int1_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet31_1Lcall_main_mask_Int1_emitted <= 5'd0;
    else
      lizzieLet31_1Lcall_main_mask_Int1_emitted <= (lizzieLet31_1Lcall_main_mask_Int1_r ? 5'd0 :
                                                    lizzieLet31_1Lcall_main_mask_Int1_done);
  
  /* destruct (Ty CTmain_mask_Int,
          Dcon Lcall_main_mask_Int2) : (lizzieLet31_1Lcall_main_mask_Int2,CTmain_mask_Int) > [(es_3_3_destruct,Pointer_QTree_Int),
                                                                                              (sc_0_12_destruct,Pointer_CTmain_mask_Int),
                                                                                              (t1a8x_2_destruct,Pointer_QTree_Int),
                                                                                              (q1a8s_2_destruct,Pointer_MaskQTree),
                                                                                              (t2a8y_2_destruct,Pointer_QTree_Int),
                                                                                              (q2a8t_2_destruct,Pointer_MaskQTree)] */
  logic [5:0] lizzieLet31_1Lcall_main_mask_Int2_emitted;
  logic [5:0] lizzieLet31_1Lcall_main_mask_Int2_done;
  assign es_3_3_destruct_d = {lizzieLet31_1Lcall_main_mask_Int2_d[19:4],
                              (lizzieLet31_1Lcall_main_mask_Int2_d[0] && (! lizzieLet31_1Lcall_main_mask_Int2_emitted[0]))};
  assign sc_0_12_destruct_d = {lizzieLet31_1Lcall_main_mask_Int2_d[35:20],
                               (lizzieLet31_1Lcall_main_mask_Int2_d[0] && (! lizzieLet31_1Lcall_main_mask_Int2_emitted[1]))};
  assign t1a8x_2_destruct_d = {lizzieLet31_1Lcall_main_mask_Int2_d[51:36],
                               (lizzieLet31_1Lcall_main_mask_Int2_d[0] && (! lizzieLet31_1Lcall_main_mask_Int2_emitted[2]))};
  assign q1a8s_2_destruct_d = {lizzieLet31_1Lcall_main_mask_Int2_d[67:52],
                               (lizzieLet31_1Lcall_main_mask_Int2_d[0] && (! lizzieLet31_1Lcall_main_mask_Int2_emitted[3]))};
  assign t2a8y_2_destruct_d = {lizzieLet31_1Lcall_main_mask_Int2_d[83:68],
                               (lizzieLet31_1Lcall_main_mask_Int2_d[0] && (! lizzieLet31_1Lcall_main_mask_Int2_emitted[4]))};
  assign q2a8t_2_destruct_d = {lizzieLet31_1Lcall_main_mask_Int2_d[99:84],
                               (lizzieLet31_1Lcall_main_mask_Int2_d[0] && (! lizzieLet31_1Lcall_main_mask_Int2_emitted[5]))};
  assign lizzieLet31_1Lcall_main_mask_Int2_done = (lizzieLet31_1Lcall_main_mask_Int2_emitted | ({q2a8t_2_destruct_d[0],
                                                                                                 t2a8y_2_destruct_d[0],
                                                                                                 q1a8s_2_destruct_d[0],
                                                                                                 t1a8x_2_destruct_d[0],
                                                                                                 sc_0_12_destruct_d[0],
                                                                                                 es_3_3_destruct_d[0]} & {q2a8t_2_destruct_r,
                                                                                                                          t2a8y_2_destruct_r,
                                                                                                                          q1a8s_2_destruct_r,
                                                                                                                          t1a8x_2_destruct_r,
                                                                                                                          sc_0_12_destruct_r,
                                                                                                                          es_3_3_destruct_r}));
  assign lizzieLet31_1Lcall_main_mask_Int2_r = (& lizzieLet31_1Lcall_main_mask_Int2_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet31_1Lcall_main_mask_Int2_emitted <= 6'd0;
    else
      lizzieLet31_1Lcall_main_mask_Int2_emitted <= (lizzieLet31_1Lcall_main_mask_Int2_r ? 6'd0 :
                                                    lizzieLet31_1Lcall_main_mask_Int2_done);
  
  /* destruct (Ty CTmain_mask_Int,
          Dcon Lcall_main_mask_Int3) : (lizzieLet31_1Lcall_main_mask_Int3,CTmain_mask_Int) > [(sc_0_11_destruct,Pointer_CTmain_mask_Int),
                                                                                              (t1a8x_1_destruct,Pointer_QTree_Int),
                                                                                              (q1a8s_1_destruct,Pointer_MaskQTree),
                                                                                              (t2a8y_1_destruct,Pointer_QTree_Int),
                                                                                              (q2a8t_1_destruct,Pointer_MaskQTree),
                                                                                              (t3a8z_1_destruct,Pointer_QTree_Int),
                                                                                              (q3a8u_1_destruct,Pointer_MaskQTree)] */
  logic [6:0] lizzieLet31_1Lcall_main_mask_Int3_emitted;
  logic [6:0] lizzieLet31_1Lcall_main_mask_Int3_done;
  assign sc_0_11_destruct_d = {lizzieLet31_1Lcall_main_mask_Int3_d[19:4],
                               (lizzieLet31_1Lcall_main_mask_Int3_d[0] && (! lizzieLet31_1Lcall_main_mask_Int3_emitted[0]))};
  assign t1a8x_1_destruct_d = {lizzieLet31_1Lcall_main_mask_Int3_d[35:20],
                               (lizzieLet31_1Lcall_main_mask_Int3_d[0] && (! lizzieLet31_1Lcall_main_mask_Int3_emitted[1]))};
  assign q1a8s_1_destruct_d = {lizzieLet31_1Lcall_main_mask_Int3_d[51:36],
                               (lizzieLet31_1Lcall_main_mask_Int3_d[0] && (! lizzieLet31_1Lcall_main_mask_Int3_emitted[2]))};
  assign t2a8y_1_destruct_d = {lizzieLet31_1Lcall_main_mask_Int3_d[67:52],
                               (lizzieLet31_1Lcall_main_mask_Int3_d[0] && (! lizzieLet31_1Lcall_main_mask_Int3_emitted[3]))};
  assign q2a8t_1_destruct_d = {lizzieLet31_1Lcall_main_mask_Int3_d[83:68],
                               (lizzieLet31_1Lcall_main_mask_Int3_d[0] && (! lizzieLet31_1Lcall_main_mask_Int3_emitted[4]))};
  assign t3a8z_1_destruct_d = {lizzieLet31_1Lcall_main_mask_Int3_d[99:84],
                               (lizzieLet31_1Lcall_main_mask_Int3_d[0] && (! lizzieLet31_1Lcall_main_mask_Int3_emitted[5]))};
  assign q3a8u_1_destruct_d = {lizzieLet31_1Lcall_main_mask_Int3_d[115:100],
                               (lizzieLet31_1Lcall_main_mask_Int3_d[0] && (! lizzieLet31_1Lcall_main_mask_Int3_emitted[6]))};
  assign lizzieLet31_1Lcall_main_mask_Int3_done = (lizzieLet31_1Lcall_main_mask_Int3_emitted | ({q3a8u_1_destruct_d[0],
                                                                                                 t3a8z_1_destruct_d[0],
                                                                                                 q2a8t_1_destruct_d[0],
                                                                                                 t2a8y_1_destruct_d[0],
                                                                                                 q1a8s_1_destruct_d[0],
                                                                                                 t1a8x_1_destruct_d[0],
                                                                                                 sc_0_11_destruct_d[0]} & {q3a8u_1_destruct_r,
                                                                                                                           t3a8z_1_destruct_r,
                                                                                                                           q2a8t_1_destruct_r,
                                                                                                                           t2a8y_1_destruct_r,
                                                                                                                           q1a8s_1_destruct_r,
                                                                                                                           t1a8x_1_destruct_r,
                                                                                                                           sc_0_11_destruct_r}));
  assign lizzieLet31_1Lcall_main_mask_Int3_r = (& lizzieLet31_1Lcall_main_mask_Int3_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet31_1Lcall_main_mask_Int3_emitted <= 7'd0;
    else
      lizzieLet31_1Lcall_main_mask_Int3_emitted <= (lizzieLet31_1Lcall_main_mask_Int3_r ? 7'd0 :
                                                    lizzieLet31_1Lcall_main_mask_Int3_done);
  
  /* demux (Ty CTmain_mask_Int,
       Ty CTmain_mask_Int) : (lizzieLet31_2,CTmain_mask_Int) (lizzieLet31_1,CTmain_mask_Int) > [(_1,CTmain_mask_Int),
                                                                                                (lizzieLet31_1Lcall_main_mask_Int3,CTmain_mask_Int),
                                                                                                (lizzieLet31_1Lcall_main_mask_Int2,CTmain_mask_Int),
                                                                                                (lizzieLet31_1Lcall_main_mask_Int1,CTmain_mask_Int),
                                                                                                (lizzieLet31_1Lcall_main_mask_Int0,CTmain_mask_Int)] */
  logic [4:0] lizzieLet31_1_onehotd;
  always_comb
    if ((lizzieLet31_2_d[0] && lizzieLet31_1_d[0]))
      unique case (lizzieLet31_2_d[3:1])
        3'd0: lizzieLet31_1_onehotd = 5'd1;
        3'd1: lizzieLet31_1_onehotd = 5'd2;
        3'd2: lizzieLet31_1_onehotd = 5'd4;
        3'd3: lizzieLet31_1_onehotd = 5'd8;
        3'd4: lizzieLet31_1_onehotd = 5'd16;
        default: lizzieLet31_1_onehotd = 5'd0;
      endcase
    else lizzieLet31_1_onehotd = 5'd0;
  assign _1_d = {lizzieLet31_1_d[115:1], lizzieLet31_1_onehotd[0]};
  assign lizzieLet31_1Lcall_main_mask_Int3_d = {lizzieLet31_1_d[115:1],
                                                lizzieLet31_1_onehotd[1]};
  assign lizzieLet31_1Lcall_main_mask_Int2_d = {lizzieLet31_1_d[115:1],
                                                lizzieLet31_1_onehotd[2]};
  assign lizzieLet31_1Lcall_main_mask_Int1_d = {lizzieLet31_1_d[115:1],
                                                lizzieLet31_1_onehotd[3]};
  assign lizzieLet31_1Lcall_main_mask_Int0_d = {lizzieLet31_1_d[115:1],
                                                lizzieLet31_1_onehotd[4]};
  assign lizzieLet31_1_r = (| (lizzieLet31_1_onehotd & {lizzieLet31_1Lcall_main_mask_Int0_r,
                                                        lizzieLet31_1Lcall_main_mask_Int1_r,
                                                        lizzieLet31_1Lcall_main_mask_Int2_r,
                                                        lizzieLet31_1Lcall_main_mask_Int3_r,
                                                        _1_r}));
  assign lizzieLet31_2_r = lizzieLet31_1_r;
  
  /* demux (Ty CTmain_mask_Int,
       Ty Go) : (lizzieLet31_3,CTmain_mask_Int) (go_12_goMux_data,Go) > [(_0,Go),
                                                                         (lizzieLet31_3Lcall_main_mask_Int3,Go),
                                                                         (lizzieLet31_3Lcall_main_mask_Int2,Go),
                                                                         (lizzieLet31_3Lcall_main_mask_Int1,Go),
                                                                         (lizzieLet31_3Lcall_main_mask_Int0,Go)] */
  logic [4:0] go_12_goMux_data_onehotd;
  always_comb
    if ((lizzieLet31_3_d[0] && go_12_goMux_data_d[0]))
      unique case (lizzieLet31_3_d[3:1])
        3'd0: go_12_goMux_data_onehotd = 5'd1;
        3'd1: go_12_goMux_data_onehotd = 5'd2;
        3'd2: go_12_goMux_data_onehotd = 5'd4;
        3'd3: go_12_goMux_data_onehotd = 5'd8;
        3'd4: go_12_goMux_data_onehotd = 5'd16;
        default: go_12_goMux_data_onehotd = 5'd0;
      endcase
    else go_12_goMux_data_onehotd = 5'd0;
  assign _0_d = go_12_goMux_data_onehotd[0];
  assign lizzieLet31_3Lcall_main_mask_Int3_d = go_12_goMux_data_onehotd[1];
  assign lizzieLet31_3Lcall_main_mask_Int2_d = go_12_goMux_data_onehotd[2];
  assign lizzieLet31_3Lcall_main_mask_Int1_d = go_12_goMux_data_onehotd[3];
  assign lizzieLet31_3Lcall_main_mask_Int0_d = go_12_goMux_data_onehotd[4];
  assign go_12_goMux_data_r = (| (go_12_goMux_data_onehotd & {lizzieLet31_3Lcall_main_mask_Int0_r,
                                                              lizzieLet31_3Lcall_main_mask_Int1_r,
                                                              lizzieLet31_3Lcall_main_mask_Int2_r,
                                                              lizzieLet31_3Lcall_main_mask_Int3_r,
                                                              _0_r}));
  assign lizzieLet31_3_r = go_12_goMux_data_r;
  
  /* buf (Ty Go) : (lizzieLet31_3Lcall_main_mask_Int0,Go) > (lizzieLet31_3Lcall_main_mask_Int0_1_argbuf,Go) */
  Go_t lizzieLet31_3Lcall_main_mask_Int0_bufchan_d;
  logic lizzieLet31_3Lcall_main_mask_Int0_bufchan_r;
  assign lizzieLet31_3Lcall_main_mask_Int0_r = ((! lizzieLet31_3Lcall_main_mask_Int0_bufchan_d[0]) || lizzieLet31_3Lcall_main_mask_Int0_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet31_3Lcall_main_mask_Int0_bufchan_d <= 1'd0;
    else
      if (lizzieLet31_3Lcall_main_mask_Int0_r)
        lizzieLet31_3Lcall_main_mask_Int0_bufchan_d <= lizzieLet31_3Lcall_main_mask_Int0_d;
  Go_t lizzieLet31_3Lcall_main_mask_Int0_bufchan_buf;
  assign lizzieLet31_3Lcall_main_mask_Int0_bufchan_r = (! lizzieLet31_3Lcall_main_mask_Int0_bufchan_buf[0]);
  assign lizzieLet31_3Lcall_main_mask_Int0_1_argbuf_d = (lizzieLet31_3Lcall_main_mask_Int0_bufchan_buf[0] ? lizzieLet31_3Lcall_main_mask_Int0_bufchan_buf :
                                                         lizzieLet31_3Lcall_main_mask_Int0_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet31_3Lcall_main_mask_Int0_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet31_3Lcall_main_mask_Int0_1_argbuf_r && lizzieLet31_3Lcall_main_mask_Int0_bufchan_buf[0]))
        lizzieLet31_3Lcall_main_mask_Int0_bufchan_buf <= 1'd0;
      else if (((! lizzieLet31_3Lcall_main_mask_Int0_1_argbuf_r) && (! lizzieLet31_3Lcall_main_mask_Int0_bufchan_buf[0])))
        lizzieLet31_3Lcall_main_mask_Int0_bufchan_buf <= lizzieLet31_3Lcall_main_mask_Int0_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet31_3Lcall_main_mask_Int1,Go) > (lizzieLet31_3Lcall_main_mask_Int1_1_argbuf,Go) */
  Go_t lizzieLet31_3Lcall_main_mask_Int1_bufchan_d;
  logic lizzieLet31_3Lcall_main_mask_Int1_bufchan_r;
  assign lizzieLet31_3Lcall_main_mask_Int1_r = ((! lizzieLet31_3Lcall_main_mask_Int1_bufchan_d[0]) || lizzieLet31_3Lcall_main_mask_Int1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet31_3Lcall_main_mask_Int1_bufchan_d <= 1'd0;
    else
      if (lizzieLet31_3Lcall_main_mask_Int1_r)
        lizzieLet31_3Lcall_main_mask_Int1_bufchan_d <= lizzieLet31_3Lcall_main_mask_Int1_d;
  Go_t lizzieLet31_3Lcall_main_mask_Int1_bufchan_buf;
  assign lizzieLet31_3Lcall_main_mask_Int1_bufchan_r = (! lizzieLet31_3Lcall_main_mask_Int1_bufchan_buf[0]);
  assign lizzieLet31_3Lcall_main_mask_Int1_1_argbuf_d = (lizzieLet31_3Lcall_main_mask_Int1_bufchan_buf[0] ? lizzieLet31_3Lcall_main_mask_Int1_bufchan_buf :
                                                         lizzieLet31_3Lcall_main_mask_Int1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet31_3Lcall_main_mask_Int1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet31_3Lcall_main_mask_Int1_1_argbuf_r && lizzieLet31_3Lcall_main_mask_Int1_bufchan_buf[0]))
        lizzieLet31_3Lcall_main_mask_Int1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet31_3Lcall_main_mask_Int1_1_argbuf_r) && (! lizzieLet31_3Lcall_main_mask_Int1_bufchan_buf[0])))
        lizzieLet31_3Lcall_main_mask_Int1_bufchan_buf <= lizzieLet31_3Lcall_main_mask_Int1_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet31_3Lcall_main_mask_Int2,Go) > (lizzieLet31_3Lcall_main_mask_Int2_1_argbuf,Go) */
  Go_t lizzieLet31_3Lcall_main_mask_Int2_bufchan_d;
  logic lizzieLet31_3Lcall_main_mask_Int2_bufchan_r;
  assign lizzieLet31_3Lcall_main_mask_Int2_r = ((! lizzieLet31_3Lcall_main_mask_Int2_bufchan_d[0]) || lizzieLet31_3Lcall_main_mask_Int2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet31_3Lcall_main_mask_Int2_bufchan_d <= 1'd0;
    else
      if (lizzieLet31_3Lcall_main_mask_Int2_r)
        lizzieLet31_3Lcall_main_mask_Int2_bufchan_d <= lizzieLet31_3Lcall_main_mask_Int2_d;
  Go_t lizzieLet31_3Lcall_main_mask_Int2_bufchan_buf;
  assign lizzieLet31_3Lcall_main_mask_Int2_bufchan_r = (! lizzieLet31_3Lcall_main_mask_Int2_bufchan_buf[0]);
  assign lizzieLet31_3Lcall_main_mask_Int2_1_argbuf_d = (lizzieLet31_3Lcall_main_mask_Int2_bufchan_buf[0] ? lizzieLet31_3Lcall_main_mask_Int2_bufchan_buf :
                                                         lizzieLet31_3Lcall_main_mask_Int2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet31_3Lcall_main_mask_Int2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet31_3Lcall_main_mask_Int2_1_argbuf_r && lizzieLet31_3Lcall_main_mask_Int2_bufchan_buf[0]))
        lizzieLet31_3Lcall_main_mask_Int2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet31_3Lcall_main_mask_Int2_1_argbuf_r) && (! lizzieLet31_3Lcall_main_mask_Int2_bufchan_buf[0])))
        lizzieLet31_3Lcall_main_mask_Int2_bufchan_buf <= lizzieLet31_3Lcall_main_mask_Int2_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet31_3Lcall_main_mask_Int3,Go) > (lizzieLet31_3Lcall_main_mask_Int3_1_argbuf,Go) */
  Go_t lizzieLet31_3Lcall_main_mask_Int3_bufchan_d;
  logic lizzieLet31_3Lcall_main_mask_Int3_bufchan_r;
  assign lizzieLet31_3Lcall_main_mask_Int3_r = ((! lizzieLet31_3Lcall_main_mask_Int3_bufchan_d[0]) || lizzieLet31_3Lcall_main_mask_Int3_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet31_3Lcall_main_mask_Int3_bufchan_d <= 1'd0;
    else
      if (lizzieLet31_3Lcall_main_mask_Int3_r)
        lizzieLet31_3Lcall_main_mask_Int3_bufchan_d <= lizzieLet31_3Lcall_main_mask_Int3_d;
  Go_t lizzieLet31_3Lcall_main_mask_Int3_bufchan_buf;
  assign lizzieLet31_3Lcall_main_mask_Int3_bufchan_r = (! lizzieLet31_3Lcall_main_mask_Int3_bufchan_buf[0]);
  assign lizzieLet31_3Lcall_main_mask_Int3_1_argbuf_d = (lizzieLet31_3Lcall_main_mask_Int3_bufchan_buf[0] ? lizzieLet31_3Lcall_main_mask_Int3_bufchan_buf :
                                                         lizzieLet31_3Lcall_main_mask_Int3_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet31_3Lcall_main_mask_Int3_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet31_3Lcall_main_mask_Int3_1_argbuf_r && lizzieLet31_3Lcall_main_mask_Int3_bufchan_buf[0]))
        lizzieLet31_3Lcall_main_mask_Int3_bufchan_buf <= 1'd0;
      else if (((! lizzieLet31_3Lcall_main_mask_Int3_1_argbuf_r) && (! lizzieLet31_3Lcall_main_mask_Int3_bufchan_buf[0])))
        lizzieLet31_3Lcall_main_mask_Int3_bufchan_buf <= lizzieLet31_3Lcall_main_mask_Int3_bufchan_d;
  
  /* demux (Ty CTmain_mask_Int,
       Ty Pointer_QTree_Int) : (lizzieLet31_4,CTmain_mask_Int) (srtarg_0_2_goMux_mux,Pointer_QTree_Int) > [(lizzieLet31_4Lmain_mask_Intsbos,Pointer_QTree_Int),
                                                                                                           (lizzieLet31_4Lcall_main_mask_Int3,Pointer_QTree_Int),
                                                                                                           (lizzieLet31_4Lcall_main_mask_Int2,Pointer_QTree_Int),
                                                                                                           (lizzieLet31_4Lcall_main_mask_Int1,Pointer_QTree_Int),
                                                                                                           (lizzieLet31_4Lcall_main_mask_Int0,Pointer_QTree_Int)] */
  logic [4:0] srtarg_0_2_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet31_4_d[0] && srtarg_0_2_goMux_mux_d[0]))
      unique case (lizzieLet31_4_d[3:1])
        3'd0: srtarg_0_2_goMux_mux_onehotd = 5'd1;
        3'd1: srtarg_0_2_goMux_mux_onehotd = 5'd2;
        3'd2: srtarg_0_2_goMux_mux_onehotd = 5'd4;
        3'd3: srtarg_0_2_goMux_mux_onehotd = 5'd8;
        3'd4: srtarg_0_2_goMux_mux_onehotd = 5'd16;
        default: srtarg_0_2_goMux_mux_onehotd = 5'd0;
      endcase
    else srtarg_0_2_goMux_mux_onehotd = 5'd0;
  assign lizzieLet31_4Lmain_mask_Intsbos_d = {srtarg_0_2_goMux_mux_d[16:1],
                                              srtarg_0_2_goMux_mux_onehotd[0]};
  assign lizzieLet31_4Lcall_main_mask_Int3_d = {srtarg_0_2_goMux_mux_d[16:1],
                                                srtarg_0_2_goMux_mux_onehotd[1]};
  assign lizzieLet31_4Lcall_main_mask_Int2_d = {srtarg_0_2_goMux_mux_d[16:1],
                                                srtarg_0_2_goMux_mux_onehotd[2]};
  assign lizzieLet31_4Lcall_main_mask_Int1_d = {srtarg_0_2_goMux_mux_d[16:1],
                                                srtarg_0_2_goMux_mux_onehotd[3]};
  assign lizzieLet31_4Lcall_main_mask_Int0_d = {srtarg_0_2_goMux_mux_d[16:1],
                                                srtarg_0_2_goMux_mux_onehotd[4]};
  assign srtarg_0_2_goMux_mux_r = (| (srtarg_0_2_goMux_mux_onehotd & {lizzieLet31_4Lcall_main_mask_Int0_r,
                                                                      lizzieLet31_4Lcall_main_mask_Int1_r,
                                                                      lizzieLet31_4Lcall_main_mask_Int2_r,
                                                                      lizzieLet31_4Lcall_main_mask_Int3_r,
                                                                      lizzieLet31_4Lmain_mask_Intsbos_r}));
  assign lizzieLet31_4_r = srtarg_0_2_goMux_mux_r;
  
  /* dcon (Ty QTree_Int,
      Dcon QNode_Int) : [(lizzieLet31_4Lcall_main_mask_Int0,Pointer_QTree_Int),
                         (es_1_1_destruct,Pointer_QTree_Int),
                         (es_2_2_destruct,Pointer_QTree_Int),
                         (es_3_5_destruct,Pointer_QTree_Int)] > (lizzieLet31_4Lcall_main_mask_Int0_1es_1_1_1es_2_2_1es_3_5_1QNode_Int,QTree_Int) */
  assign lizzieLet31_4Lcall_main_mask_Int0_1es_1_1_1es_2_2_1es_3_5_1QNode_Int_d = QNode_Int_dc((& {lizzieLet31_4Lcall_main_mask_Int0_d[0],
                                                                                                   es_1_1_destruct_d[0],
                                                                                                   es_2_2_destruct_d[0],
                                                                                                   es_3_5_destruct_d[0]}), lizzieLet31_4Lcall_main_mask_Int0_d, es_1_1_destruct_d, es_2_2_destruct_d, es_3_5_destruct_d);
  assign {lizzieLet31_4Lcall_main_mask_Int0_r,
          es_1_1_destruct_r,
          es_2_2_destruct_r,
          es_3_5_destruct_r} = {4 {(lizzieLet31_4Lcall_main_mask_Int0_1es_1_1_1es_2_2_1es_3_5_1QNode_Int_r && lizzieLet31_4Lcall_main_mask_Int0_1es_1_1_1es_2_2_1es_3_5_1QNode_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (lizzieLet31_4Lcall_main_mask_Int0_1es_1_1_1es_2_2_1es_3_5_1QNode_Int,QTree_Int) > (lizzieLet35_1_argbuf,QTree_Int) */
  QTree_Int_t lizzieLet31_4Lcall_main_mask_Int0_1es_1_1_1es_2_2_1es_3_5_1QNode_Int_bufchan_d;
  logic lizzieLet31_4Lcall_main_mask_Int0_1es_1_1_1es_2_2_1es_3_5_1QNode_Int_bufchan_r;
  assign lizzieLet31_4Lcall_main_mask_Int0_1es_1_1_1es_2_2_1es_3_5_1QNode_Int_r = ((! lizzieLet31_4Lcall_main_mask_Int0_1es_1_1_1es_2_2_1es_3_5_1QNode_Int_bufchan_d[0]) || lizzieLet31_4Lcall_main_mask_Int0_1es_1_1_1es_2_2_1es_3_5_1QNode_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet31_4Lcall_main_mask_Int0_1es_1_1_1es_2_2_1es_3_5_1QNode_Int_bufchan_d <= {66'd0,
                                                                                         1'd0};
    else
      if (lizzieLet31_4Lcall_main_mask_Int0_1es_1_1_1es_2_2_1es_3_5_1QNode_Int_r)
        lizzieLet31_4Lcall_main_mask_Int0_1es_1_1_1es_2_2_1es_3_5_1QNode_Int_bufchan_d <= lizzieLet31_4Lcall_main_mask_Int0_1es_1_1_1es_2_2_1es_3_5_1QNode_Int_d;
  QTree_Int_t lizzieLet31_4Lcall_main_mask_Int0_1es_1_1_1es_2_2_1es_3_5_1QNode_Int_bufchan_buf;
  assign lizzieLet31_4Lcall_main_mask_Int0_1es_1_1_1es_2_2_1es_3_5_1QNode_Int_bufchan_r = (! lizzieLet31_4Lcall_main_mask_Int0_1es_1_1_1es_2_2_1es_3_5_1QNode_Int_bufchan_buf[0]);
  assign lizzieLet35_1_argbuf_d = (lizzieLet31_4Lcall_main_mask_Int0_1es_1_1_1es_2_2_1es_3_5_1QNode_Int_bufchan_buf[0] ? lizzieLet31_4Lcall_main_mask_Int0_1es_1_1_1es_2_2_1es_3_5_1QNode_Int_bufchan_buf :
                                   lizzieLet31_4Lcall_main_mask_Int0_1es_1_1_1es_2_2_1es_3_5_1QNode_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet31_4Lcall_main_mask_Int0_1es_1_1_1es_2_2_1es_3_5_1QNode_Int_bufchan_buf <= {66'd0,
                                                                                           1'd0};
    else
      if ((lizzieLet35_1_argbuf_r && lizzieLet31_4Lcall_main_mask_Int0_1es_1_1_1es_2_2_1es_3_5_1QNode_Int_bufchan_buf[0]))
        lizzieLet31_4Lcall_main_mask_Int0_1es_1_1_1es_2_2_1es_3_5_1QNode_Int_bufchan_buf <= {66'd0,
                                                                                             1'd0};
      else if (((! lizzieLet35_1_argbuf_r) && (! lizzieLet31_4Lcall_main_mask_Int0_1es_1_1_1es_2_2_1es_3_5_1QNode_Int_bufchan_buf[0])))
        lizzieLet31_4Lcall_main_mask_Int0_1es_1_1_1es_2_2_1es_3_5_1QNode_Int_bufchan_buf <= lizzieLet31_4Lcall_main_mask_Int0_1es_1_1_1es_2_2_1es_3_5_1QNode_Int_bufchan_d;
  
  /* dcon (Ty CTmain_mask_Int,
      Dcon Lcall_main_mask_Int0) : [(lizzieLet31_4Lcall_main_mask_Int1,Pointer_QTree_Int),
                                    (es_2_1_destruct,Pointer_QTree_Int),
                                    (es_3_4_destruct,Pointer_QTree_Int),
                                    (sc_0_13_destruct,Pointer_CTmain_mask_Int)] > (lizzieLet31_4Lcall_main_mask_Int1_1es_2_1_1es_3_4_1sc_0_13_1Lcall_main_mask_Int0,CTmain_mask_Int) */
  assign lizzieLet31_4Lcall_main_mask_Int1_1es_2_1_1es_3_4_1sc_0_13_1Lcall_main_mask_Int0_d = Lcall_main_mask_Int0_dc((& {lizzieLet31_4Lcall_main_mask_Int1_d[0],
                                                                                                                          es_2_1_destruct_d[0],
                                                                                                                          es_3_4_destruct_d[0],
                                                                                                                          sc_0_13_destruct_d[0]}), lizzieLet31_4Lcall_main_mask_Int1_d, es_2_1_destruct_d, es_3_4_destruct_d, sc_0_13_destruct_d);
  assign {lizzieLet31_4Lcall_main_mask_Int1_r,
          es_2_1_destruct_r,
          es_3_4_destruct_r,
          sc_0_13_destruct_r} = {4 {(lizzieLet31_4Lcall_main_mask_Int1_1es_2_1_1es_3_4_1sc_0_13_1Lcall_main_mask_Int0_r && lizzieLet31_4Lcall_main_mask_Int1_1es_2_1_1es_3_4_1sc_0_13_1Lcall_main_mask_Int0_d[0])}};
  
  /* buf (Ty CTmain_mask_Int) : (lizzieLet31_4Lcall_main_mask_Int1_1es_2_1_1es_3_4_1sc_0_13_1Lcall_main_mask_Int0,CTmain_mask_Int) > (lizzieLet34_1_argbuf,CTmain_mask_Int) */
  CTmain_mask_Int_t lizzieLet31_4Lcall_main_mask_Int1_1es_2_1_1es_3_4_1sc_0_13_1Lcall_main_mask_Int0_bufchan_d;
  logic lizzieLet31_4Lcall_main_mask_Int1_1es_2_1_1es_3_4_1sc_0_13_1Lcall_main_mask_Int0_bufchan_r;
  assign lizzieLet31_4Lcall_main_mask_Int1_1es_2_1_1es_3_4_1sc_0_13_1Lcall_main_mask_Int0_r = ((! lizzieLet31_4Lcall_main_mask_Int1_1es_2_1_1es_3_4_1sc_0_13_1Lcall_main_mask_Int0_bufchan_d[0]) || lizzieLet31_4Lcall_main_mask_Int1_1es_2_1_1es_3_4_1sc_0_13_1Lcall_main_mask_Int0_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet31_4Lcall_main_mask_Int1_1es_2_1_1es_3_4_1sc_0_13_1Lcall_main_mask_Int0_bufchan_d <= {115'd0,
                                                                                                     1'd0};
    else
      if (lizzieLet31_4Lcall_main_mask_Int1_1es_2_1_1es_3_4_1sc_0_13_1Lcall_main_mask_Int0_r)
        lizzieLet31_4Lcall_main_mask_Int1_1es_2_1_1es_3_4_1sc_0_13_1Lcall_main_mask_Int0_bufchan_d <= lizzieLet31_4Lcall_main_mask_Int1_1es_2_1_1es_3_4_1sc_0_13_1Lcall_main_mask_Int0_d;
  CTmain_mask_Int_t lizzieLet31_4Lcall_main_mask_Int1_1es_2_1_1es_3_4_1sc_0_13_1Lcall_main_mask_Int0_bufchan_buf;
  assign lizzieLet31_4Lcall_main_mask_Int1_1es_2_1_1es_3_4_1sc_0_13_1Lcall_main_mask_Int0_bufchan_r = (! lizzieLet31_4Lcall_main_mask_Int1_1es_2_1_1es_3_4_1sc_0_13_1Lcall_main_mask_Int0_bufchan_buf[0]);
  assign lizzieLet34_1_argbuf_d = (lizzieLet31_4Lcall_main_mask_Int1_1es_2_1_1es_3_4_1sc_0_13_1Lcall_main_mask_Int0_bufchan_buf[0] ? lizzieLet31_4Lcall_main_mask_Int1_1es_2_1_1es_3_4_1sc_0_13_1Lcall_main_mask_Int0_bufchan_buf :
                                   lizzieLet31_4Lcall_main_mask_Int1_1es_2_1_1es_3_4_1sc_0_13_1Lcall_main_mask_Int0_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet31_4Lcall_main_mask_Int1_1es_2_1_1es_3_4_1sc_0_13_1Lcall_main_mask_Int0_bufchan_buf <= {115'd0,
                                                                                                       1'd0};
    else
      if ((lizzieLet34_1_argbuf_r && lizzieLet31_4Lcall_main_mask_Int1_1es_2_1_1es_3_4_1sc_0_13_1Lcall_main_mask_Int0_bufchan_buf[0]))
        lizzieLet31_4Lcall_main_mask_Int1_1es_2_1_1es_3_4_1sc_0_13_1Lcall_main_mask_Int0_bufchan_buf <= {115'd0,
                                                                                                         1'd0};
      else if (((! lizzieLet34_1_argbuf_r) && (! lizzieLet31_4Lcall_main_mask_Int1_1es_2_1_1es_3_4_1sc_0_13_1Lcall_main_mask_Int0_bufchan_buf[0])))
        lizzieLet31_4Lcall_main_mask_Int1_1es_2_1_1es_3_4_1sc_0_13_1Lcall_main_mask_Int0_bufchan_buf <= lizzieLet31_4Lcall_main_mask_Int1_1es_2_1_1es_3_4_1sc_0_13_1Lcall_main_mask_Int0_bufchan_d;
  
  /* dcon (Ty CTmain_mask_Int,
      Dcon Lcall_main_mask_Int1) : [(lizzieLet31_4Lcall_main_mask_Int2,Pointer_QTree_Int),
                                    (es_3_3_destruct,Pointer_QTree_Int),
                                    (sc_0_12_destruct,Pointer_CTmain_mask_Int),
                                    (t1a8x_2_destruct,Pointer_QTree_Int),
                                    (q1a8s_2_destruct,Pointer_MaskQTree)] > (lizzieLet31_4Lcall_main_mask_Int2_1es_3_3_1sc_0_12_1t1a8x_2_1q1a8s_2_1Lcall_main_mask_Int1,CTmain_mask_Int) */
  assign lizzieLet31_4Lcall_main_mask_Int2_1es_3_3_1sc_0_12_1t1a8x_2_1q1a8s_2_1Lcall_main_mask_Int1_d = Lcall_main_mask_Int1_dc((& {lizzieLet31_4Lcall_main_mask_Int2_d[0],
                                                                                                                                    es_3_3_destruct_d[0],
                                                                                                                                    sc_0_12_destruct_d[0],
                                                                                                                                    t1a8x_2_destruct_d[0],
                                                                                                                                    q1a8s_2_destruct_d[0]}), lizzieLet31_4Lcall_main_mask_Int2_d, es_3_3_destruct_d, sc_0_12_destruct_d, t1a8x_2_destruct_d, q1a8s_2_destruct_d);
  assign {lizzieLet31_4Lcall_main_mask_Int2_r,
          es_3_3_destruct_r,
          sc_0_12_destruct_r,
          t1a8x_2_destruct_r,
          q1a8s_2_destruct_r} = {5 {(lizzieLet31_4Lcall_main_mask_Int2_1es_3_3_1sc_0_12_1t1a8x_2_1q1a8s_2_1Lcall_main_mask_Int1_r && lizzieLet31_4Lcall_main_mask_Int2_1es_3_3_1sc_0_12_1t1a8x_2_1q1a8s_2_1Lcall_main_mask_Int1_d[0])}};
  
  /* buf (Ty CTmain_mask_Int) : (lizzieLet31_4Lcall_main_mask_Int2_1es_3_3_1sc_0_12_1t1a8x_2_1q1a8s_2_1Lcall_main_mask_Int1,CTmain_mask_Int) > (lizzieLet33_1_argbuf,CTmain_mask_Int) */
  CTmain_mask_Int_t lizzieLet31_4Lcall_main_mask_Int2_1es_3_3_1sc_0_12_1t1a8x_2_1q1a8s_2_1Lcall_main_mask_Int1_bufchan_d;
  logic lizzieLet31_4Lcall_main_mask_Int2_1es_3_3_1sc_0_12_1t1a8x_2_1q1a8s_2_1Lcall_main_mask_Int1_bufchan_r;
  assign lizzieLet31_4Lcall_main_mask_Int2_1es_3_3_1sc_0_12_1t1a8x_2_1q1a8s_2_1Lcall_main_mask_Int1_r = ((! lizzieLet31_4Lcall_main_mask_Int2_1es_3_3_1sc_0_12_1t1a8x_2_1q1a8s_2_1Lcall_main_mask_Int1_bufchan_d[0]) || lizzieLet31_4Lcall_main_mask_Int2_1es_3_3_1sc_0_12_1t1a8x_2_1q1a8s_2_1Lcall_main_mask_Int1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet31_4Lcall_main_mask_Int2_1es_3_3_1sc_0_12_1t1a8x_2_1q1a8s_2_1Lcall_main_mask_Int1_bufchan_d <= {115'd0,
                                                                                                               1'd0};
    else
      if (lizzieLet31_4Lcall_main_mask_Int2_1es_3_3_1sc_0_12_1t1a8x_2_1q1a8s_2_1Lcall_main_mask_Int1_r)
        lizzieLet31_4Lcall_main_mask_Int2_1es_3_3_1sc_0_12_1t1a8x_2_1q1a8s_2_1Lcall_main_mask_Int1_bufchan_d <= lizzieLet31_4Lcall_main_mask_Int2_1es_3_3_1sc_0_12_1t1a8x_2_1q1a8s_2_1Lcall_main_mask_Int1_d;
  CTmain_mask_Int_t lizzieLet31_4Lcall_main_mask_Int2_1es_3_3_1sc_0_12_1t1a8x_2_1q1a8s_2_1Lcall_main_mask_Int1_bufchan_buf;
  assign lizzieLet31_4Lcall_main_mask_Int2_1es_3_3_1sc_0_12_1t1a8x_2_1q1a8s_2_1Lcall_main_mask_Int1_bufchan_r = (! lizzieLet31_4Lcall_main_mask_Int2_1es_3_3_1sc_0_12_1t1a8x_2_1q1a8s_2_1Lcall_main_mask_Int1_bufchan_buf[0]);
  assign lizzieLet33_1_argbuf_d = (lizzieLet31_4Lcall_main_mask_Int2_1es_3_3_1sc_0_12_1t1a8x_2_1q1a8s_2_1Lcall_main_mask_Int1_bufchan_buf[0] ? lizzieLet31_4Lcall_main_mask_Int2_1es_3_3_1sc_0_12_1t1a8x_2_1q1a8s_2_1Lcall_main_mask_Int1_bufchan_buf :
                                   lizzieLet31_4Lcall_main_mask_Int2_1es_3_3_1sc_0_12_1t1a8x_2_1q1a8s_2_1Lcall_main_mask_Int1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet31_4Lcall_main_mask_Int2_1es_3_3_1sc_0_12_1t1a8x_2_1q1a8s_2_1Lcall_main_mask_Int1_bufchan_buf <= {115'd0,
                                                                                                                 1'd0};
    else
      if ((lizzieLet33_1_argbuf_r && lizzieLet31_4Lcall_main_mask_Int2_1es_3_3_1sc_0_12_1t1a8x_2_1q1a8s_2_1Lcall_main_mask_Int1_bufchan_buf[0]))
        lizzieLet31_4Lcall_main_mask_Int2_1es_3_3_1sc_0_12_1t1a8x_2_1q1a8s_2_1Lcall_main_mask_Int1_bufchan_buf <= {115'd0,
                                                                                                                   1'd0};
      else if (((! lizzieLet33_1_argbuf_r) && (! lizzieLet31_4Lcall_main_mask_Int2_1es_3_3_1sc_0_12_1t1a8x_2_1q1a8s_2_1Lcall_main_mask_Int1_bufchan_buf[0])))
        lizzieLet31_4Lcall_main_mask_Int2_1es_3_3_1sc_0_12_1t1a8x_2_1q1a8s_2_1Lcall_main_mask_Int1_bufchan_buf <= lizzieLet31_4Lcall_main_mask_Int2_1es_3_3_1sc_0_12_1t1a8x_2_1q1a8s_2_1Lcall_main_mask_Int1_bufchan_d;
  
  /* dcon (Ty CTmain_mask_Int,
      Dcon Lcall_main_mask_Int2) : [(lizzieLet31_4Lcall_main_mask_Int3,Pointer_QTree_Int),
                                    (sc_0_11_destruct,Pointer_CTmain_mask_Int),
                                    (t1a8x_1_destruct,Pointer_QTree_Int),
                                    (q1a8s_1_destruct,Pointer_MaskQTree),
                                    (t2a8y_1_destruct,Pointer_QTree_Int),
                                    (q2a8t_1_destruct,Pointer_MaskQTree)] > (lizzieLet31_4Lcall_main_mask_Int3_1sc_0_11_1t1a8x_1_1q1a8s_1_1t2a8y_1_1q2a8t_1_1Lcall_main_mask_Int2,CTmain_mask_Int) */
  assign lizzieLet31_4Lcall_main_mask_Int3_1sc_0_11_1t1a8x_1_1q1a8s_1_1t2a8y_1_1q2a8t_1_1Lcall_main_mask_Int2_d = Lcall_main_mask_Int2_dc((& {lizzieLet31_4Lcall_main_mask_Int3_d[0],
                                                                                                                                              sc_0_11_destruct_d[0],
                                                                                                                                              t1a8x_1_destruct_d[0],
                                                                                                                                              q1a8s_1_destruct_d[0],
                                                                                                                                              t2a8y_1_destruct_d[0],
                                                                                                                                              q2a8t_1_destruct_d[0]}), lizzieLet31_4Lcall_main_mask_Int3_d, sc_0_11_destruct_d, t1a8x_1_destruct_d, q1a8s_1_destruct_d, t2a8y_1_destruct_d, q2a8t_1_destruct_d);
  assign {lizzieLet31_4Lcall_main_mask_Int3_r,
          sc_0_11_destruct_r,
          t1a8x_1_destruct_r,
          q1a8s_1_destruct_r,
          t2a8y_1_destruct_r,
          q2a8t_1_destruct_r} = {6 {(lizzieLet31_4Lcall_main_mask_Int3_1sc_0_11_1t1a8x_1_1q1a8s_1_1t2a8y_1_1q2a8t_1_1Lcall_main_mask_Int2_r && lizzieLet31_4Lcall_main_mask_Int3_1sc_0_11_1t1a8x_1_1q1a8s_1_1t2a8y_1_1q2a8t_1_1Lcall_main_mask_Int2_d[0])}};
  
  /* buf (Ty CTmain_mask_Int) : (lizzieLet31_4Lcall_main_mask_Int3_1sc_0_11_1t1a8x_1_1q1a8s_1_1t2a8y_1_1q2a8t_1_1Lcall_main_mask_Int2,CTmain_mask_Int) > (lizzieLet32_1_argbuf,CTmain_mask_Int) */
  CTmain_mask_Int_t lizzieLet31_4Lcall_main_mask_Int3_1sc_0_11_1t1a8x_1_1q1a8s_1_1t2a8y_1_1q2a8t_1_1Lcall_main_mask_Int2_bufchan_d;
  logic lizzieLet31_4Lcall_main_mask_Int3_1sc_0_11_1t1a8x_1_1q1a8s_1_1t2a8y_1_1q2a8t_1_1Lcall_main_mask_Int2_bufchan_r;
  assign lizzieLet31_4Lcall_main_mask_Int3_1sc_0_11_1t1a8x_1_1q1a8s_1_1t2a8y_1_1q2a8t_1_1Lcall_main_mask_Int2_r = ((! lizzieLet31_4Lcall_main_mask_Int3_1sc_0_11_1t1a8x_1_1q1a8s_1_1t2a8y_1_1q2a8t_1_1Lcall_main_mask_Int2_bufchan_d[0]) || lizzieLet31_4Lcall_main_mask_Int3_1sc_0_11_1t1a8x_1_1q1a8s_1_1t2a8y_1_1q2a8t_1_1Lcall_main_mask_Int2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet31_4Lcall_main_mask_Int3_1sc_0_11_1t1a8x_1_1q1a8s_1_1t2a8y_1_1q2a8t_1_1Lcall_main_mask_Int2_bufchan_d <= {115'd0,
                                                                                                                         1'd0};
    else
      if (lizzieLet31_4Lcall_main_mask_Int3_1sc_0_11_1t1a8x_1_1q1a8s_1_1t2a8y_1_1q2a8t_1_1Lcall_main_mask_Int2_r)
        lizzieLet31_4Lcall_main_mask_Int3_1sc_0_11_1t1a8x_1_1q1a8s_1_1t2a8y_1_1q2a8t_1_1Lcall_main_mask_Int2_bufchan_d <= lizzieLet31_4Lcall_main_mask_Int3_1sc_0_11_1t1a8x_1_1q1a8s_1_1t2a8y_1_1q2a8t_1_1Lcall_main_mask_Int2_d;
  CTmain_mask_Int_t lizzieLet31_4Lcall_main_mask_Int3_1sc_0_11_1t1a8x_1_1q1a8s_1_1t2a8y_1_1q2a8t_1_1Lcall_main_mask_Int2_bufchan_buf;
  assign lizzieLet31_4Lcall_main_mask_Int3_1sc_0_11_1t1a8x_1_1q1a8s_1_1t2a8y_1_1q2a8t_1_1Lcall_main_mask_Int2_bufchan_r = (! lizzieLet31_4Lcall_main_mask_Int3_1sc_0_11_1t1a8x_1_1q1a8s_1_1t2a8y_1_1q2a8t_1_1Lcall_main_mask_Int2_bufchan_buf[0]);
  assign lizzieLet32_1_argbuf_d = (lizzieLet31_4Lcall_main_mask_Int3_1sc_0_11_1t1a8x_1_1q1a8s_1_1t2a8y_1_1q2a8t_1_1Lcall_main_mask_Int2_bufchan_buf[0] ? lizzieLet31_4Lcall_main_mask_Int3_1sc_0_11_1t1a8x_1_1q1a8s_1_1t2a8y_1_1q2a8t_1_1Lcall_main_mask_Int2_bufchan_buf :
                                   lizzieLet31_4Lcall_main_mask_Int3_1sc_0_11_1t1a8x_1_1q1a8s_1_1t2a8y_1_1q2a8t_1_1Lcall_main_mask_Int2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet31_4Lcall_main_mask_Int3_1sc_0_11_1t1a8x_1_1q1a8s_1_1t2a8y_1_1q2a8t_1_1Lcall_main_mask_Int2_bufchan_buf <= {115'd0,
                                                                                                                           1'd0};
    else
      if ((lizzieLet32_1_argbuf_r && lizzieLet31_4Lcall_main_mask_Int3_1sc_0_11_1t1a8x_1_1q1a8s_1_1t2a8y_1_1q2a8t_1_1Lcall_main_mask_Int2_bufchan_buf[0]))
        lizzieLet31_4Lcall_main_mask_Int3_1sc_0_11_1t1a8x_1_1q1a8s_1_1t2a8y_1_1q2a8t_1_1Lcall_main_mask_Int2_bufchan_buf <= {115'd0,
                                                                                                                             1'd0};
      else if (((! lizzieLet32_1_argbuf_r) && (! lizzieLet31_4Lcall_main_mask_Int3_1sc_0_11_1t1a8x_1_1q1a8s_1_1t2a8y_1_1q2a8t_1_1Lcall_main_mask_Int2_bufchan_buf[0])))
        lizzieLet31_4Lcall_main_mask_Int3_1sc_0_11_1t1a8x_1_1q1a8s_1_1t2a8y_1_1q2a8t_1_1Lcall_main_mask_Int2_bufchan_buf <= lizzieLet31_4Lcall_main_mask_Int3_1sc_0_11_1t1a8x_1_1q1a8s_1_1t2a8y_1_1q2a8t_1_1Lcall_main_mask_Int2_bufchan_d;
  
  /* fork (Ty Pointer_QTree_Int) : (lizzieLet31_4Lmain_mask_Intsbos,Pointer_QTree_Int) > [(lizzieLet31_4Lmain_mask_Intsbos_1_merge_merge_fork_1,Pointer_QTree_Int),
                                                                                     (lizzieLet31_4Lmain_mask_Intsbos_1_merge_merge_fork_2,Pointer_QTree_Int)] */
  logic [1:0] lizzieLet31_4Lmain_mask_Intsbos_emitted;
  logic [1:0] lizzieLet31_4Lmain_mask_Intsbos_done;
  assign lizzieLet31_4Lmain_mask_Intsbos_1_merge_merge_fork_1_d = {lizzieLet31_4Lmain_mask_Intsbos_d[16:1],
                                                                   (lizzieLet31_4Lmain_mask_Intsbos_d[0] && (! lizzieLet31_4Lmain_mask_Intsbos_emitted[0]))};
  assign lizzieLet31_4Lmain_mask_Intsbos_1_merge_merge_fork_2_d = {lizzieLet31_4Lmain_mask_Intsbos_d[16:1],
                                                                   (lizzieLet31_4Lmain_mask_Intsbos_d[0] && (! lizzieLet31_4Lmain_mask_Intsbos_emitted[1]))};
  assign lizzieLet31_4Lmain_mask_Intsbos_done = (lizzieLet31_4Lmain_mask_Intsbos_emitted | ({lizzieLet31_4Lmain_mask_Intsbos_1_merge_merge_fork_2_d[0],
                                                                                             lizzieLet31_4Lmain_mask_Intsbos_1_merge_merge_fork_1_d[0]} & {lizzieLet31_4Lmain_mask_Intsbos_1_merge_merge_fork_2_r,
                                                                                                                                                           lizzieLet31_4Lmain_mask_Intsbos_1_merge_merge_fork_1_r}));
  assign lizzieLet31_4Lmain_mask_Intsbos_r = (& lizzieLet31_4Lmain_mask_Intsbos_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet31_4Lmain_mask_Intsbos_emitted <= 2'd0;
    else
      lizzieLet31_4Lmain_mask_Intsbos_emitted <= (lizzieLet31_4Lmain_mask_Intsbos_r ? 2'd0 :
                                                  lizzieLet31_4Lmain_mask_Intsbos_done);
  
  /* togo (Ty Pointer_QTree_Int) : (lizzieLet31_4Lmain_mask_Intsbos_1_merge_merge_fork_1,Pointer_QTree_Int) > (call_main_mask_Int_goConst,Go) */
  assign call_main_mask_Int_goConst_d = lizzieLet31_4Lmain_mask_Intsbos_1_merge_merge_fork_1_d[0];
  assign lizzieLet31_4Lmain_mask_Intsbos_1_merge_merge_fork_1_r = call_main_mask_Int_goConst_r;
  
  /* buf (Ty Pointer_QTree_Int) : (lizzieLet31_4Lmain_mask_Intsbos_1_merge_merge_fork_2,Pointer_QTree_Int) > (main_mask_Int_resbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t lizzieLet31_4Lmain_mask_Intsbos_1_merge_merge_fork_2_bufchan_d;
  logic lizzieLet31_4Lmain_mask_Intsbos_1_merge_merge_fork_2_bufchan_r;
  assign lizzieLet31_4Lmain_mask_Intsbos_1_merge_merge_fork_2_r = ((! lizzieLet31_4Lmain_mask_Intsbos_1_merge_merge_fork_2_bufchan_d[0]) || lizzieLet31_4Lmain_mask_Intsbos_1_merge_merge_fork_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet31_4Lmain_mask_Intsbos_1_merge_merge_fork_2_bufchan_d <= {16'd0,
                                                                         1'd0};
    else
      if (lizzieLet31_4Lmain_mask_Intsbos_1_merge_merge_fork_2_r)
        lizzieLet31_4Lmain_mask_Intsbos_1_merge_merge_fork_2_bufchan_d <= lizzieLet31_4Lmain_mask_Intsbos_1_merge_merge_fork_2_d;
  Pointer_QTree_Int_t lizzieLet31_4Lmain_mask_Intsbos_1_merge_merge_fork_2_bufchan_buf;
  assign lizzieLet31_4Lmain_mask_Intsbos_1_merge_merge_fork_2_bufchan_r = (! lizzieLet31_4Lmain_mask_Intsbos_1_merge_merge_fork_2_bufchan_buf[0]);
  assign main_mask_Int_resbuf_d = (lizzieLet31_4Lmain_mask_Intsbos_1_merge_merge_fork_2_bufchan_buf[0] ? lizzieLet31_4Lmain_mask_Intsbos_1_merge_merge_fork_2_bufchan_buf :
                                   lizzieLet31_4Lmain_mask_Intsbos_1_merge_merge_fork_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet31_4Lmain_mask_Intsbos_1_merge_merge_fork_2_bufchan_buf <= {16'd0,
                                                                           1'd0};
    else
      if ((main_mask_Int_resbuf_r && lizzieLet31_4Lmain_mask_Intsbos_1_merge_merge_fork_2_bufchan_buf[0]))
        lizzieLet31_4Lmain_mask_Intsbos_1_merge_merge_fork_2_bufchan_buf <= {16'd0,
                                                                             1'd0};
      else if (((! main_mask_Int_resbuf_r) && (! lizzieLet31_4Lmain_mask_Intsbos_1_merge_merge_fork_2_bufchan_buf[0])))
        lizzieLet31_4Lmain_mask_Intsbos_1_merge_merge_fork_2_bufchan_buf <= lizzieLet31_4Lmain_mask_Intsbos_1_merge_merge_fork_2_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (ma8q_1,Pointer_QTree_Int) > (ma8q_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t ma8q_1_bufchan_d;
  logic ma8q_1_bufchan_r;
  assign ma8q_1_r = ((! ma8q_1_bufchan_d[0]) || ma8q_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) ma8q_1_bufchan_d <= {16'd0, 1'd0};
    else if (ma8q_1_r) ma8q_1_bufchan_d <= ma8q_1_d;
  Pointer_QTree_Int_t ma8q_1_bufchan_buf;
  assign ma8q_1_bufchan_r = (! ma8q_1_bufchan_buf[0]);
  assign ma8q_1_argbuf_d = (ma8q_1_bufchan_buf[0] ? ma8q_1_bufchan_buf :
                            ma8q_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) ma8q_1_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((ma8q_1_argbuf_r && ma8q_1_bufchan_buf[0]))
        ma8q_1_bufchan_buf <= {16'd0, 1'd0};
      else if (((! ma8q_1_argbuf_r) && (! ma8q_1_bufchan_buf[0])))
        ma8q_1_bufchan_buf <= ma8q_1_bufchan_d;
  
  /* fork (Ty Pointer_QTree_Int) : (ma8q_goMux_mux,Pointer_QTree_Int) > [(ma8q_1,Pointer_QTree_Int),
                                                                    (ma8q_2,Pointer_QTree_Int)] */
  logic [1:0] ma8q_goMux_mux_emitted;
  logic [1:0] ma8q_goMux_mux_done;
  assign ma8q_1_d = {ma8q_goMux_mux_d[16:1],
                     (ma8q_goMux_mux_d[0] && (! ma8q_goMux_mux_emitted[0]))};
  assign ma8q_2_d = {ma8q_goMux_mux_d[16:1],
                     (ma8q_goMux_mux_d[0] && (! ma8q_goMux_mux_emitted[1]))};
  assign ma8q_goMux_mux_done = (ma8q_goMux_mux_emitted | ({ma8q_2_d[0],
                                                           ma8q_1_d[0]} & {ma8q_2_r, ma8q_1_r}));
  assign ma8q_goMux_mux_r = (& ma8q_goMux_mux_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) ma8q_goMux_mux_emitted <= 2'd0;
    else
      ma8q_goMux_mux_emitted <= (ma8q_goMux_mux_r ? 2'd0 :
                                 ma8q_goMux_mux_done);
  
  /* destruct (Ty TupGo___Pointer_QTree_Int___Pointer_MaskQTree,
          Dcon TupGo___Pointer_QTree_Int___Pointer_MaskQTree) : (main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree_1,TupGo___Pointer_QTree_Int___Pointer_MaskQTree) > [(main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreego_9,Go),
                                                                                                                                                                                (main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreema8q_1,Pointer_QTree_Int),
                                                                                                                                                                                (main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreemska8r_1,Pointer_MaskQTree)] */
  logic [2:0] main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree_1_emitted;
  logic [2:0] main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree_1_done;
  assign main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreego_9_d = (main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree_1_d[0] && (! main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree_1_emitted[0]));
  assign main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreema8q_1_d = {main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree_1_d[16:1],
                                                                               (main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree_1_d[0] && (! main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree_1_emitted[1]))};
  assign main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreemska8r_1_d = {main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree_1_d[32:17],
                                                                                 (main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree_1_d[0] && (! main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree_1_emitted[2]))};
  assign main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree_1_done = (main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree_1_emitted | ({main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreemska8r_1_d[0],
                                                                                                                                                       main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreema8q_1_d[0],
                                                                                                                                                       main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreego_9_d[0]} & {main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreemska8r_1_r,
                                                                                                                                                                                                                               main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreema8q_1_r,
                                                                                                                                                                                                                               main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreego_9_r}));
  assign main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree_1_r = (& main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree_1_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree_1_emitted <= 3'd0;
    else
      main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree_1_emitted <= (main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree_1_r ? 3'd0 :
                                                                               main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree_1_done);
  
  /* fork (Ty Go) : (main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreego_9,Go) > [(go_9_1,Go),
                                                                                      (go_9_2,Go)] */
  logic [1:0] main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreego_9_emitted;
  logic [1:0] main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreego_9_done;
  assign go_9_1_d = (main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreego_9_d[0] && (! main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreego_9_emitted[0]));
  assign go_9_2_d = (main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreego_9_d[0] && (! main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreego_9_emitted[1]));
  assign main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreego_9_done = (main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreego_9_emitted | ({go_9_2_d[0],
                                                                                                                                                           go_9_1_d[0]} & {go_9_2_r,
                                                                                                                                                                           go_9_1_r}));
  assign main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreego_9_r = (& main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreego_9_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreego_9_emitted <= 2'd0;
    else
      main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreego_9_emitted <= (main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreego_9_r ? 2'd0 :
                                                                                 main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreego_9_done);
  
  /* buf (Ty Pointer_QTree_Int) : (main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreema8q_1,Pointer_QTree_Int) > (ma8q_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreema8q_1_bufchan_d;
  logic main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreema8q_1_bufchan_r;
  assign main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreema8q_1_r = ((! main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreema8q_1_bufchan_d[0]) || main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreema8q_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreema8q_1_bufchan_d <= {16'd0,
                                                                                     1'd0};
    else
      if (main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreema8q_1_r)
        main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreema8q_1_bufchan_d <= main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreema8q_1_d;
  Pointer_QTree_Int_t main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreema8q_1_bufchan_buf;
  assign main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreema8q_1_bufchan_r = (! main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreema8q_1_bufchan_buf[0]);
  assign ma8q_1_1_argbuf_d = (main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreema8q_1_bufchan_buf[0] ? main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreema8q_1_bufchan_buf :
                              main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreema8q_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreema8q_1_bufchan_buf <= {16'd0,
                                                                                       1'd0};
    else
      if ((ma8q_1_1_argbuf_r && main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreema8q_1_bufchan_buf[0]))
        main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreema8q_1_bufchan_buf <= {16'd0,
                                                                                         1'd0};
      else if (((! ma8q_1_1_argbuf_r) && (! main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreema8q_1_bufchan_buf[0])))
        main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreema8q_1_bufchan_buf <= main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreema8q_1_bufchan_d;
  
  /* buf (Ty Pointer_MaskQTree) : (main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreemska8r_1,Pointer_MaskQTree) > (mska8r_1_1_argbuf,Pointer_MaskQTree) */
  Pointer_MaskQTree_t main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreemska8r_1_bufchan_d;
  logic main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreemska8r_1_bufchan_r;
  assign main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreemska8r_1_r = ((! main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreemska8r_1_bufchan_d[0]) || main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreemska8r_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreemska8r_1_bufchan_d <= {16'd0,
                                                                                       1'd0};
    else
      if (main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreemska8r_1_r)
        main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreemska8r_1_bufchan_d <= main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreemska8r_1_d;
  Pointer_MaskQTree_t main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreemska8r_1_bufchan_buf;
  assign main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreemska8r_1_bufchan_r = (! main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreemska8r_1_bufchan_buf[0]);
  assign mska8r_1_1_argbuf_d = (main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreemska8r_1_bufchan_buf[0] ? main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreemska8r_1_bufchan_buf :
                                main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreemska8r_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreemska8r_1_bufchan_buf <= {16'd0,
                                                                                         1'd0};
    else
      if ((mska8r_1_1_argbuf_r && main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreemska8r_1_bufchan_buf[0]))
        main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreemska8r_1_bufchan_buf <= {16'd0,
                                                                                           1'd0};
      else if (((! mska8r_1_1_argbuf_r) && (! main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreemska8r_1_bufchan_buf[0])))
        main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreemska8r_1_bufchan_buf <= main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreemska8r_1_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (main_mask_Int_resbuf,Pointer_QTree_Int) > (es_0_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t main_mask_Int_resbuf_bufchan_d;
  logic main_mask_Int_resbuf_bufchan_r;
  assign main_mask_Int_resbuf_r = ((! main_mask_Int_resbuf_bufchan_d[0]) || main_mask_Int_resbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      main_mask_Int_resbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (main_mask_Int_resbuf_r)
        main_mask_Int_resbuf_bufchan_d <= main_mask_Int_resbuf_d;
  Pointer_QTree_Int_t main_mask_Int_resbuf_bufchan_buf;
  assign main_mask_Int_resbuf_bufchan_r = (! main_mask_Int_resbuf_bufchan_buf[0]);
  assign es_0_1_argbuf_d = (main_mask_Int_resbuf_bufchan_buf[0] ? main_mask_Int_resbuf_bufchan_buf :
                            main_mask_Int_resbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      main_mask_Int_resbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((es_0_1_argbuf_r && main_mask_Int_resbuf_bufchan_buf[0]))
        main_mask_Int_resbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! es_0_1_argbuf_r) && (! main_mask_Int_resbuf_bufchan_buf[0])))
        main_mask_Int_resbuf_bufchan_buf <= main_mask_Int_resbuf_bufchan_d;
  
  /* buf (Ty Pointer_MaskQTree) : (mska8r_goMux_mux,Pointer_MaskQTree) > (mska8r_1_argbuf,Pointer_MaskQTree) */
  Pointer_MaskQTree_t mska8r_goMux_mux_bufchan_d;
  logic mska8r_goMux_mux_bufchan_r;
  assign mska8r_goMux_mux_r = ((! mska8r_goMux_mux_bufchan_d[0]) || mska8r_goMux_mux_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mska8r_goMux_mux_bufchan_d <= {16'd0, 1'd0};
    else
      if (mska8r_goMux_mux_r)
        mska8r_goMux_mux_bufchan_d <= mska8r_goMux_mux_d;
  Pointer_MaskQTree_t mska8r_goMux_mux_bufchan_buf;
  assign mska8r_goMux_mux_bufchan_r = (! mska8r_goMux_mux_bufchan_buf[0]);
  assign mska8r_1_argbuf_d = (mska8r_goMux_mux_bufchan_buf[0] ? mska8r_goMux_mux_bufchan_buf :
                              mska8r_goMux_mux_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mska8r_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((mska8r_1_argbuf_r && mska8r_goMux_mux_bufchan_buf[0]))
        mska8r_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
      else if (((! mska8r_1_argbuf_r) && (! mska8r_goMux_mux_bufchan_buf[0])))
        mska8r_goMux_mux_bufchan_buf <= mska8r_goMux_mux_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (q1a8C_destruct,Pointer_QTree_Int) > (q1a8C_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t q1a8C_destruct_bufchan_d;
  logic q1a8C_destruct_bufchan_r;
  assign q1a8C_destruct_r = ((! q1a8C_destruct_bufchan_d[0]) || q1a8C_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q1a8C_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q1a8C_destruct_r) q1a8C_destruct_bufchan_d <= q1a8C_destruct_d;
  Pointer_QTree_Int_t q1a8C_destruct_bufchan_buf;
  assign q1a8C_destruct_bufchan_r = (! q1a8C_destruct_bufchan_buf[0]);
  assign q1a8C_1_argbuf_d = (q1a8C_destruct_bufchan_buf[0] ? q1a8C_destruct_bufchan_buf :
                             q1a8C_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q1a8C_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q1a8C_1_argbuf_r && q1a8C_destruct_bufchan_buf[0]))
        q1a8C_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q1a8C_1_argbuf_r) && (! q1a8C_destruct_bufchan_buf[0])))
        q1a8C_destruct_bufchan_buf <= q1a8C_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (q1a8h_3_destruct,Pointer_QTree_Int) > (q1a8h_3_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t q1a8h_3_destruct_bufchan_d;
  logic q1a8h_3_destruct_bufchan_r;
  assign q1a8h_3_destruct_r = ((! q1a8h_3_destruct_bufchan_d[0]) || q1a8h_3_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q1a8h_3_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q1a8h_3_destruct_r)
        q1a8h_3_destruct_bufchan_d <= q1a8h_3_destruct_d;
  Pointer_QTree_Int_t q1a8h_3_destruct_bufchan_buf;
  assign q1a8h_3_destruct_bufchan_r = (! q1a8h_3_destruct_bufchan_buf[0]);
  assign q1a8h_3_1_argbuf_d = (q1a8h_3_destruct_bufchan_buf[0] ? q1a8h_3_destruct_bufchan_buf :
                               q1a8h_3_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q1a8h_3_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q1a8h_3_1_argbuf_r && q1a8h_3_destruct_bufchan_buf[0]))
        q1a8h_3_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q1a8h_3_1_argbuf_r) && (! q1a8h_3_destruct_bufchan_buf[0])))
        q1a8h_3_destruct_bufchan_buf <= q1a8h_3_destruct_bufchan_d;
  
  /* buf (Ty Pointer_MaskQTree) : (q1a8s_3_destruct,Pointer_MaskQTree) > (q1a8s_3_1_argbuf,Pointer_MaskQTree) */
  Pointer_MaskQTree_t q1a8s_3_destruct_bufchan_d;
  logic q1a8s_3_destruct_bufchan_r;
  assign q1a8s_3_destruct_r = ((! q1a8s_3_destruct_bufchan_d[0]) || q1a8s_3_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q1a8s_3_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q1a8s_3_destruct_r)
        q1a8s_3_destruct_bufchan_d <= q1a8s_3_destruct_d;
  Pointer_MaskQTree_t q1a8s_3_destruct_bufchan_buf;
  assign q1a8s_3_destruct_bufchan_r = (! q1a8s_3_destruct_bufchan_buf[0]);
  assign q1a8s_3_1_argbuf_d = (q1a8s_3_destruct_bufchan_buf[0] ? q1a8s_3_destruct_bufchan_buf :
                               q1a8s_3_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q1a8s_3_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q1a8s_3_1_argbuf_r && q1a8s_3_destruct_bufchan_buf[0]))
        q1a8s_3_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q1a8s_3_1_argbuf_r) && (! q1a8s_3_destruct_bufchan_buf[0])))
        q1a8s_3_destruct_bufchan_buf <= q1a8s_3_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (q2a8D_1_destruct,Pointer_QTree_Int) > (q2a8D_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t q2a8D_1_destruct_bufchan_d;
  logic q2a8D_1_destruct_bufchan_r;
  assign q2a8D_1_destruct_r = ((! q2a8D_1_destruct_bufchan_d[0]) || q2a8D_1_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q2a8D_1_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q2a8D_1_destruct_r)
        q2a8D_1_destruct_bufchan_d <= q2a8D_1_destruct_d;
  Pointer_QTree_Int_t q2a8D_1_destruct_bufchan_buf;
  assign q2a8D_1_destruct_bufchan_r = (! q2a8D_1_destruct_bufchan_buf[0]);
  assign q2a8D_1_1_argbuf_d = (q2a8D_1_destruct_bufchan_buf[0] ? q2a8D_1_destruct_bufchan_buf :
                               q2a8D_1_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q2a8D_1_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q2a8D_1_1_argbuf_r && q2a8D_1_destruct_bufchan_buf[0]))
        q2a8D_1_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q2a8D_1_1_argbuf_r) && (! q2a8D_1_destruct_bufchan_buf[0])))
        q2a8D_1_destruct_bufchan_buf <= q2a8D_1_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (q2a8i_2_destruct,Pointer_QTree_Int) > (q2a8i_2_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t q2a8i_2_destruct_bufchan_d;
  logic q2a8i_2_destruct_bufchan_r;
  assign q2a8i_2_destruct_r = ((! q2a8i_2_destruct_bufchan_d[0]) || q2a8i_2_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q2a8i_2_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q2a8i_2_destruct_r)
        q2a8i_2_destruct_bufchan_d <= q2a8i_2_destruct_d;
  Pointer_QTree_Int_t q2a8i_2_destruct_bufchan_buf;
  assign q2a8i_2_destruct_bufchan_r = (! q2a8i_2_destruct_bufchan_buf[0]);
  assign q2a8i_2_1_argbuf_d = (q2a8i_2_destruct_bufchan_buf[0] ? q2a8i_2_destruct_bufchan_buf :
                               q2a8i_2_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q2a8i_2_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q2a8i_2_1_argbuf_r && q2a8i_2_destruct_bufchan_buf[0]))
        q2a8i_2_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q2a8i_2_1_argbuf_r) && (! q2a8i_2_destruct_bufchan_buf[0])))
        q2a8i_2_destruct_bufchan_buf <= q2a8i_2_destruct_bufchan_d;
  
  /* buf (Ty Pointer_MaskQTree) : (q2a8t_2_destruct,Pointer_MaskQTree) > (q2a8t_2_1_argbuf,Pointer_MaskQTree) */
  Pointer_MaskQTree_t q2a8t_2_destruct_bufchan_d;
  logic q2a8t_2_destruct_bufchan_r;
  assign q2a8t_2_destruct_r = ((! q2a8t_2_destruct_bufchan_d[0]) || q2a8t_2_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q2a8t_2_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q2a8t_2_destruct_r)
        q2a8t_2_destruct_bufchan_d <= q2a8t_2_destruct_d;
  Pointer_MaskQTree_t q2a8t_2_destruct_bufchan_buf;
  assign q2a8t_2_destruct_bufchan_r = (! q2a8t_2_destruct_bufchan_buf[0]);
  assign q2a8t_2_1_argbuf_d = (q2a8t_2_destruct_bufchan_buf[0] ? q2a8t_2_destruct_bufchan_buf :
                               q2a8t_2_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q2a8t_2_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q2a8t_2_1_argbuf_r && q2a8t_2_destruct_bufchan_buf[0]))
        q2a8t_2_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q2a8t_2_1_argbuf_r) && (! q2a8t_2_destruct_bufchan_buf[0])))
        q2a8t_2_destruct_bufchan_buf <= q2a8t_2_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (q3a8E_2_destruct,Pointer_QTree_Int) > (q3a8E_2_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t q3a8E_2_destruct_bufchan_d;
  logic q3a8E_2_destruct_bufchan_r;
  assign q3a8E_2_destruct_r = ((! q3a8E_2_destruct_bufchan_d[0]) || q3a8E_2_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q3a8E_2_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q3a8E_2_destruct_r)
        q3a8E_2_destruct_bufchan_d <= q3a8E_2_destruct_d;
  Pointer_QTree_Int_t q3a8E_2_destruct_bufchan_buf;
  assign q3a8E_2_destruct_bufchan_r = (! q3a8E_2_destruct_bufchan_buf[0]);
  assign q3a8E_2_1_argbuf_d = (q3a8E_2_destruct_bufchan_buf[0] ? q3a8E_2_destruct_bufchan_buf :
                               q3a8E_2_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q3a8E_2_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q3a8E_2_1_argbuf_r && q3a8E_2_destruct_bufchan_buf[0]))
        q3a8E_2_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q3a8E_2_1_argbuf_r) && (! q3a8E_2_destruct_bufchan_buf[0])))
        q3a8E_2_destruct_bufchan_buf <= q3a8E_2_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (q3a8j_1_destruct,Pointer_QTree_Int) > (q3a8j_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t q3a8j_1_destruct_bufchan_d;
  logic q3a8j_1_destruct_bufchan_r;
  assign q3a8j_1_destruct_r = ((! q3a8j_1_destruct_bufchan_d[0]) || q3a8j_1_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q3a8j_1_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q3a8j_1_destruct_r)
        q3a8j_1_destruct_bufchan_d <= q3a8j_1_destruct_d;
  Pointer_QTree_Int_t q3a8j_1_destruct_bufchan_buf;
  assign q3a8j_1_destruct_bufchan_r = (! q3a8j_1_destruct_bufchan_buf[0]);
  assign q3a8j_1_1_argbuf_d = (q3a8j_1_destruct_bufchan_buf[0] ? q3a8j_1_destruct_bufchan_buf :
                               q3a8j_1_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q3a8j_1_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q3a8j_1_1_argbuf_r && q3a8j_1_destruct_bufchan_buf[0]))
        q3a8j_1_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q3a8j_1_1_argbuf_r) && (! q3a8j_1_destruct_bufchan_buf[0])))
        q3a8j_1_destruct_bufchan_buf <= q3a8j_1_destruct_bufchan_d;
  
  /* buf (Ty Pointer_MaskQTree) : (q3a8u_1_destruct,Pointer_MaskQTree) > (q3a8u_1_1_argbuf,Pointer_MaskQTree) */
  Pointer_MaskQTree_t q3a8u_1_destruct_bufchan_d;
  logic q3a8u_1_destruct_bufchan_r;
  assign q3a8u_1_destruct_r = ((! q3a8u_1_destruct_bufchan_d[0]) || q3a8u_1_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q3a8u_1_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q3a8u_1_destruct_r)
        q3a8u_1_destruct_bufchan_d <= q3a8u_1_destruct_d;
  Pointer_MaskQTree_t q3a8u_1_destruct_bufchan_buf;
  assign q3a8u_1_destruct_bufchan_r = (! q3a8u_1_destruct_bufchan_buf[0]);
  assign q3a8u_1_1_argbuf_d = (q3a8u_1_destruct_bufchan_buf[0] ? q3a8u_1_destruct_bufchan_buf :
                               q3a8u_1_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q3a8u_1_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q3a8u_1_1_argbuf_r && q3a8u_1_destruct_bufchan_buf[0]))
        q3a8u_1_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q3a8u_1_1_argbuf_r) && (! q3a8u_1_destruct_bufchan_buf[0])))
        q3a8u_1_destruct_bufchan_buf <= q3a8u_1_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (q4a8F_3_destruct,Pointer_QTree_Int) > (q4a8F_3_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t q4a8F_3_destruct_bufchan_d;
  logic q4a8F_3_destruct_bufchan_r;
  assign q4a8F_3_destruct_r = ((! q4a8F_3_destruct_bufchan_d[0]) || q4a8F_3_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q4a8F_3_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q4a8F_3_destruct_r)
        q4a8F_3_destruct_bufchan_d <= q4a8F_3_destruct_d;
  Pointer_QTree_Int_t q4a8F_3_destruct_bufchan_buf;
  assign q4a8F_3_destruct_bufchan_r = (! q4a8F_3_destruct_bufchan_buf[0]);
  assign q4a8F_3_1_argbuf_d = (q4a8F_3_destruct_bufchan_buf[0] ? q4a8F_3_destruct_bufchan_buf :
                               q4a8F_3_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q4a8F_3_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q4a8F_3_1_argbuf_r && q4a8F_3_destruct_bufchan_buf[0]))
        q4a8F_3_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q4a8F_3_1_argbuf_r) && (! q4a8F_3_destruct_bufchan_buf[0])))
        q4a8F_3_destruct_bufchan_buf <= q4a8F_3_destruct_bufchan_d;
  
  /* buf (Ty CT$wmAdd_Int) : (readPointer_CT$wmAdd_Intscfarg_0_1_argbuf,CT$wmAdd_Int) > (readPointer_CT$wmAdd_Intscfarg_0_1_argbuf_rwb,CT$wmAdd_Int) */
  CT$wmAdd_Int_t readPointer_CT$wmAdd_Intscfarg_0_1_argbuf_bufchan_d;
  logic readPointer_CT$wmAdd_Intscfarg_0_1_argbuf_bufchan_r;
  assign readPointer_CT$wmAdd_Intscfarg_0_1_argbuf_r = ((! readPointer_CT$wmAdd_Intscfarg_0_1_argbuf_bufchan_d[0]) || readPointer_CT$wmAdd_Intscfarg_0_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_CT$wmAdd_Intscfarg_0_1_argbuf_bufchan_d <= {115'd0,
                                                              1'd0};
    else
      if (readPointer_CT$wmAdd_Intscfarg_0_1_argbuf_r)
        readPointer_CT$wmAdd_Intscfarg_0_1_argbuf_bufchan_d <= readPointer_CT$wmAdd_Intscfarg_0_1_argbuf_d;
  CT$wmAdd_Int_t readPointer_CT$wmAdd_Intscfarg_0_1_argbuf_bufchan_buf;
  assign readPointer_CT$wmAdd_Intscfarg_0_1_argbuf_bufchan_r = (! readPointer_CT$wmAdd_Intscfarg_0_1_argbuf_bufchan_buf[0]);
  assign readPointer_CT$wmAdd_Intscfarg_0_1_argbuf_rwb_d = (readPointer_CT$wmAdd_Intscfarg_0_1_argbuf_bufchan_buf[0] ? readPointer_CT$wmAdd_Intscfarg_0_1_argbuf_bufchan_buf :
                                                            readPointer_CT$wmAdd_Intscfarg_0_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_CT$wmAdd_Intscfarg_0_1_argbuf_bufchan_buf <= {115'd0,
                                                                1'd0};
    else
      if ((readPointer_CT$wmAdd_Intscfarg_0_1_argbuf_rwb_r && readPointer_CT$wmAdd_Intscfarg_0_1_argbuf_bufchan_buf[0]))
        readPointer_CT$wmAdd_Intscfarg_0_1_argbuf_bufchan_buf <= {115'd0,
                                                                  1'd0};
      else if (((! readPointer_CT$wmAdd_Intscfarg_0_1_argbuf_rwb_r) && (! readPointer_CT$wmAdd_Intscfarg_0_1_argbuf_bufchan_buf[0])))
        readPointer_CT$wmAdd_Intscfarg_0_1_argbuf_bufchan_buf <= readPointer_CT$wmAdd_Intscfarg_0_1_argbuf_bufchan_d;
  
  /* fork (Ty CT$wmAdd_Int) : (readPointer_CT$wmAdd_Intscfarg_0_1_argbuf_rwb,CT$wmAdd_Int) > [(lizzieLet22_1,CT$wmAdd_Int),
                                                                                         (lizzieLet22_2,CT$wmAdd_Int),
                                                                                         (lizzieLet22_3,CT$wmAdd_Int),
                                                                                         (lizzieLet22_4,CT$wmAdd_Int)] */
  logic [3:0] readPointer_CT$wmAdd_Intscfarg_0_1_argbuf_rwb_emitted;
  logic [3:0] readPointer_CT$wmAdd_Intscfarg_0_1_argbuf_rwb_done;
  assign lizzieLet22_1_d = {readPointer_CT$wmAdd_Intscfarg_0_1_argbuf_rwb_d[115:1],
                            (readPointer_CT$wmAdd_Intscfarg_0_1_argbuf_rwb_d[0] && (! readPointer_CT$wmAdd_Intscfarg_0_1_argbuf_rwb_emitted[0]))};
  assign lizzieLet22_2_d = {readPointer_CT$wmAdd_Intscfarg_0_1_argbuf_rwb_d[115:1],
                            (readPointer_CT$wmAdd_Intscfarg_0_1_argbuf_rwb_d[0] && (! readPointer_CT$wmAdd_Intscfarg_0_1_argbuf_rwb_emitted[1]))};
  assign lizzieLet22_3_d = {readPointer_CT$wmAdd_Intscfarg_0_1_argbuf_rwb_d[115:1],
                            (readPointer_CT$wmAdd_Intscfarg_0_1_argbuf_rwb_d[0] && (! readPointer_CT$wmAdd_Intscfarg_0_1_argbuf_rwb_emitted[2]))};
  assign lizzieLet22_4_d = {readPointer_CT$wmAdd_Intscfarg_0_1_argbuf_rwb_d[115:1],
                            (readPointer_CT$wmAdd_Intscfarg_0_1_argbuf_rwb_d[0] && (! readPointer_CT$wmAdd_Intscfarg_0_1_argbuf_rwb_emitted[3]))};
  assign readPointer_CT$wmAdd_Intscfarg_0_1_argbuf_rwb_done = (readPointer_CT$wmAdd_Intscfarg_0_1_argbuf_rwb_emitted | ({lizzieLet22_4_d[0],
                                                                                                                         lizzieLet22_3_d[0],
                                                                                                                         lizzieLet22_2_d[0],
                                                                                                                         lizzieLet22_1_d[0]} & {lizzieLet22_4_r,
                                                                                                                                                lizzieLet22_3_r,
                                                                                                                                                lizzieLet22_2_r,
                                                                                                                                                lizzieLet22_1_r}));
  assign readPointer_CT$wmAdd_Intscfarg_0_1_argbuf_rwb_r = (& readPointer_CT$wmAdd_Intscfarg_0_1_argbuf_rwb_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_CT$wmAdd_Intscfarg_0_1_argbuf_rwb_emitted <= 4'd0;
    else
      readPointer_CT$wmAdd_Intscfarg_0_1_argbuf_rwb_emitted <= (readPointer_CT$wmAdd_Intscfarg_0_1_argbuf_rwb_r ? 4'd0 :
                                                                readPointer_CT$wmAdd_Intscfarg_0_1_argbuf_rwb_done);
  
  /* buf (Ty CT$wnnz_Int) : (readPointer_CT$wnnz_Intscfarg_0_1_1_argbuf,CT$wnnz_Int) > (readPointer_CT$wnnz_Intscfarg_0_1_1_argbuf_rwb,CT$wnnz_Int) */
  CT$wnnz_Int_t readPointer_CT$wnnz_Intscfarg_0_1_1_argbuf_bufchan_d;
  logic readPointer_CT$wnnz_Intscfarg_0_1_1_argbuf_bufchan_r;
  assign readPointer_CT$wnnz_Intscfarg_0_1_1_argbuf_r = ((! readPointer_CT$wnnz_Intscfarg_0_1_1_argbuf_bufchan_d[0]) || readPointer_CT$wnnz_Intscfarg_0_1_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_CT$wnnz_Intscfarg_0_1_1_argbuf_bufchan_d <= {115'd0,
                                                               1'd0};
    else
      if (readPointer_CT$wnnz_Intscfarg_0_1_1_argbuf_r)
        readPointer_CT$wnnz_Intscfarg_0_1_1_argbuf_bufchan_d <= readPointer_CT$wnnz_Intscfarg_0_1_1_argbuf_d;
  CT$wnnz_Int_t readPointer_CT$wnnz_Intscfarg_0_1_1_argbuf_bufchan_buf;
  assign readPointer_CT$wnnz_Intscfarg_0_1_1_argbuf_bufchan_r = (! readPointer_CT$wnnz_Intscfarg_0_1_1_argbuf_bufchan_buf[0]);
  assign readPointer_CT$wnnz_Intscfarg_0_1_1_argbuf_rwb_d = (readPointer_CT$wnnz_Intscfarg_0_1_1_argbuf_bufchan_buf[0] ? readPointer_CT$wnnz_Intscfarg_0_1_1_argbuf_bufchan_buf :
                                                             readPointer_CT$wnnz_Intscfarg_0_1_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_CT$wnnz_Intscfarg_0_1_1_argbuf_bufchan_buf <= {115'd0,
                                                                 1'd0};
    else
      if ((readPointer_CT$wnnz_Intscfarg_0_1_1_argbuf_rwb_r && readPointer_CT$wnnz_Intscfarg_0_1_1_argbuf_bufchan_buf[0]))
        readPointer_CT$wnnz_Intscfarg_0_1_1_argbuf_bufchan_buf <= {115'd0,
                                                                   1'd0};
      else if (((! readPointer_CT$wnnz_Intscfarg_0_1_1_argbuf_rwb_r) && (! readPointer_CT$wnnz_Intscfarg_0_1_1_argbuf_bufchan_buf[0])))
        readPointer_CT$wnnz_Intscfarg_0_1_1_argbuf_bufchan_buf <= readPointer_CT$wnnz_Intscfarg_0_1_1_argbuf_bufchan_d;
  
  /* fork (Ty CT$wnnz_Int) : (readPointer_CT$wnnz_Intscfarg_0_1_1_argbuf_rwb,CT$wnnz_Int) > [(lizzieLet27_1,CT$wnnz_Int),
                                                                                        (lizzieLet27_2,CT$wnnz_Int),
                                                                                        (lizzieLet27_3,CT$wnnz_Int),
                                                                                        (lizzieLet27_4,CT$wnnz_Int)] */
  logic [3:0] readPointer_CT$wnnz_Intscfarg_0_1_1_argbuf_rwb_emitted;
  logic [3:0] readPointer_CT$wnnz_Intscfarg_0_1_1_argbuf_rwb_done;
  assign lizzieLet27_1_d = {readPointer_CT$wnnz_Intscfarg_0_1_1_argbuf_rwb_d[115:1],
                            (readPointer_CT$wnnz_Intscfarg_0_1_1_argbuf_rwb_d[0] && (! readPointer_CT$wnnz_Intscfarg_0_1_1_argbuf_rwb_emitted[0]))};
  assign lizzieLet27_2_d = {readPointer_CT$wnnz_Intscfarg_0_1_1_argbuf_rwb_d[115:1],
                            (readPointer_CT$wnnz_Intscfarg_0_1_1_argbuf_rwb_d[0] && (! readPointer_CT$wnnz_Intscfarg_0_1_1_argbuf_rwb_emitted[1]))};
  assign lizzieLet27_3_d = {readPointer_CT$wnnz_Intscfarg_0_1_1_argbuf_rwb_d[115:1],
                            (readPointer_CT$wnnz_Intscfarg_0_1_1_argbuf_rwb_d[0] && (! readPointer_CT$wnnz_Intscfarg_0_1_1_argbuf_rwb_emitted[2]))};
  assign lizzieLet27_4_d = {readPointer_CT$wnnz_Intscfarg_0_1_1_argbuf_rwb_d[115:1],
                            (readPointer_CT$wnnz_Intscfarg_0_1_1_argbuf_rwb_d[0] && (! readPointer_CT$wnnz_Intscfarg_0_1_1_argbuf_rwb_emitted[3]))};
  assign readPointer_CT$wnnz_Intscfarg_0_1_1_argbuf_rwb_done = (readPointer_CT$wnnz_Intscfarg_0_1_1_argbuf_rwb_emitted | ({lizzieLet27_4_d[0],
                                                                                                                           lizzieLet27_3_d[0],
                                                                                                                           lizzieLet27_2_d[0],
                                                                                                                           lizzieLet27_1_d[0]} & {lizzieLet27_4_r,
                                                                                                                                                  lizzieLet27_3_r,
                                                                                                                                                  lizzieLet27_2_r,
                                                                                                                                                  lizzieLet27_1_r}));
  assign readPointer_CT$wnnz_Intscfarg_0_1_1_argbuf_rwb_r = (& readPointer_CT$wnnz_Intscfarg_0_1_1_argbuf_rwb_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_CT$wnnz_Intscfarg_0_1_1_argbuf_rwb_emitted <= 4'd0;
    else
      readPointer_CT$wnnz_Intscfarg_0_1_1_argbuf_rwb_emitted <= (readPointer_CT$wnnz_Intscfarg_0_1_1_argbuf_rwb_r ? 4'd0 :
                                                                 readPointer_CT$wnnz_Intscfarg_0_1_1_argbuf_rwb_done);
  
  /* buf (Ty CTmain_mask_Int) : (readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf,CTmain_mask_Int) > (readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf_rwb,CTmain_mask_Int) */
  CTmain_mask_Int_t readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf_bufchan_d;
  logic readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf_bufchan_r;
  assign readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf_r = ((! readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf_bufchan_d[0]) || readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf_bufchan_d <= {115'd0,
                                                                   1'd0};
    else
      if (readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf_r)
        readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf_bufchan_d <= readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf_d;
  CTmain_mask_Int_t readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf_bufchan_buf;
  assign readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf_bufchan_r = (! readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf_bufchan_buf[0]);
  assign readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf_rwb_d = (readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf_bufchan_buf[0] ? readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf_bufchan_buf :
                                                                 readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf_bufchan_buf <= {115'd0,
                                                                     1'd0};
    else
      if ((readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf_rwb_r && readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf_bufchan_buf[0]))
        readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf_bufchan_buf <= {115'd0,
                                                                       1'd0};
      else if (((! readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf_rwb_r) && (! readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf_bufchan_buf[0])))
        readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf_bufchan_buf <= readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf_bufchan_d;
  
  /* fork (Ty CTmain_mask_Int) : (readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf_rwb,CTmain_mask_Int) > [(lizzieLet31_1,CTmain_mask_Int),
                                                                                                    (lizzieLet31_2,CTmain_mask_Int),
                                                                                                    (lizzieLet31_3,CTmain_mask_Int),
                                                                                                    (lizzieLet31_4,CTmain_mask_Int)] */
  logic [3:0] readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf_rwb_emitted;
  logic [3:0] readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf_rwb_done;
  assign lizzieLet31_1_d = {readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf_rwb_d[115:1],
                            (readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf_rwb_d[0] && (! readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf_rwb_emitted[0]))};
  assign lizzieLet31_2_d = {readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf_rwb_d[115:1],
                            (readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf_rwb_d[0] && (! readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf_rwb_emitted[1]))};
  assign lizzieLet31_3_d = {readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf_rwb_d[115:1],
                            (readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf_rwb_d[0] && (! readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf_rwb_emitted[2]))};
  assign lizzieLet31_4_d = {readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf_rwb_d[115:1],
                            (readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf_rwb_d[0] && (! readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf_rwb_emitted[3]))};
  assign readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf_rwb_done = (readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf_rwb_emitted | ({lizzieLet31_4_d[0],
                                                                                                                                   lizzieLet31_3_d[0],
                                                                                                                                   lizzieLet31_2_d[0],
                                                                                                                                   lizzieLet31_1_d[0]} & {lizzieLet31_4_r,
                                                                                                                                                          lizzieLet31_3_r,
                                                                                                                                                          lizzieLet31_2_r,
                                                                                                                                                          lizzieLet31_1_r}));
  assign readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf_rwb_r = (& readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf_rwb_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf_rwb_emitted <= 4'd0;
    else
      readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf_rwb_emitted <= (readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf_rwb_r ? 4'd0 :
                                                                     readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf_rwb_done);
  
  /* buf (Ty MaskQTree) : (readPointer_MaskQTreemska8r_1_argbuf,MaskQTree) > (readPointer_MaskQTreemska8r_1_argbuf_rwb,MaskQTree) */
  MaskQTree_t readPointer_MaskQTreemska8r_1_argbuf_bufchan_d;
  logic readPointer_MaskQTreemska8r_1_argbuf_bufchan_r;
  assign readPointer_MaskQTreemska8r_1_argbuf_r = ((! readPointer_MaskQTreemska8r_1_argbuf_bufchan_d[0]) || readPointer_MaskQTreemska8r_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_MaskQTreemska8r_1_argbuf_bufchan_d <= {66'd0, 1'd0};
    else
      if (readPointer_MaskQTreemska8r_1_argbuf_r)
        readPointer_MaskQTreemska8r_1_argbuf_bufchan_d <= readPointer_MaskQTreemska8r_1_argbuf_d;
  MaskQTree_t readPointer_MaskQTreemska8r_1_argbuf_bufchan_buf;
  assign readPointer_MaskQTreemska8r_1_argbuf_bufchan_r = (! readPointer_MaskQTreemska8r_1_argbuf_bufchan_buf[0]);
  assign readPointer_MaskQTreemska8r_1_argbuf_rwb_d = (readPointer_MaskQTreemska8r_1_argbuf_bufchan_buf[0] ? readPointer_MaskQTreemska8r_1_argbuf_bufchan_buf :
                                                       readPointer_MaskQTreemska8r_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_MaskQTreemska8r_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((readPointer_MaskQTreemska8r_1_argbuf_rwb_r && readPointer_MaskQTreemska8r_1_argbuf_bufchan_buf[0]))
        readPointer_MaskQTreemska8r_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
      else if (((! readPointer_MaskQTreemska8r_1_argbuf_rwb_r) && (! readPointer_MaskQTreemska8r_1_argbuf_bufchan_buf[0])))
        readPointer_MaskQTreemska8r_1_argbuf_bufchan_buf <= readPointer_MaskQTreemska8r_1_argbuf_bufchan_d;
  
  /* fork (Ty MaskQTree) : (readPointer_MaskQTreemska8r_1_argbuf_rwb,MaskQTree) > [(lizzieLet14_1_1,MaskQTree),
                                                                              (lizzieLet14_1_2,MaskQTree),
                                                                              (lizzieLet14_1_3,MaskQTree),
                                                                              (lizzieLet14_1_4,MaskQTree),
                                                                              (lizzieLet14_1_5,MaskQTree),
                                                                              (lizzieLet14_1_6,MaskQTree)] */
  logic [5:0] readPointer_MaskQTreemska8r_1_argbuf_rwb_emitted;
  logic [5:0] readPointer_MaskQTreemska8r_1_argbuf_rwb_done;
  assign lizzieLet14_1_1_d = {readPointer_MaskQTreemska8r_1_argbuf_rwb_d[66:1],
                              (readPointer_MaskQTreemska8r_1_argbuf_rwb_d[0] && (! readPointer_MaskQTreemska8r_1_argbuf_rwb_emitted[0]))};
  assign lizzieLet14_1_2_d = {readPointer_MaskQTreemska8r_1_argbuf_rwb_d[66:1],
                              (readPointer_MaskQTreemska8r_1_argbuf_rwb_d[0] && (! readPointer_MaskQTreemska8r_1_argbuf_rwb_emitted[1]))};
  assign lizzieLet14_1_3_d = {readPointer_MaskQTreemska8r_1_argbuf_rwb_d[66:1],
                              (readPointer_MaskQTreemska8r_1_argbuf_rwb_d[0] && (! readPointer_MaskQTreemska8r_1_argbuf_rwb_emitted[2]))};
  assign lizzieLet14_1_4_d = {readPointer_MaskQTreemska8r_1_argbuf_rwb_d[66:1],
                              (readPointer_MaskQTreemska8r_1_argbuf_rwb_d[0] && (! readPointer_MaskQTreemska8r_1_argbuf_rwb_emitted[3]))};
  assign lizzieLet14_1_5_d = {readPointer_MaskQTreemska8r_1_argbuf_rwb_d[66:1],
                              (readPointer_MaskQTreemska8r_1_argbuf_rwb_d[0] && (! readPointer_MaskQTreemska8r_1_argbuf_rwb_emitted[4]))};
  assign lizzieLet14_1_6_d = {readPointer_MaskQTreemska8r_1_argbuf_rwb_d[66:1],
                              (readPointer_MaskQTreemska8r_1_argbuf_rwb_d[0] && (! readPointer_MaskQTreemska8r_1_argbuf_rwb_emitted[5]))};
  assign readPointer_MaskQTreemska8r_1_argbuf_rwb_done = (readPointer_MaskQTreemska8r_1_argbuf_rwb_emitted | ({lizzieLet14_1_6_d[0],
                                                                                                               lizzieLet14_1_5_d[0],
                                                                                                               lizzieLet14_1_4_d[0],
                                                                                                               lizzieLet14_1_3_d[0],
                                                                                                               lizzieLet14_1_2_d[0],
                                                                                                               lizzieLet14_1_1_d[0]} & {lizzieLet14_1_6_r,
                                                                                                                                        lizzieLet14_1_5_r,
                                                                                                                                        lizzieLet14_1_4_r,
                                                                                                                                        lizzieLet14_1_3_r,
                                                                                                                                        lizzieLet14_1_2_r,
                                                                                                                                        lizzieLet14_1_1_r}));
  assign readPointer_MaskQTreemska8r_1_argbuf_rwb_r = (& readPointer_MaskQTreemska8r_1_argbuf_rwb_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_MaskQTreemska8r_1_argbuf_rwb_emitted <= 6'd0;
    else
      readPointer_MaskQTreemska8r_1_argbuf_rwb_emitted <= (readPointer_MaskQTreemska8r_1_argbuf_rwb_r ? 6'd0 :
                                                           readPointer_MaskQTreemska8r_1_argbuf_rwb_done);
  
  /* buf (Ty QTree_Int) : (readPointer_QTree_Intma8q_1_argbuf,QTree_Int) > (readPointer_QTree_Intma8q_1_argbuf_rwb,QTree_Int) */
  QTree_Int_t readPointer_QTree_Intma8q_1_argbuf_bufchan_d;
  logic readPointer_QTree_Intma8q_1_argbuf_bufchan_r;
  assign readPointer_QTree_Intma8q_1_argbuf_r = ((! readPointer_QTree_Intma8q_1_argbuf_bufchan_d[0]) || readPointer_QTree_Intma8q_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Intma8q_1_argbuf_bufchan_d <= {66'd0, 1'd0};
    else
      if (readPointer_QTree_Intma8q_1_argbuf_r)
        readPointer_QTree_Intma8q_1_argbuf_bufchan_d <= readPointer_QTree_Intma8q_1_argbuf_d;
  QTree_Int_t readPointer_QTree_Intma8q_1_argbuf_bufchan_buf;
  assign readPointer_QTree_Intma8q_1_argbuf_bufchan_r = (! readPointer_QTree_Intma8q_1_argbuf_bufchan_buf[0]);
  assign readPointer_QTree_Intma8q_1_argbuf_rwb_d = (readPointer_QTree_Intma8q_1_argbuf_bufchan_buf[0] ? readPointer_QTree_Intma8q_1_argbuf_bufchan_buf :
                                                     readPointer_QTree_Intma8q_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Intma8q_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((readPointer_QTree_Intma8q_1_argbuf_rwb_r && readPointer_QTree_Intma8q_1_argbuf_bufchan_buf[0]))
        readPointer_QTree_Intma8q_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
      else if (((! readPointer_QTree_Intma8q_1_argbuf_rwb_r) && (! readPointer_QTree_Intma8q_1_argbuf_bufchan_buf[0])))
        readPointer_QTree_Intma8q_1_argbuf_bufchan_buf <= readPointer_QTree_Intma8q_1_argbuf_bufchan_d;
  
  /* buf (Ty QTree_Int) : (readPointer_QTree_Intw1sif_1_1_argbuf,QTree_Int) > (readPointer_QTree_Intw1sif_1_1_argbuf_rwb,QTree_Int) */
  QTree_Int_t readPointer_QTree_Intw1sif_1_1_argbuf_bufchan_d;
  logic readPointer_QTree_Intw1sif_1_1_argbuf_bufchan_r;
  assign readPointer_QTree_Intw1sif_1_1_argbuf_r = ((! readPointer_QTree_Intw1sif_1_1_argbuf_bufchan_d[0]) || readPointer_QTree_Intw1sif_1_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Intw1sif_1_1_argbuf_bufchan_d <= {66'd0, 1'd0};
    else
      if (readPointer_QTree_Intw1sif_1_1_argbuf_r)
        readPointer_QTree_Intw1sif_1_1_argbuf_bufchan_d <= readPointer_QTree_Intw1sif_1_1_argbuf_d;
  QTree_Int_t readPointer_QTree_Intw1sif_1_1_argbuf_bufchan_buf;
  assign readPointer_QTree_Intw1sif_1_1_argbuf_bufchan_r = (! readPointer_QTree_Intw1sif_1_1_argbuf_bufchan_buf[0]);
  assign readPointer_QTree_Intw1sif_1_1_argbuf_rwb_d = (readPointer_QTree_Intw1sif_1_1_argbuf_bufchan_buf[0] ? readPointer_QTree_Intw1sif_1_1_argbuf_bufchan_buf :
                                                        readPointer_QTree_Intw1sif_1_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Intw1sif_1_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((readPointer_QTree_Intw1sif_1_1_argbuf_rwb_r && readPointer_QTree_Intw1sif_1_1_argbuf_bufchan_buf[0]))
        readPointer_QTree_Intw1sif_1_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
      else if (((! readPointer_QTree_Intw1sif_1_1_argbuf_rwb_r) && (! readPointer_QTree_Intw1sif_1_1_argbuf_bufchan_buf[0])))
        readPointer_QTree_Intw1sif_1_1_argbuf_bufchan_buf <= readPointer_QTree_Intw1sif_1_1_argbuf_bufchan_d;
  
  /* fork (Ty QTree_Int) : (readPointer_QTree_Intw1sif_1_1_argbuf_rwb,QTree_Int) > [(lizzieLet2_1,QTree_Int),
                                                                               (lizzieLet2_2,QTree_Int),
                                                                               (lizzieLet2_3,QTree_Int),
                                                                               (lizzieLet2_4,QTree_Int),
                                                                               (lizzieLet2_5,QTree_Int),
                                                                               (lizzieLet2_6,QTree_Int),
                                                                               (lizzieLet2_7,QTree_Int),
                                                                               (lizzieLet2_8,QTree_Int)] */
  logic [7:0] readPointer_QTree_Intw1sif_1_1_argbuf_rwb_emitted;
  logic [7:0] readPointer_QTree_Intw1sif_1_1_argbuf_rwb_done;
  assign lizzieLet2_1_d = {readPointer_QTree_Intw1sif_1_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_Intw1sif_1_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intw1sif_1_1_argbuf_rwb_emitted[0]))};
  assign lizzieLet2_2_d = {readPointer_QTree_Intw1sif_1_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_Intw1sif_1_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intw1sif_1_1_argbuf_rwb_emitted[1]))};
  assign lizzieLet2_3_d = {readPointer_QTree_Intw1sif_1_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_Intw1sif_1_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intw1sif_1_1_argbuf_rwb_emitted[2]))};
  assign lizzieLet2_4_d = {readPointer_QTree_Intw1sif_1_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_Intw1sif_1_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intw1sif_1_1_argbuf_rwb_emitted[3]))};
  assign lizzieLet2_5_d = {readPointer_QTree_Intw1sif_1_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_Intw1sif_1_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intw1sif_1_1_argbuf_rwb_emitted[4]))};
  assign lizzieLet2_6_d = {readPointer_QTree_Intw1sif_1_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_Intw1sif_1_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intw1sif_1_1_argbuf_rwb_emitted[5]))};
  assign lizzieLet2_7_d = {readPointer_QTree_Intw1sif_1_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_Intw1sif_1_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intw1sif_1_1_argbuf_rwb_emitted[6]))};
  assign lizzieLet2_8_d = {readPointer_QTree_Intw1sif_1_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_Intw1sif_1_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intw1sif_1_1_argbuf_rwb_emitted[7]))};
  assign readPointer_QTree_Intw1sif_1_1_argbuf_rwb_done = (readPointer_QTree_Intw1sif_1_1_argbuf_rwb_emitted | ({lizzieLet2_8_d[0],
                                                                                                                 lizzieLet2_7_d[0],
                                                                                                                 lizzieLet2_6_d[0],
                                                                                                                 lizzieLet2_5_d[0],
                                                                                                                 lizzieLet2_4_d[0],
                                                                                                                 lizzieLet2_3_d[0],
                                                                                                                 lizzieLet2_2_d[0],
                                                                                                                 lizzieLet2_1_d[0]} & {lizzieLet2_8_r,
                                                                                                                                       lizzieLet2_7_r,
                                                                                                                                       lizzieLet2_6_r,
                                                                                                                                       lizzieLet2_5_r,
                                                                                                                                       lizzieLet2_4_r,
                                                                                                                                       lizzieLet2_3_r,
                                                                                                                                       lizzieLet2_2_r,
                                                                                                                                       lizzieLet2_1_r}));
  assign readPointer_QTree_Intw1sif_1_1_argbuf_rwb_r = (& readPointer_QTree_Intw1sif_1_1_argbuf_rwb_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Intw1sif_1_1_argbuf_rwb_emitted <= 8'd0;
    else
      readPointer_QTree_Intw1sif_1_1_argbuf_rwb_emitted <= (readPointer_QTree_Intw1sif_1_1_argbuf_rwb_r ? 8'd0 :
                                                            readPointer_QTree_Intw1sif_1_1_argbuf_rwb_done);
  
  /* buf (Ty QTree_Int) : (readPointer_QTree_Intw2sig_1_1_argbuf,QTree_Int) > (readPointer_QTree_Intw2sig_1_1_argbuf_rwb,QTree_Int) */
  QTree_Int_t readPointer_QTree_Intw2sig_1_1_argbuf_bufchan_d;
  logic readPointer_QTree_Intw2sig_1_1_argbuf_bufchan_r;
  assign readPointer_QTree_Intw2sig_1_1_argbuf_r = ((! readPointer_QTree_Intw2sig_1_1_argbuf_bufchan_d[0]) || readPointer_QTree_Intw2sig_1_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Intw2sig_1_1_argbuf_bufchan_d <= {66'd0, 1'd0};
    else
      if (readPointer_QTree_Intw2sig_1_1_argbuf_r)
        readPointer_QTree_Intw2sig_1_1_argbuf_bufchan_d <= readPointer_QTree_Intw2sig_1_1_argbuf_d;
  QTree_Int_t readPointer_QTree_Intw2sig_1_1_argbuf_bufchan_buf;
  assign readPointer_QTree_Intw2sig_1_1_argbuf_bufchan_r = (! readPointer_QTree_Intw2sig_1_1_argbuf_bufchan_buf[0]);
  assign readPointer_QTree_Intw2sig_1_1_argbuf_rwb_d = (readPointer_QTree_Intw2sig_1_1_argbuf_bufchan_buf[0] ? readPointer_QTree_Intw2sig_1_1_argbuf_bufchan_buf :
                                                        readPointer_QTree_Intw2sig_1_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Intw2sig_1_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((readPointer_QTree_Intw2sig_1_1_argbuf_rwb_r && readPointer_QTree_Intw2sig_1_1_argbuf_bufchan_buf[0]))
        readPointer_QTree_Intw2sig_1_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
      else if (((! readPointer_QTree_Intw2sig_1_1_argbuf_rwb_r) && (! readPointer_QTree_Intw2sig_1_1_argbuf_bufchan_buf[0])))
        readPointer_QTree_Intw2sig_1_1_argbuf_bufchan_buf <= readPointer_QTree_Intw2sig_1_1_argbuf_bufchan_d;
  
  /* buf (Ty QTree_Int) : (readPointer_QTree_Intwsij_1_1_argbuf,QTree_Int) > (readPointer_QTree_Intwsij_1_1_argbuf_rwb,QTree_Int) */
  QTree_Int_t readPointer_QTree_Intwsij_1_1_argbuf_bufchan_d;
  logic readPointer_QTree_Intwsij_1_1_argbuf_bufchan_r;
  assign readPointer_QTree_Intwsij_1_1_argbuf_r = ((! readPointer_QTree_Intwsij_1_1_argbuf_bufchan_d[0]) || readPointer_QTree_Intwsij_1_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Intwsij_1_1_argbuf_bufchan_d <= {66'd0, 1'd0};
    else
      if (readPointer_QTree_Intwsij_1_1_argbuf_r)
        readPointer_QTree_Intwsij_1_1_argbuf_bufchan_d <= readPointer_QTree_Intwsij_1_1_argbuf_d;
  QTree_Int_t readPointer_QTree_Intwsij_1_1_argbuf_bufchan_buf;
  assign readPointer_QTree_Intwsij_1_1_argbuf_bufchan_r = (! readPointer_QTree_Intwsij_1_1_argbuf_bufchan_buf[0]);
  assign readPointer_QTree_Intwsij_1_1_argbuf_rwb_d = (readPointer_QTree_Intwsij_1_1_argbuf_bufchan_buf[0] ? readPointer_QTree_Intwsij_1_1_argbuf_bufchan_buf :
                                                       readPointer_QTree_Intwsij_1_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Intwsij_1_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((readPointer_QTree_Intwsij_1_1_argbuf_rwb_r && readPointer_QTree_Intwsij_1_1_argbuf_bufchan_buf[0]))
        readPointer_QTree_Intwsij_1_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
      else if (((! readPointer_QTree_Intwsij_1_1_argbuf_rwb_r) && (! readPointer_QTree_Intwsij_1_1_argbuf_bufchan_buf[0])))
        readPointer_QTree_Intwsij_1_1_argbuf_bufchan_buf <= readPointer_QTree_Intwsij_1_1_argbuf_bufchan_d;
  
  /* fork (Ty QTree_Int) : (readPointer_QTree_Intwsij_1_1_argbuf_rwb,QTree_Int) > [(lizzieLet12_1_1,QTree_Int),
                                                                              (lizzieLet12_1_2,QTree_Int),
                                                                              (lizzieLet12_1_3,QTree_Int),
                                                                              (lizzieLet12_1_4,QTree_Int)] */
  logic [3:0] readPointer_QTree_Intwsij_1_1_argbuf_rwb_emitted;
  logic [3:0] readPointer_QTree_Intwsij_1_1_argbuf_rwb_done;
  assign lizzieLet12_1_1_d = {readPointer_QTree_Intwsij_1_1_argbuf_rwb_d[66:1],
                              (readPointer_QTree_Intwsij_1_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intwsij_1_1_argbuf_rwb_emitted[0]))};
  assign lizzieLet12_1_2_d = {readPointer_QTree_Intwsij_1_1_argbuf_rwb_d[66:1],
                              (readPointer_QTree_Intwsij_1_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intwsij_1_1_argbuf_rwb_emitted[1]))};
  assign lizzieLet12_1_3_d = {readPointer_QTree_Intwsij_1_1_argbuf_rwb_d[66:1],
                              (readPointer_QTree_Intwsij_1_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intwsij_1_1_argbuf_rwb_emitted[2]))};
  assign lizzieLet12_1_4_d = {readPointer_QTree_Intwsij_1_1_argbuf_rwb_d[66:1],
                              (readPointer_QTree_Intwsij_1_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intwsij_1_1_argbuf_rwb_emitted[3]))};
  assign readPointer_QTree_Intwsij_1_1_argbuf_rwb_done = (readPointer_QTree_Intwsij_1_1_argbuf_rwb_emitted | ({lizzieLet12_1_4_d[0],
                                                                                                               lizzieLet12_1_3_d[0],
                                                                                                               lizzieLet12_1_2_d[0],
                                                                                                               lizzieLet12_1_1_d[0]} & {lizzieLet12_1_4_r,
                                                                                                                                        lizzieLet12_1_3_r,
                                                                                                                                        lizzieLet12_1_2_r,
                                                                                                                                        lizzieLet12_1_1_r}));
  assign readPointer_QTree_Intwsij_1_1_argbuf_rwb_r = (& readPointer_QTree_Intwsij_1_1_argbuf_rwb_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Intwsij_1_1_argbuf_rwb_emitted <= 4'd0;
    else
      readPointer_QTree_Intwsij_1_1_argbuf_rwb_emitted <= (readPointer_QTree_Intwsij_1_1_argbuf_rwb_r ? 4'd0 :
                                                           readPointer_QTree_Intwsij_1_1_argbuf_rwb_done);
  
  /* buf (Ty Pointer_CT$wnnz_Int) : (sc_0_10_destruct,Pointer_CT$wnnz_Int) > (sc_0_10_1_argbuf,Pointer_CT$wnnz_Int) */
  Pointer_CT$wnnz_Int_t sc_0_10_destruct_bufchan_d;
  logic sc_0_10_destruct_bufchan_r;
  assign sc_0_10_destruct_r = ((! sc_0_10_destruct_bufchan_d[0]) || sc_0_10_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) sc_0_10_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (sc_0_10_destruct_r)
        sc_0_10_destruct_bufchan_d <= sc_0_10_destruct_d;
  Pointer_CT$wnnz_Int_t sc_0_10_destruct_bufchan_buf;
  assign sc_0_10_destruct_bufchan_r = (! sc_0_10_destruct_bufchan_buf[0]);
  assign sc_0_10_1_argbuf_d = (sc_0_10_destruct_bufchan_buf[0] ? sc_0_10_destruct_bufchan_buf :
                               sc_0_10_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) sc_0_10_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((sc_0_10_1_argbuf_r && sc_0_10_destruct_bufchan_buf[0]))
        sc_0_10_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! sc_0_10_1_argbuf_r) && (! sc_0_10_destruct_bufchan_buf[0])))
        sc_0_10_destruct_bufchan_buf <= sc_0_10_destruct_bufchan_d;
  
  /* buf (Ty Pointer_CTmain_mask_Int) : (sc_0_14_destruct,Pointer_CTmain_mask_Int) > (sc_0_14_1_argbuf,Pointer_CTmain_mask_Int) */
  Pointer_CTmain_mask_Int_t sc_0_14_destruct_bufchan_d;
  logic sc_0_14_destruct_bufchan_r;
  assign sc_0_14_destruct_r = ((! sc_0_14_destruct_bufchan_d[0]) || sc_0_14_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) sc_0_14_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (sc_0_14_destruct_r)
        sc_0_14_destruct_bufchan_d <= sc_0_14_destruct_d;
  Pointer_CTmain_mask_Int_t sc_0_14_destruct_bufchan_buf;
  assign sc_0_14_destruct_bufchan_r = (! sc_0_14_destruct_bufchan_buf[0]);
  assign sc_0_14_1_argbuf_d = (sc_0_14_destruct_bufchan_buf[0] ? sc_0_14_destruct_bufchan_buf :
                               sc_0_14_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) sc_0_14_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((sc_0_14_1_argbuf_r && sc_0_14_destruct_bufchan_buf[0]))
        sc_0_14_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! sc_0_14_1_argbuf_r) && (! sc_0_14_destruct_bufchan_buf[0])))
        sc_0_14_destruct_bufchan_buf <= sc_0_14_destruct_bufchan_d;
  
  /* buf (Ty Pointer_CT$wmAdd_Int) : (sc_0_6_destruct,Pointer_CT$wmAdd_Int) > (sc_0_6_1_argbuf,Pointer_CT$wmAdd_Int) */
  Pointer_CT$wmAdd_Int_t sc_0_6_destruct_bufchan_d;
  logic sc_0_6_destruct_bufchan_r;
  assign sc_0_6_destruct_r = ((! sc_0_6_destruct_bufchan_d[0]) || sc_0_6_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) sc_0_6_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (sc_0_6_destruct_r)
        sc_0_6_destruct_bufchan_d <= sc_0_6_destruct_d;
  Pointer_CT$wmAdd_Int_t sc_0_6_destruct_bufchan_buf;
  assign sc_0_6_destruct_bufchan_r = (! sc_0_6_destruct_bufchan_buf[0]);
  assign sc_0_6_1_argbuf_d = (sc_0_6_destruct_bufchan_buf[0] ? sc_0_6_destruct_bufchan_buf :
                              sc_0_6_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) sc_0_6_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((sc_0_6_1_argbuf_r && sc_0_6_destruct_bufchan_buf[0]))
        sc_0_6_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! sc_0_6_1_argbuf_r) && (! sc_0_6_destruct_bufchan_buf[0])))
        sc_0_6_destruct_bufchan_buf <= sc_0_6_destruct_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz_Int) : (scfarg_0_1_goMux_mux,Pointer_CT$wnnz_Int) > (scfarg_0_1_1_argbuf,Pointer_CT$wnnz_Int) */
  Pointer_CT$wnnz_Int_t scfarg_0_1_goMux_mux_bufchan_d;
  logic scfarg_0_1_goMux_mux_bufchan_r;
  assign scfarg_0_1_goMux_mux_r = ((! scfarg_0_1_goMux_mux_bufchan_d[0]) || scfarg_0_1_goMux_mux_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      scfarg_0_1_goMux_mux_bufchan_d <= {16'd0, 1'd0};
    else
      if (scfarg_0_1_goMux_mux_r)
        scfarg_0_1_goMux_mux_bufchan_d <= scfarg_0_1_goMux_mux_d;
  Pointer_CT$wnnz_Int_t scfarg_0_1_goMux_mux_bufchan_buf;
  assign scfarg_0_1_goMux_mux_bufchan_r = (! scfarg_0_1_goMux_mux_bufchan_buf[0]);
  assign scfarg_0_1_1_argbuf_d = (scfarg_0_1_goMux_mux_bufchan_buf[0] ? scfarg_0_1_goMux_mux_bufchan_buf :
                                  scfarg_0_1_goMux_mux_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      scfarg_0_1_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((scfarg_0_1_1_argbuf_r && scfarg_0_1_goMux_mux_bufchan_buf[0]))
        scfarg_0_1_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
      else if (((! scfarg_0_1_1_argbuf_r) && (! scfarg_0_1_goMux_mux_bufchan_buf[0])))
        scfarg_0_1_goMux_mux_bufchan_buf <= scfarg_0_1_goMux_mux_bufchan_d;
  
  /* buf (Ty Pointer_CTmain_mask_Int) : (scfarg_0_2_goMux_mux,Pointer_CTmain_mask_Int) > (scfarg_0_2_1_argbuf,Pointer_CTmain_mask_Int) */
  Pointer_CTmain_mask_Int_t scfarg_0_2_goMux_mux_bufchan_d;
  logic scfarg_0_2_goMux_mux_bufchan_r;
  assign scfarg_0_2_goMux_mux_r = ((! scfarg_0_2_goMux_mux_bufchan_d[0]) || scfarg_0_2_goMux_mux_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      scfarg_0_2_goMux_mux_bufchan_d <= {16'd0, 1'd0};
    else
      if (scfarg_0_2_goMux_mux_r)
        scfarg_0_2_goMux_mux_bufchan_d <= scfarg_0_2_goMux_mux_d;
  Pointer_CTmain_mask_Int_t scfarg_0_2_goMux_mux_bufchan_buf;
  assign scfarg_0_2_goMux_mux_bufchan_r = (! scfarg_0_2_goMux_mux_bufchan_buf[0]);
  assign scfarg_0_2_1_argbuf_d = (scfarg_0_2_goMux_mux_bufchan_buf[0] ? scfarg_0_2_goMux_mux_bufchan_buf :
                                  scfarg_0_2_goMux_mux_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      scfarg_0_2_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((scfarg_0_2_1_argbuf_r && scfarg_0_2_goMux_mux_bufchan_buf[0]))
        scfarg_0_2_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
      else if (((! scfarg_0_2_1_argbuf_r) && (! scfarg_0_2_goMux_mux_bufchan_buf[0])))
        scfarg_0_2_goMux_mux_bufchan_buf <= scfarg_0_2_goMux_mux_bufchan_d;
  
  /* buf (Ty Pointer_CT$wmAdd_Int) : (scfarg_0_goMux_mux,Pointer_CT$wmAdd_Int) > (scfarg_0_1_argbuf,Pointer_CT$wmAdd_Int) */
  Pointer_CT$wmAdd_Int_t scfarg_0_goMux_mux_bufchan_d;
  logic scfarg_0_goMux_mux_bufchan_r;
  assign scfarg_0_goMux_mux_r = ((! scfarg_0_goMux_mux_bufchan_d[0]) || scfarg_0_goMux_mux_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) scfarg_0_goMux_mux_bufchan_d <= {16'd0, 1'd0};
    else
      if (scfarg_0_goMux_mux_r)
        scfarg_0_goMux_mux_bufchan_d <= scfarg_0_goMux_mux_d;
  Pointer_CT$wmAdd_Int_t scfarg_0_goMux_mux_bufchan_buf;
  assign scfarg_0_goMux_mux_bufchan_r = (! scfarg_0_goMux_mux_bufchan_buf[0]);
  assign scfarg_0_1_argbuf_d = (scfarg_0_goMux_mux_bufchan_buf[0] ? scfarg_0_goMux_mux_bufchan_buf :
                                scfarg_0_goMux_mux_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      scfarg_0_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((scfarg_0_1_argbuf_r && scfarg_0_goMux_mux_bufchan_buf[0]))
        scfarg_0_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
      else if (((! scfarg_0_1_argbuf_r) && (! scfarg_0_goMux_mux_bufchan_buf[0])))
        scfarg_0_goMux_mux_bufchan_buf <= scfarg_0_goMux_mux_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (t1a8m_3_destruct,Pointer_QTree_Int) > (t1a8m_3_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t t1a8m_3_destruct_bufchan_d;
  logic t1a8m_3_destruct_bufchan_r;
  assign t1a8m_3_destruct_r = ((! t1a8m_3_destruct_bufchan_d[0]) || t1a8m_3_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t1a8m_3_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (t1a8m_3_destruct_r)
        t1a8m_3_destruct_bufchan_d <= t1a8m_3_destruct_d;
  Pointer_QTree_Int_t t1a8m_3_destruct_bufchan_buf;
  assign t1a8m_3_destruct_bufchan_r = (! t1a8m_3_destruct_bufchan_buf[0]);
  assign t1a8m_3_1_argbuf_d = (t1a8m_3_destruct_bufchan_buf[0] ? t1a8m_3_destruct_bufchan_buf :
                               t1a8m_3_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t1a8m_3_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((t1a8m_3_1_argbuf_r && t1a8m_3_destruct_bufchan_buf[0]))
        t1a8m_3_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! t1a8m_3_1_argbuf_r) && (! t1a8m_3_destruct_bufchan_buf[0])))
        t1a8m_3_destruct_bufchan_buf <= t1a8m_3_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (t1a8x_3_destruct,Pointer_QTree_Int) > (t1a8x_3_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t t1a8x_3_destruct_bufchan_d;
  logic t1a8x_3_destruct_bufchan_r;
  assign t1a8x_3_destruct_r = ((! t1a8x_3_destruct_bufchan_d[0]) || t1a8x_3_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t1a8x_3_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (t1a8x_3_destruct_r)
        t1a8x_3_destruct_bufchan_d <= t1a8x_3_destruct_d;
  Pointer_QTree_Int_t t1a8x_3_destruct_bufchan_buf;
  assign t1a8x_3_destruct_bufchan_r = (! t1a8x_3_destruct_bufchan_buf[0]);
  assign t1a8x_3_1_argbuf_d = (t1a8x_3_destruct_bufchan_buf[0] ? t1a8x_3_destruct_bufchan_buf :
                               t1a8x_3_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t1a8x_3_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((t1a8x_3_1_argbuf_r && t1a8x_3_destruct_bufchan_buf[0]))
        t1a8x_3_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! t1a8x_3_1_argbuf_r) && (! t1a8x_3_destruct_bufchan_buf[0])))
        t1a8x_3_destruct_bufchan_buf <= t1a8x_3_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (t2a8n_2_destruct,Pointer_QTree_Int) > (t2a8n_2_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t t2a8n_2_destruct_bufchan_d;
  logic t2a8n_2_destruct_bufchan_r;
  assign t2a8n_2_destruct_r = ((! t2a8n_2_destruct_bufchan_d[0]) || t2a8n_2_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t2a8n_2_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (t2a8n_2_destruct_r)
        t2a8n_2_destruct_bufchan_d <= t2a8n_2_destruct_d;
  Pointer_QTree_Int_t t2a8n_2_destruct_bufchan_buf;
  assign t2a8n_2_destruct_bufchan_r = (! t2a8n_2_destruct_bufchan_buf[0]);
  assign t2a8n_2_1_argbuf_d = (t2a8n_2_destruct_bufchan_buf[0] ? t2a8n_2_destruct_bufchan_buf :
                               t2a8n_2_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t2a8n_2_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((t2a8n_2_1_argbuf_r && t2a8n_2_destruct_bufchan_buf[0]))
        t2a8n_2_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! t2a8n_2_1_argbuf_r) && (! t2a8n_2_destruct_bufchan_buf[0])))
        t2a8n_2_destruct_bufchan_buf <= t2a8n_2_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (t2a8y_2_destruct,Pointer_QTree_Int) > (t2a8y_2_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t t2a8y_2_destruct_bufchan_d;
  logic t2a8y_2_destruct_bufchan_r;
  assign t2a8y_2_destruct_r = ((! t2a8y_2_destruct_bufchan_d[0]) || t2a8y_2_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t2a8y_2_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (t2a8y_2_destruct_r)
        t2a8y_2_destruct_bufchan_d <= t2a8y_2_destruct_d;
  Pointer_QTree_Int_t t2a8y_2_destruct_bufchan_buf;
  assign t2a8y_2_destruct_bufchan_r = (! t2a8y_2_destruct_bufchan_buf[0]);
  assign t2a8y_2_1_argbuf_d = (t2a8y_2_destruct_bufchan_buf[0] ? t2a8y_2_destruct_bufchan_buf :
                               t2a8y_2_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t2a8y_2_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((t2a8y_2_1_argbuf_r && t2a8y_2_destruct_bufchan_buf[0]))
        t2a8y_2_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! t2a8y_2_1_argbuf_r) && (! t2a8y_2_destruct_bufchan_buf[0])))
        t2a8y_2_destruct_bufchan_buf <= t2a8y_2_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (t3a8o_1_destruct,Pointer_QTree_Int) > (t3a8o_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t t3a8o_1_destruct_bufchan_d;
  logic t3a8o_1_destruct_bufchan_r;
  assign t3a8o_1_destruct_r = ((! t3a8o_1_destruct_bufchan_d[0]) || t3a8o_1_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t3a8o_1_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (t3a8o_1_destruct_r)
        t3a8o_1_destruct_bufchan_d <= t3a8o_1_destruct_d;
  Pointer_QTree_Int_t t3a8o_1_destruct_bufchan_buf;
  assign t3a8o_1_destruct_bufchan_r = (! t3a8o_1_destruct_bufchan_buf[0]);
  assign t3a8o_1_1_argbuf_d = (t3a8o_1_destruct_bufchan_buf[0] ? t3a8o_1_destruct_bufchan_buf :
                               t3a8o_1_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t3a8o_1_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((t3a8o_1_1_argbuf_r && t3a8o_1_destruct_bufchan_buf[0]))
        t3a8o_1_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! t3a8o_1_1_argbuf_r) && (! t3a8o_1_destruct_bufchan_buf[0])))
        t3a8o_1_destruct_bufchan_buf <= t3a8o_1_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (t3a8z_1_destruct,Pointer_QTree_Int) > (t3a8z_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t t3a8z_1_destruct_bufchan_d;
  logic t3a8z_1_destruct_bufchan_r;
  assign t3a8z_1_destruct_r = ((! t3a8z_1_destruct_bufchan_d[0]) || t3a8z_1_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t3a8z_1_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (t3a8z_1_destruct_r)
        t3a8z_1_destruct_bufchan_d <= t3a8z_1_destruct_d;
  Pointer_QTree_Int_t t3a8z_1_destruct_bufchan_buf;
  assign t3a8z_1_destruct_bufchan_r = (! t3a8z_1_destruct_bufchan_buf[0]);
  assign t3a8z_1_1_argbuf_d = (t3a8z_1_destruct_bufchan_buf[0] ? t3a8z_1_destruct_bufchan_buf :
                               t3a8z_1_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t3a8z_1_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((t3a8z_1_1_argbuf_r && t3a8z_1_destruct_bufchan_buf[0]))
        t3a8z_1_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! t3a8z_1_1_argbuf_r) && (! t3a8z_1_destruct_bufchan_buf[0])))
        t3a8z_1_destruct_bufchan_buf <= t3a8z_1_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (t4a8A_destruct,Pointer_QTree_Int) > (t4a8A_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t t4a8A_destruct_bufchan_d;
  logic t4a8A_destruct_bufchan_r;
  assign t4a8A_destruct_r = ((! t4a8A_destruct_bufchan_d[0]) || t4a8A_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t4a8A_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (t4a8A_destruct_r) t4a8A_destruct_bufchan_d <= t4a8A_destruct_d;
  Pointer_QTree_Int_t t4a8A_destruct_bufchan_buf;
  assign t4a8A_destruct_bufchan_r = (! t4a8A_destruct_bufchan_buf[0]);
  assign t4a8A_1_argbuf_d = (t4a8A_destruct_bufchan_buf[0] ? t4a8A_destruct_bufchan_buf :
                             t4a8A_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t4a8A_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((t4a8A_1_argbuf_r && t4a8A_destruct_bufchan_buf[0]))
        t4a8A_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! t4a8A_1_argbuf_r) && (! t4a8A_destruct_bufchan_buf[0])))
        t4a8A_destruct_bufchan_buf <= t4a8A_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (t4a8p_destruct,Pointer_QTree_Int) > (t4a8p_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t t4a8p_destruct_bufchan_d;
  logic t4a8p_destruct_bufchan_r;
  assign t4a8p_destruct_r = ((! t4a8p_destruct_bufchan_d[0]) || t4a8p_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t4a8p_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (t4a8p_destruct_r) t4a8p_destruct_bufchan_d <= t4a8p_destruct_d;
  Pointer_QTree_Int_t t4a8p_destruct_bufchan_buf;
  assign t4a8p_destruct_bufchan_r = (! t4a8p_destruct_bufchan_buf[0]);
  assign t4a8p_1_argbuf_d = (t4a8p_destruct_bufchan_buf[0] ? t4a8p_destruct_bufchan_buf :
                             t4a8p_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t4a8p_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((t4a8p_1_argbuf_r && t4a8p_destruct_bufchan_buf[0]))
        t4a8p_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! t4a8p_1_argbuf_r) && (! t4a8p_destruct_bufchan_buf[0])))
        t4a8p_destruct_bufchan_buf <= t4a8p_destruct_bufchan_d;
  
  /* buf (Ty Int) : (va8c_destruct,Int) > (va8c_1_argbuf,Int) */
  Int_t va8c_destruct_bufchan_d;
  logic va8c_destruct_bufchan_r;
  assign va8c_destruct_r = ((! va8c_destruct_bufchan_d[0]) || va8c_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) va8c_destruct_bufchan_d <= {32'd0, 1'd0};
    else
      if (va8c_destruct_r) va8c_destruct_bufchan_d <= va8c_destruct_d;
  Int_t va8c_destruct_bufchan_buf;
  assign va8c_destruct_bufchan_r = (! va8c_destruct_bufchan_buf[0]);
  assign va8c_1_argbuf_d = (va8c_destruct_bufchan_buf[0] ? va8c_destruct_bufchan_buf :
                            va8c_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) va8c_destruct_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((va8c_1_argbuf_r && va8c_destruct_bufchan_buf[0]))
        va8c_destruct_bufchan_buf <= {32'd0, 1'd0};
      else if (((! va8c_1_argbuf_r) && (! va8c_destruct_bufchan_buf[0])))
        va8c_destruct_bufchan_buf <= va8c_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (w1sif_1_1,Pointer_QTree_Int) > (w1sif_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t w1sif_1_1_bufchan_d;
  logic w1sif_1_1_bufchan_r;
  assign w1sif_1_1_r = ((! w1sif_1_1_bufchan_d[0]) || w1sif_1_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) w1sif_1_1_bufchan_d <= {16'd0, 1'd0};
    else if (w1sif_1_1_r) w1sif_1_1_bufchan_d <= w1sif_1_1_d;
  Pointer_QTree_Int_t w1sif_1_1_bufchan_buf;
  assign w1sif_1_1_bufchan_r = (! w1sif_1_1_bufchan_buf[0]);
  assign w1sif_1_1_argbuf_d = (w1sif_1_1_bufchan_buf[0] ? w1sif_1_1_bufchan_buf :
                               w1sif_1_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) w1sif_1_1_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((w1sif_1_1_argbuf_r && w1sif_1_1_bufchan_buf[0]))
        w1sif_1_1_bufchan_buf <= {16'd0, 1'd0};
      else if (((! w1sif_1_1_argbuf_r) && (! w1sif_1_1_bufchan_buf[0])))
        w1sif_1_1_bufchan_buf <= w1sif_1_1_bufchan_d;
  
  /* fork (Ty Pointer_QTree_Int) : (w1sif_1_goMux_mux,Pointer_QTree_Int) > [(w1sif_1_1,Pointer_QTree_Int),
                                                                       (w1sif_1_2,Pointer_QTree_Int)] */
  logic [1:0] w1sif_1_goMux_mux_emitted;
  logic [1:0] w1sif_1_goMux_mux_done;
  assign w1sif_1_1_d = {w1sif_1_goMux_mux_d[16:1],
                        (w1sif_1_goMux_mux_d[0] && (! w1sif_1_goMux_mux_emitted[0]))};
  assign w1sif_1_2_d = {w1sif_1_goMux_mux_d[16:1],
                        (w1sif_1_goMux_mux_d[0] && (! w1sif_1_goMux_mux_emitted[1]))};
  assign w1sif_1_goMux_mux_done = (w1sif_1_goMux_mux_emitted | ({w1sif_1_2_d[0],
                                                                 w1sif_1_1_d[0]} & {w1sif_1_2_r,
                                                                                    w1sif_1_1_r}));
  assign w1sif_1_goMux_mux_r = (& w1sif_1_goMux_mux_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) w1sif_1_goMux_mux_emitted <= 2'd0;
    else
      w1sif_1_goMux_mux_emitted <= (w1sif_1_goMux_mux_r ? 2'd0 :
                                    w1sif_1_goMux_mux_done);
  
  /* buf (Ty Pointer_QTree_Int) : (w2sig_1_1,Pointer_QTree_Int) > (w2sig_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t w2sig_1_1_bufchan_d;
  logic w2sig_1_1_bufchan_r;
  assign w2sig_1_1_r = ((! w2sig_1_1_bufchan_d[0]) || w2sig_1_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) w2sig_1_1_bufchan_d <= {16'd0, 1'd0};
    else if (w2sig_1_1_r) w2sig_1_1_bufchan_d <= w2sig_1_1_d;
  Pointer_QTree_Int_t w2sig_1_1_bufchan_buf;
  assign w2sig_1_1_bufchan_r = (! w2sig_1_1_bufchan_buf[0]);
  assign w2sig_1_1_argbuf_d = (w2sig_1_1_bufchan_buf[0] ? w2sig_1_1_bufchan_buf :
                               w2sig_1_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) w2sig_1_1_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((w2sig_1_1_argbuf_r && w2sig_1_1_bufchan_buf[0]))
        w2sig_1_1_bufchan_buf <= {16'd0, 1'd0};
      else if (((! w2sig_1_1_argbuf_r) && (! w2sig_1_1_bufchan_buf[0])))
        w2sig_1_1_bufchan_buf <= w2sig_1_1_bufchan_d;
  
  /* fork (Ty Pointer_QTree_Int) : (w2sig_1_goMux_mux,Pointer_QTree_Int) > [(w2sig_1_1,Pointer_QTree_Int),
                                                                       (w2sig_1_2,Pointer_QTree_Int)] */
  logic [1:0] w2sig_1_goMux_mux_emitted;
  logic [1:0] w2sig_1_goMux_mux_done;
  assign w2sig_1_1_d = {w2sig_1_goMux_mux_d[16:1],
                        (w2sig_1_goMux_mux_d[0] && (! w2sig_1_goMux_mux_emitted[0]))};
  assign w2sig_1_2_d = {w2sig_1_goMux_mux_d[16:1],
                        (w2sig_1_goMux_mux_d[0] && (! w2sig_1_goMux_mux_emitted[1]))};
  assign w2sig_1_goMux_mux_done = (w2sig_1_goMux_mux_emitted | ({w2sig_1_2_d[0],
                                                                 w2sig_1_1_d[0]} & {w2sig_1_2_r,
                                                                                    w2sig_1_1_r}));
  assign w2sig_1_goMux_mux_r = (& w2sig_1_goMux_mux_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) w2sig_1_goMux_mux_emitted <= 2'd0;
    else
      w2sig_1_goMux_mux_emitted <= (w2sig_1_goMux_mux_r ? 2'd0 :
                                    w2sig_1_goMux_mux_done);
  
  /* buf (Ty Pointer_CT$wmAdd_Int) : (writeCT$wmAdd_IntlizzieLet0_1_argbuf,Pointer_CT$wmAdd_Int) > (writeCT$wmAdd_IntlizzieLet0_1_argbuf_rwb,Pointer_CT$wmAdd_Int) */
  Pointer_CT$wmAdd_Int_t writeCT$wmAdd_IntlizzieLet0_1_argbuf_bufchan_d;
  logic writeCT$wmAdd_IntlizzieLet0_1_argbuf_bufchan_r;
  assign writeCT$wmAdd_IntlizzieLet0_1_argbuf_r = ((! writeCT$wmAdd_IntlizzieLet0_1_argbuf_bufchan_d[0]) || writeCT$wmAdd_IntlizzieLet0_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wmAdd_IntlizzieLet0_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCT$wmAdd_IntlizzieLet0_1_argbuf_r)
        writeCT$wmAdd_IntlizzieLet0_1_argbuf_bufchan_d <= writeCT$wmAdd_IntlizzieLet0_1_argbuf_d;
  Pointer_CT$wmAdd_Int_t writeCT$wmAdd_IntlizzieLet0_1_argbuf_bufchan_buf;
  assign writeCT$wmAdd_IntlizzieLet0_1_argbuf_bufchan_r = (! writeCT$wmAdd_IntlizzieLet0_1_argbuf_bufchan_buf[0]);
  assign writeCT$wmAdd_IntlizzieLet0_1_argbuf_rwb_d = (writeCT$wmAdd_IntlizzieLet0_1_argbuf_bufchan_buf[0] ? writeCT$wmAdd_IntlizzieLet0_1_argbuf_bufchan_buf :
                                                       writeCT$wmAdd_IntlizzieLet0_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wmAdd_IntlizzieLet0_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeCT$wmAdd_IntlizzieLet0_1_argbuf_rwb_r && writeCT$wmAdd_IntlizzieLet0_1_argbuf_bufchan_buf[0]))
        writeCT$wmAdd_IntlizzieLet0_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeCT$wmAdd_IntlizzieLet0_1_argbuf_rwb_r) && (! writeCT$wmAdd_IntlizzieLet0_1_argbuf_bufchan_buf[0])))
        writeCT$wmAdd_IntlizzieLet0_1_argbuf_bufchan_buf <= writeCT$wmAdd_IntlizzieLet0_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CT$wmAdd_Int) : (writeCT$wmAdd_IntlizzieLet0_1_argbuf_rwb,Pointer_CT$wmAdd_Int) > (lizzieLet14_1_argbuf,Pointer_CT$wmAdd_Int) */
  Pointer_CT$wmAdd_Int_t writeCT$wmAdd_IntlizzieLet0_1_argbuf_rwb_bufchan_d;
  logic writeCT$wmAdd_IntlizzieLet0_1_argbuf_rwb_bufchan_r;
  assign writeCT$wmAdd_IntlizzieLet0_1_argbuf_rwb_r = ((! writeCT$wmAdd_IntlizzieLet0_1_argbuf_rwb_bufchan_d[0]) || writeCT$wmAdd_IntlizzieLet0_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wmAdd_IntlizzieLet0_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                             1'd0};
    else
      if (writeCT$wmAdd_IntlizzieLet0_1_argbuf_rwb_r)
        writeCT$wmAdd_IntlizzieLet0_1_argbuf_rwb_bufchan_d <= writeCT$wmAdd_IntlizzieLet0_1_argbuf_rwb_d;
  Pointer_CT$wmAdd_Int_t writeCT$wmAdd_IntlizzieLet0_1_argbuf_rwb_bufchan_buf;
  assign writeCT$wmAdd_IntlizzieLet0_1_argbuf_rwb_bufchan_r = (! writeCT$wmAdd_IntlizzieLet0_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet14_1_argbuf_d = (writeCT$wmAdd_IntlizzieLet0_1_argbuf_rwb_bufchan_buf[0] ? writeCT$wmAdd_IntlizzieLet0_1_argbuf_rwb_bufchan_buf :
                                   writeCT$wmAdd_IntlizzieLet0_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wmAdd_IntlizzieLet0_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
    else
      if ((lizzieLet14_1_argbuf_r && writeCT$wmAdd_IntlizzieLet0_1_argbuf_rwb_bufchan_buf[0]))
        writeCT$wmAdd_IntlizzieLet0_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                 1'd0};
      else if (((! lizzieLet14_1_argbuf_r) && (! writeCT$wmAdd_IntlizzieLet0_1_argbuf_rwb_bufchan_buf[0])))
        writeCT$wmAdd_IntlizzieLet0_1_argbuf_rwb_bufchan_buf <= writeCT$wmAdd_IntlizzieLet0_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CT$wmAdd_Int) : (writeCT$wmAdd_IntlizzieLet23_1_argbuf,Pointer_CT$wmAdd_Int) > (writeCT$wmAdd_IntlizzieLet23_1_argbuf_rwb,Pointer_CT$wmAdd_Int) */
  Pointer_CT$wmAdd_Int_t writeCT$wmAdd_IntlizzieLet23_1_argbuf_bufchan_d;
  logic writeCT$wmAdd_IntlizzieLet23_1_argbuf_bufchan_r;
  assign writeCT$wmAdd_IntlizzieLet23_1_argbuf_r = ((! writeCT$wmAdd_IntlizzieLet23_1_argbuf_bufchan_d[0]) || writeCT$wmAdd_IntlizzieLet23_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wmAdd_IntlizzieLet23_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCT$wmAdd_IntlizzieLet23_1_argbuf_r)
        writeCT$wmAdd_IntlizzieLet23_1_argbuf_bufchan_d <= writeCT$wmAdd_IntlizzieLet23_1_argbuf_d;
  Pointer_CT$wmAdd_Int_t writeCT$wmAdd_IntlizzieLet23_1_argbuf_bufchan_buf;
  assign writeCT$wmAdd_IntlizzieLet23_1_argbuf_bufchan_r = (! writeCT$wmAdd_IntlizzieLet23_1_argbuf_bufchan_buf[0]);
  assign writeCT$wmAdd_IntlizzieLet23_1_argbuf_rwb_d = (writeCT$wmAdd_IntlizzieLet23_1_argbuf_bufchan_buf[0] ? writeCT$wmAdd_IntlizzieLet23_1_argbuf_bufchan_buf :
                                                        writeCT$wmAdd_IntlizzieLet23_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wmAdd_IntlizzieLet23_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeCT$wmAdd_IntlizzieLet23_1_argbuf_rwb_r && writeCT$wmAdd_IntlizzieLet23_1_argbuf_bufchan_buf[0]))
        writeCT$wmAdd_IntlizzieLet23_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeCT$wmAdd_IntlizzieLet23_1_argbuf_rwb_r) && (! writeCT$wmAdd_IntlizzieLet23_1_argbuf_bufchan_buf[0])))
        writeCT$wmAdd_IntlizzieLet23_1_argbuf_bufchan_buf <= writeCT$wmAdd_IntlizzieLet23_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CT$wmAdd_Int) : (writeCT$wmAdd_IntlizzieLet23_1_argbuf_rwb,Pointer_CT$wmAdd_Int) > (sca2_1_argbuf,Pointer_CT$wmAdd_Int) */
  Pointer_CT$wmAdd_Int_t writeCT$wmAdd_IntlizzieLet23_1_argbuf_rwb_bufchan_d;
  logic writeCT$wmAdd_IntlizzieLet23_1_argbuf_rwb_bufchan_r;
  assign writeCT$wmAdd_IntlizzieLet23_1_argbuf_rwb_r = ((! writeCT$wmAdd_IntlizzieLet23_1_argbuf_rwb_bufchan_d[0]) || writeCT$wmAdd_IntlizzieLet23_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wmAdd_IntlizzieLet23_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                              1'd0};
    else
      if (writeCT$wmAdd_IntlizzieLet23_1_argbuf_rwb_r)
        writeCT$wmAdd_IntlizzieLet23_1_argbuf_rwb_bufchan_d <= writeCT$wmAdd_IntlizzieLet23_1_argbuf_rwb_d;
  Pointer_CT$wmAdd_Int_t writeCT$wmAdd_IntlizzieLet23_1_argbuf_rwb_bufchan_buf;
  assign writeCT$wmAdd_IntlizzieLet23_1_argbuf_rwb_bufchan_r = (! writeCT$wmAdd_IntlizzieLet23_1_argbuf_rwb_bufchan_buf[0]);
  assign sca2_1_argbuf_d = (writeCT$wmAdd_IntlizzieLet23_1_argbuf_rwb_bufchan_buf[0] ? writeCT$wmAdd_IntlizzieLet23_1_argbuf_rwb_bufchan_buf :
                            writeCT$wmAdd_IntlizzieLet23_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wmAdd_IntlizzieLet23_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
    else
      if ((sca2_1_argbuf_r && writeCT$wmAdd_IntlizzieLet23_1_argbuf_rwb_bufchan_buf[0]))
        writeCT$wmAdd_IntlizzieLet23_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                  1'd0};
      else if (((! sca2_1_argbuf_r) && (! writeCT$wmAdd_IntlizzieLet23_1_argbuf_rwb_bufchan_buf[0])))
        writeCT$wmAdd_IntlizzieLet23_1_argbuf_rwb_bufchan_buf <= writeCT$wmAdd_IntlizzieLet23_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CT$wmAdd_Int) : (writeCT$wmAdd_IntlizzieLet24_1_argbuf,Pointer_CT$wmAdd_Int) > (writeCT$wmAdd_IntlizzieLet24_1_argbuf_rwb,Pointer_CT$wmAdd_Int) */
  Pointer_CT$wmAdd_Int_t writeCT$wmAdd_IntlizzieLet24_1_argbuf_bufchan_d;
  logic writeCT$wmAdd_IntlizzieLet24_1_argbuf_bufchan_r;
  assign writeCT$wmAdd_IntlizzieLet24_1_argbuf_r = ((! writeCT$wmAdd_IntlizzieLet24_1_argbuf_bufchan_d[0]) || writeCT$wmAdd_IntlizzieLet24_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wmAdd_IntlizzieLet24_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCT$wmAdd_IntlizzieLet24_1_argbuf_r)
        writeCT$wmAdd_IntlizzieLet24_1_argbuf_bufchan_d <= writeCT$wmAdd_IntlizzieLet24_1_argbuf_d;
  Pointer_CT$wmAdd_Int_t writeCT$wmAdd_IntlizzieLet24_1_argbuf_bufchan_buf;
  assign writeCT$wmAdd_IntlizzieLet24_1_argbuf_bufchan_r = (! writeCT$wmAdd_IntlizzieLet24_1_argbuf_bufchan_buf[0]);
  assign writeCT$wmAdd_IntlizzieLet24_1_argbuf_rwb_d = (writeCT$wmAdd_IntlizzieLet24_1_argbuf_bufchan_buf[0] ? writeCT$wmAdd_IntlizzieLet24_1_argbuf_bufchan_buf :
                                                        writeCT$wmAdd_IntlizzieLet24_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wmAdd_IntlizzieLet24_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeCT$wmAdd_IntlizzieLet24_1_argbuf_rwb_r && writeCT$wmAdd_IntlizzieLet24_1_argbuf_bufchan_buf[0]))
        writeCT$wmAdd_IntlizzieLet24_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeCT$wmAdd_IntlizzieLet24_1_argbuf_rwb_r) && (! writeCT$wmAdd_IntlizzieLet24_1_argbuf_bufchan_buf[0])))
        writeCT$wmAdd_IntlizzieLet24_1_argbuf_bufchan_buf <= writeCT$wmAdd_IntlizzieLet24_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CT$wmAdd_Int) : (writeCT$wmAdd_IntlizzieLet24_1_argbuf_rwb,Pointer_CT$wmAdd_Int) > (sca1_1_argbuf,Pointer_CT$wmAdd_Int) */
  Pointer_CT$wmAdd_Int_t writeCT$wmAdd_IntlizzieLet24_1_argbuf_rwb_bufchan_d;
  logic writeCT$wmAdd_IntlizzieLet24_1_argbuf_rwb_bufchan_r;
  assign writeCT$wmAdd_IntlizzieLet24_1_argbuf_rwb_r = ((! writeCT$wmAdd_IntlizzieLet24_1_argbuf_rwb_bufchan_d[0]) || writeCT$wmAdd_IntlizzieLet24_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wmAdd_IntlizzieLet24_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                              1'd0};
    else
      if (writeCT$wmAdd_IntlizzieLet24_1_argbuf_rwb_r)
        writeCT$wmAdd_IntlizzieLet24_1_argbuf_rwb_bufchan_d <= writeCT$wmAdd_IntlizzieLet24_1_argbuf_rwb_d;
  Pointer_CT$wmAdd_Int_t writeCT$wmAdd_IntlizzieLet24_1_argbuf_rwb_bufchan_buf;
  assign writeCT$wmAdd_IntlizzieLet24_1_argbuf_rwb_bufchan_r = (! writeCT$wmAdd_IntlizzieLet24_1_argbuf_rwb_bufchan_buf[0]);
  assign sca1_1_argbuf_d = (writeCT$wmAdd_IntlizzieLet24_1_argbuf_rwb_bufchan_buf[0] ? writeCT$wmAdd_IntlizzieLet24_1_argbuf_rwb_bufchan_buf :
                            writeCT$wmAdd_IntlizzieLet24_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wmAdd_IntlizzieLet24_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
    else
      if ((sca1_1_argbuf_r && writeCT$wmAdd_IntlizzieLet24_1_argbuf_rwb_bufchan_buf[0]))
        writeCT$wmAdd_IntlizzieLet24_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                  1'd0};
      else if (((! sca1_1_argbuf_r) && (! writeCT$wmAdd_IntlizzieLet24_1_argbuf_rwb_bufchan_buf[0])))
        writeCT$wmAdd_IntlizzieLet24_1_argbuf_rwb_bufchan_buf <= writeCT$wmAdd_IntlizzieLet24_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CT$wmAdd_Int) : (writeCT$wmAdd_IntlizzieLet25_1_argbuf,Pointer_CT$wmAdd_Int) > (writeCT$wmAdd_IntlizzieLet25_1_argbuf_rwb,Pointer_CT$wmAdd_Int) */
  Pointer_CT$wmAdd_Int_t writeCT$wmAdd_IntlizzieLet25_1_argbuf_bufchan_d;
  logic writeCT$wmAdd_IntlizzieLet25_1_argbuf_bufchan_r;
  assign writeCT$wmAdd_IntlizzieLet25_1_argbuf_r = ((! writeCT$wmAdd_IntlizzieLet25_1_argbuf_bufchan_d[0]) || writeCT$wmAdd_IntlizzieLet25_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wmAdd_IntlizzieLet25_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCT$wmAdd_IntlizzieLet25_1_argbuf_r)
        writeCT$wmAdd_IntlizzieLet25_1_argbuf_bufchan_d <= writeCT$wmAdd_IntlizzieLet25_1_argbuf_d;
  Pointer_CT$wmAdd_Int_t writeCT$wmAdd_IntlizzieLet25_1_argbuf_bufchan_buf;
  assign writeCT$wmAdd_IntlizzieLet25_1_argbuf_bufchan_r = (! writeCT$wmAdd_IntlizzieLet25_1_argbuf_bufchan_buf[0]);
  assign writeCT$wmAdd_IntlizzieLet25_1_argbuf_rwb_d = (writeCT$wmAdd_IntlizzieLet25_1_argbuf_bufchan_buf[0] ? writeCT$wmAdd_IntlizzieLet25_1_argbuf_bufchan_buf :
                                                        writeCT$wmAdd_IntlizzieLet25_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wmAdd_IntlizzieLet25_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeCT$wmAdd_IntlizzieLet25_1_argbuf_rwb_r && writeCT$wmAdd_IntlizzieLet25_1_argbuf_bufchan_buf[0]))
        writeCT$wmAdd_IntlizzieLet25_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeCT$wmAdd_IntlizzieLet25_1_argbuf_rwb_r) && (! writeCT$wmAdd_IntlizzieLet25_1_argbuf_bufchan_buf[0])))
        writeCT$wmAdd_IntlizzieLet25_1_argbuf_bufchan_buf <= writeCT$wmAdd_IntlizzieLet25_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CT$wmAdd_Int) : (writeCT$wmAdd_IntlizzieLet25_1_argbuf_rwb,Pointer_CT$wmAdd_Int) > (sca0_1_argbuf,Pointer_CT$wmAdd_Int) */
  Pointer_CT$wmAdd_Int_t writeCT$wmAdd_IntlizzieLet25_1_argbuf_rwb_bufchan_d;
  logic writeCT$wmAdd_IntlizzieLet25_1_argbuf_rwb_bufchan_r;
  assign writeCT$wmAdd_IntlizzieLet25_1_argbuf_rwb_r = ((! writeCT$wmAdd_IntlizzieLet25_1_argbuf_rwb_bufchan_d[0]) || writeCT$wmAdd_IntlizzieLet25_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wmAdd_IntlizzieLet25_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                              1'd0};
    else
      if (writeCT$wmAdd_IntlizzieLet25_1_argbuf_rwb_r)
        writeCT$wmAdd_IntlizzieLet25_1_argbuf_rwb_bufchan_d <= writeCT$wmAdd_IntlizzieLet25_1_argbuf_rwb_d;
  Pointer_CT$wmAdd_Int_t writeCT$wmAdd_IntlizzieLet25_1_argbuf_rwb_bufchan_buf;
  assign writeCT$wmAdd_IntlizzieLet25_1_argbuf_rwb_bufchan_r = (! writeCT$wmAdd_IntlizzieLet25_1_argbuf_rwb_bufchan_buf[0]);
  assign sca0_1_argbuf_d = (writeCT$wmAdd_IntlizzieLet25_1_argbuf_rwb_bufchan_buf[0] ? writeCT$wmAdd_IntlizzieLet25_1_argbuf_rwb_bufchan_buf :
                            writeCT$wmAdd_IntlizzieLet25_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wmAdd_IntlizzieLet25_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
    else
      if ((sca0_1_argbuf_r && writeCT$wmAdd_IntlizzieLet25_1_argbuf_rwb_bufchan_buf[0]))
        writeCT$wmAdd_IntlizzieLet25_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                  1'd0};
      else if (((! sca0_1_argbuf_r) && (! writeCT$wmAdd_IntlizzieLet25_1_argbuf_rwb_bufchan_buf[0])))
        writeCT$wmAdd_IntlizzieLet25_1_argbuf_rwb_bufchan_buf <= writeCT$wmAdd_IntlizzieLet25_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CT$wmAdd_Int) : (writeCT$wmAdd_IntlizzieLet9_1_1_argbuf,Pointer_CT$wmAdd_Int) > (writeCT$wmAdd_IntlizzieLet9_1_1_argbuf_rwb,Pointer_CT$wmAdd_Int) */
  Pointer_CT$wmAdd_Int_t writeCT$wmAdd_IntlizzieLet9_1_1_argbuf_bufchan_d;
  logic writeCT$wmAdd_IntlizzieLet9_1_1_argbuf_bufchan_r;
  assign writeCT$wmAdd_IntlizzieLet9_1_1_argbuf_r = ((! writeCT$wmAdd_IntlizzieLet9_1_1_argbuf_bufchan_d[0]) || writeCT$wmAdd_IntlizzieLet9_1_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wmAdd_IntlizzieLet9_1_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCT$wmAdd_IntlizzieLet9_1_1_argbuf_r)
        writeCT$wmAdd_IntlizzieLet9_1_1_argbuf_bufchan_d <= writeCT$wmAdd_IntlizzieLet9_1_1_argbuf_d;
  Pointer_CT$wmAdd_Int_t writeCT$wmAdd_IntlizzieLet9_1_1_argbuf_bufchan_buf;
  assign writeCT$wmAdd_IntlizzieLet9_1_1_argbuf_bufchan_r = (! writeCT$wmAdd_IntlizzieLet9_1_1_argbuf_bufchan_buf[0]);
  assign writeCT$wmAdd_IntlizzieLet9_1_1_argbuf_rwb_d = (writeCT$wmAdd_IntlizzieLet9_1_1_argbuf_bufchan_buf[0] ? writeCT$wmAdd_IntlizzieLet9_1_1_argbuf_bufchan_buf :
                                                         writeCT$wmAdd_IntlizzieLet9_1_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wmAdd_IntlizzieLet9_1_1_argbuf_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((writeCT$wmAdd_IntlizzieLet9_1_1_argbuf_rwb_r && writeCT$wmAdd_IntlizzieLet9_1_1_argbuf_bufchan_buf[0]))
        writeCT$wmAdd_IntlizzieLet9_1_1_argbuf_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! writeCT$wmAdd_IntlizzieLet9_1_1_argbuf_rwb_r) && (! writeCT$wmAdd_IntlizzieLet9_1_1_argbuf_bufchan_buf[0])))
        writeCT$wmAdd_IntlizzieLet9_1_1_argbuf_bufchan_buf <= writeCT$wmAdd_IntlizzieLet9_1_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CT$wmAdd_Int) : (writeCT$wmAdd_IntlizzieLet9_1_1_argbuf_rwb,Pointer_CT$wmAdd_Int) > (sca3_1_argbuf,Pointer_CT$wmAdd_Int) */
  Pointer_CT$wmAdd_Int_t writeCT$wmAdd_IntlizzieLet9_1_1_argbuf_rwb_bufchan_d;
  logic writeCT$wmAdd_IntlizzieLet9_1_1_argbuf_rwb_bufchan_r;
  assign writeCT$wmAdd_IntlizzieLet9_1_1_argbuf_rwb_r = ((! writeCT$wmAdd_IntlizzieLet9_1_1_argbuf_rwb_bufchan_d[0]) || writeCT$wmAdd_IntlizzieLet9_1_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wmAdd_IntlizzieLet9_1_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                               1'd0};
    else
      if (writeCT$wmAdd_IntlizzieLet9_1_1_argbuf_rwb_r)
        writeCT$wmAdd_IntlizzieLet9_1_1_argbuf_rwb_bufchan_d <= writeCT$wmAdd_IntlizzieLet9_1_1_argbuf_rwb_d;
  Pointer_CT$wmAdd_Int_t writeCT$wmAdd_IntlizzieLet9_1_1_argbuf_rwb_bufchan_buf;
  assign writeCT$wmAdd_IntlizzieLet9_1_1_argbuf_rwb_bufchan_r = (! writeCT$wmAdd_IntlizzieLet9_1_1_argbuf_rwb_bufchan_buf[0]);
  assign sca3_1_argbuf_d = (writeCT$wmAdd_IntlizzieLet9_1_1_argbuf_rwb_bufchan_buf[0] ? writeCT$wmAdd_IntlizzieLet9_1_1_argbuf_rwb_bufchan_buf :
                            writeCT$wmAdd_IntlizzieLet9_1_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wmAdd_IntlizzieLet9_1_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                 1'd0};
    else
      if ((sca3_1_argbuf_r && writeCT$wmAdd_IntlizzieLet9_1_1_argbuf_rwb_bufchan_buf[0]))
        writeCT$wmAdd_IntlizzieLet9_1_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                   1'd0};
      else if (((! sca3_1_argbuf_r) && (! writeCT$wmAdd_IntlizzieLet9_1_1_argbuf_rwb_bufchan_buf[0])))
        writeCT$wmAdd_IntlizzieLet9_1_1_argbuf_rwb_bufchan_buf <= writeCT$wmAdd_IntlizzieLet9_1_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz_Int) : (writeCT$wnnz_IntlizzieLet13_1_1_argbuf,Pointer_CT$wnnz_Int) > (writeCT$wnnz_IntlizzieLet13_1_1_argbuf_rwb,Pointer_CT$wnnz_Int) */
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet13_1_1_argbuf_bufchan_d;
  logic writeCT$wnnz_IntlizzieLet13_1_1_argbuf_bufchan_r;
  assign writeCT$wnnz_IntlizzieLet13_1_1_argbuf_r = ((! writeCT$wnnz_IntlizzieLet13_1_1_argbuf_bufchan_d[0]) || writeCT$wnnz_IntlizzieLet13_1_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnz_IntlizzieLet13_1_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCT$wnnz_IntlizzieLet13_1_1_argbuf_r)
        writeCT$wnnz_IntlizzieLet13_1_1_argbuf_bufchan_d <= writeCT$wnnz_IntlizzieLet13_1_1_argbuf_d;
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet13_1_1_argbuf_bufchan_buf;
  assign writeCT$wnnz_IntlizzieLet13_1_1_argbuf_bufchan_r = (! writeCT$wnnz_IntlizzieLet13_1_1_argbuf_bufchan_buf[0]);
  assign writeCT$wnnz_IntlizzieLet13_1_1_argbuf_rwb_d = (writeCT$wnnz_IntlizzieLet13_1_1_argbuf_bufchan_buf[0] ? writeCT$wnnz_IntlizzieLet13_1_1_argbuf_bufchan_buf :
                                                         writeCT$wnnz_IntlizzieLet13_1_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnz_IntlizzieLet13_1_1_argbuf_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((writeCT$wnnz_IntlizzieLet13_1_1_argbuf_rwb_r && writeCT$wnnz_IntlizzieLet13_1_1_argbuf_bufchan_buf[0]))
        writeCT$wnnz_IntlizzieLet13_1_1_argbuf_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! writeCT$wnnz_IntlizzieLet13_1_1_argbuf_rwb_r) && (! writeCT$wnnz_IntlizzieLet13_1_1_argbuf_bufchan_buf[0])))
        writeCT$wnnz_IntlizzieLet13_1_1_argbuf_bufchan_buf <= writeCT$wnnz_IntlizzieLet13_1_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz_Int) : (writeCT$wnnz_IntlizzieLet13_1_1_argbuf_rwb,Pointer_CT$wnnz_Int) > (sca3_1_1_argbuf,Pointer_CT$wnnz_Int) */
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet13_1_1_argbuf_rwb_bufchan_d;
  logic writeCT$wnnz_IntlizzieLet13_1_1_argbuf_rwb_bufchan_r;
  assign writeCT$wnnz_IntlizzieLet13_1_1_argbuf_rwb_r = ((! writeCT$wnnz_IntlizzieLet13_1_1_argbuf_rwb_bufchan_d[0]) || writeCT$wnnz_IntlizzieLet13_1_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnz_IntlizzieLet13_1_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                               1'd0};
    else
      if (writeCT$wnnz_IntlizzieLet13_1_1_argbuf_rwb_r)
        writeCT$wnnz_IntlizzieLet13_1_1_argbuf_rwb_bufchan_d <= writeCT$wnnz_IntlizzieLet13_1_1_argbuf_rwb_d;
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet13_1_1_argbuf_rwb_bufchan_buf;
  assign writeCT$wnnz_IntlizzieLet13_1_1_argbuf_rwb_bufchan_r = (! writeCT$wnnz_IntlizzieLet13_1_1_argbuf_rwb_bufchan_buf[0]);
  assign sca3_1_1_argbuf_d = (writeCT$wnnz_IntlizzieLet13_1_1_argbuf_rwb_bufchan_buf[0] ? writeCT$wnnz_IntlizzieLet13_1_1_argbuf_rwb_bufchan_buf :
                              writeCT$wnnz_IntlizzieLet13_1_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnz_IntlizzieLet13_1_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                 1'd0};
    else
      if ((sca3_1_1_argbuf_r && writeCT$wnnz_IntlizzieLet13_1_1_argbuf_rwb_bufchan_buf[0]))
        writeCT$wnnz_IntlizzieLet13_1_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                   1'd0};
      else if (((! sca3_1_1_argbuf_r) && (! writeCT$wnnz_IntlizzieLet13_1_1_argbuf_rwb_bufchan_buf[0])))
        writeCT$wnnz_IntlizzieLet13_1_1_argbuf_rwb_bufchan_buf <= writeCT$wnnz_IntlizzieLet13_1_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz_Int) : (writeCT$wnnz_IntlizzieLet1_1_argbuf,Pointer_CT$wnnz_Int) > (writeCT$wnnz_IntlizzieLet1_1_argbuf_rwb,Pointer_CT$wnnz_Int) */
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet1_1_argbuf_bufchan_d;
  logic writeCT$wnnz_IntlizzieLet1_1_argbuf_bufchan_r;
  assign writeCT$wnnz_IntlizzieLet1_1_argbuf_r = ((! writeCT$wnnz_IntlizzieLet1_1_argbuf_bufchan_d[0]) || writeCT$wnnz_IntlizzieLet1_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnz_IntlizzieLet1_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCT$wnnz_IntlizzieLet1_1_argbuf_r)
        writeCT$wnnz_IntlizzieLet1_1_argbuf_bufchan_d <= writeCT$wnnz_IntlizzieLet1_1_argbuf_d;
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet1_1_argbuf_bufchan_buf;
  assign writeCT$wnnz_IntlizzieLet1_1_argbuf_bufchan_r = (! writeCT$wnnz_IntlizzieLet1_1_argbuf_bufchan_buf[0]);
  assign writeCT$wnnz_IntlizzieLet1_1_argbuf_rwb_d = (writeCT$wnnz_IntlizzieLet1_1_argbuf_bufchan_buf[0] ? writeCT$wnnz_IntlizzieLet1_1_argbuf_bufchan_buf :
                                                      writeCT$wnnz_IntlizzieLet1_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnz_IntlizzieLet1_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeCT$wnnz_IntlizzieLet1_1_argbuf_rwb_r && writeCT$wnnz_IntlizzieLet1_1_argbuf_bufchan_buf[0]))
        writeCT$wnnz_IntlizzieLet1_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeCT$wnnz_IntlizzieLet1_1_argbuf_rwb_r) && (! writeCT$wnnz_IntlizzieLet1_1_argbuf_bufchan_buf[0])))
        writeCT$wnnz_IntlizzieLet1_1_argbuf_bufchan_buf <= writeCT$wnnz_IntlizzieLet1_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz_Int) : (writeCT$wnnz_IntlizzieLet1_1_argbuf_rwb,Pointer_CT$wnnz_Int) > (lizzieLet7_1_argbuf,Pointer_CT$wnnz_Int) */
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet1_1_argbuf_rwb_bufchan_d;
  logic writeCT$wnnz_IntlizzieLet1_1_argbuf_rwb_bufchan_r;
  assign writeCT$wnnz_IntlizzieLet1_1_argbuf_rwb_r = ((! writeCT$wnnz_IntlizzieLet1_1_argbuf_rwb_bufchan_d[0]) || writeCT$wnnz_IntlizzieLet1_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnz_IntlizzieLet1_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCT$wnnz_IntlizzieLet1_1_argbuf_rwb_r)
        writeCT$wnnz_IntlizzieLet1_1_argbuf_rwb_bufchan_d <= writeCT$wnnz_IntlizzieLet1_1_argbuf_rwb_d;
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet1_1_argbuf_rwb_bufchan_buf;
  assign writeCT$wnnz_IntlizzieLet1_1_argbuf_rwb_bufchan_r = (! writeCT$wnnz_IntlizzieLet1_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet7_1_argbuf_d = (writeCT$wnnz_IntlizzieLet1_1_argbuf_rwb_bufchan_buf[0] ? writeCT$wnnz_IntlizzieLet1_1_argbuf_rwb_bufchan_buf :
                                  writeCT$wnnz_IntlizzieLet1_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnz_IntlizzieLet1_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                              1'd0};
    else
      if ((lizzieLet7_1_argbuf_r && writeCT$wnnz_IntlizzieLet1_1_argbuf_rwb_bufchan_buf[0]))
        writeCT$wnnz_IntlizzieLet1_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
      else if (((! lizzieLet7_1_argbuf_r) && (! writeCT$wnnz_IntlizzieLet1_1_argbuf_rwb_bufchan_buf[0])))
        writeCT$wnnz_IntlizzieLet1_1_argbuf_rwb_bufchan_buf <= writeCT$wnnz_IntlizzieLet1_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz_Int) : (writeCT$wnnz_IntlizzieLet28_1_argbuf,Pointer_CT$wnnz_Int) > (writeCT$wnnz_IntlizzieLet28_1_argbuf_rwb,Pointer_CT$wnnz_Int) */
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet28_1_argbuf_bufchan_d;
  logic writeCT$wnnz_IntlizzieLet28_1_argbuf_bufchan_r;
  assign writeCT$wnnz_IntlizzieLet28_1_argbuf_r = ((! writeCT$wnnz_IntlizzieLet28_1_argbuf_bufchan_d[0]) || writeCT$wnnz_IntlizzieLet28_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnz_IntlizzieLet28_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCT$wnnz_IntlizzieLet28_1_argbuf_r)
        writeCT$wnnz_IntlizzieLet28_1_argbuf_bufchan_d <= writeCT$wnnz_IntlizzieLet28_1_argbuf_d;
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet28_1_argbuf_bufchan_buf;
  assign writeCT$wnnz_IntlizzieLet28_1_argbuf_bufchan_r = (! writeCT$wnnz_IntlizzieLet28_1_argbuf_bufchan_buf[0]);
  assign writeCT$wnnz_IntlizzieLet28_1_argbuf_rwb_d = (writeCT$wnnz_IntlizzieLet28_1_argbuf_bufchan_buf[0] ? writeCT$wnnz_IntlizzieLet28_1_argbuf_bufchan_buf :
                                                       writeCT$wnnz_IntlizzieLet28_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnz_IntlizzieLet28_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeCT$wnnz_IntlizzieLet28_1_argbuf_rwb_r && writeCT$wnnz_IntlizzieLet28_1_argbuf_bufchan_buf[0]))
        writeCT$wnnz_IntlizzieLet28_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeCT$wnnz_IntlizzieLet28_1_argbuf_rwb_r) && (! writeCT$wnnz_IntlizzieLet28_1_argbuf_bufchan_buf[0])))
        writeCT$wnnz_IntlizzieLet28_1_argbuf_bufchan_buf <= writeCT$wnnz_IntlizzieLet28_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz_Int) : (writeCT$wnnz_IntlizzieLet28_1_argbuf_rwb,Pointer_CT$wnnz_Int) > (sca2_1_1_argbuf,Pointer_CT$wnnz_Int) */
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet28_1_argbuf_rwb_bufchan_d;
  logic writeCT$wnnz_IntlizzieLet28_1_argbuf_rwb_bufchan_r;
  assign writeCT$wnnz_IntlizzieLet28_1_argbuf_rwb_r = ((! writeCT$wnnz_IntlizzieLet28_1_argbuf_rwb_bufchan_d[0]) || writeCT$wnnz_IntlizzieLet28_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnz_IntlizzieLet28_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                             1'd0};
    else
      if (writeCT$wnnz_IntlizzieLet28_1_argbuf_rwb_r)
        writeCT$wnnz_IntlizzieLet28_1_argbuf_rwb_bufchan_d <= writeCT$wnnz_IntlizzieLet28_1_argbuf_rwb_d;
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet28_1_argbuf_rwb_bufchan_buf;
  assign writeCT$wnnz_IntlizzieLet28_1_argbuf_rwb_bufchan_r = (! writeCT$wnnz_IntlizzieLet28_1_argbuf_rwb_bufchan_buf[0]);
  assign sca2_1_1_argbuf_d = (writeCT$wnnz_IntlizzieLet28_1_argbuf_rwb_bufchan_buf[0] ? writeCT$wnnz_IntlizzieLet28_1_argbuf_rwb_bufchan_buf :
                              writeCT$wnnz_IntlizzieLet28_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnz_IntlizzieLet28_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
    else
      if ((sca2_1_1_argbuf_r && writeCT$wnnz_IntlizzieLet28_1_argbuf_rwb_bufchan_buf[0]))
        writeCT$wnnz_IntlizzieLet28_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                 1'd0};
      else if (((! sca2_1_1_argbuf_r) && (! writeCT$wnnz_IntlizzieLet28_1_argbuf_rwb_bufchan_buf[0])))
        writeCT$wnnz_IntlizzieLet28_1_argbuf_rwb_bufchan_buf <= writeCT$wnnz_IntlizzieLet28_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz_Int) : (writeCT$wnnz_IntlizzieLet29_1_argbuf,Pointer_CT$wnnz_Int) > (writeCT$wnnz_IntlizzieLet29_1_argbuf_rwb,Pointer_CT$wnnz_Int) */
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet29_1_argbuf_bufchan_d;
  logic writeCT$wnnz_IntlizzieLet29_1_argbuf_bufchan_r;
  assign writeCT$wnnz_IntlizzieLet29_1_argbuf_r = ((! writeCT$wnnz_IntlizzieLet29_1_argbuf_bufchan_d[0]) || writeCT$wnnz_IntlizzieLet29_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnz_IntlizzieLet29_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCT$wnnz_IntlizzieLet29_1_argbuf_r)
        writeCT$wnnz_IntlizzieLet29_1_argbuf_bufchan_d <= writeCT$wnnz_IntlizzieLet29_1_argbuf_d;
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet29_1_argbuf_bufchan_buf;
  assign writeCT$wnnz_IntlizzieLet29_1_argbuf_bufchan_r = (! writeCT$wnnz_IntlizzieLet29_1_argbuf_bufchan_buf[0]);
  assign writeCT$wnnz_IntlizzieLet29_1_argbuf_rwb_d = (writeCT$wnnz_IntlizzieLet29_1_argbuf_bufchan_buf[0] ? writeCT$wnnz_IntlizzieLet29_1_argbuf_bufchan_buf :
                                                       writeCT$wnnz_IntlizzieLet29_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnz_IntlizzieLet29_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeCT$wnnz_IntlizzieLet29_1_argbuf_rwb_r && writeCT$wnnz_IntlizzieLet29_1_argbuf_bufchan_buf[0]))
        writeCT$wnnz_IntlizzieLet29_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeCT$wnnz_IntlizzieLet29_1_argbuf_rwb_r) && (! writeCT$wnnz_IntlizzieLet29_1_argbuf_bufchan_buf[0])))
        writeCT$wnnz_IntlizzieLet29_1_argbuf_bufchan_buf <= writeCT$wnnz_IntlizzieLet29_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz_Int) : (writeCT$wnnz_IntlizzieLet29_1_argbuf_rwb,Pointer_CT$wnnz_Int) > (sca1_1_1_argbuf,Pointer_CT$wnnz_Int) */
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet29_1_argbuf_rwb_bufchan_d;
  logic writeCT$wnnz_IntlizzieLet29_1_argbuf_rwb_bufchan_r;
  assign writeCT$wnnz_IntlizzieLet29_1_argbuf_rwb_r = ((! writeCT$wnnz_IntlizzieLet29_1_argbuf_rwb_bufchan_d[0]) || writeCT$wnnz_IntlizzieLet29_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnz_IntlizzieLet29_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                             1'd0};
    else
      if (writeCT$wnnz_IntlizzieLet29_1_argbuf_rwb_r)
        writeCT$wnnz_IntlizzieLet29_1_argbuf_rwb_bufchan_d <= writeCT$wnnz_IntlizzieLet29_1_argbuf_rwb_d;
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet29_1_argbuf_rwb_bufchan_buf;
  assign writeCT$wnnz_IntlizzieLet29_1_argbuf_rwb_bufchan_r = (! writeCT$wnnz_IntlizzieLet29_1_argbuf_rwb_bufchan_buf[0]);
  assign sca1_1_1_argbuf_d = (writeCT$wnnz_IntlizzieLet29_1_argbuf_rwb_bufchan_buf[0] ? writeCT$wnnz_IntlizzieLet29_1_argbuf_rwb_bufchan_buf :
                              writeCT$wnnz_IntlizzieLet29_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnz_IntlizzieLet29_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
    else
      if ((sca1_1_1_argbuf_r && writeCT$wnnz_IntlizzieLet29_1_argbuf_rwb_bufchan_buf[0]))
        writeCT$wnnz_IntlizzieLet29_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                 1'd0};
      else if (((! sca1_1_1_argbuf_r) && (! writeCT$wnnz_IntlizzieLet29_1_argbuf_rwb_bufchan_buf[0])))
        writeCT$wnnz_IntlizzieLet29_1_argbuf_rwb_bufchan_buf <= writeCT$wnnz_IntlizzieLet29_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz_Int) : (writeCT$wnnz_IntlizzieLet30_1_argbuf,Pointer_CT$wnnz_Int) > (writeCT$wnnz_IntlizzieLet30_1_argbuf_rwb,Pointer_CT$wnnz_Int) */
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet30_1_argbuf_bufchan_d;
  logic writeCT$wnnz_IntlizzieLet30_1_argbuf_bufchan_r;
  assign writeCT$wnnz_IntlizzieLet30_1_argbuf_r = ((! writeCT$wnnz_IntlizzieLet30_1_argbuf_bufchan_d[0]) || writeCT$wnnz_IntlizzieLet30_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnz_IntlizzieLet30_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCT$wnnz_IntlizzieLet30_1_argbuf_r)
        writeCT$wnnz_IntlizzieLet30_1_argbuf_bufchan_d <= writeCT$wnnz_IntlizzieLet30_1_argbuf_d;
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet30_1_argbuf_bufchan_buf;
  assign writeCT$wnnz_IntlizzieLet30_1_argbuf_bufchan_r = (! writeCT$wnnz_IntlizzieLet30_1_argbuf_bufchan_buf[0]);
  assign writeCT$wnnz_IntlizzieLet30_1_argbuf_rwb_d = (writeCT$wnnz_IntlizzieLet30_1_argbuf_bufchan_buf[0] ? writeCT$wnnz_IntlizzieLet30_1_argbuf_bufchan_buf :
                                                       writeCT$wnnz_IntlizzieLet30_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnz_IntlizzieLet30_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeCT$wnnz_IntlizzieLet30_1_argbuf_rwb_r && writeCT$wnnz_IntlizzieLet30_1_argbuf_bufchan_buf[0]))
        writeCT$wnnz_IntlizzieLet30_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeCT$wnnz_IntlizzieLet30_1_argbuf_rwb_r) && (! writeCT$wnnz_IntlizzieLet30_1_argbuf_bufchan_buf[0])))
        writeCT$wnnz_IntlizzieLet30_1_argbuf_bufchan_buf <= writeCT$wnnz_IntlizzieLet30_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz_Int) : (writeCT$wnnz_IntlizzieLet30_1_argbuf_rwb,Pointer_CT$wnnz_Int) > (sca0_1_1_argbuf,Pointer_CT$wnnz_Int) */
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet30_1_argbuf_rwb_bufchan_d;
  logic writeCT$wnnz_IntlizzieLet30_1_argbuf_rwb_bufchan_r;
  assign writeCT$wnnz_IntlizzieLet30_1_argbuf_rwb_r = ((! writeCT$wnnz_IntlizzieLet30_1_argbuf_rwb_bufchan_d[0]) || writeCT$wnnz_IntlizzieLet30_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnz_IntlizzieLet30_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                             1'd0};
    else
      if (writeCT$wnnz_IntlizzieLet30_1_argbuf_rwb_r)
        writeCT$wnnz_IntlizzieLet30_1_argbuf_rwb_bufchan_d <= writeCT$wnnz_IntlizzieLet30_1_argbuf_rwb_d;
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet30_1_argbuf_rwb_bufchan_buf;
  assign writeCT$wnnz_IntlizzieLet30_1_argbuf_rwb_bufchan_r = (! writeCT$wnnz_IntlizzieLet30_1_argbuf_rwb_bufchan_buf[0]);
  assign sca0_1_1_argbuf_d = (writeCT$wnnz_IntlizzieLet30_1_argbuf_rwb_bufchan_buf[0] ? writeCT$wnnz_IntlizzieLet30_1_argbuf_rwb_bufchan_buf :
                              writeCT$wnnz_IntlizzieLet30_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnz_IntlizzieLet30_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
    else
      if ((sca0_1_1_argbuf_r && writeCT$wnnz_IntlizzieLet30_1_argbuf_rwb_bufchan_buf[0]))
        writeCT$wnnz_IntlizzieLet30_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                 1'd0};
      else if (((! sca0_1_1_argbuf_r) && (! writeCT$wnnz_IntlizzieLet30_1_argbuf_rwb_bufchan_buf[0])))
        writeCT$wnnz_IntlizzieLet30_1_argbuf_rwb_bufchan_buf <= writeCT$wnnz_IntlizzieLet30_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CTmain_mask_Int) : (writeCTmain_mask_IntlizzieLet19_1_argbuf,Pointer_CTmain_mask_Int) > (writeCTmain_mask_IntlizzieLet19_1_argbuf_rwb,Pointer_CTmain_mask_Int) */
  Pointer_CTmain_mask_Int_t writeCTmain_mask_IntlizzieLet19_1_argbuf_bufchan_d;
  logic writeCTmain_mask_IntlizzieLet19_1_argbuf_bufchan_r;
  assign writeCTmain_mask_IntlizzieLet19_1_argbuf_r = ((! writeCTmain_mask_IntlizzieLet19_1_argbuf_bufchan_d[0]) || writeCTmain_mask_IntlizzieLet19_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTmain_mask_IntlizzieLet19_1_argbuf_bufchan_d <= {16'd0,
                                                             1'd0};
    else
      if (writeCTmain_mask_IntlizzieLet19_1_argbuf_r)
        writeCTmain_mask_IntlizzieLet19_1_argbuf_bufchan_d <= writeCTmain_mask_IntlizzieLet19_1_argbuf_d;
  Pointer_CTmain_mask_Int_t writeCTmain_mask_IntlizzieLet19_1_argbuf_bufchan_buf;
  assign writeCTmain_mask_IntlizzieLet19_1_argbuf_bufchan_r = (! writeCTmain_mask_IntlizzieLet19_1_argbuf_bufchan_buf[0]);
  assign writeCTmain_mask_IntlizzieLet19_1_argbuf_rwb_d = (writeCTmain_mask_IntlizzieLet19_1_argbuf_bufchan_buf[0] ? writeCTmain_mask_IntlizzieLet19_1_argbuf_bufchan_buf :
                                                           writeCTmain_mask_IntlizzieLet19_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTmain_mask_IntlizzieLet19_1_argbuf_bufchan_buf <= {16'd0,
                                                               1'd0};
    else
      if ((writeCTmain_mask_IntlizzieLet19_1_argbuf_rwb_r && writeCTmain_mask_IntlizzieLet19_1_argbuf_bufchan_buf[0]))
        writeCTmain_mask_IntlizzieLet19_1_argbuf_bufchan_buf <= {16'd0,
                                                                 1'd0};
      else if (((! writeCTmain_mask_IntlizzieLet19_1_argbuf_rwb_r) && (! writeCTmain_mask_IntlizzieLet19_1_argbuf_bufchan_buf[0])))
        writeCTmain_mask_IntlizzieLet19_1_argbuf_bufchan_buf <= writeCTmain_mask_IntlizzieLet19_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CTmain_mask_Int) : (writeCTmain_mask_IntlizzieLet19_1_argbuf_rwb,Pointer_CTmain_mask_Int) > (sca3_2_1_argbuf,Pointer_CTmain_mask_Int) */
  Pointer_CTmain_mask_Int_t writeCTmain_mask_IntlizzieLet19_1_argbuf_rwb_bufchan_d;
  logic writeCTmain_mask_IntlizzieLet19_1_argbuf_rwb_bufchan_r;
  assign writeCTmain_mask_IntlizzieLet19_1_argbuf_rwb_r = ((! writeCTmain_mask_IntlizzieLet19_1_argbuf_rwb_bufchan_d[0]) || writeCTmain_mask_IntlizzieLet19_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTmain_mask_IntlizzieLet19_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                                 1'd0};
    else
      if (writeCTmain_mask_IntlizzieLet19_1_argbuf_rwb_r)
        writeCTmain_mask_IntlizzieLet19_1_argbuf_rwb_bufchan_d <= writeCTmain_mask_IntlizzieLet19_1_argbuf_rwb_d;
  Pointer_CTmain_mask_Int_t writeCTmain_mask_IntlizzieLet19_1_argbuf_rwb_bufchan_buf;
  assign writeCTmain_mask_IntlizzieLet19_1_argbuf_rwb_bufchan_r = (! writeCTmain_mask_IntlizzieLet19_1_argbuf_rwb_bufchan_buf[0]);
  assign sca3_2_1_argbuf_d = (writeCTmain_mask_IntlizzieLet19_1_argbuf_rwb_bufchan_buf[0] ? writeCTmain_mask_IntlizzieLet19_1_argbuf_rwb_bufchan_buf :
                              writeCTmain_mask_IntlizzieLet19_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTmain_mask_IntlizzieLet19_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                   1'd0};
    else
      if ((sca3_2_1_argbuf_r && writeCTmain_mask_IntlizzieLet19_1_argbuf_rwb_bufchan_buf[0]))
        writeCTmain_mask_IntlizzieLet19_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                     1'd0};
      else if (((! sca3_2_1_argbuf_r) && (! writeCTmain_mask_IntlizzieLet19_1_argbuf_rwb_bufchan_buf[0])))
        writeCTmain_mask_IntlizzieLet19_1_argbuf_rwb_bufchan_buf <= writeCTmain_mask_IntlizzieLet19_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CTmain_mask_Int) : (writeCTmain_mask_IntlizzieLet21_1_argbuf,Pointer_CTmain_mask_Int) > (writeCTmain_mask_IntlizzieLet21_1_argbuf_rwb,Pointer_CTmain_mask_Int) */
  Pointer_CTmain_mask_Int_t writeCTmain_mask_IntlizzieLet21_1_argbuf_bufchan_d;
  logic writeCTmain_mask_IntlizzieLet21_1_argbuf_bufchan_r;
  assign writeCTmain_mask_IntlizzieLet21_1_argbuf_r = ((! writeCTmain_mask_IntlizzieLet21_1_argbuf_bufchan_d[0]) || writeCTmain_mask_IntlizzieLet21_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTmain_mask_IntlizzieLet21_1_argbuf_bufchan_d <= {16'd0,
                                                             1'd0};
    else
      if (writeCTmain_mask_IntlizzieLet21_1_argbuf_r)
        writeCTmain_mask_IntlizzieLet21_1_argbuf_bufchan_d <= writeCTmain_mask_IntlizzieLet21_1_argbuf_d;
  Pointer_CTmain_mask_Int_t writeCTmain_mask_IntlizzieLet21_1_argbuf_bufchan_buf;
  assign writeCTmain_mask_IntlizzieLet21_1_argbuf_bufchan_r = (! writeCTmain_mask_IntlizzieLet21_1_argbuf_bufchan_buf[0]);
  assign writeCTmain_mask_IntlizzieLet21_1_argbuf_rwb_d = (writeCTmain_mask_IntlizzieLet21_1_argbuf_bufchan_buf[0] ? writeCTmain_mask_IntlizzieLet21_1_argbuf_bufchan_buf :
                                                           writeCTmain_mask_IntlizzieLet21_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTmain_mask_IntlizzieLet21_1_argbuf_bufchan_buf <= {16'd0,
                                                               1'd0};
    else
      if ((writeCTmain_mask_IntlizzieLet21_1_argbuf_rwb_r && writeCTmain_mask_IntlizzieLet21_1_argbuf_bufchan_buf[0]))
        writeCTmain_mask_IntlizzieLet21_1_argbuf_bufchan_buf <= {16'd0,
                                                                 1'd0};
      else if (((! writeCTmain_mask_IntlizzieLet21_1_argbuf_rwb_r) && (! writeCTmain_mask_IntlizzieLet21_1_argbuf_bufchan_buf[0])))
        writeCTmain_mask_IntlizzieLet21_1_argbuf_bufchan_buf <= writeCTmain_mask_IntlizzieLet21_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CTmain_mask_Int) : (writeCTmain_mask_IntlizzieLet21_1_argbuf_rwb,Pointer_CTmain_mask_Int) > (lizzieLet4_1_1_argbuf,Pointer_CTmain_mask_Int) */
  Pointer_CTmain_mask_Int_t writeCTmain_mask_IntlizzieLet21_1_argbuf_rwb_bufchan_d;
  logic writeCTmain_mask_IntlizzieLet21_1_argbuf_rwb_bufchan_r;
  assign writeCTmain_mask_IntlizzieLet21_1_argbuf_rwb_r = ((! writeCTmain_mask_IntlizzieLet21_1_argbuf_rwb_bufchan_d[0]) || writeCTmain_mask_IntlizzieLet21_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTmain_mask_IntlizzieLet21_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                                 1'd0};
    else
      if (writeCTmain_mask_IntlizzieLet21_1_argbuf_rwb_r)
        writeCTmain_mask_IntlizzieLet21_1_argbuf_rwb_bufchan_d <= writeCTmain_mask_IntlizzieLet21_1_argbuf_rwb_d;
  Pointer_CTmain_mask_Int_t writeCTmain_mask_IntlizzieLet21_1_argbuf_rwb_bufchan_buf;
  assign writeCTmain_mask_IntlizzieLet21_1_argbuf_rwb_bufchan_r = (! writeCTmain_mask_IntlizzieLet21_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet4_1_1_argbuf_d = (writeCTmain_mask_IntlizzieLet21_1_argbuf_rwb_bufchan_buf[0] ? writeCTmain_mask_IntlizzieLet21_1_argbuf_rwb_bufchan_buf :
                                    writeCTmain_mask_IntlizzieLet21_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTmain_mask_IntlizzieLet21_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                   1'd0};
    else
      if ((lizzieLet4_1_1_argbuf_r && writeCTmain_mask_IntlizzieLet21_1_argbuf_rwb_bufchan_buf[0]))
        writeCTmain_mask_IntlizzieLet21_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                     1'd0};
      else if (((! lizzieLet4_1_1_argbuf_r) && (! writeCTmain_mask_IntlizzieLet21_1_argbuf_rwb_bufchan_buf[0])))
        writeCTmain_mask_IntlizzieLet21_1_argbuf_rwb_bufchan_buf <= writeCTmain_mask_IntlizzieLet21_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CTmain_mask_Int) : (writeCTmain_mask_IntlizzieLet32_1_argbuf,Pointer_CTmain_mask_Int) > (writeCTmain_mask_IntlizzieLet32_1_argbuf_rwb,Pointer_CTmain_mask_Int) */
  Pointer_CTmain_mask_Int_t writeCTmain_mask_IntlizzieLet32_1_argbuf_bufchan_d;
  logic writeCTmain_mask_IntlizzieLet32_1_argbuf_bufchan_r;
  assign writeCTmain_mask_IntlizzieLet32_1_argbuf_r = ((! writeCTmain_mask_IntlizzieLet32_1_argbuf_bufchan_d[0]) || writeCTmain_mask_IntlizzieLet32_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTmain_mask_IntlizzieLet32_1_argbuf_bufchan_d <= {16'd0,
                                                             1'd0};
    else
      if (writeCTmain_mask_IntlizzieLet32_1_argbuf_r)
        writeCTmain_mask_IntlizzieLet32_1_argbuf_bufchan_d <= writeCTmain_mask_IntlizzieLet32_1_argbuf_d;
  Pointer_CTmain_mask_Int_t writeCTmain_mask_IntlizzieLet32_1_argbuf_bufchan_buf;
  assign writeCTmain_mask_IntlizzieLet32_1_argbuf_bufchan_r = (! writeCTmain_mask_IntlizzieLet32_1_argbuf_bufchan_buf[0]);
  assign writeCTmain_mask_IntlizzieLet32_1_argbuf_rwb_d = (writeCTmain_mask_IntlizzieLet32_1_argbuf_bufchan_buf[0] ? writeCTmain_mask_IntlizzieLet32_1_argbuf_bufchan_buf :
                                                           writeCTmain_mask_IntlizzieLet32_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTmain_mask_IntlizzieLet32_1_argbuf_bufchan_buf <= {16'd0,
                                                               1'd0};
    else
      if ((writeCTmain_mask_IntlizzieLet32_1_argbuf_rwb_r && writeCTmain_mask_IntlizzieLet32_1_argbuf_bufchan_buf[0]))
        writeCTmain_mask_IntlizzieLet32_1_argbuf_bufchan_buf <= {16'd0,
                                                                 1'd0};
      else if (((! writeCTmain_mask_IntlizzieLet32_1_argbuf_rwb_r) && (! writeCTmain_mask_IntlizzieLet32_1_argbuf_bufchan_buf[0])))
        writeCTmain_mask_IntlizzieLet32_1_argbuf_bufchan_buf <= writeCTmain_mask_IntlizzieLet32_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CTmain_mask_Int) : (writeCTmain_mask_IntlizzieLet32_1_argbuf_rwb,Pointer_CTmain_mask_Int) > (sca2_2_1_argbuf,Pointer_CTmain_mask_Int) */
  Pointer_CTmain_mask_Int_t writeCTmain_mask_IntlizzieLet32_1_argbuf_rwb_bufchan_d;
  logic writeCTmain_mask_IntlizzieLet32_1_argbuf_rwb_bufchan_r;
  assign writeCTmain_mask_IntlizzieLet32_1_argbuf_rwb_r = ((! writeCTmain_mask_IntlizzieLet32_1_argbuf_rwb_bufchan_d[0]) || writeCTmain_mask_IntlizzieLet32_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTmain_mask_IntlizzieLet32_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                                 1'd0};
    else
      if (writeCTmain_mask_IntlizzieLet32_1_argbuf_rwb_r)
        writeCTmain_mask_IntlizzieLet32_1_argbuf_rwb_bufchan_d <= writeCTmain_mask_IntlizzieLet32_1_argbuf_rwb_d;
  Pointer_CTmain_mask_Int_t writeCTmain_mask_IntlizzieLet32_1_argbuf_rwb_bufchan_buf;
  assign writeCTmain_mask_IntlizzieLet32_1_argbuf_rwb_bufchan_r = (! writeCTmain_mask_IntlizzieLet32_1_argbuf_rwb_bufchan_buf[0]);
  assign sca2_2_1_argbuf_d = (writeCTmain_mask_IntlizzieLet32_1_argbuf_rwb_bufchan_buf[0] ? writeCTmain_mask_IntlizzieLet32_1_argbuf_rwb_bufchan_buf :
                              writeCTmain_mask_IntlizzieLet32_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTmain_mask_IntlizzieLet32_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                   1'd0};
    else
      if ((sca2_2_1_argbuf_r && writeCTmain_mask_IntlizzieLet32_1_argbuf_rwb_bufchan_buf[0]))
        writeCTmain_mask_IntlizzieLet32_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                     1'd0};
      else if (((! sca2_2_1_argbuf_r) && (! writeCTmain_mask_IntlizzieLet32_1_argbuf_rwb_bufchan_buf[0])))
        writeCTmain_mask_IntlizzieLet32_1_argbuf_rwb_bufchan_buf <= writeCTmain_mask_IntlizzieLet32_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CTmain_mask_Int) : (writeCTmain_mask_IntlizzieLet33_1_argbuf,Pointer_CTmain_mask_Int) > (writeCTmain_mask_IntlizzieLet33_1_argbuf_rwb,Pointer_CTmain_mask_Int) */
  Pointer_CTmain_mask_Int_t writeCTmain_mask_IntlizzieLet33_1_argbuf_bufchan_d;
  logic writeCTmain_mask_IntlizzieLet33_1_argbuf_bufchan_r;
  assign writeCTmain_mask_IntlizzieLet33_1_argbuf_r = ((! writeCTmain_mask_IntlizzieLet33_1_argbuf_bufchan_d[0]) || writeCTmain_mask_IntlizzieLet33_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTmain_mask_IntlizzieLet33_1_argbuf_bufchan_d <= {16'd0,
                                                             1'd0};
    else
      if (writeCTmain_mask_IntlizzieLet33_1_argbuf_r)
        writeCTmain_mask_IntlizzieLet33_1_argbuf_bufchan_d <= writeCTmain_mask_IntlizzieLet33_1_argbuf_d;
  Pointer_CTmain_mask_Int_t writeCTmain_mask_IntlizzieLet33_1_argbuf_bufchan_buf;
  assign writeCTmain_mask_IntlizzieLet33_1_argbuf_bufchan_r = (! writeCTmain_mask_IntlizzieLet33_1_argbuf_bufchan_buf[0]);
  assign writeCTmain_mask_IntlizzieLet33_1_argbuf_rwb_d = (writeCTmain_mask_IntlizzieLet33_1_argbuf_bufchan_buf[0] ? writeCTmain_mask_IntlizzieLet33_1_argbuf_bufchan_buf :
                                                           writeCTmain_mask_IntlizzieLet33_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTmain_mask_IntlizzieLet33_1_argbuf_bufchan_buf <= {16'd0,
                                                               1'd0};
    else
      if ((writeCTmain_mask_IntlizzieLet33_1_argbuf_rwb_r && writeCTmain_mask_IntlizzieLet33_1_argbuf_bufchan_buf[0]))
        writeCTmain_mask_IntlizzieLet33_1_argbuf_bufchan_buf <= {16'd0,
                                                                 1'd0};
      else if (((! writeCTmain_mask_IntlizzieLet33_1_argbuf_rwb_r) && (! writeCTmain_mask_IntlizzieLet33_1_argbuf_bufchan_buf[0])))
        writeCTmain_mask_IntlizzieLet33_1_argbuf_bufchan_buf <= writeCTmain_mask_IntlizzieLet33_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CTmain_mask_Int) : (writeCTmain_mask_IntlizzieLet33_1_argbuf_rwb,Pointer_CTmain_mask_Int) > (sca1_2_1_argbuf,Pointer_CTmain_mask_Int) */
  Pointer_CTmain_mask_Int_t writeCTmain_mask_IntlizzieLet33_1_argbuf_rwb_bufchan_d;
  logic writeCTmain_mask_IntlizzieLet33_1_argbuf_rwb_bufchan_r;
  assign writeCTmain_mask_IntlizzieLet33_1_argbuf_rwb_r = ((! writeCTmain_mask_IntlizzieLet33_1_argbuf_rwb_bufchan_d[0]) || writeCTmain_mask_IntlizzieLet33_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTmain_mask_IntlizzieLet33_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                                 1'd0};
    else
      if (writeCTmain_mask_IntlizzieLet33_1_argbuf_rwb_r)
        writeCTmain_mask_IntlizzieLet33_1_argbuf_rwb_bufchan_d <= writeCTmain_mask_IntlizzieLet33_1_argbuf_rwb_d;
  Pointer_CTmain_mask_Int_t writeCTmain_mask_IntlizzieLet33_1_argbuf_rwb_bufchan_buf;
  assign writeCTmain_mask_IntlizzieLet33_1_argbuf_rwb_bufchan_r = (! writeCTmain_mask_IntlizzieLet33_1_argbuf_rwb_bufchan_buf[0]);
  assign sca1_2_1_argbuf_d = (writeCTmain_mask_IntlizzieLet33_1_argbuf_rwb_bufchan_buf[0] ? writeCTmain_mask_IntlizzieLet33_1_argbuf_rwb_bufchan_buf :
                              writeCTmain_mask_IntlizzieLet33_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTmain_mask_IntlizzieLet33_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                   1'd0};
    else
      if ((sca1_2_1_argbuf_r && writeCTmain_mask_IntlizzieLet33_1_argbuf_rwb_bufchan_buf[0]))
        writeCTmain_mask_IntlizzieLet33_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                     1'd0};
      else if (((! sca1_2_1_argbuf_r) && (! writeCTmain_mask_IntlizzieLet33_1_argbuf_rwb_bufchan_buf[0])))
        writeCTmain_mask_IntlizzieLet33_1_argbuf_rwb_bufchan_buf <= writeCTmain_mask_IntlizzieLet33_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CTmain_mask_Int) : (writeCTmain_mask_IntlizzieLet34_1_argbuf,Pointer_CTmain_mask_Int) > (writeCTmain_mask_IntlizzieLet34_1_argbuf_rwb,Pointer_CTmain_mask_Int) */
  Pointer_CTmain_mask_Int_t writeCTmain_mask_IntlizzieLet34_1_argbuf_bufchan_d;
  logic writeCTmain_mask_IntlizzieLet34_1_argbuf_bufchan_r;
  assign writeCTmain_mask_IntlizzieLet34_1_argbuf_r = ((! writeCTmain_mask_IntlizzieLet34_1_argbuf_bufchan_d[0]) || writeCTmain_mask_IntlizzieLet34_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTmain_mask_IntlizzieLet34_1_argbuf_bufchan_d <= {16'd0,
                                                             1'd0};
    else
      if (writeCTmain_mask_IntlizzieLet34_1_argbuf_r)
        writeCTmain_mask_IntlizzieLet34_1_argbuf_bufchan_d <= writeCTmain_mask_IntlizzieLet34_1_argbuf_d;
  Pointer_CTmain_mask_Int_t writeCTmain_mask_IntlizzieLet34_1_argbuf_bufchan_buf;
  assign writeCTmain_mask_IntlizzieLet34_1_argbuf_bufchan_r = (! writeCTmain_mask_IntlizzieLet34_1_argbuf_bufchan_buf[0]);
  assign writeCTmain_mask_IntlizzieLet34_1_argbuf_rwb_d = (writeCTmain_mask_IntlizzieLet34_1_argbuf_bufchan_buf[0] ? writeCTmain_mask_IntlizzieLet34_1_argbuf_bufchan_buf :
                                                           writeCTmain_mask_IntlizzieLet34_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTmain_mask_IntlizzieLet34_1_argbuf_bufchan_buf <= {16'd0,
                                                               1'd0};
    else
      if ((writeCTmain_mask_IntlizzieLet34_1_argbuf_rwb_r && writeCTmain_mask_IntlizzieLet34_1_argbuf_bufchan_buf[0]))
        writeCTmain_mask_IntlizzieLet34_1_argbuf_bufchan_buf <= {16'd0,
                                                                 1'd0};
      else if (((! writeCTmain_mask_IntlizzieLet34_1_argbuf_rwb_r) && (! writeCTmain_mask_IntlizzieLet34_1_argbuf_bufchan_buf[0])))
        writeCTmain_mask_IntlizzieLet34_1_argbuf_bufchan_buf <= writeCTmain_mask_IntlizzieLet34_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CTmain_mask_Int) : (writeCTmain_mask_IntlizzieLet34_1_argbuf_rwb,Pointer_CTmain_mask_Int) > (sca0_2_1_argbuf,Pointer_CTmain_mask_Int) */
  Pointer_CTmain_mask_Int_t writeCTmain_mask_IntlizzieLet34_1_argbuf_rwb_bufchan_d;
  logic writeCTmain_mask_IntlizzieLet34_1_argbuf_rwb_bufchan_r;
  assign writeCTmain_mask_IntlizzieLet34_1_argbuf_rwb_r = ((! writeCTmain_mask_IntlizzieLet34_1_argbuf_rwb_bufchan_d[0]) || writeCTmain_mask_IntlizzieLet34_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTmain_mask_IntlizzieLet34_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                                 1'd0};
    else
      if (writeCTmain_mask_IntlizzieLet34_1_argbuf_rwb_r)
        writeCTmain_mask_IntlizzieLet34_1_argbuf_rwb_bufchan_d <= writeCTmain_mask_IntlizzieLet34_1_argbuf_rwb_d;
  Pointer_CTmain_mask_Int_t writeCTmain_mask_IntlizzieLet34_1_argbuf_rwb_bufchan_buf;
  assign writeCTmain_mask_IntlizzieLet34_1_argbuf_rwb_bufchan_r = (! writeCTmain_mask_IntlizzieLet34_1_argbuf_rwb_bufchan_buf[0]);
  assign sca0_2_1_argbuf_d = (writeCTmain_mask_IntlizzieLet34_1_argbuf_rwb_bufchan_buf[0] ? writeCTmain_mask_IntlizzieLet34_1_argbuf_rwb_bufchan_buf :
                              writeCTmain_mask_IntlizzieLet34_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTmain_mask_IntlizzieLet34_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                   1'd0};
    else
      if ((sca0_2_1_argbuf_r && writeCTmain_mask_IntlizzieLet34_1_argbuf_rwb_bufchan_buf[0]))
        writeCTmain_mask_IntlizzieLet34_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                     1'd0};
      else if (((! sca0_2_1_argbuf_r) && (! writeCTmain_mask_IntlizzieLet34_1_argbuf_rwb_bufchan_buf[0])))
        writeCTmain_mask_IntlizzieLet34_1_argbuf_rwb_bufchan_buf <= writeCTmain_mask_IntlizzieLet34_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet10_1_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet10_1_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet10_1_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet10_1_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet10_1_1_argbuf_r = ((! writeQTree_IntlizzieLet10_1_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet10_1_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet10_1_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet10_1_1_argbuf_r)
        writeQTree_IntlizzieLet10_1_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet10_1_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet10_1_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet10_1_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet10_1_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet10_1_1_argbuf_rwb_d = (writeQTree_IntlizzieLet10_1_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet10_1_1_argbuf_bufchan_buf :
                                                       writeQTree_IntlizzieLet10_1_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet10_1_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet10_1_1_argbuf_rwb_r && writeQTree_IntlizzieLet10_1_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet10_1_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet10_1_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet10_1_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet10_1_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet10_1_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet10_1_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet12_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet10_1_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet10_1_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet10_1_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet10_1_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet10_1_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet10_1_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                             1'd0};
    else
      if (writeQTree_IntlizzieLet10_1_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet10_1_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet10_1_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet10_1_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet10_1_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet10_1_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet12_1_argbuf_d = (writeQTree_IntlizzieLet10_1_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet10_1_1_argbuf_rwb_bufchan_buf :
                                   writeQTree_IntlizzieLet10_1_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet10_1_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
    else
      if ((lizzieLet12_1_argbuf_r && writeQTree_IntlizzieLet10_1_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet10_1_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                 1'd0};
      else if (((! lizzieLet12_1_argbuf_r) && (! writeQTree_IntlizzieLet10_1_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet10_1_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet10_1_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet11_1_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet11_1_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet11_1_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet11_1_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet11_1_1_argbuf_r = ((! writeQTree_IntlizzieLet11_1_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet11_1_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet11_1_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet11_1_1_argbuf_r)
        writeQTree_IntlizzieLet11_1_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet11_1_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet11_1_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet11_1_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet11_1_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet11_1_1_argbuf_rwb_d = (writeQTree_IntlizzieLet11_1_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet11_1_1_argbuf_bufchan_buf :
                                                       writeQTree_IntlizzieLet11_1_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet11_1_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet11_1_1_argbuf_rwb_r && writeQTree_IntlizzieLet11_1_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet11_1_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet11_1_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet11_1_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet11_1_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet11_1_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet11_1_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet13_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet11_1_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet11_1_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet11_1_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet11_1_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet11_1_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet11_1_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                             1'd0};
    else
      if (writeQTree_IntlizzieLet11_1_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet11_1_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet11_1_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet11_1_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet11_1_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet11_1_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet13_1_argbuf_d = (writeQTree_IntlizzieLet11_1_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet11_1_1_argbuf_rwb_bufchan_buf :
                                   writeQTree_IntlizzieLet11_1_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet11_1_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
    else
      if ((lizzieLet13_1_argbuf_r && writeQTree_IntlizzieLet11_1_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet11_1_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                 1'd0};
      else if (((! lizzieLet13_1_argbuf_r) && (! writeQTree_IntlizzieLet11_1_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet11_1_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet11_1_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet15_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet15_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet15_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet15_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet15_1_argbuf_r = ((! writeQTree_IntlizzieLet15_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet15_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet15_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet15_1_argbuf_r)
        writeQTree_IntlizzieLet15_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet15_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet15_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet15_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet15_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet15_1_argbuf_rwb_d = (writeQTree_IntlizzieLet15_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet15_1_argbuf_bufchan_buf :
                                                     writeQTree_IntlizzieLet15_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet15_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet15_1_argbuf_rwb_r && writeQTree_IntlizzieLet15_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet15_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet15_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet15_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet15_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet15_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet15_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet0_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet15_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet15_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet15_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet15_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet15_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet15_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet15_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet15_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet15_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet15_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet15_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet15_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet0_1_1_argbuf_d = (writeQTree_IntlizzieLet15_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet15_1_argbuf_rwb_bufchan_buf :
                                    writeQTree_IntlizzieLet15_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet15_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((lizzieLet0_1_1_argbuf_r && writeQTree_IntlizzieLet15_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet15_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! lizzieLet0_1_1_argbuf_r) && (! writeQTree_IntlizzieLet15_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet15_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet15_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet17_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet17_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet17_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet17_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet17_1_argbuf_r = ((! writeQTree_IntlizzieLet17_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet17_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet17_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet17_1_argbuf_r)
        writeQTree_IntlizzieLet17_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet17_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet17_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet17_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet17_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet17_1_argbuf_rwb_d = (writeQTree_IntlizzieLet17_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet17_1_argbuf_bufchan_buf :
                                                     writeQTree_IntlizzieLet17_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet17_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet17_1_argbuf_rwb_r && writeQTree_IntlizzieLet17_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet17_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet17_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet17_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet17_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet17_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet17_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet1_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet17_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet17_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet17_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet17_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet17_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet17_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet17_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet17_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet17_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet17_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet17_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet17_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet1_1_1_argbuf_d = (writeQTree_IntlizzieLet17_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet17_1_argbuf_rwb_bufchan_buf :
                                    writeQTree_IntlizzieLet17_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet17_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((lizzieLet1_1_1_argbuf_r && writeQTree_IntlizzieLet17_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet17_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! lizzieLet1_1_1_argbuf_r) && (! writeQTree_IntlizzieLet17_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet17_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet17_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet18_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet18_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet18_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet18_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet18_1_argbuf_r = ((! writeQTree_IntlizzieLet18_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet18_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet18_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet18_1_argbuf_r)
        writeQTree_IntlizzieLet18_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet18_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet18_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet18_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet18_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet18_1_argbuf_rwb_d = (writeQTree_IntlizzieLet18_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet18_1_argbuf_bufchan_buf :
                                                     writeQTree_IntlizzieLet18_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet18_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet18_1_argbuf_rwb_r && writeQTree_IntlizzieLet18_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet18_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet18_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet18_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet18_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet18_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet18_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet2_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet18_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet18_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet18_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet18_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet18_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet18_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet18_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet18_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet18_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet18_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet18_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet18_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet2_1_1_argbuf_d = (writeQTree_IntlizzieLet18_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet18_1_argbuf_rwb_bufchan_buf :
                                    writeQTree_IntlizzieLet18_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet18_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((lizzieLet2_1_1_argbuf_r && writeQTree_IntlizzieLet18_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet18_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! lizzieLet2_1_1_argbuf_r) && (! writeQTree_IntlizzieLet18_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet18_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet18_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet20_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet20_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet20_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet20_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet20_1_argbuf_r = ((! writeQTree_IntlizzieLet20_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet20_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet20_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet20_1_argbuf_r)
        writeQTree_IntlizzieLet20_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet20_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet20_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet20_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet20_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet20_1_argbuf_rwb_d = (writeQTree_IntlizzieLet20_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet20_1_argbuf_bufchan_buf :
                                                     writeQTree_IntlizzieLet20_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet20_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet20_1_argbuf_rwb_r && writeQTree_IntlizzieLet20_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet20_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet20_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet20_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet20_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet20_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet20_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet3_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet20_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet20_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet20_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet20_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet20_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet20_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet20_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet20_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet20_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet20_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet20_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet20_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet3_1_1_argbuf_d = (writeQTree_IntlizzieLet20_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet20_1_argbuf_rwb_bufchan_buf :
                                    writeQTree_IntlizzieLet20_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet20_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((lizzieLet3_1_1_argbuf_r && writeQTree_IntlizzieLet20_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet20_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! lizzieLet3_1_1_argbuf_r) && (! writeQTree_IntlizzieLet20_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet20_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet20_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet26_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet26_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet26_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet26_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet26_1_argbuf_r = ((! writeQTree_IntlizzieLet26_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet26_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet26_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet26_1_argbuf_r)
        writeQTree_IntlizzieLet26_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet26_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet26_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet26_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet26_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet26_1_argbuf_rwb_d = (writeQTree_IntlizzieLet26_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet26_1_argbuf_bufchan_buf :
                                                     writeQTree_IntlizzieLet26_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet26_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet26_1_argbuf_rwb_r && writeQTree_IntlizzieLet26_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet26_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet26_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet26_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet26_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet26_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet26_1_argbuf_rwb,Pointer_QTree_Int) > (contRet_0_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet26_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet26_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet26_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet26_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet26_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet26_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet26_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet26_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet26_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet26_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet26_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet26_1_argbuf_rwb_bufchan_buf[0]);
  assign contRet_0_1_argbuf_d = (writeQTree_IntlizzieLet26_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet26_1_argbuf_rwb_bufchan_buf :
                                 writeQTree_IntlizzieLet26_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet26_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((contRet_0_1_argbuf_r && writeQTree_IntlizzieLet26_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet26_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! contRet_0_1_argbuf_r) && (! writeQTree_IntlizzieLet26_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet26_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet26_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet35_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet35_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet35_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet35_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet35_1_argbuf_r = ((! writeQTree_IntlizzieLet35_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet35_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet35_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet35_1_argbuf_r)
        writeQTree_IntlizzieLet35_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet35_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet35_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet35_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet35_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet35_1_argbuf_rwb_d = (writeQTree_IntlizzieLet35_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet35_1_argbuf_bufchan_buf :
                                                     writeQTree_IntlizzieLet35_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet35_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet35_1_argbuf_rwb_r && writeQTree_IntlizzieLet35_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet35_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet35_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet35_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet35_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet35_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet35_1_argbuf_rwb,Pointer_QTree_Int) > (contRet_0_2_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet35_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet35_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet35_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet35_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet35_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet35_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet35_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet35_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet35_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet35_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet35_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet35_1_argbuf_rwb_bufchan_buf[0]);
  assign contRet_0_2_1_argbuf_d = (writeQTree_IntlizzieLet35_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet35_1_argbuf_rwb_bufchan_buf :
                                   writeQTree_IntlizzieLet35_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet35_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((contRet_0_2_1_argbuf_r && writeQTree_IntlizzieLet35_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet35_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! contRet_0_2_1_argbuf_r) && (! writeQTree_IntlizzieLet35_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet35_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet35_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet4_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet4_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet4_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet4_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet4_1_argbuf_r = ((! writeQTree_IntlizzieLet4_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet4_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet4_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet4_1_argbuf_r)
        writeQTree_IntlizzieLet4_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet4_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet4_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet4_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet4_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet4_1_argbuf_rwb_d = (writeQTree_IntlizzieLet4_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet4_1_argbuf_bufchan_buf :
                                                    writeQTree_IntlizzieLet4_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet4_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet4_1_argbuf_rwb_r && writeQTree_IntlizzieLet4_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet4_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet4_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet4_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet4_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet4_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet4_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet8_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet4_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet4_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet4_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet4_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet4_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet4_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet4_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet4_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet4_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet4_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet4_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet4_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet8_1_argbuf_d = (writeQTree_IntlizzieLet4_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet4_1_argbuf_rwb_bufchan_buf :
                                  writeQTree_IntlizzieLet4_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet4_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet8_1_argbuf_r && writeQTree_IntlizzieLet4_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet4_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet8_1_argbuf_r) && (! writeQTree_IntlizzieLet4_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet4_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet4_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet5_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet5_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet5_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet5_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet5_1_argbuf_r = ((! writeQTree_IntlizzieLet5_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet5_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet5_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet5_1_argbuf_r)
        writeQTree_IntlizzieLet5_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet5_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet5_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet5_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet5_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet5_1_argbuf_rwb_d = (writeQTree_IntlizzieLet5_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet5_1_argbuf_bufchan_buf :
                                                    writeQTree_IntlizzieLet5_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet5_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet5_1_argbuf_rwb_r && writeQTree_IntlizzieLet5_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet5_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet5_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet5_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet5_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet5_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet5_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet9_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet5_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet5_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet5_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet5_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet5_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet5_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet5_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet5_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet5_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet5_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet5_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet5_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet9_1_argbuf_d = (writeQTree_IntlizzieLet5_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet5_1_argbuf_rwb_bufchan_buf :
                                  writeQTree_IntlizzieLet5_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet5_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet9_1_argbuf_r && writeQTree_IntlizzieLet5_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet5_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet9_1_argbuf_r) && (! writeQTree_IntlizzieLet5_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet5_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet5_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet6_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet6_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet6_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet6_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet6_1_argbuf_r = ((! writeQTree_IntlizzieLet6_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet6_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet6_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet6_1_argbuf_r)
        writeQTree_IntlizzieLet6_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet6_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet6_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet6_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet6_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet6_1_argbuf_rwb_d = (writeQTree_IntlizzieLet6_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet6_1_argbuf_bufchan_buf :
                                                    writeQTree_IntlizzieLet6_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet6_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet6_1_argbuf_rwb_r && writeQTree_IntlizzieLet6_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet6_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet6_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet6_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet6_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet6_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet6_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet10_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet6_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet6_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet6_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet6_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet6_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet6_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet6_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet6_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet6_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet6_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet6_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet6_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet10_1_argbuf_d = (writeQTree_IntlizzieLet6_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet6_1_argbuf_rwb_bufchan_buf :
                                   writeQTree_IntlizzieLet6_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet6_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet10_1_argbuf_r && writeQTree_IntlizzieLet6_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet6_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet10_1_argbuf_r) && (! writeQTree_IntlizzieLet6_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet6_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet6_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet8_1_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet8_1_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet8_1_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet8_1_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet8_1_1_argbuf_r = ((! writeQTree_IntlizzieLet8_1_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet8_1_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet8_1_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet8_1_1_argbuf_r)
        writeQTree_IntlizzieLet8_1_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet8_1_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet8_1_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet8_1_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet8_1_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet8_1_1_argbuf_rwb_d = (writeQTree_IntlizzieLet8_1_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet8_1_1_argbuf_bufchan_buf :
                                                      writeQTree_IntlizzieLet8_1_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet8_1_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet8_1_1_argbuf_rwb_r && writeQTree_IntlizzieLet8_1_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet8_1_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet8_1_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet8_1_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet8_1_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet8_1_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet8_1_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet11_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet8_1_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet8_1_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet8_1_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet8_1_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet8_1_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet8_1_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet8_1_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet8_1_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet8_1_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet8_1_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet8_1_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet8_1_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet11_1_argbuf_d = (writeQTree_IntlizzieLet8_1_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet8_1_1_argbuf_rwb_bufchan_buf :
                                   writeQTree_IntlizzieLet8_1_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet8_1_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                              1'd0};
    else
      if ((lizzieLet11_1_argbuf_r && writeQTree_IntlizzieLet8_1_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet8_1_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
      else if (((! lizzieLet11_1_argbuf_r) && (! writeQTree_IntlizzieLet8_1_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet8_1_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet8_1_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty MyDTInt_Int_Int) : (wsie_2_2,MyDTInt_Int_Int) > (wsie_2_2_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t wsie_2_2_bufchan_d;
  logic wsie_2_2_bufchan_r;
  assign wsie_2_2_r = ((! wsie_2_2_bufchan_d[0]) || wsie_2_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) wsie_2_2_bufchan_d <= 1'd0;
    else if (wsie_2_2_r) wsie_2_2_bufchan_d <= wsie_2_2_d;
  MyDTInt_Int_Int_t wsie_2_2_bufchan_buf;
  assign wsie_2_2_bufchan_r = (! wsie_2_2_bufchan_buf[0]);
  assign wsie_2_2_argbuf_d = (wsie_2_2_bufchan_buf[0] ? wsie_2_2_bufchan_buf :
                              wsie_2_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) wsie_2_2_bufchan_buf <= 1'd0;
    else
      if ((wsie_2_2_argbuf_r && wsie_2_2_bufchan_buf[0]))
        wsie_2_2_bufchan_buf <= 1'd0;
      else if (((! wsie_2_2_argbuf_r) && (! wsie_2_2_bufchan_buf[0])))
        wsie_2_2_bufchan_buf <= wsie_2_2_bufchan_d;
  
  /* fork (Ty MyDTInt_Int_Int) : (wsie_2_destruct,MyDTInt_Int_Int) > [(wsie_2_1,MyDTInt_Int_Int),
                                                                 (wsie_2_2,MyDTInt_Int_Int)] */
  logic [1:0] wsie_2_destruct_emitted;
  logic [1:0] wsie_2_destruct_done;
  assign wsie_2_1_d = (wsie_2_destruct_d[0] && (! wsie_2_destruct_emitted[0]));
  assign wsie_2_2_d = (wsie_2_destruct_d[0] && (! wsie_2_destruct_emitted[1]));
  assign wsie_2_destruct_done = (wsie_2_destruct_emitted | ({wsie_2_2_d[0],
                                                             wsie_2_1_d[0]} & {wsie_2_2_r,
                                                                               wsie_2_1_r}));
  assign wsie_2_destruct_r = (& wsie_2_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) wsie_2_destruct_emitted <= 2'd0;
    else
      wsie_2_destruct_emitted <= (wsie_2_destruct_r ? 2'd0 :
                                  wsie_2_destruct_done);
  
  /* buf (Ty MyDTInt_Int_Int) : (wsie_3_2,MyDTInt_Int_Int) > (wsie_3_2_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t wsie_3_2_bufchan_d;
  logic wsie_3_2_bufchan_r;
  assign wsie_3_2_r = ((! wsie_3_2_bufchan_d[0]) || wsie_3_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) wsie_3_2_bufchan_d <= 1'd0;
    else if (wsie_3_2_r) wsie_3_2_bufchan_d <= wsie_3_2_d;
  MyDTInt_Int_Int_t wsie_3_2_bufchan_buf;
  assign wsie_3_2_bufchan_r = (! wsie_3_2_bufchan_buf[0]);
  assign wsie_3_2_argbuf_d = (wsie_3_2_bufchan_buf[0] ? wsie_3_2_bufchan_buf :
                              wsie_3_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) wsie_3_2_bufchan_buf <= 1'd0;
    else
      if ((wsie_3_2_argbuf_r && wsie_3_2_bufchan_buf[0]))
        wsie_3_2_bufchan_buf <= 1'd0;
      else if (((! wsie_3_2_argbuf_r) && (! wsie_3_2_bufchan_buf[0])))
        wsie_3_2_bufchan_buf <= wsie_3_2_bufchan_d;
  
  /* fork (Ty MyDTInt_Int_Int) : (wsie_3_destruct,MyDTInt_Int_Int) > [(wsie_3_1,MyDTInt_Int_Int),
                                                                 (wsie_3_2,MyDTInt_Int_Int)] */
  logic [1:0] wsie_3_destruct_emitted;
  logic [1:0] wsie_3_destruct_done;
  assign wsie_3_1_d = (wsie_3_destruct_d[0] && (! wsie_3_destruct_emitted[0]));
  assign wsie_3_2_d = (wsie_3_destruct_d[0] && (! wsie_3_destruct_emitted[1]));
  assign wsie_3_destruct_done = (wsie_3_destruct_emitted | ({wsie_3_2_d[0],
                                                             wsie_3_1_d[0]} & {wsie_3_2_r,
                                                                               wsie_3_1_r}));
  assign wsie_3_destruct_r = (& wsie_3_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) wsie_3_destruct_emitted <= 2'd0;
    else
      wsie_3_destruct_emitted <= (wsie_3_destruct_r ? 2'd0 :
                                  wsie_3_destruct_done);
  
  /* buf (Ty MyDTInt_Int_Int) : (wsie_4_destruct,MyDTInt_Int_Int) > (wsie_4_1_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t wsie_4_destruct_bufchan_d;
  logic wsie_4_destruct_bufchan_r;
  assign wsie_4_destruct_r = ((! wsie_4_destruct_bufchan_d[0]) || wsie_4_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) wsie_4_destruct_bufchan_d <= 1'd0;
    else
      if (wsie_4_destruct_r)
        wsie_4_destruct_bufchan_d <= wsie_4_destruct_d;
  MyDTInt_Int_Int_t wsie_4_destruct_bufchan_buf;
  assign wsie_4_destruct_bufchan_r = (! wsie_4_destruct_bufchan_buf[0]);
  assign wsie_4_1_argbuf_d = (wsie_4_destruct_bufchan_buf[0] ? wsie_4_destruct_bufchan_buf :
                              wsie_4_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) wsie_4_destruct_bufchan_buf <= 1'd0;
    else
      if ((wsie_4_1_argbuf_r && wsie_4_destruct_bufchan_buf[0]))
        wsie_4_destruct_bufchan_buf <= 1'd0;
      else if (((! wsie_4_1_argbuf_r) && (! wsie_4_destruct_bufchan_buf[0])))
        wsie_4_destruct_bufchan_buf <= wsie_4_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (wsij_1_goMux_mux,Pointer_QTree_Int) > (wsij_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t wsij_1_goMux_mux_bufchan_d;
  logic wsij_1_goMux_mux_bufchan_r;
  assign wsij_1_goMux_mux_r = ((! wsij_1_goMux_mux_bufchan_d[0]) || wsij_1_goMux_mux_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) wsij_1_goMux_mux_bufchan_d <= {16'd0, 1'd0};
    else
      if (wsij_1_goMux_mux_r)
        wsij_1_goMux_mux_bufchan_d <= wsij_1_goMux_mux_d;
  Pointer_QTree_Int_t wsij_1_goMux_mux_bufchan_buf;
  assign wsij_1_goMux_mux_bufchan_r = (! wsij_1_goMux_mux_bufchan_buf[0]);
  assign wsij_1_1_argbuf_d = (wsij_1_goMux_mux_bufchan_buf[0] ? wsij_1_goMux_mux_bufchan_buf :
                              wsij_1_goMux_mux_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) wsij_1_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((wsij_1_1_argbuf_r && wsij_1_goMux_mux_bufchan_buf[0]))
        wsij_1_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
      else if (((! wsij_1_1_argbuf_r) && (! wsij_1_goMux_mux_bufchan_buf[0])))
        wsij_1_goMux_mux_bufchan_buf <= wsij_1_goMux_mux_bufchan_d;
  
  /* buf (Ty CT$wnnz_Int) : (wwsim_2_1lizzieLet27_4Lcall_$wnnz_Int2_1sc_0_8_1q4a8F_2_1Lcall_$wnnz_Int1,CT$wnnz_Int) > (lizzieLet29_1_argbuf,CT$wnnz_Int) */
  CT$wnnz_Int_t wwsim_2_1lizzieLet27_4Lcall_$wnnz_Int2_1sc_0_8_1q4a8F_2_1Lcall_$wnnz_Int1_bufchan_d;
  logic wwsim_2_1lizzieLet27_4Lcall_$wnnz_Int2_1sc_0_8_1q4a8F_2_1Lcall_$wnnz_Int1_bufchan_r;
  assign wwsim_2_1lizzieLet27_4Lcall_$wnnz_Int2_1sc_0_8_1q4a8F_2_1Lcall_$wnnz_Int1_r = ((! wwsim_2_1lizzieLet27_4Lcall_$wnnz_Int2_1sc_0_8_1q4a8F_2_1Lcall_$wnnz_Int1_bufchan_d[0]) || wwsim_2_1lizzieLet27_4Lcall_$wnnz_Int2_1sc_0_8_1q4a8F_2_1Lcall_$wnnz_Int1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      wwsim_2_1lizzieLet27_4Lcall_$wnnz_Int2_1sc_0_8_1q4a8F_2_1Lcall_$wnnz_Int1_bufchan_d <= {115'd0,
                                                                                              1'd0};
    else
      if (wwsim_2_1lizzieLet27_4Lcall_$wnnz_Int2_1sc_0_8_1q4a8F_2_1Lcall_$wnnz_Int1_r)
        wwsim_2_1lizzieLet27_4Lcall_$wnnz_Int2_1sc_0_8_1q4a8F_2_1Lcall_$wnnz_Int1_bufchan_d <= wwsim_2_1lizzieLet27_4Lcall_$wnnz_Int2_1sc_0_8_1q4a8F_2_1Lcall_$wnnz_Int1_d;
  CT$wnnz_Int_t wwsim_2_1lizzieLet27_4Lcall_$wnnz_Int2_1sc_0_8_1q4a8F_2_1Lcall_$wnnz_Int1_bufchan_buf;
  assign wwsim_2_1lizzieLet27_4Lcall_$wnnz_Int2_1sc_0_8_1q4a8F_2_1Lcall_$wnnz_Int1_bufchan_r = (! wwsim_2_1lizzieLet27_4Lcall_$wnnz_Int2_1sc_0_8_1q4a8F_2_1Lcall_$wnnz_Int1_bufchan_buf[0]);
  assign lizzieLet29_1_argbuf_d = (wwsim_2_1lizzieLet27_4Lcall_$wnnz_Int2_1sc_0_8_1q4a8F_2_1Lcall_$wnnz_Int1_bufchan_buf[0] ? wwsim_2_1lizzieLet27_4Lcall_$wnnz_Int2_1sc_0_8_1q4a8F_2_1Lcall_$wnnz_Int1_bufchan_buf :
                                   wwsim_2_1lizzieLet27_4Lcall_$wnnz_Int2_1sc_0_8_1q4a8F_2_1Lcall_$wnnz_Int1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      wwsim_2_1lizzieLet27_4Lcall_$wnnz_Int2_1sc_0_8_1q4a8F_2_1Lcall_$wnnz_Int1_bufchan_buf <= {115'd0,
                                                                                                1'd0};
    else
      if ((lizzieLet29_1_argbuf_r && wwsim_2_1lizzieLet27_4Lcall_$wnnz_Int2_1sc_0_8_1q4a8F_2_1Lcall_$wnnz_Int1_bufchan_buf[0]))
        wwsim_2_1lizzieLet27_4Lcall_$wnnz_Int2_1sc_0_8_1q4a8F_2_1Lcall_$wnnz_Int1_bufchan_buf <= {115'd0,
                                                                                                  1'd0};
      else if (((! lizzieLet29_1_argbuf_r) && (! wwsim_2_1lizzieLet27_4Lcall_$wnnz_Int2_1sc_0_8_1q4a8F_2_1Lcall_$wnnz_Int1_bufchan_buf[0])))
        wwsim_2_1lizzieLet27_4Lcall_$wnnz_Int2_1sc_0_8_1q4a8F_2_1Lcall_$wnnz_Int1_bufchan_buf <= wwsim_2_1lizzieLet27_4Lcall_$wnnz_Int2_1sc_0_8_1q4a8F_2_1Lcall_$wnnz_Int1_bufchan_d;
  
  /* dcon (Ty CT$wnnz_Int,
      Dcon Lcall_$wnnz_Int1) : [(wwsim_2_destruct,Int#),
                                (lizzieLet27_4Lcall_$wnnz_Int2,Int#),
                                (sc_0_8_destruct,Pointer_CT$wnnz_Int),
                                (q4a8F_2_destruct,Pointer_QTree_Int)] > (wwsim_2_1lizzieLet27_4Lcall_$wnnz_Int2_1sc_0_8_1q4a8F_2_1Lcall_$wnnz_Int1,CT$wnnz_Int) */
  assign wwsim_2_1lizzieLet27_4Lcall_$wnnz_Int2_1sc_0_8_1q4a8F_2_1Lcall_$wnnz_Int1_d = Lcall_$wnnz_Int1_dc((& {wwsim_2_destruct_d[0],
                                                                                                               lizzieLet27_4Lcall_$wnnz_Int2_d[0],
                                                                                                               sc_0_8_destruct_d[0],
                                                                                                               q4a8F_2_destruct_d[0]}), wwsim_2_destruct_d, lizzieLet27_4Lcall_$wnnz_Int2_d, sc_0_8_destruct_d, q4a8F_2_destruct_d);
  assign {wwsim_2_destruct_r,
          lizzieLet27_4Lcall_$wnnz_Int2_r,
          sc_0_8_destruct_r,
          q4a8F_2_destruct_r} = {4 {(wwsim_2_1lizzieLet27_4Lcall_$wnnz_Int2_1sc_0_8_1q4a8F_2_1Lcall_$wnnz_Int1_r && wwsim_2_1lizzieLet27_4Lcall_$wnnz_Int2_1sc_0_8_1q4a8F_2_1Lcall_$wnnz_Int1_d[0])}};
  
  /* buf (Ty CT$wnnz_Int) : (wwsim_3_1ww1XiS_1_1lizzieLet27_4Lcall_$wnnz_Int1_1sc_0_9_1Lcall_$wnnz_Int0,CT$wnnz_Int) > (lizzieLet30_1_argbuf,CT$wnnz_Int) */
  CT$wnnz_Int_t wwsim_3_1ww1XiS_1_1lizzieLet27_4Lcall_$wnnz_Int1_1sc_0_9_1Lcall_$wnnz_Int0_bufchan_d;
  logic wwsim_3_1ww1XiS_1_1lizzieLet27_4Lcall_$wnnz_Int1_1sc_0_9_1Lcall_$wnnz_Int0_bufchan_r;
  assign wwsim_3_1ww1XiS_1_1lizzieLet27_4Lcall_$wnnz_Int1_1sc_0_9_1Lcall_$wnnz_Int0_r = ((! wwsim_3_1ww1XiS_1_1lizzieLet27_4Lcall_$wnnz_Int1_1sc_0_9_1Lcall_$wnnz_Int0_bufchan_d[0]) || wwsim_3_1ww1XiS_1_1lizzieLet27_4Lcall_$wnnz_Int1_1sc_0_9_1Lcall_$wnnz_Int0_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      wwsim_3_1ww1XiS_1_1lizzieLet27_4Lcall_$wnnz_Int1_1sc_0_9_1Lcall_$wnnz_Int0_bufchan_d <= {115'd0,
                                                                                               1'd0};
    else
      if (wwsim_3_1ww1XiS_1_1lizzieLet27_4Lcall_$wnnz_Int1_1sc_0_9_1Lcall_$wnnz_Int0_r)
        wwsim_3_1ww1XiS_1_1lizzieLet27_4Lcall_$wnnz_Int1_1sc_0_9_1Lcall_$wnnz_Int0_bufchan_d <= wwsim_3_1ww1XiS_1_1lizzieLet27_4Lcall_$wnnz_Int1_1sc_0_9_1Lcall_$wnnz_Int0_d;
  CT$wnnz_Int_t wwsim_3_1ww1XiS_1_1lizzieLet27_4Lcall_$wnnz_Int1_1sc_0_9_1Lcall_$wnnz_Int0_bufchan_buf;
  assign wwsim_3_1ww1XiS_1_1lizzieLet27_4Lcall_$wnnz_Int1_1sc_0_9_1Lcall_$wnnz_Int0_bufchan_r = (! wwsim_3_1ww1XiS_1_1lizzieLet27_4Lcall_$wnnz_Int1_1sc_0_9_1Lcall_$wnnz_Int0_bufchan_buf[0]);
  assign lizzieLet30_1_argbuf_d = (wwsim_3_1ww1XiS_1_1lizzieLet27_4Lcall_$wnnz_Int1_1sc_0_9_1Lcall_$wnnz_Int0_bufchan_buf[0] ? wwsim_3_1ww1XiS_1_1lizzieLet27_4Lcall_$wnnz_Int1_1sc_0_9_1Lcall_$wnnz_Int0_bufchan_buf :
                                   wwsim_3_1ww1XiS_1_1lizzieLet27_4Lcall_$wnnz_Int1_1sc_0_9_1Lcall_$wnnz_Int0_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      wwsim_3_1ww1XiS_1_1lizzieLet27_4Lcall_$wnnz_Int1_1sc_0_9_1Lcall_$wnnz_Int0_bufchan_buf <= {115'd0,
                                                                                                 1'd0};
    else
      if ((lizzieLet30_1_argbuf_r && wwsim_3_1ww1XiS_1_1lizzieLet27_4Lcall_$wnnz_Int1_1sc_0_9_1Lcall_$wnnz_Int0_bufchan_buf[0]))
        wwsim_3_1ww1XiS_1_1lizzieLet27_4Lcall_$wnnz_Int1_1sc_0_9_1Lcall_$wnnz_Int0_bufchan_buf <= {115'd0,
                                                                                                   1'd0};
      else if (((! lizzieLet30_1_argbuf_r) && (! wwsim_3_1ww1XiS_1_1lizzieLet27_4Lcall_$wnnz_Int1_1sc_0_9_1Lcall_$wnnz_Int0_bufchan_buf[0])))
        wwsim_3_1ww1XiS_1_1lizzieLet27_4Lcall_$wnnz_Int1_1sc_0_9_1Lcall_$wnnz_Int0_bufchan_buf <= wwsim_3_1ww1XiS_1_1lizzieLet27_4Lcall_$wnnz_Int1_1sc_0_9_1Lcall_$wnnz_Int0_bufchan_d;
  
  /* dcon (Ty CT$wnnz_Int,
      Dcon Lcall_$wnnz_Int0) : [(wwsim_3_destruct,Int#),
                                (ww1XiS_1_destruct,Int#),
                                (lizzieLet27_4Lcall_$wnnz_Int1,Int#),
                                (sc_0_9_destruct,Pointer_CT$wnnz_Int)] > (wwsim_3_1ww1XiS_1_1lizzieLet27_4Lcall_$wnnz_Int1_1sc_0_9_1Lcall_$wnnz_Int0,CT$wnnz_Int) */
  assign wwsim_3_1ww1XiS_1_1lizzieLet27_4Lcall_$wnnz_Int1_1sc_0_9_1Lcall_$wnnz_Int0_d = Lcall_$wnnz_Int0_dc((& {wwsim_3_destruct_d[0],
                                                                                                                ww1XiS_1_destruct_d[0],
                                                                                                                lizzieLet27_4Lcall_$wnnz_Int1_d[0],
                                                                                                                sc_0_9_destruct_d[0]}), wwsim_3_destruct_d, ww1XiS_1_destruct_d, lizzieLet27_4Lcall_$wnnz_Int1_d, sc_0_9_destruct_d);
  assign {wwsim_3_destruct_r,
          ww1XiS_1_destruct_r,
          lizzieLet27_4Lcall_$wnnz_Int1_r,
          sc_0_9_destruct_r} = {4 {(wwsim_3_1ww1XiS_1_1lizzieLet27_4Lcall_$wnnz_Int1_1sc_0_9_1Lcall_$wnnz_Int0_r && wwsim_3_1ww1XiS_1_1lizzieLet27_4Lcall_$wnnz_Int1_1sc_0_9_1Lcall_$wnnz_Int0_d[0])}};
  
  /* op_add (Ty Int#) : (wwsim_4_1ww1XiS_2_1_Add32,Int#) (ww2XiV_1_destruct,Int#) > (es_6_1_1ww2XiV_1_1_Add32,Int#) */
  assign es_6_1_1ww2XiV_1_1_Add32_d = {(wwsim_4_1ww1XiS_2_1_Add32_d[32:1] + ww2XiV_1_destruct_d[32:1]),
                                       (wwsim_4_1ww1XiS_2_1_Add32_d[0] && ww2XiV_1_destruct_d[0])};
  assign {wwsim_4_1ww1XiS_2_1_Add32_r,
          ww2XiV_1_destruct_r} = {2 {(es_6_1_1ww2XiV_1_1_Add32_r && es_6_1_1ww2XiV_1_1_Add32_d[0])}};
  
  /* op_add (Ty Int#) : (wwsim_4_destruct,Int#) (ww1XiS_2_destruct,Int#) > (wwsim_4_1ww1XiS_2_1_Add32,Int#) */
  assign wwsim_4_1ww1XiS_2_1_Add32_d = {(wwsim_4_destruct_d[32:1] + ww1XiS_2_destruct_d[32:1]),
                                        (wwsim_4_destruct_d[0] && ww1XiS_2_destruct_d[0])};
  assign {wwsim_4_destruct_r,
          ww1XiS_2_destruct_r} = {2 {(wwsim_4_1ww1XiS_2_1_Add32_r && wwsim_4_1ww1XiS_2_1_Add32_d[0])}};
endmodule