`timescale 1ns/1ns
import mMapAdd_package::*;

module mMapAdd(
  input logic clk,
  input logic reset,
  input Go_t \\QTree_Int_src_d ,
  output logic \\QTree_Int_src_r ,
  input QTree_Int_t dummy_write_QTree_Int_d,
  output logic dummy_write_QTree_Int_r,
  input Go_t sourceGo_d,
  output logic sourceGo_r,
  input Pointer_QTree_Int_t m1aey_0_d,
  output logic m1aey_0_r,
  input Pointer_QTree_Int_t m2aez_1_d,
  output logic m2aez_1_r,
  output \Word16#_t  forkHP1_QTree_Int_snk_dout,
  input logic forkHP1_QTree_Int_snk_rout,
  output Pointer_QTree_Int_t dummy_write_QTree_Int_sink_dout,
  input logic dummy_write_QTree_Int_sink_rout,
  output Int_t \es_7_1I#_dout ,
  input logic \es_7_1I#_rout 
  );
  /* --define=INPUTS=((__05CQTree_Int_src, 0, 1, Go), (dummy_write_QTree_Int, 66, 73786976294838206464, QTree_Int), (sourceGo, 0, 1, Go), (m1aey_0, 16, 65536, Pointer_QTree_Int), (m2aez_1, 16, 65536, Pointer_QTree_Int)) */
  /* --define=TAPS=() */
  /* --define=OUTPUTS=((forkHP1_QTree_Int_snk, 16, 65536, Word16__023), (dummy_write_QTree_Int_sink, 16, 65536, Pointer_QTree_Int), (es_7_1I__023, 32, 4294967296, Int)) */
  /* TYPE_START
CT__024wnnz 16 3 (0,[0]) (1,[16p,16p,16p,16p]) (2,[32,16p,16p,16p]) (3,[32,32,16p,16p]) (4,[32,32,32,16p])
CTf__027__027__027__027__027__027__027__027_f__027__027__027__027__027__027__027__027_Int_Int 16 3 (0,[0]) (1,[16p,16p,0,0,16p,16p]) (2,[16p,16p,16p,0,0,16p]) (3,[16p,16p,16p,16p,0,0]) (4,[16p,16p,16p,16p])
QTree_Int 16 2 (0,[0]) (1,[32]) (2,[16p,16p,16p,16p]) (3,[0])
CTf_f_Int_Int 16 3 (0,[0]) (1,[16p,16p,16p,0,0,0,0,16p,16p,16p,16p]) (2,[16p,16p,16p,16p,0,0,0,0,16p,16p]) (3,[16p,16p,16p,16p,16p,0,0,0,0]) (4,[16p,16p,16p,16p])
TupGo___Pointer_QTree_Int 16 0 (0,[0,16p])
TupGo___Pointer_QTree_Int___Pointer_CT__024wnnz 16 0 (0,[0,16p,16p])
TupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf__027__027__027__027__027__027__027__027_f__027__027__027__027__027__027__027__027_Int_Int 16 0 (0,[0,16p,0,0,16p])
TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Int 16 0 (0,[0,16p,16p,0,0,0,0,16p])
TupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int 16 0 (0,[0,16p,0,0])
TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int 16 0 (0,[0,16p,16p,0,0,0,0])
TYPE_END */
  /*  */
  /*  */
  Go_t go_1_d;
  logic go_1_r;
  Go_t go_2_d;
  logic go_2_r;
  Go_t go_3_d;
  logic go_3_r;
  Go_t go_4_d;
  logic go_4_r;
  Go_t go_5_d;
  logic go_5_r;
  Go_t go_6_d;
  logic go_6_r;
  Go_t go__7_d;
  logic go__7_r;
  Go_t go__8_d;
  logic go__8_r;
  Go_t go__9_d;
  logic go__9_r;
  Go_t go__10_d;
  logic go__10_r;
  Go_t go__11_d;
  logic go__11_r;
  Go_t go__12_d;
  logic go__12_r;
  \Word16#_t  initHP_CT$wnnz_d;
  logic initHP_CT$wnnz_r;
  \Word16#_t  incrHP_CT$wnnz_d;
  logic incrHP_CT$wnnz_r;
  Go_t incrHP_mergeCT$wnnz_d;
  logic incrHP_mergeCT$wnnz_r;
  Go_t incrHP_CT$wnnz1_d;
  logic incrHP_CT$wnnz1_r;
  Go_t incrHP_CT$wnnz2_d;
  logic incrHP_CT$wnnz2_r;
  \Word16#_t  addHP_CT$wnnz_d;
  logic addHP_CT$wnnz_r;
  \Word16#_t  mergeHP_CT$wnnz_d;
  logic mergeHP_CT$wnnz_r;
  Go_t incrHP_mergeCT$wnnz_buf_d;
  logic incrHP_mergeCT$wnnz_buf_r;
  \Word16#_t  mergeHP_CT$wnnz_buf_d;
  logic mergeHP_CT$wnnz_buf_r;
  \Word16#_t  forkHP1_CT$wnnz_d;
  logic forkHP1_CT$wnnz_r;
  \Word16#_t  forkHP1_CT$wnn2_d;
  logic forkHP1_CT$wnn2_r;
  \Word16#_t  forkHP1_CT$wnn3_d;
  logic forkHP1_CT$wnn3_r;
  C2_t memMergeChoice_CT$wnnz_d;
  logic memMergeChoice_CT$wnnz_r;
  MemIn_CT$wnnz_t memMergeIn_CT$wnnz_d;
  logic memMergeIn_CT$wnnz_r;
  MemOut_CT$wnnz_t memOut_CT$wnnz_d;
  logic memOut_CT$wnnz_r;
  MemOut_CT$wnnz_t memReadOut_CT$wnnz_d;
  logic memReadOut_CT$wnnz_r;
  MemOut_CT$wnnz_t memWriteOut_CT$wnnz_d;
  logic memWriteOut_CT$wnnz_r;
  MemIn_CT$wnnz_t memMergeIn_CT$wnnz_dbuf_d;
  logic memMergeIn_CT$wnnz_dbuf_r;
  MemIn_CT$wnnz_t memMergeIn_CT$wnnz_rbuf_d;
  logic memMergeIn_CT$wnnz_rbuf_r;
  MemOut_CT$wnnz_t memOut_CT$wnnz_dbuf_d;
  logic memOut_CT$wnnz_dbuf_r;
  MemOut_CT$wnnz_t memOut_CT$wnnz_rbuf_d;
  logic memOut_CT$wnnz_rbuf_r;
  \Word16#_t  destructReadIn_CT$wnnz_d;
  logic destructReadIn_CT$wnnz_r;
  MemIn_CT$wnnz_t dconReadIn_CT$wnnz_d;
  logic dconReadIn_CT$wnnz_r;
  CT$wnnz_t readPointer_CT$wnnzscfarg_0_1_argbuf_d;
  logic readPointer_CT$wnnzscfarg_0_1_argbuf_r;
  C5_t writeMerge_choice_CT$wnnz_d;
  logic writeMerge_choice_CT$wnnz_r;
  CT$wnnz_t writeMerge_data_CT$wnnz_d;
  logic writeMerge_data_CT$wnnz_r;
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet0_1_argbuf_d;
  logic writeCT$wnnzlizzieLet0_1_argbuf_r;
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet36_1_argbuf_d;
  logic writeCT$wnnzlizzieLet36_1_argbuf_r;
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet37_1_argbuf_d;
  logic writeCT$wnnzlizzieLet37_1_argbuf_r;
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet38_1_argbuf_d;
  logic writeCT$wnnzlizzieLet38_1_argbuf_r;
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet5_1_argbuf_d;
  logic writeCT$wnnzlizzieLet5_1_argbuf_r;
  MemIn_CT$wnnz_t dconWriteIn_CT$wnnz_d;
  logic dconWriteIn_CT$wnnz_r;
  Pointer_CT$wnnz_t dconPtr_CT$wnnz_d;
  logic dconPtr_CT$wnnz_r;
  Pointer_CT$wnnz_t _84_d;
  logic _84_r;
  assign _84_r = 1'd1;
  Pointer_CT$wnnz_t demuxWriteResult_CT$wnnz_d;
  logic demuxWriteResult_CT$wnnz_r;
  \Word16#_t  \initHP_CTf''''''''_f''''''''_Int_Int_d ;
  logic \initHP_CTf''''''''_f''''''''_Int_Int_r ;
  \Word16#_t  \incrHP_CTf''''''''_f''''''''_Int_Int_d ;
  logic \incrHP_CTf''''''''_f''''''''_Int_Int_r ;
  Go_t \incrHP_mergeCTf''''''''_f''''''''_Int_Int_d ;
  logic \incrHP_mergeCTf''''''''_f''''''''_Int_Int_r ;
  Go_t \incrHP_CTf''''''''_f''''''''_Int_Int1_d ;
  logic \incrHP_CTf''''''''_f''''''''_Int_Int1_r ;
  Go_t \incrHP_CTf''''''''_f''''''''_Int_Int2_d ;
  logic \incrHP_CTf''''''''_f''''''''_Int_Int2_r ;
  \Word16#_t  \addHP_CTf''''''''_f''''''''_Int_Int_d ;
  logic \addHP_CTf''''''''_f''''''''_Int_Int_r ;
  \Word16#_t  \mergeHP_CTf''''''''_f''''''''_Int_Int_d ;
  logic \mergeHP_CTf''''''''_f''''''''_Int_Int_r ;
  Go_t \incrHP_mergeCTf''''''''_f''''''''_Int_Int_buf_d ;
  logic \incrHP_mergeCTf''''''''_f''''''''_Int_Int_buf_r ;
  \Word16#_t  \mergeHP_CTf''''''''_f''''''''_Int_Int_buf_d ;
  logic \mergeHP_CTf''''''''_f''''''''_Int_Int_buf_r ;
  \Word16#_t  \forkHP1_CTf''''''''_f''''''''_Int_Int_d ;
  logic \forkHP1_CTf''''''''_f''''''''_Int_Int_r ;
  \Word16#_t  \forkHP1_CTf''''''''_f''''''''_Int_In2_d ;
  logic \forkHP1_CTf''''''''_f''''''''_Int_In2_r ;
  \Word16#_t  \forkHP1_CTf''''''''_f''''''''_Int_In3_d ;
  logic \forkHP1_CTf''''''''_f''''''''_Int_In3_r ;
  C2_t \memMergeChoice_CTf''''''''_f''''''''_Int_Int_d ;
  logic \memMergeChoice_CTf''''''''_f''''''''_Int_Int_r ;
  \MemIn_CTf''''''''_f''''''''_Int_Int_t  \memMergeIn_CTf''''''''_f''''''''_Int_Int_d ;
  logic \memMergeIn_CTf''''''''_f''''''''_Int_Int_r ;
  \MemOut_CTf''''''''_f''''''''_Int_Int_t  \memOut_CTf''''''''_f''''''''_Int_Int_d ;
  logic \memOut_CTf''''''''_f''''''''_Int_Int_r ;
  \MemOut_CTf''''''''_f''''''''_Int_Int_t  \memReadOut_CTf''''''''_f''''''''_Int_Int_d ;
  logic \memReadOut_CTf''''''''_f''''''''_Int_Int_r ;
  \MemOut_CTf''''''''_f''''''''_Int_Int_t  \memWriteOut_CTf''''''''_f''''''''_Int_Int_d ;
  logic \memWriteOut_CTf''''''''_f''''''''_Int_Int_r ;
  \MemIn_CTf''''''''_f''''''''_Int_Int_t  \memMergeIn_CTf''''''''_f''''''''_Int_Int_dbuf_d ;
  logic \memMergeIn_CTf''''''''_f''''''''_Int_Int_dbuf_r ;
  \MemIn_CTf''''''''_f''''''''_Int_Int_t  \memMergeIn_CTf''''''''_f''''''''_Int_Int_rbuf_d ;
  logic \memMergeIn_CTf''''''''_f''''''''_Int_Int_rbuf_r ;
  \MemOut_CTf''''''''_f''''''''_Int_Int_t  \memOut_CTf''''''''_f''''''''_Int_Int_dbuf_d ;
  logic \memOut_CTf''''''''_f''''''''_Int_Int_dbuf_r ;
  \MemOut_CTf''''''''_f''''''''_Int_Int_t  \memOut_CTf''''''''_f''''''''_Int_Int_rbuf_d ;
  logic \memOut_CTf''''''''_f''''''''_Int_Int_rbuf_r ;
  \Word16#_t  \destructReadIn_CTf''''''''_f''''''''_Int_Int_d ;
  logic \destructReadIn_CTf''''''''_f''''''''_Int_Int_r ;
  \MemIn_CTf''''''''_f''''''''_Int_Int_t  \dconReadIn_CTf''''''''_f''''''''_Int_Int_d ;
  logic \dconReadIn_CTf''''''''_f''''''''_Int_Int_r ;
  \CTf''''''''_f''''''''_Int_Int_t  \readPointer_CTf''''''''_f''''''''_Int_Intscfarg_0_1_1_argbuf_d ;
  logic \readPointer_CTf''''''''_f''''''''_Int_Intscfarg_0_1_1_argbuf_r ;
  C5_t \writeMerge_choice_CTf''''''''_f''''''''_Int_Int_d ;
  logic \writeMerge_choice_CTf''''''''_f''''''''_Int_Int_r ;
  \CTf''''''''_f''''''''_Int_Int_t  \writeMerge_data_CTf''''''''_f''''''''_Int_Int_d ;
  logic \writeMerge_data_CTf''''''''_f''''''''_Int_Int_r ;
  \Pointer_CTf''''''''_f''''''''_Int_Int_t  \writeCTf''''''''_f''''''''_Int_IntlizzieLet10_1_argbuf_d ;
  logic \writeCTf''''''''_f''''''''_Int_IntlizzieLet10_1_argbuf_r ;
  \Pointer_CTf''''''''_f''''''''_Int_Int_t  \writeCTf''''''''_f''''''''_Int_IntlizzieLet33_1_argbuf_d ;
  logic \writeCTf''''''''_f''''''''_Int_IntlizzieLet33_1_argbuf_r ;
  \Pointer_CTf''''''''_f''''''''_Int_Int_t  \writeCTf''''''''_f''''''''_Int_IntlizzieLet40_1_argbuf_d ;
  logic \writeCTf''''''''_f''''''''_Int_IntlizzieLet40_1_argbuf_r ;
  \Pointer_CTf''''''''_f''''''''_Int_Int_t  \writeCTf''''''''_f''''''''_Int_IntlizzieLet41_1_argbuf_d ;
  logic \writeCTf''''''''_f''''''''_Int_IntlizzieLet41_1_argbuf_r ;
  \Pointer_CTf''''''''_f''''''''_Int_Int_t  \writeCTf''''''''_f''''''''_Int_IntlizzieLet42_1_argbuf_d ;
  logic \writeCTf''''''''_f''''''''_Int_IntlizzieLet42_1_argbuf_r ;
  \MemIn_CTf''''''''_f''''''''_Int_Int_t  \dconWriteIn_CTf''''''''_f''''''''_Int_Int_d ;
  logic \dconWriteIn_CTf''''''''_f''''''''_Int_Int_r ;
  \Pointer_CTf''''''''_f''''''''_Int_Int_t  \dconPtr_CTf''''''''_f''''''''_Int_Int_d ;
  logic \dconPtr_CTf''''''''_f''''''''_Int_Int_r ;
  \Pointer_CTf''''''''_f''''''''_Int_Int_t  _83_d;
  logic _83_r;
  assign _83_r = 1'd1;
  \Pointer_CTf''''''''_f''''''''_Int_Int_t  \demuxWriteResult_CTf''''''''_f''''''''_Int_Int_d ;
  logic \demuxWriteResult_CTf''''''''_f''''''''_Int_Int_r ;
  \Word16#_t  initHP_QTree_Int_d;
  logic initHP_QTree_Int_r;
  \Word16#_t  incrHP_QTree_Int_d;
  logic incrHP_QTree_Int_r;
  Go_t incrHP_mergeQTree_Int_d;
  logic incrHP_mergeQTree_Int_r;
  Go_t incrHP_QTree_Int1_d;
  logic incrHP_QTree_Int1_r;
  Go_t incrHP_QTree_Int2_d;
  logic incrHP_QTree_Int2_r;
  \Word16#_t  addHP_QTree_Int_d;
  logic addHP_QTree_Int_r;
  \Word16#_t  mergeHP_QTree_Int_d;
  logic mergeHP_QTree_Int_r;
  Go_t incrHP_mergeQTree_Int_buf_d;
  logic incrHP_mergeQTree_Int_buf_r;
  \Word16#_t  mergeHP_QTree_Int_buf_d;
  logic mergeHP_QTree_Int_buf_r;
  Go_t go_1_dummy_write_QTree_Int_d;
  logic go_1_dummy_write_QTree_Int_r;
  Go_t go_2_dummy_write_QTree_Int_d;
  logic go_2_dummy_write_QTree_Int_r;
  \Word16#_t  forkHP1_QTree_Int_d;
  logic forkHP1_QTree_Int_r;
  \Word16#_t  forkHP1_QTree_Int_snk_d;
  logic forkHP1_QTree_Int_snk_r;
  \Word16#_t  forkHP1_QTree_In3_d;
  logic forkHP1_QTree_In3_r;
  \Word16#_t  forkHP1_QTree_In4_d;
  logic forkHP1_QTree_In4_r;
  C2_t memMergeChoice_QTree_Int_d;
  logic memMergeChoice_QTree_Int_r;
  MemIn_QTree_Int_t memMergeIn_QTree_Int_d;
  logic memMergeIn_QTree_Int_r;
  MemOut_QTree_Int_t memOut_QTree_Int_d;
  logic memOut_QTree_Int_r;
  MemOut_QTree_Int_t memReadOut_QTree_Int_d;
  logic memReadOut_QTree_Int_r;
  MemOut_QTree_Int_t memWriteOut_QTree_Int_d;
  logic memWriteOut_QTree_Int_r;
  MemIn_QTree_Int_t memMergeIn_QTree_Int_dbuf_d;
  logic memMergeIn_QTree_Int_dbuf_r;
  MemIn_QTree_Int_t memMergeIn_QTree_Int_rbuf_d;
  logic memMergeIn_QTree_Int_rbuf_r;
  MemOut_QTree_Int_t memOut_QTree_Int_dbuf_d;
  logic memOut_QTree_Int_dbuf_r;
  MemOut_QTree_Int_t memOut_QTree_Int_rbuf_d;
  logic memOut_QTree_Int_rbuf_r;
  C4_t readMerge_choice_QTree_Int_d;
  logic readMerge_choice_QTree_Int_r;
  Pointer_QTree_Int_t readMerge_data_QTree_Int_d;
  logic readMerge_data_QTree_Int_r;
  QTree_Int_t readPointer_QTree_Intm1a8C_1_argbuf_d;
  logic readPointer_QTree_Intm1a8C_1_argbuf_r;
  QTree_Int_t readPointer_QTree_Intm2a8D_1_argbuf_d;
  logic readPointer_QTree_Intm2a8D_1_argbuf_r;
  QTree_Int_t readPointer_QTree_Intq4a8u_1_argbuf_d;
  logic readPointer_QTree_Intq4a8u_1_argbuf_r;
  QTree_Int_t readPointer_QTree_IntwsiX_1_1_argbuf_d;
  logic readPointer_QTree_IntwsiX_1_1_argbuf_r;
  \Word16#_t  destructReadIn_QTree_Int_d;
  logic destructReadIn_QTree_Int_r;
  MemIn_QTree_Int_t dconReadIn_QTree_Int_d;
  logic dconReadIn_QTree_Int_r;
  QTree_Int_t destructReadOut_QTree_Int_d;
  logic destructReadOut_QTree_Int_r;
  C23_t writeMerge_choice_QTree_Int_d;
  logic writeMerge_choice_QTree_Int_r;
  QTree_Int_t writeMerge_data_QTree_Int_d;
  logic writeMerge_data_QTree_Int_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet11_1_argbuf_d;
  logic writeQTree_IntlizzieLet11_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet14_1_argbuf_d;
  logic writeQTree_IntlizzieLet14_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet15_1_argbuf_d;
  logic writeQTree_IntlizzieLet15_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet16_1_argbuf_d;
  logic writeQTree_IntlizzieLet16_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet17_1_argbuf_d;
  logic writeQTree_IntlizzieLet17_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet18_1_argbuf_d;
  logic writeQTree_IntlizzieLet18_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet20_1_argbuf_d;
  logic writeQTree_IntlizzieLet20_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet21_1_argbuf_d;
  logic writeQTree_IntlizzieLet21_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet22_1_argbuf_d;
  logic writeQTree_IntlizzieLet22_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet23_2_1_argbuf_d;
  logic writeQTree_IntlizzieLet23_2_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet24_1_1_argbuf_d;
  logic writeQTree_IntlizzieLet24_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet25_1_1_argbuf_d;
  logic writeQTree_IntlizzieLet25_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet26_1_argbuf_d;
  logic writeQTree_IntlizzieLet26_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet28_1_argbuf_d;
  logic writeQTree_IntlizzieLet28_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet29_1_argbuf_d;
  logic writeQTree_IntlizzieLet29_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet31_1_argbuf_d;
  logic writeQTree_IntlizzieLet31_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet32_1_argbuf_d;
  logic writeQTree_IntlizzieLet32_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet43_1_argbuf_d;
  logic writeQTree_IntlizzieLet43_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet48_1_argbuf_d;
  logic writeQTree_IntlizzieLet48_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet7_1_argbuf_d;
  logic writeQTree_IntlizzieLet7_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet8_1_argbuf_d;
  logic writeQTree_IntlizzieLet8_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet9_1_argbuf_d;
  logic writeQTree_IntlizzieLet9_1_argbuf_r;
  Pointer_QTree_Int_t dummy_write_QTree_Int_sink_d;
  logic dummy_write_QTree_Int_sink_r;
  MemIn_QTree_Int_t dconWriteIn_QTree_Int_d;
  logic dconWriteIn_QTree_Int_r;
  Pointer_QTree_Int_t dconPtr_QTree_Int_d;
  logic dconPtr_QTree_Int_r;
  Pointer_QTree_Int_t _82_d;
  logic _82_r;
  assign _82_r = 1'd1;
  Pointer_QTree_Int_t demuxWriteResult_QTree_Int_d;
  logic demuxWriteResult_QTree_Int_r;
  \Word16#_t  initHP_CTf_f_Int_Int_d;
  logic initHP_CTf_f_Int_Int_r;
  \Word16#_t  incrHP_CTf_f_Int_Int_d;
  logic incrHP_CTf_f_Int_Int_r;
  Go_t incrHP_mergeCTf_f_Int_Int_d;
  logic incrHP_mergeCTf_f_Int_Int_r;
  Go_t incrHP_CTf_f_Int_Int1_d;
  logic incrHP_CTf_f_Int_Int1_r;
  Go_t incrHP_CTf_f_Int_Int2_d;
  logic incrHP_CTf_f_Int_Int2_r;
  \Word16#_t  addHP_CTf_f_Int_Int_d;
  logic addHP_CTf_f_Int_Int_r;
  \Word16#_t  mergeHP_CTf_f_Int_Int_d;
  logic mergeHP_CTf_f_Int_Int_r;
  Go_t incrHP_mergeCTf_f_Int_Int_buf_d;
  logic incrHP_mergeCTf_f_Int_Int_buf_r;
  \Word16#_t  mergeHP_CTf_f_Int_Int_buf_d;
  logic mergeHP_CTf_f_Int_Int_buf_r;
  \Word16#_t  forkHP1_CTf_f_Int_Int_d;
  logic forkHP1_CTf_f_Int_Int_r;
  \Word16#_t  forkHP1_CTf_f_Int_In2_d;
  logic forkHP1_CTf_f_Int_In2_r;
  \Word16#_t  forkHP1_CTf_f_Int_In3_d;
  logic forkHP1_CTf_f_Int_In3_r;
  C2_t memMergeChoice_CTf_f_Int_Int_d;
  logic memMergeChoice_CTf_f_Int_Int_r;
  MemIn_CTf_f_Int_Int_t memMergeIn_CTf_f_Int_Int_d;
  logic memMergeIn_CTf_f_Int_Int_r;
  MemOut_CTf_f_Int_Int_t memOut_CTf_f_Int_Int_d;
  logic memOut_CTf_f_Int_Int_r;
  MemOut_CTf_f_Int_Int_t memReadOut_CTf_f_Int_Int_d;
  logic memReadOut_CTf_f_Int_Int_r;
  MemOut_CTf_f_Int_Int_t memWriteOut_CTf_f_Int_Int_d;
  logic memWriteOut_CTf_f_Int_Int_r;
  MemIn_CTf_f_Int_Int_t memMergeIn_CTf_f_Int_Int_dbuf_d;
  logic memMergeIn_CTf_f_Int_Int_dbuf_r;
  MemIn_CTf_f_Int_Int_t memMergeIn_CTf_f_Int_Int_rbuf_d;
  logic memMergeIn_CTf_f_Int_Int_rbuf_r;
  MemOut_CTf_f_Int_Int_t memOut_CTf_f_Int_Int_dbuf_d;
  logic memOut_CTf_f_Int_Int_dbuf_r;
  MemOut_CTf_f_Int_Int_t memOut_CTf_f_Int_Int_rbuf_d;
  logic memOut_CTf_f_Int_Int_rbuf_r;
  \Word16#_t  destructReadIn_CTf_f_Int_Int_d;
  logic destructReadIn_CTf_f_Int_Int_r;
  MemIn_CTf_f_Int_Int_t dconReadIn_CTf_f_Int_Int_d;
  logic dconReadIn_CTf_f_Int_Int_r;
  CTf_f_Int_Int_t readPointer_CTf_f_Int_Intscfarg_0_2_1_argbuf_d;
  logic readPointer_CTf_f_Int_Intscfarg_0_2_1_argbuf_r;
  C5_t writeMerge_choice_CTf_f_Int_Int_d;
  logic writeMerge_choice_CTf_f_Int_Int_r;
  CTf_f_Int_Int_t writeMerge_data_CTf_f_Int_Int_d;
  logic writeMerge_data_CTf_f_Int_Int_r;
  Pointer_CTf_f_Int_Int_t writeCTf_f_Int_IntlizzieLet30_1_argbuf_d;
  logic writeCTf_f_Int_IntlizzieLet30_1_argbuf_r;
  Pointer_CTf_f_Int_Int_t writeCTf_f_Int_IntlizzieLet34_1_argbuf_d;
  logic writeCTf_f_Int_IntlizzieLet34_1_argbuf_r;
  Pointer_CTf_f_Int_Int_t writeCTf_f_Int_IntlizzieLet45_1_argbuf_d;
  logic writeCTf_f_Int_IntlizzieLet45_1_argbuf_r;
  Pointer_CTf_f_Int_Int_t writeCTf_f_Int_IntlizzieLet46_1_argbuf_d;
  logic writeCTf_f_Int_IntlizzieLet46_1_argbuf_r;
  Pointer_CTf_f_Int_Int_t writeCTf_f_Int_IntlizzieLet47_1_argbuf_d;
  logic writeCTf_f_Int_IntlizzieLet47_1_argbuf_r;
  MemIn_CTf_f_Int_Int_t dconWriteIn_CTf_f_Int_Int_d;
  logic dconWriteIn_CTf_f_Int_Int_r;
  Pointer_CTf_f_Int_Int_t dconPtr_CTf_f_Int_Int_d;
  logic dconPtr_CTf_f_Int_Int_r;
  Pointer_CTf_f_Int_Int_t _81_d;
  logic _81_r;
  assign _81_r = 1'd1;
  Pointer_CTf_f_Int_Int_t demuxWriteResult_CTf_f_Int_Int_d;
  logic demuxWriteResult_CTf_f_Int_Int_r;
  Go_t \$wnnzTupGo___Pointer_QTree_Intgo_7_d ;
  logic \$wnnzTupGo___Pointer_QTree_Intgo_7_r ;
  Pointer_QTree_Int_t \$wnnzTupGo___Pointer_QTree_IntwsiX_d ;
  logic \$wnnzTupGo___Pointer_QTree_IntwsiX_r ;
  Go_t go_7_1_d;
  logic go_7_1_r;
  Go_t go_7_2_d;
  logic go_7_2_r;
  Pointer_QTree_Int_t wsiX_1_argbuf_d;
  logic wsiX_1_argbuf_r;
  Int_t \es_7_1I#_d ;
  logic \es_7_1I#_r ;
  C5_t applyfnInt_Bool_5_choice_d;
  logic applyfnInt_Bool_5_choice_r;
  TupGo___MyDTInt_Bool___Int_t applyfnInt_Bool_5_data_d;
  logic applyfnInt_Bool_5_data_r;
  MyDTInt_Bool_t arg0_1_d;
  logic arg0_1_r;
  MyDTInt_Bool_t arg0_2_d;
  logic arg0_2_r;
  MyDTInt_Bool_t arg0_3_d;
  logic arg0_3_r;
  MyBool_t applyfnInt_Bool_5_resbuf_d;
  logic applyfnInt_Bool_5_resbuf_r;
  MyBool_t applyfnInt_Bool_5_2_argbuf_d;
  logic applyfnInt_Bool_5_2_argbuf_r;
  MyBool_t es_2_1_d;
  logic es_2_1_r;
  MyBool_t es_2_2_d;
  logic es_2_2_r;
  MyBool_t es_2_3_d;
  logic es_2_3_r;
  MyBool_t es_2_4_d;
  logic es_2_4_r;
  MyBool_t applyfnInt_Bool_5_3_argbuf_d;
  logic applyfnInt_Bool_5_3_argbuf_r;
  MyBool_t es_10_1_d;
  logic es_10_1_r;
  MyBool_t es_10_2_d;
  logic es_10_2_r;
  MyBool_t es_10_3_d;
  logic es_10_3_r;
  MyBool_t es_10_4_d;
  logic es_10_4_r;
  MyBool_t applyfnInt_Bool_5_4_argbuf_d;
  logic applyfnInt_Bool_5_4_argbuf_r;
  MyBool_t es_14_1_d;
  logic es_14_1_r;
  MyBool_t es_14_2_d;
  logic es_14_2_r;
  MyBool_t es_14_3_d;
  logic es_14_3_r;
  MyBool_t es_14_4_d;
  logic es_14_4_r;
  MyBool_t es_14_5_d;
  logic es_14_5_r;
  MyBool_t es_14_6_d;
  logic es_14_6_r;
  MyBool_t es_14_7_d;
  logic es_14_7_r;
  MyBool_t applyfnInt_Bool_5_5_argbuf_d;
  logic applyfnInt_Bool_5_5_argbuf_r;
  MyBool_t es_19_1_d;
  logic es_19_1_r;
  MyBool_t es_19_2_d;
  logic es_19_2_r;
  MyBool_t es_19_3_d;
  logic es_19_3_r;
  MyBool_t es_19_4_d;
  logic es_19_4_r;
  MyBool_t es_19_5_d;
  logic es_19_5_r;
  MyBool_t es_19_6_d;
  logic es_19_6_r;
  MyBool_t applyfnInt_Bool_5_1_d;
  logic applyfnInt_Bool_5_1_r;
  MyBool_t applyfnInt_Bool_5_2_d;
  logic applyfnInt_Bool_5_2_r;
  MyBool_t applyfnInt_Bool_5_3_d;
  logic applyfnInt_Bool_5_3_r;
  MyBool_t applyfnInt_Bool_5_4_d;
  logic applyfnInt_Bool_5_4_r;
  MyBool_t applyfnInt_Bool_5_5_d;
  logic applyfnInt_Bool_5_5_r;
  Go_t applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intgo_8_d;
  logic applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intgo_8_r;
  MyDTInt_Bool_t applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_d;
  logic applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_r;
  Int_t applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg1_d;
  logic applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg1_r;
  MyBool_t es_2_1_1_d;
  logic es_2_1_1_r;
  MyBool_t es_2_1_2_d;
  logic es_2_1_2_r;
  MyBool_t es_2_1_3_d;
  logic es_2_1_3_r;
  MyBool_t es_2_1_4_d;
  logic es_2_1_4_r;
  C8_t applyfnInt_Int_5_choice_d;
  logic applyfnInt_Int_5_choice_r;
  TupGo___MyDTInt_Int___Int_t applyfnInt_Int_5_data_d;
  logic applyfnInt_Int_5_data_r;
  MyDTInt_Int_t arg0_2_1_d;
  logic arg0_2_1_r;
  MyDTInt_Int_t arg0_2_2_d;
  logic arg0_2_2_r;
  MyDTInt_Int_t arg0_2_3_d;
  logic arg0_2_3_r;
  Int_t applyfnInt_Int_5_resbuf_d;
  logic applyfnInt_Int_5_resbuf_r;
  Int_t applyfnInt_Int_5_2_argbuf_d;
  logic applyfnInt_Int_5_2_argbuf_r;
  QTree_Int_t es_3_2_1QVal_Int_d;
  logic es_3_2_1QVal_Int_r;
  Int_t applyfnInt_Int_5_3_argbuf_d;
  logic applyfnInt_Int_5_3_argbuf_r;
  Int_t es_1_1_argbuf_d;
  logic es_1_1_argbuf_r;
  Int_t applyfnInt_Int_5_4_argbuf_d;
  logic applyfnInt_Int_5_4_argbuf_r;
  QTree_Int_t es_3_1_1QVal_Int_d;
  logic es_3_1_1QVal_Int_r;
  Int_t applyfnInt_Int_5_5_argbuf_d;
  logic applyfnInt_Int_5_5_argbuf_r;
  Int_t es_9_1_argbuf_d;
  logic es_9_1_argbuf_r;
  Int_t applyfnInt_Int_5_6_argbuf_d;
  logic applyfnInt_Int_5_6_argbuf_r;
  QTree_Int_t es_11_1QVal_Int_d;
  logic es_11_1QVal_Int_r;
  Int_t applyfnInt_Int_5_7_argbuf_d;
  logic applyfnInt_Int_5_7_argbuf_r;
  Int_t es_16_1_argbuf_d;
  logic es_16_1_argbuf_r;
  Int_t applyfnInt_Int_5_8_argbuf_d;
  logic applyfnInt_Int_5_8_argbuf_r;
  QTree_Int_t es_20_1QVal_Int_d;
  logic es_20_1QVal_Int_r;
  Int_t applyfnInt_Int_5_1_d;
  logic applyfnInt_Int_5_1_r;
  Int_t applyfnInt_Int_5_2_d;
  logic applyfnInt_Int_5_2_r;
  Int_t applyfnInt_Int_5_3_d;
  logic applyfnInt_Int_5_3_r;
  Int_t applyfnInt_Int_5_4_d;
  logic applyfnInt_Int_5_4_r;
  Int_t applyfnInt_Int_5_5_d;
  logic applyfnInt_Int_5_5_r;
  Int_t applyfnInt_Int_5_6_d;
  logic applyfnInt_Int_5_6_r;
  Int_t applyfnInt_Int_5_7_d;
  logic applyfnInt_Int_5_7_r;
  Int_t applyfnInt_Int_5_8_d;
  logic applyfnInt_Int_5_8_r;
  Go_t applyfnInt_Int_5TupGo___MyDTInt_Int___Intgo_9_d;
  logic applyfnInt_Int_5TupGo___MyDTInt_Int___Intgo_9_r;
  MyDTInt_Int_t applyfnInt_Int_5TupGo___MyDTInt_Int___Intarg0_2_d;
  logic applyfnInt_Int_5TupGo___MyDTInt_Int___Intarg0_2_r;
  Int_t applyfnInt_Int_5TupGo___MyDTInt_Int___Intarg1_1_d;
  logic applyfnInt_Int_5TupGo___MyDTInt_Int___Intarg1_1_r;
  Int_t es_1_1_1_argbuf_d;
  logic es_1_1_1_argbuf_r;
  C3_t applyfnInt_Int_Int_5_choice_d;
  logic applyfnInt_Int_Int_5_choice_r;
  TupMyDTInt_Int_Int___Int___Int_t applyfnInt_Int_Int_5_data_d;
  logic applyfnInt_Int_Int_5_data_r;
  MyDTInt_Int_Int_t arg0_4_1_d;
  logic arg0_4_1_r;
  MyDTInt_Int_Int_t arg0_4_2_d;
  logic arg0_4_2_r;
  MyDTInt_Int_Int_t arg0_4_3_d;
  logic arg0_4_3_r;
  Int_t applyfnInt_Int_Int_5_resbuf_d;
  logic applyfnInt_Int_Int_5_resbuf_r;
  Int_t applyfnInt_Int_Int_5_2_argbuf_d;
  logic applyfnInt_Int_Int_5_2_argbuf_r;
  Int_t es_18_1_argbuf_d;
  logic es_18_1_argbuf_r;
  Int_t applyfnInt_Int_Int_5_3_argbuf_d;
  logic applyfnInt_Int_Int_5_3_argbuf_r;
  Int_t es_22_1_argbuf_d;
  logic es_22_1_argbuf_r;
  Int_t applyfnInt_Int_Int_5_1_d;
  logic applyfnInt_Int_Int_5_1_r;
  Int_t applyfnInt_Int_Int_5_2_d;
  logic applyfnInt_Int_Int_5_2_r;
  Int_t applyfnInt_Int_Int_5_3_d;
  logic applyfnInt_Int_Int_5_3_r;
  MyDTInt_Int_Int_t applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_4_d;
  logic applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_4_r;
  Int_t applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg2_d;
  logic applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg2_r;
  Int_t applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg1_2_d;
  logic applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg1_2_r;
  Int_t es_13_1_argbuf_d;
  logic es_13_1_argbuf_r;
  Int_t arg0_1Dcon_is_z_1_d;
  logic arg0_1Dcon_is_z_1_r;
  Int_t arg0_1Dcon_is_z_1_1_d;
  logic arg0_1Dcon_is_z_1_1_r;
  Int_t arg0_1Dcon_is_z_1_2_d;
  logic arg0_1Dcon_is_z_1_2_r;
  Int_t arg0_1Dcon_is_z_1_3_d;
  logic arg0_1Dcon_is_z_1_3_r;
  Int_t arg0_1Dcon_is_z_1_4_d;
  logic arg0_1Dcon_is_z_1_4_r;
  \Int#_t  x1ah2_destruct_d;
  logic x1ah2_destruct_r;
  Int_t \arg0_1Dcon_is_z_1_1I#_d ;
  logic \arg0_1Dcon_is_z_1_1I#_r ;
  Go_t \arg0_1Dcon_is_z_1_3I#_d ;
  logic \arg0_1Dcon_is_z_1_3I#_r ;
  Go_t \arg0_1Dcon_is_z_1_3I#_1_d ;
  logic \arg0_1Dcon_is_z_1_3I#_1_r ;
  Go_t \arg0_1Dcon_is_z_1_3I#_2_d ;
  logic \arg0_1Dcon_is_z_1_3I#_2_r ;
  Go_t \arg0_1Dcon_is_z_1_3I#_3_d ;
  logic \arg0_1Dcon_is_z_1_3I#_3_r ;
  Go_t \arg0_1Dcon_is_z_1_3I#_1_argbuf_d ;
  logic \arg0_1Dcon_is_z_1_3I#_1_argbuf_r ;
  \Int#_t  \arg0_1Dcon_is_z_1_3I#_1_argbuf_0_d ;
  logic \arg0_1Dcon_is_z_1_3I#_1_argbuf_0_r ;
  Bool_t lizzieLet1_1wild1Xr_1_Eq_d;
  logic lizzieLet1_1wild1Xr_1_Eq_r;
  Go_t \arg0_1Dcon_is_z_1_3I#_2_argbuf_d ;
  logic \arg0_1Dcon_is_z_1_3I#_2_argbuf_r ;
  TupGo___Bool_t boolConvert_1TupGo___Bool_1_d;
  logic boolConvert_1TupGo___Bool_1_r;
  MyBool_t lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_d;
  logic lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_r;
  Go_t arg0_2Dcon_is_z_1_d;
  logic arg0_2Dcon_is_z_1_r;
  Int_t arg0_2_1Dcon_main1_d;
  logic arg0_2_1Dcon_main1_r;
  Int_t arg0_2_1Dcon_main1_1_d;
  logic arg0_2_1Dcon_main1_1_r;
  Int_t arg0_2_1Dcon_main1_2_d;
  logic arg0_2_1Dcon_main1_2_r;
  Int_t arg0_2_1Dcon_main1_3_d;
  logic arg0_2_1Dcon_main1_3_r;
  Int_t arg0_2_1Dcon_main1_4_d;
  logic arg0_2_1Dcon_main1_4_r;
  \Int#_t  x1agS_destruct_d;
  logic x1agS_destruct_r;
  Int_t \arg0_2_1Dcon_main1_1I#_d ;
  logic \arg0_2_1Dcon_main1_1I#_r ;
  Go_t \arg0_2_1Dcon_main1_3I#_d ;
  logic \arg0_2_1Dcon_main1_3I#_r ;
  Go_t \arg0_2_1Dcon_main1_3I#_1_argbuf_d ;
  logic \arg0_2_1Dcon_main1_3I#_1_argbuf_r ;
  \Int#_t  \arg0_2_1Dcon_main1_3I#_1_argbuf_2_d ;
  logic \arg0_2_1Dcon_main1_3I#_1_argbuf_2_r ;
  Int_t \es_0_1_1I#_mux_d ;
  logic \es_0_1_1I#_mux_r ;
  Go_t arg0_2_2Dcon_main1_d;
  logic arg0_2_2Dcon_main1_r;
  Int_t \es_0_1_1I#_mux_mux_d ;
  logic \es_0_1_1I#_mux_mux_r ;
  MyBool_t lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_d;
  logic lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_r;
  Int_t \arg0_4_1Dcon_$fNumInt_$c+_d ;
  logic \arg0_4_1Dcon_$fNumInt_$c+_r ;
  Int_t \arg0_4_2Dcon_$fNumInt_$c+_d ;
  logic \arg0_4_2Dcon_$fNumInt_$c+_r ;
  Int_t \arg0_4_2Dcon_$fNumInt_$c+_1_d ;
  logic \arg0_4_2Dcon_$fNumInt_$c+_1_r ;
  Int_t \arg0_4_2Dcon_$fNumInt_$c+_2_d ;
  logic \arg0_4_2Dcon_$fNumInt_$c+_2_r ;
  Int_t \arg0_4_2Dcon_$fNumInt_$c+_3_d ;
  logic \arg0_4_2Dcon_$fNumInt_$c+_3_r ;
  Int_t \arg0_4_2Dcon_$fNumInt_$c+_4_d ;
  logic \arg0_4_2Dcon_$fNumInt_$c+_4_r ;
  \Int#_t  xa1lV_destruct_d;
  logic xa1lV_destruct_r;
  Int_t \arg0_4_2Dcon_$fNumInt_$c+_1I#_d ;
  logic \arg0_4_2Dcon_$fNumInt_$c+_1I#_r ;
  Int_t \arg0_4_2Dcon_$fNumInt_$c+_3I#_d ;
  logic \arg0_4_2Dcon_$fNumInt_$c+_3I#_r ;
  Int_t \arg0_4_2Dcon_$fNumInt_$c+_3I#_1_d ;
  logic \arg0_4_2Dcon_$fNumInt_$c+_3I#_1_r ;
  Int_t \arg0_4_2Dcon_$fNumInt_$c+_3I#_2_d ;
  logic \arg0_4_2Dcon_$fNumInt_$c+_3I#_2_r ;
  Int_t \arg0_4_2Dcon_$fNumInt_$c+_3I#_3_d ;
  logic \arg0_4_2Dcon_$fNumInt_$c+_3I#_3_r ;
  Int_t \arg0_4_2Dcon_$fNumInt_$c+_3I#_4_d ;
  logic \arg0_4_2Dcon_$fNumInt_$c+_3I#_4_r ;
  \Int#_t  ya1lW_destruct_d;
  logic ya1lW_destruct_r;
  Int_t \arg0_4_2Dcon_$fNumInt_$c+_3I#_1I#_d ;
  logic \arg0_4_2Dcon_$fNumInt_$c+_3I#_1I#_r ;
  \Int#_t  \arg0_4_2Dcon_$fNumInt_$c+_3I#_3I#_d ;
  logic \arg0_4_2Dcon_$fNumInt_$c+_3I#_3I#_r ;
  \Int#_t  \arg0_4_2Dcon_$fNumInt_$c+_3I#_3I#_1ya1lW_1_Add32_d ;
  logic \arg0_4_2Dcon_$fNumInt_$c+_3I#_3I#_1ya1lW_1_Add32_r ;
  Int_t \es_0_2_1I#_d ;
  logic \es_0_2_1I#_r ;
  Int_t \es_0_2_1I#_mux_d ;
  logic \es_0_2_1I#_mux_r ;
  Int_t \es_0_2_1I#_mux_mux_d ;
  logic \es_0_2_1I#_mux_mux_r ;
  Int_t \es_0_2_1I#_mux_mux_mux_d ;
  logic \es_0_2_1I#_mux_mux_mux_r ;
  Pointer_QTree_Int_t bla8A_1_1_argbuf_d;
  logic bla8A_1_1_argbuf_r;
  Pointer_QTree_Int_t bla8L_1_argbuf_d;
  logic bla8L_1_argbuf_r;
  Go_t boolConvert_1TupGo___Boolgo_1_d;
  logic boolConvert_1TupGo___Boolgo_1_r;
  Bool_t boolConvert_1TupGo___Boolbool_d;
  logic boolConvert_1TupGo___Boolbool_r;
  Bool_t bool_1_d;
  logic bool_1_r;
  Bool_t bool_2_d;
  logic bool_2_r;
  MyBool_t lizzieLet3_1_d;
  logic lizzieLet3_1_r;
  MyBool_t lizzieLet3_2_d;
  logic lizzieLet3_2_r;
  Go_t bool_1False_d;
  logic bool_1False_r;
  Go_t bool_1True_d;
  logic bool_1True_r;
  MyBool_t bool_1False_1MyFalse_d;
  logic bool_1False_1MyFalse_r;
  MyBool_t boolConvert_1_resbuf_d;
  logic boolConvert_1_resbuf_r;
  MyBool_t bool_1True_1MyTrue_d;
  logic bool_1True_1MyTrue_r;
  MyBool_t bool_1False_1MyFalsebool_1True_1MyTrue_mux_d;
  logic bool_1False_1MyFalsebool_1True_1MyTrue_mux_r;
  Pointer_QTree_Int_t bra8B_1_argbuf_d;
  logic bra8B_1_argbuf_r;
  Pointer_QTree_Int_t bra8M_1_argbuf_d;
  logic bra8M_1_argbuf_r;
  Go_t call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnzgo_10_d;
  logic call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnzgo_10_r;
  Pointer_QTree_Int_t call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnzwsiX_1_d;
  logic call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnzwsiX_1_r;
  Pointer_CT$wnnz_t call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnzsc_0_d;
  logic call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnzsc_0_r;
  Go_t call_$wnnz_initBufi_d;
  logic call_$wnnz_initBufi_r;
  C5_t go_10_goMux_choice_d;
  logic go_10_goMux_choice_r;
  Go_t go_10_goMux_data_d;
  logic go_10_goMux_data_r;
  Go_t call_$wnnz_unlockFork1_d;
  logic call_$wnnz_unlockFork1_r;
  Go_t call_$wnnz_unlockFork2_d;
  logic call_$wnnz_unlockFork2_r;
  Go_t call_$wnnz_unlockFork3_d;
  logic call_$wnnz_unlockFork3_r;
  Go_t call_$wnnz_initBuf_d;
  logic call_$wnnz_initBuf_r;
  Go_t call_$wnnz_goMux1_d;
  logic call_$wnnz_goMux1_r;
  Pointer_QTree_Int_t call_$wnnz_goMux2_d;
  logic call_$wnnz_goMux2_r;
  Pointer_CT$wnnz_t call_$wnnz_goMux3_d;
  logic call_$wnnz_goMux3_r;
  Go_t \call_f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf''''''''_f''''''''_Int_Intgo_11_d ;
  logic \call_f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf''''''''_f''''''''_Int_Intgo_11_r ;
  Pointer_QTree_Int_t \call_f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf''''''''_f''''''''_Int_Intq4a8u_d ;
  logic \call_f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf''''''''_f''''''''_Int_Intq4a8u_r ;
  MyDTInt_Bool_t \call_f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf''''''''_f''''''''_Int_Intis_z_mapa8v_d ;
  logic \call_f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf''''''''_f''''''''_Int_Intis_z_mapa8v_r ;
  MyDTInt_Int_t \call_f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf''''''''_f''''''''_Int_Intop_mapa8w_d ;
  logic \call_f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf''''''''_f''''''''_Int_Intop_mapa8w_r ;
  \Pointer_CTf''''''''_f''''''''_Int_Int_t  \call_f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf''''''''_f''''''''_Int_Intsc_0_1_d ;
  logic \call_f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf''''''''_f''''''''_Int_Intsc_0_1_r ;
  Go_t \call_f''''''''_f''''''''_Int_Int_initBufi_d ;
  logic \call_f''''''''_f''''''''_Int_Int_initBufi_r ;
  C5_t go_11_goMux_choice_d;
  logic go_11_goMux_choice_r;
  Go_t go_11_goMux_data_d;
  logic go_11_goMux_data_r;
  Go_t \call_f''''''''_f''''''''_Int_Int_unlockFork1_d ;
  logic \call_f''''''''_f''''''''_Int_Int_unlockFork1_r ;
  Go_t \call_f''''''''_f''''''''_Int_Int_unlockFork2_d ;
  logic \call_f''''''''_f''''''''_Int_Int_unlockFork2_r ;
  Go_t \call_f''''''''_f''''''''_Int_Int_unlockFork3_d ;
  logic \call_f''''''''_f''''''''_Int_Int_unlockFork3_r ;
  Go_t \call_f''''''''_f''''''''_Int_Int_unlockFork4_d ;
  logic \call_f''''''''_f''''''''_Int_Int_unlockFork4_r ;
  Go_t \call_f''''''''_f''''''''_Int_Int_unlockFork5_d ;
  logic \call_f''''''''_f''''''''_Int_Int_unlockFork5_r ;
  Go_t \call_f''''''''_f''''''''_Int_Int_initBuf_d ;
  logic \call_f''''''''_f''''''''_Int_Int_initBuf_r ;
  Go_t \call_f''''''''_f''''''''_Int_Int_goMux1_d ;
  logic \call_f''''''''_f''''''''_Int_Int_goMux1_r ;
  Pointer_QTree_Int_t \call_f''''''''_f''''''''_Int_Int_goMux2_d ;
  logic \call_f''''''''_f''''''''_Int_Int_goMux2_r ;
  MyDTInt_Bool_t \call_f''''''''_f''''''''_Int_Int_goMux3_d ;
  logic \call_f''''''''_f''''''''_Int_Int_goMux3_r ;
  MyDTInt_Int_t \call_f''''''''_f''''''''_Int_Int_goMux4_d ;
  logic \call_f''''''''_f''''''''_Int_Int_goMux4_r ;
  \Pointer_CTf''''''''_f''''''''_Int_Int_t  \call_f''''''''_f''''''''_Int_Int_goMux5_d ;
  logic \call_f''''''''_f''''''''_Int_Int_goMux5_r ;
  Go_t call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Intgo_12_d;
  logic call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Intgo_12_r;
  Pointer_QTree_Int_t call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Intm1a8C_d;
  logic call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Intm1a8C_r;
  Pointer_QTree_Int_t call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Intm2a8D_d;
  logic call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Intm2a8D_r;
  MyDTInt_Bool_t call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Intis_z_mapa8E_d;
  logic call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Intis_z_mapa8E_r;
  MyDTInt_Int_t call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Intop_mapa8F_d;
  logic call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Intop_mapa8F_r;
  MyDTInt_Bool_t call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Intis_z_adda8G_d;
  logic call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Intis_z_adda8G_r;
  MyDTInt_Int_Int_t call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Intop_adda8H_d;
  logic call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Intop_adda8H_r;
  Pointer_CTf_f_Int_Int_t call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Intsc_0_2_d;
  logic call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Intsc_0_2_r;
  Go_t call_f_f_Int_Int_initBufi_d;
  logic call_f_f_Int_Int_initBufi_r;
  C5_t go_12_goMux_choice_d;
  logic go_12_goMux_choice_r;
  Go_t go_12_goMux_data_d;
  logic go_12_goMux_data_r;
  Go_t call_f_f_Int_Int_unlockFork1_d;
  logic call_f_f_Int_Int_unlockFork1_r;
  Go_t call_f_f_Int_Int_unlockFork2_d;
  logic call_f_f_Int_Int_unlockFork2_r;
  Go_t call_f_f_Int_Int_unlockFork3_d;
  logic call_f_f_Int_Int_unlockFork3_r;
  Go_t call_f_f_Int_Int_unlockFork4_d;
  logic call_f_f_Int_Int_unlockFork4_r;
  Go_t call_f_f_Int_Int_unlockFork5_d;
  logic call_f_f_Int_Int_unlockFork5_r;
  Go_t call_f_f_Int_Int_unlockFork6_d;
  logic call_f_f_Int_Int_unlockFork6_r;
  Go_t call_f_f_Int_Int_unlockFork7_d;
  logic call_f_f_Int_Int_unlockFork7_r;
  Go_t call_f_f_Int_Int_unlockFork8_d;
  logic call_f_f_Int_Int_unlockFork8_r;
  Go_t call_f_f_Int_Int_initBuf_d;
  logic call_f_f_Int_Int_initBuf_r;
  Go_t call_f_f_Int_Int_goMux1_d;
  logic call_f_f_Int_Int_goMux1_r;
  Pointer_QTree_Int_t call_f_f_Int_Int_goMux2_d;
  logic call_f_f_Int_Int_goMux2_r;
  Pointer_QTree_Int_t call_f_f_Int_Int_goMux3_d;
  logic call_f_f_Int_Int_goMux3_r;
  MyDTInt_Bool_t call_f_f_Int_Int_goMux4_d;
  logic call_f_f_Int_Int_goMux4_r;
  MyDTInt_Int_t call_f_f_Int_Int_goMux5_d;
  logic call_f_f_Int_Int_goMux5_r;
  MyDTInt_Bool_t call_f_f_Int_Int_goMux6_d;
  logic call_f_f_Int_Int_goMux6_r;
  MyDTInt_Int_Int_t call_f_f_Int_Int_goMux7_d;
  logic call_f_f_Int_Int_goMux7_r;
  Pointer_CTf_f_Int_Int_t call_f_f_Int_Int_goMux8_d;
  logic call_f_f_Int_Int_goMux8_r;
  Go_t es_10_1MyFalse_d;
  logic es_10_1MyFalse_r;
  Go_t es_10_1MyTrue_d;
  logic es_10_1MyTrue_r;
  Go_t es_10_1MyFalse_1_d;
  logic es_10_1MyFalse_1_r;
  Go_t es_10_1MyFalse_2_d;
  logic es_10_1MyFalse_2_r;
  Go_t es_10_1MyFalse_1_argbuf_d;
  logic es_10_1MyFalse_1_argbuf_r;
  TupGo___MyDTInt_Int___Int_t applyfnInt_Int_5TupGo___MyDTInt_Int___Int6_d;
  logic applyfnInt_Int_5TupGo___MyDTInt_Int___Int6_r;
  Go_t es_10_1MyFalse_2_argbuf_d;
  logic es_10_1MyFalse_2_argbuf_r;
  Go_t es_10_1MyTrue_1_d;
  logic es_10_1MyTrue_1_r;
  Go_t es_10_1MyTrue_2_d;
  logic es_10_1MyTrue_2_r;
  QTree_Int_t es_10_1MyTrue_1QNone_Int_d;
  logic es_10_1MyTrue_1QNone_Int_r;
  QTree_Int_t lizzieLet21_1_argbuf_d;
  logic lizzieLet21_1_argbuf_r;
  Go_t es_10_1MyTrue_2_argbuf_d;
  logic es_10_1MyTrue_2_argbuf_r;
  MyDTInt_Int_t es_10_2MyFalse_d;
  logic es_10_2MyFalse_r;
  MyDTInt_Int_t _80_d;
  logic _80_r;
  assign _80_r = 1'd1;
  MyDTInt_Int_t es_10_2MyFalse_1_argbuf_d;
  logic es_10_2MyFalse_1_argbuf_r;
  Pointer_CTf_f_Int_Int_t es_10_3MyFalse_d;
  logic es_10_3MyFalse_r;
  Pointer_CTf_f_Int_Int_t es_10_3MyTrue_d;
  logic es_10_3MyTrue_r;
  Pointer_CTf_f_Int_Int_t es_10_3MyFalse_1_argbuf_d;
  logic es_10_3MyFalse_1_argbuf_r;
  Pointer_CTf_f_Int_Int_t es_10_3MyTrue_1_argbuf_d;
  logic es_10_3MyTrue_1_argbuf_r;
  Int_t es_10_4MyFalse_d;
  logic es_10_4MyFalse_r;
  Int_t _79_d;
  logic _79_r;
  assign _79_r = 1'd1;
  Int_t es_10_4MyFalse_1_argbuf_d;
  logic es_10_4MyFalse_1_argbuf_r;
  QTree_Int_t lizzieLet20_1_argbuf_d;
  logic lizzieLet20_1_argbuf_r;
  Go_t es_14_1MyFalse_d;
  logic es_14_1MyFalse_r;
  Go_t es_14_1MyTrue_d;
  logic es_14_1MyTrue_r;
  Go_t es_14_1MyFalse_1_d;
  logic es_14_1MyFalse_1_r;
  Go_t es_14_1MyFalse_2_d;
  logic es_14_1MyFalse_2_r;
  Go_t es_14_1MyFalse_3_d;
  logic es_14_1MyFalse_3_r;
  Go_t es_14_1MyFalse_1_argbuf_d;
  logic es_14_1MyFalse_1_argbuf_r;
  TupGo___MyDTInt_Int___Int_t applyfnInt_Int_5TupGo___MyDTInt_Int___Int7_d;
  logic applyfnInt_Int_5TupGo___MyDTInt_Int___Int7_r;
  Go_t es_14_1MyFalse_2_argbuf_d;
  logic es_14_1MyFalse_2_argbuf_r;
  TupGo___MyDTInt_Bool___Int_t applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int5_d;
  logic applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int5_r;
  Go_t es_14_1MyTrue_1_d;
  logic es_14_1MyTrue_1_r;
  Go_t es_14_1MyTrue_2_d;
  logic es_14_1MyTrue_2_r;
  QTree_Int_t es_14_1MyTrue_1QNone_Int_d;
  logic es_14_1MyTrue_1QNone_Int_r;
  QTree_Int_t lizzieLet24_1_1_argbuf_d;
  logic lizzieLet24_1_1_argbuf_r;
  Go_t es_14_1MyTrue_2_argbuf_d;
  logic es_14_1MyTrue_2_argbuf_r;
  MyDTInt_Bool_t es_14_2MyFalse_d;
  logic es_14_2MyFalse_r;
  MyDTInt_Bool_t _78_d;
  logic _78_r;
  assign _78_r = 1'd1;
  MyDTInt_Bool_t es_14_2MyFalse_1_argbuf_d;
  logic es_14_2MyFalse_1_argbuf_r;
  MyDTInt_Int_Int_t es_14_3MyFalse_d;
  logic es_14_3MyFalse_r;
  MyDTInt_Int_Int_t _77_d;
  logic _77_r;
  assign _77_r = 1'd1;
  MyDTInt_Int_Int_t es_14_3MyFalse_1_d;
  logic es_14_3MyFalse_1_r;
  MyDTInt_Int_Int_t es_14_3MyFalse_2_d;
  logic es_14_3MyFalse_2_r;
  MyDTInt_Int_Int_t es_14_3MyFalse_1_argbuf_d;
  logic es_14_3MyFalse_1_argbuf_r;
  TupMyDTInt_Int_Int___Int___Int_t applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int2_d;
  logic applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int2_r;
  MyDTInt_Int_t es_14_4MyFalse_d;
  logic es_14_4MyFalse_r;
  MyDTInt_Int_t _76_d;
  logic _76_r;
  assign _76_r = 1'd1;
  MyDTInt_Int_t es_14_4MyFalse_1_d;
  logic es_14_4MyFalse_1_r;
  MyDTInt_Int_t es_14_4MyFalse_2_d;
  logic es_14_4MyFalse_2_r;
  MyDTInt_Int_t es_14_4MyFalse_1_argbuf_d;
  logic es_14_4MyFalse_1_argbuf_r;
  Pointer_CTf_f_Int_Int_t es_14_5MyFalse_d;
  logic es_14_5MyFalse_r;
  Pointer_CTf_f_Int_Int_t es_14_5MyTrue_d;
  logic es_14_5MyTrue_r;
  Pointer_CTf_f_Int_Int_t es_14_5MyTrue_1_argbuf_d;
  logic es_14_5MyTrue_1_argbuf_r;
  Int_t es_14_6MyFalse_d;
  logic es_14_6MyFalse_r;
  Int_t _75_d;
  logic _75_r;
  assign _75_r = 1'd1;
  Int_t es_14_6MyFalse_1_d;
  logic es_14_6MyFalse_1_r;
  Int_t es_14_6MyFalse_2_d;
  logic es_14_6MyFalse_2_r;
  Int_t es_14_6MyFalse_1_argbuf_d;
  logic es_14_6MyFalse_1_argbuf_r;
  Int_t es_14_7MyFalse_d;
  logic es_14_7MyFalse_r;
  Int_t _74_d;
  logic _74_r;
  assign _74_r = 1'd1;
  Int_t es_14_7MyFalse_1_d;
  logic es_14_7MyFalse_1_r;
  Int_t es_14_7MyFalse_2_d;
  logic es_14_7MyFalse_2_r;
  Int_t es_14_7MyFalse_1_argbuf_d;
  logic es_14_7MyFalse_1_argbuf_r;
  Go_t es_19_1MyFalse_d;
  logic es_19_1MyFalse_r;
  Go_t es_19_1MyTrue_d;
  logic es_19_1MyTrue_r;
  Go_t es_19_1MyFalse_1_d;
  logic es_19_1MyFalse_1_r;
  Go_t es_19_1MyFalse_2_d;
  logic es_19_1MyFalse_2_r;
  Go_t es_19_1MyFalse_1_argbuf_d;
  logic es_19_1MyFalse_1_argbuf_r;
  TupGo___MyDTInt_Int___Int_t applyfnInt_Int_5TupGo___MyDTInt_Int___Int8_d;
  logic applyfnInt_Int_5TupGo___MyDTInt_Int___Int8_r;
  Go_t es_19_1MyFalse_2_argbuf_d;
  logic es_19_1MyFalse_2_argbuf_r;
  Go_t es_19_1MyTrue_1_d;
  logic es_19_1MyTrue_1_r;
  Go_t es_19_1MyTrue_2_d;
  logic es_19_1MyTrue_2_r;
  QTree_Int_t es_19_1MyTrue_1QNone_Int_d;
  logic es_19_1MyTrue_1QNone_Int_r;
  QTree_Int_t lizzieLet23_2_1_argbuf_d;
  logic lizzieLet23_2_1_argbuf_r;
  Go_t es_19_1MyTrue_2_argbuf_d;
  logic es_19_1MyTrue_2_argbuf_r;
  MyDTInt_Int_Int_t es_19_2MyFalse_d;
  logic es_19_2MyFalse_r;
  MyDTInt_Int_Int_t _73_d;
  logic _73_r;
  assign _73_r = 1'd1;
  MyDTInt_Int_Int_t es_19_2MyFalse_1_argbuf_d;
  logic es_19_2MyFalse_1_argbuf_r;
  TupMyDTInt_Int_Int___Int___Int_t applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int3_d;
  logic applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int3_r;
  MyDTInt_Int_t es_19_3MyFalse_d;
  logic es_19_3MyFalse_r;
  MyDTInt_Int_t _72_d;
  logic _72_r;
  assign _72_r = 1'd1;
  MyDTInt_Int_t es_19_3MyFalse_1_argbuf_d;
  logic es_19_3MyFalse_1_argbuf_r;
  Pointer_CTf_f_Int_Int_t es_19_4MyFalse_d;
  logic es_19_4MyFalse_r;
  Pointer_CTf_f_Int_Int_t es_19_4MyTrue_d;
  logic es_19_4MyTrue_r;
  Pointer_CTf_f_Int_Int_t es_19_4MyFalse_1_argbuf_d;
  logic es_19_4MyFalse_1_argbuf_r;
  Pointer_CTf_f_Int_Int_t es_19_4MyTrue_1_argbuf_d;
  logic es_19_4MyTrue_1_argbuf_r;
  Int_t es_19_5MyFalse_d;
  logic es_19_5MyFalse_r;
  Int_t _71_d;
  logic _71_r;
  assign _71_r = 1'd1;
  Int_t es_19_5MyFalse_1_argbuf_d;
  logic es_19_5MyFalse_1_argbuf_r;
  Int_t es_19_6MyFalse_d;
  logic es_19_6MyFalse_r;
  Int_t _70_d;
  logic _70_r;
  assign _70_r = 1'd1;
  Int_t es_19_6MyFalse_1_argbuf_d;
  logic es_19_6MyFalse_1_argbuf_r;
  QTree_Int_t lizzieLet22_1_argbuf_d;
  logic lizzieLet22_1_argbuf_r;
  QTree_Int_t lizzieLet28_1_argbuf_d;
  logic lizzieLet28_1_argbuf_r;
  Go_t es_2_1MyFalse_d;
  logic es_2_1MyFalse_r;
  Go_t es_2_1MyTrue_d;
  logic es_2_1MyTrue_r;
  Go_t es_2_1MyFalse_1_d;
  logic es_2_1MyFalse_1_r;
  Go_t es_2_1MyFalse_2_d;
  logic es_2_1MyFalse_2_r;
  Go_t es_2_1MyFalse_1_argbuf_d;
  logic es_2_1MyFalse_1_argbuf_r;
  TupGo___MyDTInt_Int___Int_t applyfnInt_Int_5TupGo___MyDTInt_Int___Int4_d;
  logic applyfnInt_Int_5TupGo___MyDTInt_Int___Int4_r;
  Go_t es_2_1MyFalse_2_argbuf_d;
  logic es_2_1MyFalse_2_argbuf_r;
  Go_t es_2_1MyTrue_1_d;
  logic es_2_1MyTrue_1_r;
  Go_t es_2_1MyTrue_2_d;
  logic es_2_1MyTrue_2_r;
  QTree_Int_t es_2_1MyTrue_1QNone_Int_d;
  logic es_2_1MyTrue_1QNone_Int_r;
  QTree_Int_t lizzieLet9_1_argbuf_d;
  logic lizzieLet9_1_argbuf_r;
  Go_t es_2_1MyTrue_2_argbuf_d;
  logic es_2_1MyTrue_2_argbuf_r;
  Go_t es_2_1_1MyFalse_d;
  logic es_2_1_1MyFalse_r;
  Go_t es_2_1_1MyTrue_d;
  logic es_2_1_1MyTrue_r;
  Go_t es_2_1_1MyFalse_1_d;
  logic es_2_1_1MyFalse_1_r;
  Go_t es_2_1_1MyFalse_2_d;
  logic es_2_1_1MyFalse_2_r;
  Go_t es_2_1_1MyFalse_1_argbuf_d;
  logic es_2_1_1MyFalse_1_argbuf_r;
  TupGo___MyDTInt_Int___Int_t applyfnInt_Int_5TupGo___MyDTInt_Int___Int2_d;
  logic applyfnInt_Int_5TupGo___MyDTInt_Int___Int2_r;
  Go_t es_2_1_1MyFalse_2_argbuf_d;
  logic es_2_1_1MyFalse_2_argbuf_r;
  Go_t es_2_1_1MyTrue_1_d;
  logic es_2_1_1MyTrue_1_r;
  Go_t es_2_1_1MyTrue_2_d;
  logic es_2_1_1MyTrue_2_r;
  QTree_Int_t es_2_1_1MyTrue_1QNone_Int_d;
  logic es_2_1_1MyTrue_1QNone_Int_r;
  QTree_Int_t lizzieLet16_1_argbuf_d;
  logic lizzieLet16_1_argbuf_r;
  Go_t es_2_1_1MyTrue_2_argbuf_d;
  logic es_2_1_1MyTrue_2_argbuf_r;
  MyDTInt_Int_t es_2_1_2MyFalse_d;
  logic es_2_1_2MyFalse_r;
  MyDTInt_Int_t _69_d;
  logic _69_r;
  assign _69_r = 1'd1;
  MyDTInt_Int_t es_2_1_2MyFalse_1_argbuf_d;
  logic es_2_1_2MyFalse_1_argbuf_r;
  Pointer_CTf_f_Int_Int_t es_2_1_3MyFalse_d;
  logic es_2_1_3MyFalse_r;
  Pointer_CTf_f_Int_Int_t es_2_1_3MyTrue_d;
  logic es_2_1_3MyTrue_r;
  Pointer_CTf_f_Int_Int_t es_2_1_3MyFalse_1_argbuf_d;
  logic es_2_1_3MyFalse_1_argbuf_r;
  Pointer_CTf_f_Int_Int_t es_2_1_3MyTrue_1_argbuf_d;
  logic es_2_1_3MyTrue_1_argbuf_r;
  Int_t es_2_1_4MyFalse_d;
  logic es_2_1_4MyFalse_r;
  Int_t _68_d;
  logic _68_r;
  assign _68_r = 1'd1;
  Int_t es_2_1_4MyFalse_1_argbuf_d;
  logic es_2_1_4MyFalse_1_argbuf_r;
  MyDTInt_Int_t es_2_2MyFalse_d;
  logic es_2_2MyFalse_r;
  MyDTInt_Int_t _67_d;
  logic _67_r;
  assign _67_r = 1'd1;
  MyDTInt_Int_t es_2_2MyFalse_1_argbuf_d;
  logic es_2_2MyFalse_1_argbuf_r;
  \Pointer_CTf''''''''_f''''''''_Int_Int_t  es_2_3MyFalse_d;
  logic es_2_3MyFalse_r;
  \Pointer_CTf''''''''_f''''''''_Int_Int_t  es_2_3MyTrue_d;
  logic es_2_3MyTrue_r;
  \Pointer_CTf''''''''_f''''''''_Int_Int_t  es_2_3MyFalse_1_argbuf_d;
  logic es_2_3MyFalse_1_argbuf_r;
  \Pointer_CTf''''''''_f''''''''_Int_Int_t  es_2_3MyTrue_1_argbuf_d;
  logic es_2_3MyTrue_1_argbuf_r;
  Int_t es_2_4MyFalse_d;
  logic es_2_4MyFalse_r;
  Int_t _66_d;
  logic _66_r;
  assign _66_r = 1'd1;
  Int_t es_2_4MyFalse_1_argbuf_d;
  logic es_2_4MyFalse_1_argbuf_r;
  QTree_Int_t lizzieLet8_1_argbuf_d;
  logic lizzieLet8_1_argbuf_r;
  QTree_Int_t lizzieLet15_1_argbuf_d;
  logic lizzieLet15_1_argbuf_r;
  QTree_Int_t lizzieLet17_1_argbuf_d;
  logic lizzieLet17_1_argbuf_r;
  \Int#_t  contRet_0_1_argbuf_d;
  logic contRet_0_1_argbuf_r;
  \Int#_t  es_4_2_1lizzieLet35_4Lcall_$wnnz0_1_Add32_d;
  logic es_4_2_1lizzieLet35_4Lcall_$wnnz0_1_Add32_r;
  C8_t \f''''''''_f''''''''_Int_Int_choice_d ;
  logic \f''''''''_f''''''''_Int_Int_choice_r ;
  TupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_t \f''''''''_f''''''''_Int_Int_data_d ;
  logic \f''''''''_f''''''''_Int_Int_data_r ;
  Go_t go_13_1_d;
  logic go_13_1_r;
  Go_t go_13_2_d;
  logic go_13_2_r;
  MyDTInt_Bool_t is_z_mapa8v_1_1_argbuf_d;
  logic is_z_mapa8v_1_1_argbuf_r;
  MyDTInt_Int_t op_mapa8w_1_1_argbuf_d;
  logic op_mapa8w_1_1_argbuf_r;
  Pointer_QTree_Int_t q4a8u_1_1_argbuf_d;
  logic q4a8u_1_1_argbuf_r;
  Pointer_QTree_Int_t \f''''''''_f''''''''_Int_Int_resbuf_d ;
  logic \f''''''''_f''''''''_Int_Int_resbuf_r ;
  Pointer_QTree_Int_t \f''''''''_f''''''''_Int_Int_2_argbuf_d ;
  logic \f''''''''_f''''''''_Int_Int_2_argbuf_r ;
  Pointer_QTree_Int_t \f''''''''_f''''''''_Int_Int_3_argbuf_d ;
  logic \f''''''''_f''''''''_Int_Int_3_argbuf_r ;
  Pointer_QTree_Int_t \f''''''''_f''''''''_Int_Int_4_argbuf_d ;
  logic \f''''''''_f''''''''_Int_Int_4_argbuf_r ;
  QTree_Int_t es_4_1_1es_5_1_1es_6_1_1es_7_1_1QNode_Int_d;
  logic es_4_1_1es_5_1_1es_6_1_1es_7_1_1QNode_Int_r;
  Pointer_QTree_Int_t \f''''''''_f''''''''_Int_Int_5_argbuf_d ;
  logic \f''''''''_f''''''''_Int_Int_5_argbuf_r ;
  Pointer_QTree_Int_t \f''''''''_f''''''''_Int_Int_6_argbuf_d ;
  logic \f''''''''_f''''''''_Int_Int_6_argbuf_r ;
  Pointer_QTree_Int_t \f''''''''_f''''''''_Int_Int_7_argbuf_d ;
  logic \f''''''''_f''''''''_Int_Int_7_argbuf_r ;
  Pointer_QTree_Int_t \f''''''''_f''''''''_Int_Int_8_argbuf_d ;
  logic \f''''''''_f''''''''_Int_Int_8_argbuf_r ;
  QTree_Int_t es_23_1es_24_1es_25_1es_26_1QNode_Int_d;
  logic es_23_1es_24_1es_25_1es_26_1QNode_Int_r;
  Pointer_QTree_Int_t \f''''''''_f''''''''_Int_Int_1_d ;
  logic \f''''''''_f''''''''_Int_Int_1_r ;
  Pointer_QTree_Int_t \f''''''''_f''''''''_Int_Int_2_d ;
  logic \f''''''''_f''''''''_Int_Int_2_r ;
  Pointer_QTree_Int_t \f''''''''_f''''''''_Int_Int_3_d ;
  logic \f''''''''_f''''''''_Int_Int_3_r ;
  Pointer_QTree_Int_t \f''''''''_f''''''''_Int_Int_4_d ;
  logic \f''''''''_f''''''''_Int_Int_4_r ;
  Pointer_QTree_Int_t \f''''''''_f''''''''_Int_Int_5_d ;
  logic \f''''''''_f''''''''_Int_Int_5_r ;
  Pointer_QTree_Int_t \f''''''''_f''''''''_Int_Int_6_d ;
  logic \f''''''''_f''''''''_Int_Int_6_r ;
  Pointer_QTree_Int_t \f''''''''_f''''''''_Int_Int_7_d ;
  logic \f''''''''_f''''''''_Int_Int_7_r ;
  Pointer_QTree_Int_t \f''''''''_f''''''''_Int_Int_8_d ;
  logic \f''''''''_f''''''''_Int_Int_8_r ;
  Go_t \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Intgo_13_d ;
  logic \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Intgo_13_r ;
  Pointer_QTree_Int_t \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Intq4a8u_1_d ;
  logic \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Intq4a8u_1_r ;
  MyDTInt_Bool_t \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Intis_z_mapa8v_1_d ;
  logic \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Intis_z_mapa8v_1_r ;
  MyDTInt_Int_t \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Intop_mapa8w_1_d ;
  logic \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Intop_mapa8w_1_r ;
  Go_t f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intgo_14_d;
  logic f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intgo_14_r;
  Pointer_QTree_Int_t f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intm1a8C_1_d;
  logic f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intm1a8C_1_r;
  Pointer_QTree_Int_t f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intm2a8D_1_d;
  logic f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intm2a8D_1_r;
  MyDTInt_Bool_t f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intis_z_mapa8E_1_d;
  logic f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intis_z_mapa8E_1_r;
  MyDTInt_Int_t f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intop_mapa8F_1_d;
  logic f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intop_mapa8F_1_r;
  MyDTInt_Bool_t f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intis_z_adda8G_1_d;
  logic f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intis_z_adda8G_1_r;
  MyDTInt_Int_Int_t f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intop_adda8H_1_d;
  logic f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intop_adda8H_1_r;
  Go_t go_14_1_d;
  logic go_14_1_r;
  Go_t go_14_2_d;
  logic go_14_2_r;
  MyDTInt_Bool_t is_z_adda8G_1_1_argbuf_d;
  logic is_z_adda8G_1_1_argbuf_r;
  MyDTInt_Bool_t is_z_mapa8E_1_1_argbuf_d;
  logic is_z_mapa8E_1_1_argbuf_r;
  Pointer_QTree_Int_t m1a8C_1_1_argbuf_d;
  logic m1a8C_1_1_argbuf_r;
  Pointer_QTree_Int_t m2a8D_1_1_argbuf_d;
  logic m2a8D_1_1_argbuf_r;
  MyDTInt_Int_Int_t op_adda8H_1_1_argbuf_d;
  logic op_adda8H_1_1_argbuf_r;
  MyDTInt_Int_t op_mapa8F_1_1_argbuf_d;
  logic op_mapa8F_1_1_argbuf_r;
  Pointer_QTree_Int_t es_0_1_argbuf_d;
  logic es_0_1_argbuf_r;
  MyDTInt_Int_Int_t \go_1Dcon_$fNumInt_$c+_d ;
  logic \go_1Dcon_$fNumInt_$c+_r ;
  C5_t go_10_goMux_choice_1_d;
  logic go_10_goMux_choice_1_r;
  C5_t go_10_goMux_choice_2_d;
  logic go_10_goMux_choice_2_r;
  Pointer_QTree_Int_t wsiX_1_goMux_mux_d;
  logic wsiX_1_goMux_mux_r;
  Pointer_CT$wnnz_t sc_0_goMux_mux_d;
  logic sc_0_goMux_mux_r;
  C5_t go_11_goMux_choice_1_d;
  logic go_11_goMux_choice_1_r;
  C5_t go_11_goMux_choice_2_d;
  logic go_11_goMux_choice_2_r;
  C5_t go_11_goMux_choice_3_d;
  logic go_11_goMux_choice_3_r;
  C5_t go_11_goMux_choice_4_d;
  logic go_11_goMux_choice_4_r;
  Pointer_QTree_Int_t q4a8u_goMux_mux_d;
  logic q4a8u_goMux_mux_r;
  MyDTInt_Bool_t is_z_mapa8v_goMux_mux_d;
  logic is_z_mapa8v_goMux_mux_r;
  MyDTInt_Int_t op_mapa8w_goMux_mux_d;
  logic op_mapa8w_goMux_mux_r;
  \Pointer_CTf''''''''_f''''''''_Int_Int_t  sc_0_1_goMux_mux_d;
  logic sc_0_1_goMux_mux_r;
  C5_t go_12_goMux_choice_1_d;
  logic go_12_goMux_choice_1_r;
  C5_t go_12_goMux_choice_2_d;
  logic go_12_goMux_choice_2_r;
  C5_t go_12_goMux_choice_3_d;
  logic go_12_goMux_choice_3_r;
  C5_t go_12_goMux_choice_4_d;
  logic go_12_goMux_choice_4_r;
  C5_t go_12_goMux_choice_5_d;
  logic go_12_goMux_choice_5_r;
  C5_t go_12_goMux_choice_6_d;
  logic go_12_goMux_choice_6_r;
  C5_t go_12_goMux_choice_7_d;
  logic go_12_goMux_choice_7_r;
  Pointer_QTree_Int_t m1a8C_goMux_mux_d;
  logic m1a8C_goMux_mux_r;
  Pointer_QTree_Int_t m2a8D_goMux_mux_d;
  logic m2a8D_goMux_mux_r;
  MyDTInt_Bool_t is_z_mapa8E_goMux_mux_d;
  logic is_z_mapa8E_goMux_mux_r;
  MyDTInt_Int_t op_mapa8F_goMux_mux_d;
  logic op_mapa8F_goMux_mux_r;
  MyDTInt_Bool_t is_z_adda8G_goMux_mux_d;
  logic is_z_adda8G_goMux_mux_r;
  MyDTInt_Int_Int_t op_adda8H_goMux_mux_d;
  logic op_adda8H_goMux_mux_r;
  Pointer_CTf_f_Int_Int_t sc_0_2_goMux_mux_d;
  logic sc_0_2_goMux_mux_r;
  \CTf''''''''_f''''''''_Int_Int_t  \go_13_1Lf''''''''_f''''''''_Int_Intsbos_d ;
  logic \go_13_1Lf''''''''_f''''''''_Int_Intsbos_r ;
  \CTf''''''''_f''''''''_Int_Int_t  lizzieLet33_1_argbuf_d;
  logic lizzieLet33_1_argbuf_r;
  Go_t go_13_2_argbuf_d;
  logic go_13_2_argbuf_r;
  \TupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf''''''''_f''''''''_Int_Int_t  \call_f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf''''''''_f''''''''_Int_Int_1_d ;
  logic \call_f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf''''''''_f''''''''_Int_Int_1_r ;
  CTf_f_Int_Int_t go_14_1Lf_f_Int_Intsbos_d;
  logic go_14_1Lf_f_Int_Intsbos_r;
  CTf_f_Int_Int_t lizzieLet34_1_argbuf_d;
  logic lizzieLet34_1_argbuf_r;
  Go_t go_14_2_argbuf_d;
  logic go_14_2_argbuf_r;
  TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Int_t call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Int_1_d;
  logic call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Int_1_r;
  C4_t go_15_goMux_choice_1_d;
  logic go_15_goMux_choice_1_r;
  C4_t go_15_goMux_choice_2_d;
  logic go_15_goMux_choice_2_r;
  \Int#_t  srtarg_0_goMux_mux_d;
  logic srtarg_0_goMux_mux_r;
  Pointer_CT$wnnz_t scfarg_0_goMux_mux_d;
  logic scfarg_0_goMux_mux_r;
  C5_t go_16_goMux_choice_1_d;
  logic go_16_goMux_choice_1_r;
  C5_t go_16_goMux_choice_2_d;
  logic go_16_goMux_choice_2_r;
  Pointer_QTree_Int_t srtarg_0_1_goMux_mux_d;
  logic srtarg_0_1_goMux_mux_r;
  \Pointer_CTf''''''''_f''''''''_Int_Int_t  scfarg_0_1_goMux_mux_d;
  logic scfarg_0_1_goMux_mux_r;
  C17_t go_17_goMux_choice_1_d;
  logic go_17_goMux_choice_1_r;
  C17_t go_17_goMux_choice_2_d;
  logic go_17_goMux_choice_2_r;
  Pointer_QTree_Int_t srtarg_0_2_goMux_mux_d;
  logic srtarg_0_2_goMux_mux_r;
  Pointer_CTf_f_Int_Int_t scfarg_0_2_goMux_mux_d;
  logic scfarg_0_2_goMux_mux_r;
  MyDTInt_Int_Int_t es_6_1_argbuf_d;
  logic es_6_1_argbuf_r;
  MyDTInt_Bool_t go_2Dcon_is_z_1_d;
  logic go_2Dcon_is_z_1_r;
  MyDTInt_Bool_t es_5_1_argbuf_d;
  logic es_5_1_argbuf_r;
  MyDTInt_Int_t go_3Dcon_main1_d;
  logic go_3Dcon_main1_r;
  MyDTInt_Int_t es_4_1_argbuf_d;
  logic es_4_1_argbuf_r;
  MyDTInt_Bool_t go_4Dcon_is_z_1_d;
  logic go_4Dcon_is_z_1_r;
  MyDTInt_Bool_t es_3_1_argbuf_d;
  logic es_3_1_argbuf_r;
  Go_t go_5_argbuf_d;
  logic go_5_argbuf_r;
  TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int_t f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_d;
  logic f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_r;
  Go_t go_6_argbuf_d;
  logic go_6_argbuf_r;
  TupGo___Pointer_QTree_Int_t \$wnnzTupGo___Pointer_QTree_Int_1_d ;
  logic \$wnnzTupGo___Pointer_QTree_Int_1_r ;
  CT$wnnz_t go_7_1L$wnnzsbos_d;
  logic go_7_1L$wnnzsbos_r;
  CT$wnnz_t lizzieLet0_1_argbuf_d;
  logic lizzieLet0_1_argbuf_r;
  Go_t go_7_2_argbuf_d;
  logic go_7_2_argbuf_r;
  TupGo___Pointer_QTree_Int___Pointer_CT$wnnz_t call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_1_d;
  logic call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_1_r;
  MyDTInt_Bool_t is_z_adda8G_2_2_argbuf_d;
  logic is_z_adda8G_2_2_argbuf_r;
  MyDTInt_Bool_t is_z_adda8G_2_1_d;
  logic is_z_adda8G_2_1_r;
  MyDTInt_Bool_t is_z_adda8G_2_2_d;
  logic is_z_adda8G_2_2_r;
  MyDTInt_Bool_t is_z_adda8G_3_2_argbuf_d;
  logic is_z_adda8G_3_2_argbuf_r;
  MyDTInt_Bool_t is_z_adda8G_3_1_d;
  logic is_z_adda8G_3_1_r;
  MyDTInt_Bool_t is_z_adda8G_3_2_d;
  logic is_z_adda8G_3_2_r;
  MyDTInt_Bool_t is_z_adda8G_4_1_argbuf_d;
  logic is_z_adda8G_4_1_argbuf_r;
  MyDTInt_Bool_t is_z_mapa8E_2_2_argbuf_d;
  logic is_z_mapa8E_2_2_argbuf_r;
  MyDTInt_Bool_t is_z_mapa8E_2_1_d;
  logic is_z_mapa8E_2_1_r;
  MyDTInt_Bool_t is_z_mapa8E_2_2_d;
  logic is_z_mapa8E_2_2_r;
  MyDTInt_Bool_t is_z_mapa8E_3_2_argbuf_d;
  logic is_z_mapa8E_3_2_argbuf_r;
  MyDTInt_Bool_t is_z_mapa8E_3_1_d;
  logic is_z_mapa8E_3_1_r;
  MyDTInt_Bool_t is_z_mapa8E_3_2_d;
  logic is_z_mapa8E_3_2_r;
  MyDTInt_Bool_t is_z_mapa8E_4_1_argbuf_d;
  logic is_z_mapa8E_4_1_argbuf_r;
  MyDTInt_Bool_t is_z_mapa8v_2_2_argbuf_d;
  logic is_z_mapa8v_2_2_argbuf_r;
  MyDTInt_Bool_t is_z_mapa8v_2_1_d;
  logic is_z_mapa8v_2_1_r;
  MyDTInt_Bool_t is_z_mapa8v_2_2_d;
  logic is_z_mapa8v_2_2_r;
  MyDTInt_Bool_t is_z_mapa8v_3_2_argbuf_d;
  logic is_z_mapa8v_3_2_argbuf_r;
  MyDTInt_Bool_t is_z_mapa8v_3_1_d;
  logic is_z_mapa8v_3_1_r;
  MyDTInt_Bool_t is_z_mapa8v_3_2_d;
  logic is_z_mapa8v_3_2_r;
  MyDTInt_Bool_t is_z_mapa8v_4_1_argbuf_d;
  logic is_z_mapa8v_4_1_argbuf_r;
  Pointer_QTree_Int_t q1a8T_destruct_d;
  logic q1a8T_destruct_r;
  Pointer_QTree_Int_t q2a8U_destruct_d;
  logic q2a8U_destruct_r;
  Pointer_QTree_Int_t q3a8V_destruct_d;
  logic q3a8V_destruct_r;
  Pointer_QTree_Int_t q4a8W_destruct_d;
  logic q4a8W_destruct_r;
  Int_t v1a8N_destruct_d;
  logic v1a8N_destruct_r;
  QTree_Int_t _65_d;
  logic _65_r;
  assign _65_r = 1'd1;
  QTree_Int_t lizzieLet12_1QVal_Int_d;
  logic lizzieLet12_1QVal_Int_r;
  QTree_Int_t lizzieLet12_1QNode_Int_d;
  logic lizzieLet12_1QNode_Int_r;
  QTree_Int_t _64_d;
  logic _64_r;
  assign _64_r = 1'd1;
  Go_t lizzieLet12_3QNone_Int_d;
  logic lizzieLet12_3QNone_Int_r;
  Go_t lizzieLet12_3QVal_Int_d;
  logic lizzieLet12_3QVal_Int_r;
  Go_t lizzieLet12_3QNode_Int_d;
  logic lizzieLet12_3QNode_Int_r;
  Go_t lizzieLet12_3QError_Int_d;
  logic lizzieLet12_3QError_Int_r;
  Go_t lizzieLet12_3QError_Int_1_d;
  logic lizzieLet12_3QError_Int_1_r;
  Go_t lizzieLet12_3QError_Int_2_d;
  logic lizzieLet12_3QError_Int_2_r;
  QTree_Int_t lizzieLet12_3QError_Int_1QError_Int_d;
  logic lizzieLet12_3QError_Int_1QError_Int_r;
  QTree_Int_t lizzieLet32_1_argbuf_d;
  logic lizzieLet32_1_argbuf_r;
  Go_t lizzieLet12_3QError_Int_2_argbuf_d;
  logic lizzieLet12_3QError_Int_2_argbuf_r;
  MyDTInt_Bool_t _63_d;
  logic _63_r;
  assign _63_r = 1'd1;
  MyDTInt_Bool_t lizzieLet12_4QVal_Int_d;
  logic lizzieLet12_4QVal_Int_r;
  MyDTInt_Bool_t lizzieLet12_4QNode_Int_d;
  logic lizzieLet12_4QNode_Int_r;
  MyDTInt_Bool_t _62_d;
  logic _62_r;
  assign _62_r = 1'd1;
  MyDTInt_Bool_t lizzieLet12_5QNone_Int_d;
  logic lizzieLet12_5QNone_Int_r;
  MyDTInt_Bool_t lizzieLet12_5QVal_Int_d;
  logic lizzieLet12_5QVal_Int_r;
  MyDTInt_Bool_t lizzieLet12_5QNode_Int_d;
  logic lizzieLet12_5QNode_Int_r;
  MyDTInt_Bool_t _61_d;
  logic _61_r;
  assign _61_r = 1'd1;
  QTree_Int_t lizzieLet12_6QNone_Int_d;
  logic lizzieLet12_6QNone_Int_r;
  QTree_Int_t lizzieLet12_6QVal_Int_d;
  logic lizzieLet12_6QVal_Int_r;
  QTree_Int_t lizzieLet12_6QNode_Int_d;
  logic lizzieLet12_6QNode_Int_r;
  QTree_Int_t _60_d;
  logic _60_r;
  assign _60_r = 1'd1;
  QTree_Int_t lizzieLet12_6QNode_Int_1_d;
  logic lizzieLet12_6QNode_Int_1_r;
  QTree_Int_t lizzieLet12_6QNode_Int_2_d;
  logic lizzieLet12_6QNode_Int_2_r;
  QTree_Int_t lizzieLet12_6QNode_Int_3_d;
  logic lizzieLet12_6QNode_Int_3_r;
  QTree_Int_t lizzieLet12_6QNode_Int_4_d;
  logic lizzieLet12_6QNode_Int_4_r;
  QTree_Int_t lizzieLet12_6QNode_Int_5_d;
  logic lizzieLet12_6QNode_Int_5_r;
  QTree_Int_t lizzieLet12_6QNode_Int_6_d;
  logic lizzieLet12_6QNode_Int_6_r;
  QTree_Int_t lizzieLet12_6QNode_Int_7_d;
  logic lizzieLet12_6QNode_Int_7_r;
  QTree_Int_t lizzieLet12_6QNode_Int_8_d;
  logic lizzieLet12_6QNode_Int_8_r;
  QTree_Int_t lizzieLet12_6QNode_Int_9_d;
  logic lizzieLet12_6QNode_Int_9_r;
  QTree_Int_t lizzieLet12_6QNode_Int_10_d;
  logic lizzieLet12_6QNode_Int_10_r;
  QTree_Int_t lizzieLet12_6QNode_Int_11_d;
  logic lizzieLet12_6QNode_Int_11_r;
  QTree_Int_t lizzieLet12_6QNode_Int_12_d;
  logic lizzieLet12_6QNode_Int_12_r;
  Pointer_QTree_Int_t lizzieLet12_6QNode_Int_10QNone_Int_d;
  logic lizzieLet12_6QNode_Int_10QNone_Int_r;
  Pointer_QTree_Int_t _59_d;
  logic _59_r;
  assign _59_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet12_6QNode_Int_10QNode_Int_d;
  logic lizzieLet12_6QNode_Int_10QNode_Int_r;
  Pointer_QTree_Int_t _58_d;
  logic _58_r;
  assign _58_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet12_6QNode_Int_10QNone_Int_1_argbuf_d;
  logic lizzieLet12_6QNode_Int_10QNone_Int_1_argbuf_r;
  Pointer_QTree_Int_t lizzieLet12_6QNode_Int_11QNone_Int_d;
  logic lizzieLet12_6QNode_Int_11QNone_Int_r;
  Pointer_QTree_Int_t _57_d;
  logic _57_r;
  assign _57_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet12_6QNode_Int_11QNode_Int_d;
  logic lizzieLet12_6QNode_Int_11QNode_Int_r;
  Pointer_QTree_Int_t _56_d;
  logic _56_r;
  assign _56_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet12_6QNode_Int_11QNone_Int_1_argbuf_d;
  logic lizzieLet12_6QNode_Int_11QNone_Int_1_argbuf_r;
  Pointer_QTree_Int_t lizzieLet12_6QNode_Int_12QNone_Int_d;
  logic lizzieLet12_6QNode_Int_12QNone_Int_r;
  Pointer_QTree_Int_t _55_d;
  logic _55_r;
  assign _55_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet12_6QNode_Int_12QNode_Int_d;
  logic lizzieLet12_6QNode_Int_12QNode_Int_r;
  Pointer_QTree_Int_t _54_d;
  logic _54_r;
  assign _54_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet12_6QNode_Int_12QNode_Int_1_argbuf_d;
  logic lizzieLet12_6QNode_Int_12QNode_Int_1_argbuf_r;
  Pointer_QTree_Int_t lizzieLet12_6QNode_Int_12QNone_Int_1_argbuf_d;
  logic lizzieLet12_6QNode_Int_12QNone_Int_1_argbuf_r;
  Pointer_QTree_Int_t t1a8Y_destruct_d;
  logic t1a8Y_destruct_r;
  Pointer_QTree_Int_t t2a8Z_destruct_d;
  logic t2a8Z_destruct_r;
  Pointer_QTree_Int_t t3a90_destruct_d;
  logic t3a90_destruct_r;
  Pointer_QTree_Int_t t4a91_destruct_d;
  logic t4a91_destruct_r;
  QTree_Int_t _53_d;
  logic _53_r;
  assign _53_r = 1'd1;
  QTree_Int_t _52_d;
  logic _52_r;
  assign _52_r = 1'd1;
  QTree_Int_t lizzieLet12_6QNode_Int_1QNode_Int_d;
  logic lizzieLet12_6QNode_Int_1QNode_Int_r;
  QTree_Int_t _51_d;
  logic _51_r;
  assign _51_r = 1'd1;
  Go_t lizzieLet12_6QNode_Int_3QNone_Int_d;
  logic lizzieLet12_6QNode_Int_3QNone_Int_r;
  Go_t lizzieLet12_6QNode_Int_3QVal_Int_d;
  logic lizzieLet12_6QNode_Int_3QVal_Int_r;
  Go_t lizzieLet12_6QNode_Int_3QNode_Int_d;
  logic lizzieLet12_6QNode_Int_3QNode_Int_r;
  Go_t lizzieLet12_6QNode_Int_3QError_Int_d;
  logic lizzieLet12_6QNode_Int_3QError_Int_r;
  Go_t lizzieLet12_6QNode_Int_3QError_Int_1_d;
  logic lizzieLet12_6QNode_Int_3QError_Int_1_r;
  Go_t lizzieLet12_6QNode_Int_3QError_Int_2_d;
  logic lizzieLet12_6QNode_Int_3QError_Int_2_r;
  QTree_Int_t lizzieLet12_6QNode_Int_3QError_Int_1QError_Int_d;
  logic lizzieLet12_6QNode_Int_3QError_Int_1QError_Int_r;
  QTree_Int_t lizzieLet31_1_argbuf_d;
  logic lizzieLet31_1_argbuf_r;
  Go_t lizzieLet12_6QNode_Int_3QError_Int_2_argbuf_d;
  logic lizzieLet12_6QNode_Int_3QError_Int_2_argbuf_r;
  Go_t lizzieLet12_6QNode_Int_3QNode_Int_1_argbuf_d;
  logic lizzieLet12_6QNode_Int_3QNode_Int_1_argbuf_r;
  Go_t lizzieLet12_6QNode_Int_3QNone_Int_1_d;
  logic lizzieLet12_6QNode_Int_3QNone_Int_1_r;
  Go_t lizzieLet12_6QNode_Int_3QNone_Int_2_d;
  logic lizzieLet12_6QNode_Int_3QNone_Int_2_r;
  Go_t lizzieLet12_6QNode_Int_3QNone_Int_3_d;
  logic lizzieLet12_6QNode_Int_3QNone_Int_3_r;
  Go_t lizzieLet12_6QNode_Int_3QNone_Int_4_d;
  logic lizzieLet12_6QNode_Int_3QNone_Int_4_r;
  Go_t lizzieLet12_6QNode_Int_3QNone_Int_5_d;
  logic lizzieLet12_6QNode_Int_3QNone_Int_5_r;
  Go_t lizzieLet12_6QNode_Int_3QNone_Int_1_argbuf_d;
  logic lizzieLet12_6QNode_Int_3QNone_Int_1_argbuf_r;
  TupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_t \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int5_d ;
  logic \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int5_r ;
  Go_t lizzieLet12_6QNode_Int_3QNone_Int_2_argbuf_d;
  logic lizzieLet12_6QNode_Int_3QNone_Int_2_argbuf_r;
  TupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_t \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int6_d ;
  logic \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int6_r ;
  Go_t lizzieLet12_6QNode_Int_3QNone_Int_3_argbuf_d;
  logic lizzieLet12_6QNode_Int_3QNone_Int_3_argbuf_r;
  TupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_t \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int7_d ;
  logic \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int7_r ;
  Go_t lizzieLet12_6QNode_Int_3QNone_Int_4_argbuf_d;
  logic lizzieLet12_6QNode_Int_3QNone_Int_4_argbuf_r;
  TupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_t \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int8_d ;
  logic \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int8_r ;
  Go_t lizzieLet12_6QNode_Int_3QNone_Int_5_argbuf_d;
  logic lizzieLet12_6QNode_Int_3QNone_Int_5_argbuf_r;
  Go_t lizzieLet12_6QNode_Int_3QVal_Int_1_d;
  logic lizzieLet12_6QNode_Int_3QVal_Int_1_r;
  Go_t lizzieLet12_6QNode_Int_3QVal_Int_2_d;
  logic lizzieLet12_6QNode_Int_3QVal_Int_2_r;
  QTree_Int_t lizzieLet12_6QNode_Int_3QVal_Int_1QError_Int_d;
  logic lizzieLet12_6QNode_Int_3QVal_Int_1QError_Int_r;
  QTree_Int_t lizzieLet29_1_argbuf_d;
  logic lizzieLet29_1_argbuf_r;
  Go_t lizzieLet12_6QNode_Int_3QVal_Int_2_argbuf_d;
  logic lizzieLet12_6QNode_Int_3QVal_Int_2_argbuf_r;
  MyDTInt_Bool_t _50_d;
  logic _50_r;
  assign _50_r = 1'd1;
  MyDTInt_Bool_t _49_d;
  logic _49_r;
  assign _49_r = 1'd1;
  MyDTInt_Bool_t lizzieLet12_6QNode_Int_4QNode_Int_d;
  logic lizzieLet12_6QNode_Int_4QNode_Int_r;
  MyDTInt_Bool_t _48_d;
  logic _48_r;
  assign _48_r = 1'd1;
  MyDTInt_Bool_t lizzieLet12_6QNode_Int_4QNode_Int_1_d;
  logic lizzieLet12_6QNode_Int_4QNode_Int_1_r;
  MyDTInt_Bool_t lizzieLet12_6QNode_Int_4QNode_Int_2_d;
  logic lizzieLet12_6QNode_Int_4QNode_Int_2_r;
  MyDTInt_Bool_t lizzieLet12_6QNode_Int_4QNode_Int_2_argbuf_d;
  logic lizzieLet12_6QNode_Int_4QNode_Int_2_argbuf_r;
  MyDTInt_Bool_t lizzieLet12_6QNode_Int_5QNone_Int_d;
  logic lizzieLet12_6QNode_Int_5QNone_Int_r;
  MyDTInt_Bool_t _47_d;
  logic _47_r;
  assign _47_r = 1'd1;
  MyDTInt_Bool_t lizzieLet12_6QNode_Int_5QNode_Int_d;
  logic lizzieLet12_6QNode_Int_5QNode_Int_r;
  MyDTInt_Bool_t _46_d;
  logic _46_r;
  assign _46_r = 1'd1;
  MyDTInt_Bool_t lizzieLet12_6QNode_Int_5QNode_Int_1_d;
  logic lizzieLet12_6QNode_Int_5QNode_Int_1_r;
  MyDTInt_Bool_t lizzieLet12_6QNode_Int_5QNode_Int_2_d;
  logic lizzieLet12_6QNode_Int_5QNode_Int_2_r;
  MyDTInt_Bool_t lizzieLet12_6QNode_Int_5QNode_Int_2_argbuf_d;
  logic lizzieLet12_6QNode_Int_5QNode_Int_2_argbuf_r;
  MyDTInt_Bool_t lizzieLet12_6QNode_Int_5QNone_Int_1_d;
  logic lizzieLet12_6QNode_Int_5QNone_Int_1_r;
  MyDTInt_Bool_t lizzieLet12_6QNode_Int_5QNone_Int_2_d;
  logic lizzieLet12_6QNode_Int_5QNone_Int_2_r;
  MyDTInt_Bool_t lizzieLet12_6QNode_Int_5QNone_Int_3_d;
  logic lizzieLet12_6QNode_Int_5QNone_Int_3_r;
  MyDTInt_Bool_t lizzieLet12_6QNode_Int_5QNone_Int_4_d;
  logic lizzieLet12_6QNode_Int_5QNone_Int_4_r;
  MyDTInt_Bool_t lizzieLet12_6QNode_Int_5QNone_Int_1_argbuf_d;
  logic lizzieLet12_6QNode_Int_5QNone_Int_1_argbuf_r;
  MyDTInt_Bool_t lizzieLet12_6QNode_Int_5QNone_Int_2_argbuf_d;
  logic lizzieLet12_6QNode_Int_5QNone_Int_2_argbuf_r;
  MyDTInt_Bool_t lizzieLet12_6QNode_Int_5QNone_Int_3_argbuf_d;
  logic lizzieLet12_6QNode_Int_5QNone_Int_3_argbuf_r;
  MyDTInt_Bool_t lizzieLet12_6QNode_Int_5QNone_Int_4_argbuf_d;
  logic lizzieLet12_6QNode_Int_5QNone_Int_4_argbuf_r;
  MyDTInt_Int_Int_t _45_d;
  logic _45_r;
  assign _45_r = 1'd1;
  MyDTInt_Int_Int_t _44_d;
  logic _44_r;
  assign _44_r = 1'd1;
  MyDTInt_Int_Int_t lizzieLet12_6QNode_Int_6QNode_Int_d;
  logic lizzieLet12_6QNode_Int_6QNode_Int_r;
  MyDTInt_Int_Int_t _43_d;
  logic _43_r;
  assign _43_r = 1'd1;
  MyDTInt_Int_Int_t lizzieLet12_6QNode_Int_6QNode_Int_1_d;
  logic lizzieLet12_6QNode_Int_6QNode_Int_1_r;
  MyDTInt_Int_Int_t lizzieLet12_6QNode_Int_6QNode_Int_2_d;
  logic lizzieLet12_6QNode_Int_6QNode_Int_2_r;
  MyDTInt_Int_Int_t lizzieLet12_6QNode_Int_6QNode_Int_2_argbuf_d;
  logic lizzieLet12_6QNode_Int_6QNode_Int_2_argbuf_r;
  MyDTInt_Int_t lizzieLet12_6QNode_Int_7QNone_Int_d;
  logic lizzieLet12_6QNode_Int_7QNone_Int_r;
  MyDTInt_Int_t _42_d;
  logic _42_r;
  assign _42_r = 1'd1;
  MyDTInt_Int_t lizzieLet12_6QNode_Int_7QNode_Int_d;
  logic lizzieLet12_6QNode_Int_7QNode_Int_r;
  MyDTInt_Int_t _41_d;
  logic _41_r;
  assign _41_r = 1'd1;
  MyDTInt_Int_t lizzieLet12_6QNode_Int_7QNode_Int_1_d;
  logic lizzieLet12_6QNode_Int_7QNode_Int_1_r;
  MyDTInt_Int_t lizzieLet12_6QNode_Int_7QNode_Int_2_d;
  logic lizzieLet12_6QNode_Int_7QNode_Int_2_r;
  MyDTInt_Int_t lizzieLet12_6QNode_Int_7QNode_Int_2_argbuf_d;
  logic lizzieLet12_6QNode_Int_7QNode_Int_2_argbuf_r;
  MyDTInt_Int_t lizzieLet12_6QNode_Int_7QNone_Int_1_d;
  logic lizzieLet12_6QNode_Int_7QNone_Int_1_r;
  MyDTInt_Int_t lizzieLet12_6QNode_Int_7QNone_Int_2_d;
  logic lizzieLet12_6QNode_Int_7QNone_Int_2_r;
  MyDTInt_Int_t lizzieLet12_6QNode_Int_7QNone_Int_3_d;
  logic lizzieLet12_6QNode_Int_7QNone_Int_3_r;
  MyDTInt_Int_t lizzieLet12_6QNode_Int_7QNone_Int_4_d;
  logic lizzieLet12_6QNode_Int_7QNone_Int_4_r;
  MyDTInt_Int_t lizzieLet12_6QNode_Int_7QNone_Int_1_argbuf_d;
  logic lizzieLet12_6QNode_Int_7QNone_Int_1_argbuf_r;
  MyDTInt_Int_t lizzieLet12_6QNode_Int_7QNone_Int_2_argbuf_d;
  logic lizzieLet12_6QNode_Int_7QNone_Int_2_argbuf_r;
  MyDTInt_Int_t lizzieLet12_6QNode_Int_7QNone_Int_3_argbuf_d;
  logic lizzieLet12_6QNode_Int_7QNone_Int_3_argbuf_r;
  MyDTInt_Int_t lizzieLet12_6QNode_Int_7QNone_Int_4_argbuf_d;
  logic lizzieLet12_6QNode_Int_7QNone_Int_4_argbuf_r;
  Pointer_CTf_f_Int_Int_t lizzieLet12_6QNode_Int_8QNone_Int_d;
  logic lizzieLet12_6QNode_Int_8QNone_Int_r;
  Pointer_CTf_f_Int_Int_t lizzieLet12_6QNode_Int_8QVal_Int_d;
  logic lizzieLet12_6QNode_Int_8QVal_Int_r;
  Pointer_CTf_f_Int_Int_t lizzieLet12_6QNode_Int_8QNode_Int_d;
  logic lizzieLet12_6QNode_Int_8QNode_Int_r;
  Pointer_CTf_f_Int_Int_t lizzieLet12_6QNode_Int_8QError_Int_d;
  logic lizzieLet12_6QNode_Int_8QError_Int_r;
  Pointer_CTf_f_Int_Int_t lizzieLet12_6QNode_Int_8QError_Int_1_argbuf_d;
  logic lizzieLet12_6QNode_Int_8QError_Int_1_argbuf_r;
  CTf_f_Int_Int_t lizzieLet12_6QNode_Int_8QNode_Int_1lizzieLet12_6QNode_Int_9QNode_Int_1t1a8Y_1lizzieLet12_6QNode_Int_5QNode_Int_1lizzieLet12_6QNode_Int_7QNode_Int_1lizzieLet12_6QNode_Int_4QNode_Int_1lizzieLet12_6QNode_Int_6QNode_Int_1lizzieLet12_6QNode_Int_10QNode_Int_1t2a8Z_1lizzieLet12_6QNode_Int_11QNode_Int_1t3a90_1Lcall_f_f_Int_Int3_d;
  logic lizzieLet12_6QNode_Int_8QNode_Int_1lizzieLet12_6QNode_Int_9QNode_Int_1t1a8Y_1lizzieLet12_6QNode_Int_5QNode_Int_1lizzieLet12_6QNode_Int_7QNode_Int_1lizzieLet12_6QNode_Int_4QNode_Int_1lizzieLet12_6QNode_Int_6QNode_Int_1lizzieLet12_6QNode_Int_10QNode_Int_1t2a8Z_1lizzieLet12_6QNode_Int_11QNode_Int_1t3a90_1Lcall_f_f_Int_Int3_r;
  CTf_f_Int_Int_t lizzieLet30_1_argbuf_d;
  logic lizzieLet30_1_argbuf_r;
  Pointer_CTf_f_Int_Int_t lizzieLet12_6QNode_Int_8QNone_Int_1_argbuf_d;
  logic lizzieLet12_6QNode_Int_8QNone_Int_1_argbuf_r;
  Pointer_CTf_f_Int_Int_t lizzieLet12_6QNode_Int_8QVal_Int_1_argbuf_d;
  logic lizzieLet12_6QNode_Int_8QVal_Int_1_argbuf_r;
  Pointer_QTree_Int_t lizzieLet12_6QNode_Int_9QNone_Int_d;
  logic lizzieLet12_6QNode_Int_9QNone_Int_r;
  Pointer_QTree_Int_t _40_d;
  logic _40_r;
  assign _40_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet12_6QNode_Int_9QNode_Int_d;
  logic lizzieLet12_6QNode_Int_9QNode_Int_r;
  Pointer_QTree_Int_t _39_d;
  logic _39_r;
  assign _39_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet12_6QNode_Int_9QNone_Int_1_argbuf_d;
  logic lizzieLet12_6QNode_Int_9QNone_Int_1_argbuf_r;
  QTree_Int_t lizzieLet12_6QNone_Int_1_d;
  logic lizzieLet12_6QNone_Int_1_r;
  QTree_Int_t lizzieLet12_6QNone_Int_2_d;
  logic lizzieLet12_6QNone_Int_2_r;
  QTree_Int_t lizzieLet12_6QNone_Int_3_d;
  logic lizzieLet12_6QNone_Int_3_r;
  QTree_Int_t lizzieLet12_6QNone_Int_4_d;
  logic lizzieLet12_6QNone_Int_4_r;
  QTree_Int_t lizzieLet12_6QNone_Int_5_d;
  logic lizzieLet12_6QNone_Int_5_r;
  QTree_Int_t lizzieLet12_6QNone_Int_6_d;
  logic lizzieLet12_6QNone_Int_6_r;
  Pointer_QTree_Int_t tla8J_destruct_d;
  logic tla8J_destruct_r;
  Pointer_QTree_Int_t tra8K_destruct_d;
  logic tra8K_destruct_r;
  Pointer_QTree_Int_t bla8L_destruct_d;
  logic bla8L_destruct_r;
  Pointer_QTree_Int_t bra8M_destruct_d;
  logic bra8M_destruct_r;
  Int_t va8I_destruct_d;
  logic va8I_destruct_r;
  QTree_Int_t _38_d;
  logic _38_r;
  assign _38_r = 1'd1;
  QTree_Int_t lizzieLet12_6QNone_Int_1QVal_Int_d;
  logic lizzieLet12_6QNone_Int_1QVal_Int_r;
  QTree_Int_t lizzieLet12_6QNone_Int_1QNode_Int_d;
  logic lizzieLet12_6QNone_Int_1QNode_Int_r;
  QTree_Int_t _37_d;
  logic _37_r;
  assign _37_r = 1'd1;
  Go_t lizzieLet12_6QNone_Int_3QNone_Int_d;
  logic lizzieLet12_6QNone_Int_3QNone_Int_r;
  Go_t lizzieLet12_6QNone_Int_3QVal_Int_d;
  logic lizzieLet12_6QNone_Int_3QVal_Int_r;
  Go_t lizzieLet12_6QNone_Int_3QNode_Int_d;
  logic lizzieLet12_6QNone_Int_3QNode_Int_r;
  Go_t lizzieLet12_6QNone_Int_3QError_Int_d;
  logic lizzieLet12_6QNone_Int_3QError_Int_r;
  Go_t lizzieLet12_6QNone_Int_3QError_Int_1_d;
  logic lizzieLet12_6QNone_Int_3QError_Int_1_r;
  Go_t lizzieLet12_6QNone_Int_3QError_Int_2_d;
  logic lizzieLet12_6QNone_Int_3QError_Int_2_r;
  QTree_Int_t lizzieLet12_6QNone_Int_3QError_Int_1QError_Int_d;
  logic lizzieLet12_6QNone_Int_3QError_Int_1QError_Int_r;
  QTree_Int_t lizzieLet18_1_argbuf_d;
  logic lizzieLet18_1_argbuf_r;
  Go_t lizzieLet12_6QNone_Int_3QError_Int_2_argbuf_d;
  logic lizzieLet12_6QNone_Int_3QError_Int_2_argbuf_r;
  Go_t lizzieLet12_6QNone_Int_3QNode_Int_1_d;
  logic lizzieLet12_6QNone_Int_3QNode_Int_1_r;
  Go_t lizzieLet12_6QNone_Int_3QNode_Int_2_d;
  logic lizzieLet12_6QNone_Int_3QNode_Int_2_r;
  Go_t lizzieLet12_6QNone_Int_3QNode_Int_3_d;
  logic lizzieLet12_6QNone_Int_3QNode_Int_3_r;
  Go_t lizzieLet12_6QNone_Int_3QNode_Int_4_d;
  logic lizzieLet12_6QNone_Int_3QNode_Int_4_r;
  Go_t lizzieLet12_6QNone_Int_3QNode_Int_5_d;
  logic lizzieLet12_6QNone_Int_3QNode_Int_5_r;
  Go_t lizzieLet12_6QNone_Int_3QNode_Int_1_argbuf_d;
  logic lizzieLet12_6QNone_Int_3QNode_Int_1_argbuf_r;
  TupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_t \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_1_d ;
  logic \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_1_r ;
  Go_t lizzieLet12_6QNone_Int_3QNode_Int_2_argbuf_d;
  logic lizzieLet12_6QNone_Int_3QNode_Int_2_argbuf_r;
  TupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_t \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int2_d ;
  logic \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int2_r ;
  Go_t lizzieLet12_6QNone_Int_3QNode_Int_3_argbuf_d;
  logic lizzieLet12_6QNone_Int_3QNode_Int_3_argbuf_r;
  TupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_t \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int3_d ;
  logic \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int3_r ;
  Go_t lizzieLet12_6QNone_Int_3QNode_Int_4_argbuf_d;
  logic lizzieLet12_6QNone_Int_3QNode_Int_4_argbuf_r;
  TupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_t \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int4_d ;
  logic \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int4_r ;
  Go_t lizzieLet12_6QNone_Int_3QNode_Int_5_argbuf_d;
  logic lizzieLet12_6QNone_Int_3QNode_Int_5_argbuf_r;
  Go_t lizzieLet12_6QNone_Int_3QNone_Int_1_d;
  logic lizzieLet12_6QNone_Int_3QNone_Int_1_r;
  Go_t lizzieLet12_6QNone_Int_3QNone_Int_2_d;
  logic lizzieLet12_6QNone_Int_3QNone_Int_2_r;
  QTree_Int_t lizzieLet12_6QNone_Int_3QNone_Int_1QNone_Int_d;
  logic lizzieLet12_6QNone_Int_3QNone_Int_1QNone_Int_r;
  QTree_Int_t lizzieLet14_1_argbuf_d;
  logic lizzieLet14_1_argbuf_r;
  Go_t lizzieLet12_6QNone_Int_3QNone_Int_2_argbuf_d;
  logic lizzieLet12_6QNone_Int_3QNone_Int_2_argbuf_r;
  C17_t go_17_goMux_choice_d;
  logic go_17_goMux_choice_r;
  Go_t go_17_goMux_data_d;
  logic go_17_goMux_data_r;
  Go_t lizzieLet12_6QNone_Int_3QVal_Int_1_d;
  logic lizzieLet12_6QNone_Int_3QVal_Int_1_r;
  Go_t lizzieLet12_6QNone_Int_3QVal_Int_2_d;
  logic lizzieLet12_6QNone_Int_3QVal_Int_2_r;
  Go_t lizzieLet12_6QNone_Int_3QVal_Int_3_d;
  logic lizzieLet12_6QNone_Int_3QVal_Int_3_r;
  Go_t lizzieLet12_6QNone_Int_3QVal_Int_1_argbuf_d;
  logic lizzieLet12_6QNone_Int_3QVal_Int_1_argbuf_r;
  TupGo___MyDTInt_Int___Int_t applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_d;
  logic applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_r;
  Go_t lizzieLet12_6QNone_Int_3QVal_Int_2_argbuf_d;
  logic lizzieLet12_6QNone_Int_3QVal_Int_2_argbuf_r;
  TupGo___MyDTInt_Bool___Int_t applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_d;
  logic applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_r;
  MyDTInt_Bool_t _36_d;
  logic _36_r;
  assign _36_r = 1'd1;
  MyDTInt_Bool_t lizzieLet12_6QNone_Int_4QVal_Int_d;
  logic lizzieLet12_6QNone_Int_4QVal_Int_r;
  MyDTInt_Bool_t lizzieLet12_6QNone_Int_4QNode_Int_d;
  logic lizzieLet12_6QNone_Int_4QNode_Int_r;
  MyDTInt_Bool_t _35_d;
  logic _35_r;
  assign _35_r = 1'd1;
  MyDTInt_Bool_t lizzieLet12_6QNone_Int_4QNode_Int_1_d;
  logic lizzieLet12_6QNone_Int_4QNode_Int_1_r;
  MyDTInt_Bool_t lizzieLet12_6QNone_Int_4QNode_Int_2_d;
  logic lizzieLet12_6QNone_Int_4QNode_Int_2_r;
  MyDTInt_Bool_t lizzieLet12_6QNone_Int_4QNode_Int_3_d;
  logic lizzieLet12_6QNone_Int_4QNode_Int_3_r;
  MyDTInt_Bool_t lizzieLet12_6QNone_Int_4QNode_Int_4_d;
  logic lizzieLet12_6QNone_Int_4QNode_Int_4_r;
  MyDTInt_Bool_t lizzieLet12_6QNone_Int_4QNode_Int_1_argbuf_d;
  logic lizzieLet12_6QNone_Int_4QNode_Int_1_argbuf_r;
  MyDTInt_Bool_t lizzieLet12_6QNone_Int_4QNode_Int_2_argbuf_d;
  logic lizzieLet12_6QNone_Int_4QNode_Int_2_argbuf_r;
  MyDTInt_Bool_t lizzieLet12_6QNone_Int_4QNode_Int_3_argbuf_d;
  logic lizzieLet12_6QNone_Int_4QNode_Int_3_argbuf_r;
  MyDTInt_Bool_t lizzieLet12_6QNone_Int_4QNode_Int_4_argbuf_d;
  logic lizzieLet12_6QNone_Int_4QNode_Int_4_argbuf_r;
  MyDTInt_Bool_t lizzieLet12_6QNone_Int_4QVal_Int_1_argbuf_d;
  logic lizzieLet12_6QNone_Int_4QVal_Int_1_argbuf_r;
  MyDTInt_Int_t _34_d;
  logic _34_r;
  assign _34_r = 1'd1;
  MyDTInt_Int_t lizzieLet12_6QNone_Int_5QVal_Int_d;
  logic lizzieLet12_6QNone_Int_5QVal_Int_r;
  MyDTInt_Int_t lizzieLet12_6QNone_Int_5QNode_Int_d;
  logic lizzieLet12_6QNone_Int_5QNode_Int_r;
  MyDTInt_Int_t _33_d;
  logic _33_r;
  assign _33_r = 1'd1;
  MyDTInt_Int_t lizzieLet12_6QNone_Int_5QNode_Int_1_d;
  logic lizzieLet12_6QNone_Int_5QNode_Int_1_r;
  MyDTInt_Int_t lizzieLet12_6QNone_Int_5QNode_Int_2_d;
  logic lizzieLet12_6QNone_Int_5QNode_Int_2_r;
  MyDTInt_Int_t lizzieLet12_6QNone_Int_5QNode_Int_3_d;
  logic lizzieLet12_6QNone_Int_5QNode_Int_3_r;
  MyDTInt_Int_t lizzieLet12_6QNone_Int_5QNode_Int_4_d;
  logic lizzieLet12_6QNone_Int_5QNode_Int_4_r;
  MyDTInt_Int_t lizzieLet12_6QNone_Int_5QNode_Int_1_argbuf_d;
  logic lizzieLet12_6QNone_Int_5QNode_Int_1_argbuf_r;
  MyDTInt_Int_t lizzieLet12_6QNone_Int_5QNode_Int_2_argbuf_d;
  logic lizzieLet12_6QNone_Int_5QNode_Int_2_argbuf_r;
  MyDTInt_Int_t lizzieLet12_6QNone_Int_5QNode_Int_3_argbuf_d;
  logic lizzieLet12_6QNone_Int_5QNode_Int_3_argbuf_r;
  MyDTInt_Int_t lizzieLet12_6QNone_Int_5QNode_Int_4_argbuf_d;
  logic lizzieLet12_6QNone_Int_5QNode_Int_4_argbuf_r;
  MyDTInt_Int_t lizzieLet12_6QNone_Int_5QVal_Int_1_d;
  logic lizzieLet12_6QNone_Int_5QVal_Int_1_r;
  MyDTInt_Int_t lizzieLet12_6QNone_Int_5QVal_Int_2_d;
  logic lizzieLet12_6QNone_Int_5QVal_Int_2_r;
  MyDTInt_Int_t lizzieLet12_6QNone_Int_5QVal_Int_1_argbuf_d;
  logic lizzieLet12_6QNone_Int_5QVal_Int_1_argbuf_r;
  Pointer_CTf_f_Int_Int_t lizzieLet12_6QNone_Int_6QNone_Int_d;
  logic lizzieLet12_6QNone_Int_6QNone_Int_r;
  Pointer_CTf_f_Int_Int_t lizzieLet12_6QNone_Int_6QVal_Int_d;
  logic lizzieLet12_6QNone_Int_6QVal_Int_r;
  Pointer_CTf_f_Int_Int_t lizzieLet12_6QNone_Int_6QNode_Int_d;
  logic lizzieLet12_6QNone_Int_6QNode_Int_r;
  Pointer_CTf_f_Int_Int_t lizzieLet12_6QNone_Int_6QError_Int_d;
  logic lizzieLet12_6QNone_Int_6QError_Int_r;
  Pointer_CTf_f_Int_Int_t lizzieLet12_6QNone_Int_6QError_Int_1_argbuf_d;
  logic lizzieLet12_6QNone_Int_6QError_Int_1_argbuf_r;
  Pointer_CTf_f_Int_Int_t lizzieLet12_6QNone_Int_6QNode_Int_1_argbuf_d;
  logic lizzieLet12_6QNone_Int_6QNode_Int_1_argbuf_r;
  Pointer_CTf_f_Int_Int_t lizzieLet12_6QNone_Int_6QNone_Int_1_argbuf_d;
  logic lizzieLet12_6QNone_Int_6QNone_Int_1_argbuf_r;
  QTree_Int_t lizzieLet12_6QVal_Int_1_d;
  logic lizzieLet12_6QVal_Int_1_r;
  QTree_Int_t lizzieLet12_6QVal_Int_2_d;
  logic lizzieLet12_6QVal_Int_2_r;
  QTree_Int_t lizzieLet12_6QVal_Int_3_d;
  logic lizzieLet12_6QVal_Int_3_r;
  QTree_Int_t lizzieLet12_6QVal_Int_4_d;
  logic lizzieLet12_6QVal_Int_4_r;
  QTree_Int_t lizzieLet12_6QVal_Int_5_d;
  logic lizzieLet12_6QVal_Int_5_r;
  QTree_Int_t lizzieLet12_6QVal_Int_6_d;
  logic lizzieLet12_6QVal_Int_6_r;
  QTree_Int_t lizzieLet12_6QVal_Int_7_d;
  logic lizzieLet12_6QVal_Int_7_r;
  QTree_Int_t lizzieLet12_6QVal_Int_8_d;
  logic lizzieLet12_6QVal_Int_8_r;
  QTree_Int_t lizzieLet12_6QVal_Int_9_d;
  logic lizzieLet12_6QVal_Int_9_r;
  Int_t va8O_destruct_d;
  logic va8O_destruct_r;
  QTree_Int_t _32_d;
  logic _32_r;
  assign _32_r = 1'd1;
  QTree_Int_t lizzieLet12_6QVal_Int_1QVal_Int_d;
  logic lizzieLet12_6QVal_Int_1QVal_Int_r;
  QTree_Int_t _31_d;
  logic _31_r;
  assign _31_r = 1'd1;
  QTree_Int_t _30_d;
  logic _30_r;
  assign _30_r = 1'd1;
  Go_t lizzieLet12_6QVal_Int_3QNone_Int_d;
  logic lizzieLet12_6QVal_Int_3QNone_Int_r;
  Go_t lizzieLet12_6QVal_Int_3QVal_Int_d;
  logic lizzieLet12_6QVal_Int_3QVal_Int_r;
  Go_t lizzieLet12_6QVal_Int_3QNode_Int_d;
  logic lizzieLet12_6QVal_Int_3QNode_Int_r;
  Go_t lizzieLet12_6QVal_Int_3QError_Int_d;
  logic lizzieLet12_6QVal_Int_3QError_Int_r;
  Go_t lizzieLet12_6QVal_Int_3QError_Int_1_d;
  logic lizzieLet12_6QVal_Int_3QError_Int_1_r;
  Go_t lizzieLet12_6QVal_Int_3QError_Int_2_d;
  logic lizzieLet12_6QVal_Int_3QError_Int_2_r;
  QTree_Int_t lizzieLet12_6QVal_Int_3QError_Int_1QError_Int_d;
  logic lizzieLet12_6QVal_Int_3QError_Int_1QError_Int_r;
  QTree_Int_t lizzieLet26_1_argbuf_d;
  logic lizzieLet26_1_argbuf_r;
  Go_t lizzieLet12_6QVal_Int_3QError_Int_2_argbuf_d;
  logic lizzieLet12_6QVal_Int_3QError_Int_2_argbuf_r;
  Go_t lizzieLet12_6QVal_Int_3QNode_Int_1_d;
  logic lizzieLet12_6QVal_Int_3QNode_Int_1_r;
  Go_t lizzieLet12_6QVal_Int_3QNode_Int_2_d;
  logic lizzieLet12_6QVal_Int_3QNode_Int_2_r;
  QTree_Int_t lizzieLet12_6QVal_Int_3QNode_Int_1QError_Int_d;
  logic lizzieLet12_6QVal_Int_3QNode_Int_1QError_Int_r;
  QTree_Int_t lizzieLet25_1_1_argbuf_d;
  logic lizzieLet25_1_1_argbuf_r;
  Go_t lizzieLet12_6QVal_Int_3QNode_Int_2_argbuf_d;
  logic lizzieLet12_6QVal_Int_3QNode_Int_2_argbuf_r;
  Go_t lizzieLet12_6QVal_Int_3QNone_Int_1_d;
  logic lizzieLet12_6QVal_Int_3QNone_Int_1_r;
  Go_t lizzieLet12_6QVal_Int_3QNone_Int_2_d;
  logic lizzieLet12_6QVal_Int_3QNone_Int_2_r;
  Go_t lizzieLet12_6QVal_Int_3QNone_Int_3_d;
  logic lizzieLet12_6QVal_Int_3QNone_Int_3_r;
  Go_t lizzieLet12_6QVal_Int_3QNone_Int_1_argbuf_d;
  logic lizzieLet12_6QVal_Int_3QNone_Int_1_argbuf_r;
  TupGo___MyDTInt_Int___Int_t applyfnInt_Int_5TupGo___MyDTInt_Int___Int5_d;
  logic applyfnInt_Int_5TupGo___MyDTInt_Int___Int5_r;
  Go_t lizzieLet12_6QVal_Int_3QNone_Int_2_argbuf_d;
  logic lizzieLet12_6QVal_Int_3QNone_Int_2_argbuf_r;
  TupGo___MyDTInt_Bool___Int_t applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int3_d;
  logic applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int3_r;
  Go_t lizzieLet12_6QVal_Int_3QVal_Int_1_d;
  logic lizzieLet12_6QVal_Int_3QVal_Int_1_r;
  Go_t lizzieLet12_6QVal_Int_3QVal_Int_2_d;
  logic lizzieLet12_6QVal_Int_3QVal_Int_2_r;
  Go_t lizzieLet12_6QVal_Int_3QVal_Int_1_argbuf_d;
  logic lizzieLet12_6QVal_Int_3QVal_Int_1_argbuf_r;
  TupGo___MyDTInt_Bool___Int_t applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int4_d;
  logic applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int4_r;
  MyDTInt_Bool_t _29_d;
  logic _29_r;
  assign _29_r = 1'd1;
  MyDTInt_Bool_t lizzieLet12_6QVal_Int_4QVal_Int_d;
  logic lizzieLet12_6QVal_Int_4QVal_Int_r;
  MyDTInt_Bool_t _28_d;
  logic _28_r;
  assign _28_r = 1'd1;
  MyDTInt_Bool_t _27_d;
  logic _27_r;
  assign _27_r = 1'd1;
  MyDTInt_Bool_t lizzieLet12_6QVal_Int_4QVal_Int_1_argbuf_d;
  logic lizzieLet12_6QVal_Int_4QVal_Int_1_argbuf_r;
  MyDTInt_Bool_t lizzieLet12_6QVal_Int_5QNone_Int_d;
  logic lizzieLet12_6QVal_Int_5QNone_Int_r;
  MyDTInt_Bool_t lizzieLet12_6QVal_Int_5QVal_Int_d;
  logic lizzieLet12_6QVal_Int_5QVal_Int_r;
  MyDTInt_Bool_t _26_d;
  logic _26_r;
  assign _26_r = 1'd1;
  MyDTInt_Bool_t _25_d;
  logic _25_r;
  assign _25_r = 1'd1;
  MyDTInt_Bool_t lizzieLet12_6QVal_Int_5QNone_Int_1_argbuf_d;
  logic lizzieLet12_6QVal_Int_5QNone_Int_1_argbuf_r;
  MyDTInt_Int_Int_t _24_d;
  logic _24_r;
  assign _24_r = 1'd1;
  MyDTInt_Int_Int_t lizzieLet12_6QVal_Int_6QVal_Int_d;
  logic lizzieLet12_6QVal_Int_6QVal_Int_r;
  MyDTInt_Int_Int_t _23_d;
  logic _23_r;
  assign _23_r = 1'd1;
  MyDTInt_Int_Int_t _22_d;
  logic _22_r;
  assign _22_r = 1'd1;
  MyDTInt_Int_Int_t lizzieLet12_6QVal_Int_6QVal_Int_1_d;
  logic lizzieLet12_6QVal_Int_6QVal_Int_1_r;
  MyDTInt_Int_Int_t lizzieLet12_6QVal_Int_6QVal_Int_2_d;
  logic lizzieLet12_6QVal_Int_6QVal_Int_2_r;
  MyDTInt_Int_Int_t lizzieLet12_6QVal_Int_6QVal_Int_1_argbuf_d;
  logic lizzieLet12_6QVal_Int_6QVal_Int_1_argbuf_r;
  TupMyDTInt_Int_Int___Int___Int_t applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_d;
  logic applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_r;
  MyDTInt_Int_t lizzieLet12_6QVal_Int_7QNone_Int_d;
  logic lizzieLet12_6QVal_Int_7QNone_Int_r;
  MyDTInt_Int_t lizzieLet12_6QVal_Int_7QVal_Int_d;
  logic lizzieLet12_6QVal_Int_7QVal_Int_r;
  MyDTInt_Int_t _21_d;
  logic _21_r;
  assign _21_r = 1'd1;
  MyDTInt_Int_t _20_d;
  logic _20_r;
  assign _20_r = 1'd1;
  MyDTInt_Int_t lizzieLet12_6QVal_Int_7QNone_Int_1_d;
  logic lizzieLet12_6QVal_Int_7QNone_Int_1_r;
  MyDTInt_Int_t lizzieLet12_6QVal_Int_7QNone_Int_2_d;
  logic lizzieLet12_6QVal_Int_7QNone_Int_2_r;
  MyDTInt_Int_t lizzieLet12_6QVal_Int_7QNone_Int_1_argbuf_d;
  logic lizzieLet12_6QVal_Int_7QNone_Int_1_argbuf_r;
  Pointer_CTf_f_Int_Int_t lizzieLet12_6QVal_Int_8QNone_Int_d;
  logic lizzieLet12_6QVal_Int_8QNone_Int_r;
  Pointer_CTf_f_Int_Int_t lizzieLet12_6QVal_Int_8QVal_Int_d;
  logic lizzieLet12_6QVal_Int_8QVal_Int_r;
  Pointer_CTf_f_Int_Int_t lizzieLet12_6QVal_Int_8QNode_Int_d;
  logic lizzieLet12_6QVal_Int_8QNode_Int_r;
  Pointer_CTf_f_Int_Int_t lizzieLet12_6QVal_Int_8QError_Int_d;
  logic lizzieLet12_6QVal_Int_8QError_Int_r;
  Pointer_CTf_f_Int_Int_t lizzieLet12_6QVal_Int_8QError_Int_1_argbuf_d;
  logic lizzieLet12_6QVal_Int_8QError_Int_1_argbuf_r;
  Pointer_CTf_f_Int_Int_t lizzieLet12_6QVal_Int_8QNode_Int_1_argbuf_d;
  logic lizzieLet12_6QVal_Int_8QNode_Int_1_argbuf_r;
  Int_t lizzieLet12_6QVal_Int_9QNone_Int_d;
  logic lizzieLet12_6QVal_Int_9QNone_Int_r;
  Int_t lizzieLet12_6QVal_Int_9QVal_Int_d;
  logic lizzieLet12_6QVal_Int_9QVal_Int_r;
  Int_t _19_d;
  logic _19_r;
  assign _19_r = 1'd1;
  Int_t _18_d;
  logic _18_r;
  assign _18_r = 1'd1;
  Int_t lizzieLet12_6QVal_Int_9QNone_Int_1_d;
  logic lizzieLet12_6QVal_Int_9QNone_Int_1_r;
  Int_t lizzieLet12_6QVal_Int_9QNone_Int_2_d;
  logic lizzieLet12_6QVal_Int_9QNone_Int_2_r;
  Int_t lizzieLet12_6QVal_Int_9QNone_Int_1_argbuf_d;
  logic lizzieLet12_6QVal_Int_9QNone_Int_1_argbuf_r;
  Int_t lizzieLet12_6QVal_Int_9QVal_Int_1_d;
  logic lizzieLet12_6QVal_Int_9QVal_Int_1_r;
  Int_t lizzieLet12_6QVal_Int_9QVal_Int_2_d;
  logic lizzieLet12_6QVal_Int_9QVal_Int_2_r;
  Int_t lizzieLet12_6QVal_Int_9QVal_Int_1_argbuf_d;
  logic lizzieLet12_6QVal_Int_9QVal_Int_1_argbuf_r;
  MyDTInt_Int_Int_t _17_d;
  logic _17_r;
  assign _17_r = 1'd1;
  MyDTInt_Int_Int_t lizzieLet12_7QVal_Int_d;
  logic lizzieLet12_7QVal_Int_r;
  MyDTInt_Int_Int_t lizzieLet12_7QNode_Int_d;
  logic lizzieLet12_7QNode_Int_r;
  MyDTInt_Int_Int_t _16_d;
  logic _16_r;
  assign _16_r = 1'd1;
  MyDTInt_Int_t lizzieLet12_8QNone_Int_d;
  logic lizzieLet12_8QNone_Int_r;
  MyDTInt_Int_t lizzieLet12_8QVal_Int_d;
  logic lizzieLet12_8QVal_Int_r;
  MyDTInt_Int_t lizzieLet12_8QNode_Int_d;
  logic lizzieLet12_8QNode_Int_r;
  MyDTInt_Int_t _15_d;
  logic _15_r;
  assign _15_r = 1'd1;
  Pointer_CTf_f_Int_Int_t lizzieLet12_9QNone_Int_d;
  logic lizzieLet12_9QNone_Int_r;
  Pointer_CTf_f_Int_Int_t lizzieLet12_9QVal_Int_d;
  logic lizzieLet12_9QVal_Int_r;
  Pointer_CTf_f_Int_Int_t lizzieLet12_9QNode_Int_d;
  logic lizzieLet12_9QNode_Int_r;
  Pointer_CTf_f_Int_Int_t lizzieLet12_9QError_Int_d;
  logic lizzieLet12_9QError_Int_r;
  Pointer_CTf_f_Int_Int_t lizzieLet12_9QError_Int_1_argbuf_d;
  logic lizzieLet12_9QError_Int_1_argbuf_r;
  Bool_t lizzieLet2_1_argbuf_d;
  logic lizzieLet2_1_argbuf_r;
  \Int#_t  wwsj0_4_destruct_d;
  logic wwsj0_4_destruct_r;
  \Int#_t  ww1Xju_2_destruct_d;
  logic ww1Xju_2_destruct_r;
  \Int#_t  ww2Xjx_1_destruct_d;
  logic ww2Xjx_1_destruct_r;
  Pointer_CT$wnnz_t sc_0_6_destruct_d;
  logic sc_0_6_destruct_r;
  \Int#_t  wwsj0_3_destruct_d;
  logic wwsj0_3_destruct_r;
  \Int#_t  ww1Xju_1_destruct_d;
  logic ww1Xju_1_destruct_r;
  Pointer_CT$wnnz_t sc_0_5_destruct_d;
  logic sc_0_5_destruct_r;
  Pointer_QTree_Int_t q4a87_3_destruct_d;
  logic q4a87_3_destruct_r;
  \Int#_t  wwsj0_2_destruct_d;
  logic wwsj0_2_destruct_r;
  Pointer_CT$wnnz_t sc_0_4_destruct_d;
  logic sc_0_4_destruct_r;
  Pointer_QTree_Int_t q4a87_2_destruct_d;
  logic q4a87_2_destruct_r;
  Pointer_QTree_Int_t q3a86_2_destruct_d;
  logic q3a86_2_destruct_r;
  Pointer_CT$wnnz_t sc_0_3_destruct_d;
  logic sc_0_3_destruct_r;
  Pointer_QTree_Int_t q4a87_1_destruct_d;
  logic q4a87_1_destruct_r;
  Pointer_QTree_Int_t q3a86_1_destruct_d;
  logic q3a86_1_destruct_r;
  Pointer_QTree_Int_t q2a85_1_destruct_d;
  logic q2a85_1_destruct_r;
  CT$wnnz_t _14_d;
  logic _14_r;
  assign _14_r = 1'd1;
  CT$wnnz_t lizzieLet35_1Lcall_$wnnz3_d;
  logic lizzieLet35_1Lcall_$wnnz3_r;
  CT$wnnz_t lizzieLet35_1Lcall_$wnnz2_d;
  logic lizzieLet35_1Lcall_$wnnz2_r;
  CT$wnnz_t lizzieLet35_1Lcall_$wnnz1_d;
  logic lizzieLet35_1Lcall_$wnnz1_r;
  CT$wnnz_t lizzieLet35_1Lcall_$wnnz0_d;
  logic lizzieLet35_1Lcall_$wnnz0_r;
  Go_t _13_d;
  logic _13_r;
  assign _13_r = 1'd1;
  Go_t lizzieLet35_3Lcall_$wnnz3_d;
  logic lizzieLet35_3Lcall_$wnnz3_r;
  Go_t lizzieLet35_3Lcall_$wnnz2_d;
  logic lizzieLet35_3Lcall_$wnnz2_r;
  Go_t lizzieLet35_3Lcall_$wnnz1_d;
  logic lizzieLet35_3Lcall_$wnnz1_r;
  Go_t lizzieLet35_3Lcall_$wnnz0_d;
  logic lizzieLet35_3Lcall_$wnnz0_r;
  Go_t lizzieLet35_3Lcall_$wnnz0_1_argbuf_d;
  logic lizzieLet35_3Lcall_$wnnz0_1_argbuf_r;
  Go_t lizzieLet35_3Lcall_$wnnz1_1_argbuf_d;
  logic lizzieLet35_3Lcall_$wnnz1_1_argbuf_r;
  Go_t lizzieLet35_3Lcall_$wnnz2_1_argbuf_d;
  logic lizzieLet35_3Lcall_$wnnz2_1_argbuf_r;
  Go_t lizzieLet35_3Lcall_$wnnz3_1_argbuf_d;
  logic lizzieLet35_3Lcall_$wnnz3_1_argbuf_r;
  \Int#_t  lizzieLet35_4L$wnnzsbos_d;
  logic lizzieLet35_4L$wnnzsbos_r;
  \Int#_t  lizzieLet35_4Lcall_$wnnz3_d;
  logic lizzieLet35_4Lcall_$wnnz3_r;
  \Int#_t  lizzieLet35_4Lcall_$wnnz2_d;
  logic lizzieLet35_4Lcall_$wnnz2_r;
  \Int#_t  lizzieLet35_4Lcall_$wnnz1_d;
  logic lizzieLet35_4Lcall_$wnnz1_r;
  \Int#_t  lizzieLet35_4Lcall_$wnnz0_d;
  logic lizzieLet35_4Lcall_$wnnz0_r;
  \Int#_t  lizzieLet35_4L$wnnzsbos_1_merge_merge_fork_1_d;
  logic lizzieLet35_4L$wnnzsbos_1_merge_merge_fork_1_r;
  \Int#_t  lizzieLet35_4L$wnnzsbos_1_merge_merge_fork_2_d;
  logic lizzieLet35_4L$wnnzsbos_1_merge_merge_fork_2_r;
  Go_t call_$wnnz_goConst_d;
  logic call_$wnnz_goConst_r;
  \Int#_t  \$wnnz_resbuf_d ;
  logic \$wnnz_resbuf_r ;
  CT$wnnz_t lizzieLet35_4Lcall_$wnnz3_1sc_0_3_1q4a87_1_1q3a86_1_1Lcall_$wnnz2_d;
  logic lizzieLet35_4Lcall_$wnnz3_1sc_0_3_1q4a87_1_1q3a86_1_1Lcall_$wnnz2_r;
  CT$wnnz_t lizzieLet36_1_argbuf_d;
  logic lizzieLet36_1_argbuf_r;
  Pointer_QTree_Int_t es_5_2_destruct_d;
  logic es_5_2_destruct_r;
  Pointer_QTree_Int_t es_6_4_destruct_d;
  logic es_6_4_destruct_r;
  Pointer_QTree_Int_t es_7_4_destruct_d;
  logic es_7_4_destruct_r;
  \Pointer_CTf''''''''_f''''''''_Int_Int_t  sc_0_10_destruct_d;
  logic sc_0_10_destruct_r;
  Pointer_QTree_Int_t es_6_3_destruct_d;
  logic es_6_3_destruct_r;
  Pointer_QTree_Int_t es_7_3_destruct_d;
  logic es_7_3_destruct_r;
  \Pointer_CTf''''''''_f''''''''_Int_Int_t  sc_0_9_destruct_d;
  logic sc_0_9_destruct_r;
  Pointer_QTree_Int_t tla8y_3_destruct_d;
  logic tla8y_3_destruct_r;
  MyDTInt_Bool_t is_z_mapa8v_4_destruct_d;
  logic is_z_mapa8v_4_destruct_r;
  MyDTInt_Int_t op_mapa8w_4_destruct_d;
  logic op_mapa8w_4_destruct_r;
  Pointer_QTree_Int_t es_7_2_destruct_d;
  logic es_7_2_destruct_r;
  \Pointer_CTf''''''''_f''''''''_Int_Int_t  sc_0_8_destruct_d;
  logic sc_0_8_destruct_r;
  Pointer_QTree_Int_t tla8y_2_destruct_d;
  logic tla8y_2_destruct_r;
  MyDTInt_Bool_t is_z_mapa8v_3_destruct_d;
  logic is_z_mapa8v_3_destruct_r;
  MyDTInt_Int_t op_mapa8w_3_destruct_d;
  logic op_mapa8w_3_destruct_r;
  Pointer_QTree_Int_t tra8z_2_destruct_d;
  logic tra8z_2_destruct_r;
  \Pointer_CTf''''''''_f''''''''_Int_Int_t  sc_0_7_destruct_d;
  logic sc_0_7_destruct_r;
  Pointer_QTree_Int_t tla8y_1_destruct_d;
  logic tla8y_1_destruct_r;
  MyDTInt_Bool_t is_z_mapa8v_2_destruct_d;
  logic is_z_mapa8v_2_destruct_r;
  MyDTInt_Int_t op_mapa8w_2_destruct_d;
  logic op_mapa8w_2_destruct_r;
  Pointer_QTree_Int_t tra8z_1_destruct_d;
  logic tra8z_1_destruct_r;
  Pointer_QTree_Int_t bla8A_1_destruct_d;
  logic bla8A_1_destruct_r;
  \CTf''''''''_f''''''''_Int_Int_t  _12_d;
  logic _12_r;
  assign _12_r = 1'd1;
  \CTf''''''''_f''''''''_Int_Int_t  \lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int3_d ;
  logic \lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int3_r ;
  \CTf''''''''_f''''''''_Int_Int_t  \lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int2_d ;
  logic \lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int2_r ;
  \CTf''''''''_f''''''''_Int_Int_t  \lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int1_d ;
  logic \lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int1_r ;
  \CTf''''''''_f''''''''_Int_Int_t  \lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int0_d ;
  logic \lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int0_r ;
  Go_t _11_d;
  logic _11_r;
  assign _11_r = 1'd1;
  Go_t \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int3_d ;
  logic \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int3_r ;
  Go_t \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int2_d ;
  logic \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int2_r ;
  Go_t \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int1_d ;
  logic \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int1_r ;
  Go_t \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int0_d ;
  logic \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int0_r ;
  Go_t \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int0_1_argbuf_d ;
  logic \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int0_1_argbuf_r ;
  Go_t \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int1_1_argbuf_d ;
  logic \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int1_1_argbuf_r ;
  Go_t \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int2_1_argbuf_d ;
  logic \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int2_1_argbuf_r ;
  Go_t \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int3_1_argbuf_d ;
  logic \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int3_1_argbuf_r ;
  Pointer_QTree_Int_t \lizzieLet39_4Lf''''''''_f''''''''_Int_Intsbos_d ;
  logic \lizzieLet39_4Lf''''''''_f''''''''_Int_Intsbos_r ;
  Pointer_QTree_Int_t \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int3_d ;
  logic \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int3_r ;
  Pointer_QTree_Int_t \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int2_d ;
  logic \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int2_r ;
  Pointer_QTree_Int_t \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int1_d ;
  logic \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int1_r ;
  Pointer_QTree_Int_t \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int0_d ;
  logic \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int0_r ;
  QTree_Int_t \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int0_1es_5_2_1es_6_4_1es_7_4_1QNode_Int_d ;
  logic \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int0_1es_5_2_1es_6_4_1es_7_4_1QNode_Int_r ;
  QTree_Int_t lizzieLet43_1_argbuf_d;
  logic lizzieLet43_1_argbuf_r;
  \CTf''''''''_f''''''''_Int_Int_t  \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int1_1es_6_3_1es_7_3_1sc_0_9_1Lcall_f''''''''_f''''''''_Int_Int0_d ;
  logic \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int1_1es_6_3_1es_7_3_1sc_0_9_1Lcall_f''''''''_f''''''''_Int_Int0_r ;
  \CTf''''''''_f''''''''_Int_Int_t  lizzieLet42_1_argbuf_d;
  logic lizzieLet42_1_argbuf_r;
  \CTf''''''''_f''''''''_Int_Int_t  \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int2_1es_7_2_1sc_0_8_1tla8y_2_1is_z_mapa8v_3_1op_mapa8w_3_1Lcall_f''''''''_f''''''''_Int_Int1_d ;
  logic \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int2_1es_7_2_1sc_0_8_1tla8y_2_1is_z_mapa8v_3_1op_mapa8w_3_1Lcall_f''''''''_f''''''''_Int_Int1_r ;
  \CTf''''''''_f''''''''_Int_Int_t  lizzieLet41_1_argbuf_d;
  logic lizzieLet41_1_argbuf_r;
  \CTf''''''''_f''''''''_Int_Int_t  \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int3_1sc_0_7_1tla8y_1_1is_z_mapa8v_2_1op_mapa8w_2_1tra8z_1_1Lcall_f''''''''_f''''''''_Int_Int2_d ;
  logic \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int3_1sc_0_7_1tla8y_1_1is_z_mapa8v_2_1op_mapa8w_2_1tra8z_1_1Lcall_f''''''''_f''''''''_Int_Int2_r ;
  \CTf''''''''_f''''''''_Int_Int_t  lizzieLet40_1_argbuf_d;
  logic lizzieLet40_1_argbuf_r;
  Pointer_QTree_Int_t \lizzieLet39_4Lf''''''''_f''''''''_Int_Intsbos_1_merge_merge_fork_1_d ;
  logic \lizzieLet39_4Lf''''''''_f''''''''_Int_Intsbos_1_merge_merge_fork_1_r ;
  Pointer_QTree_Int_t \lizzieLet39_4Lf''''''''_f''''''''_Int_Intsbos_1_merge_merge_fork_2_d ;
  logic \lizzieLet39_4Lf''''''''_f''''''''_Int_Intsbos_1_merge_merge_fork_2_r ;
  Go_t \call_f''''''''_f''''''''_Int_Int_goConst_d ;
  logic \call_f''''''''_f''''''''_Int_Int_goConst_r ;
  Go_t lizzieLet3_1MyFalse_d;
  logic lizzieLet3_1MyFalse_r;
  Go_t lizzieLet3_1MyTrue_d;
  logic lizzieLet3_1MyTrue_r;
  MyBool_t lizzieLet3_1MyFalse_1MyFalse_d;
  logic lizzieLet3_1MyFalse_1MyFalse_r;
  MyBool_t lizzieLet3_1MyTrue_1MyTrue_d;
  logic lizzieLet3_1MyTrue_1MyTrue_r;
  MyBool_t lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_d;
  logic lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_r;
  Pointer_QTree_Int_t es_28_destruct_d;
  logic es_28_destruct_r;
  Pointer_QTree_Int_t es_29_1_destruct_d;
  logic es_29_1_destruct_r;
  Pointer_QTree_Int_t es_30_2_destruct_d;
  logic es_30_2_destruct_r;
  Pointer_CTf_f_Int_Int_t sc_0_14_destruct_d;
  logic sc_0_14_destruct_r;
  Pointer_QTree_Int_t es_29_destruct_d;
  logic es_29_destruct_r;
  Pointer_QTree_Int_t es_30_1_destruct_d;
  logic es_30_1_destruct_r;
  Pointer_CTf_f_Int_Int_t sc_0_13_destruct_d;
  logic sc_0_13_destruct_r;
  Pointer_QTree_Int_t q1a8T_3_destruct_d;
  logic q1a8T_3_destruct_r;
  Pointer_QTree_Int_t t1a8Y_3_destruct_d;
  logic t1a8Y_3_destruct_r;
  MyDTInt_Bool_t is_z_mapa8E_4_destruct_d;
  logic is_z_mapa8E_4_destruct_r;
  MyDTInt_Int_t op_mapa8F_4_destruct_d;
  logic op_mapa8F_4_destruct_r;
  MyDTInt_Bool_t is_z_adda8G_4_destruct_d;
  logic is_z_adda8G_4_destruct_r;
  MyDTInt_Int_Int_t op_adda8H_4_destruct_d;
  logic op_adda8H_4_destruct_r;
  Pointer_QTree_Int_t es_30_destruct_d;
  logic es_30_destruct_r;
  Pointer_CTf_f_Int_Int_t sc_0_12_destruct_d;
  logic sc_0_12_destruct_r;
  Pointer_QTree_Int_t q1a8T_2_destruct_d;
  logic q1a8T_2_destruct_r;
  Pointer_QTree_Int_t t1a8Y_2_destruct_d;
  logic t1a8Y_2_destruct_r;
  MyDTInt_Bool_t is_z_mapa8E_3_destruct_d;
  logic is_z_mapa8E_3_destruct_r;
  MyDTInt_Int_t op_mapa8F_3_destruct_d;
  logic op_mapa8F_3_destruct_r;
  MyDTInt_Bool_t is_z_adda8G_3_destruct_d;
  logic is_z_adda8G_3_destruct_r;
  MyDTInt_Int_Int_t op_adda8H_3_destruct_d;
  logic op_adda8H_3_destruct_r;
  Pointer_QTree_Int_t q2a8U_2_destruct_d;
  logic q2a8U_2_destruct_r;
  Pointer_QTree_Int_t t2a8Z_2_destruct_d;
  logic t2a8Z_2_destruct_r;
  Pointer_CTf_f_Int_Int_t sc_0_11_destruct_d;
  logic sc_0_11_destruct_r;
  Pointer_QTree_Int_t q1a8T_1_destruct_d;
  logic q1a8T_1_destruct_r;
  Pointer_QTree_Int_t t1a8Y_1_destruct_d;
  logic t1a8Y_1_destruct_r;
  MyDTInt_Bool_t is_z_mapa8E_2_destruct_d;
  logic is_z_mapa8E_2_destruct_r;
  MyDTInt_Int_t op_mapa8F_2_destruct_d;
  logic op_mapa8F_2_destruct_r;
  MyDTInt_Bool_t is_z_adda8G_2_destruct_d;
  logic is_z_adda8G_2_destruct_r;
  MyDTInt_Int_Int_t op_adda8H_2_destruct_d;
  logic op_adda8H_2_destruct_r;
  Pointer_QTree_Int_t q2a8U_1_destruct_d;
  logic q2a8U_1_destruct_r;
  Pointer_QTree_Int_t t2a8Z_1_destruct_d;
  logic t2a8Z_1_destruct_r;
  Pointer_QTree_Int_t q3a8V_1_destruct_d;
  logic q3a8V_1_destruct_r;
  Pointer_QTree_Int_t t3a90_1_destruct_d;
  logic t3a90_1_destruct_r;
  CTf_f_Int_Int_t _10_d;
  logic _10_r;
  assign _10_r = 1'd1;
  CTf_f_Int_Int_t lizzieLet44_1Lcall_f_f_Int_Int3_d;
  logic lizzieLet44_1Lcall_f_f_Int_Int3_r;
  CTf_f_Int_Int_t lizzieLet44_1Lcall_f_f_Int_Int2_d;
  logic lizzieLet44_1Lcall_f_f_Int_Int2_r;
  CTf_f_Int_Int_t lizzieLet44_1Lcall_f_f_Int_Int1_d;
  logic lizzieLet44_1Lcall_f_f_Int_Int1_r;
  CTf_f_Int_Int_t lizzieLet44_1Lcall_f_f_Int_Int0_d;
  logic lizzieLet44_1Lcall_f_f_Int_Int0_r;
  Go_t _9_d;
  logic _9_r;
  assign _9_r = 1'd1;
  Go_t lizzieLet44_3Lcall_f_f_Int_Int3_d;
  logic lizzieLet44_3Lcall_f_f_Int_Int3_r;
  Go_t lizzieLet44_3Lcall_f_f_Int_Int2_d;
  logic lizzieLet44_3Lcall_f_f_Int_Int2_r;
  Go_t lizzieLet44_3Lcall_f_f_Int_Int1_d;
  logic lizzieLet44_3Lcall_f_f_Int_Int1_r;
  Go_t lizzieLet44_3Lcall_f_f_Int_Int0_d;
  logic lizzieLet44_3Lcall_f_f_Int_Int0_r;
  Go_t lizzieLet44_3Lcall_f_f_Int_Int0_1_argbuf_d;
  logic lizzieLet44_3Lcall_f_f_Int_Int0_1_argbuf_r;
  Go_t lizzieLet44_3Lcall_f_f_Int_Int1_1_argbuf_d;
  logic lizzieLet44_3Lcall_f_f_Int_Int1_1_argbuf_r;
  Go_t lizzieLet44_3Lcall_f_f_Int_Int2_1_argbuf_d;
  logic lizzieLet44_3Lcall_f_f_Int_Int2_1_argbuf_r;
  Go_t lizzieLet44_3Lcall_f_f_Int_Int3_1_argbuf_d;
  logic lizzieLet44_3Lcall_f_f_Int_Int3_1_argbuf_r;
  Pointer_QTree_Int_t lizzieLet44_4Lf_f_Int_Intsbos_d;
  logic lizzieLet44_4Lf_f_Int_Intsbos_r;
  Pointer_QTree_Int_t lizzieLet44_4Lcall_f_f_Int_Int3_d;
  logic lizzieLet44_4Lcall_f_f_Int_Int3_r;
  Pointer_QTree_Int_t lizzieLet44_4Lcall_f_f_Int_Int2_d;
  logic lizzieLet44_4Lcall_f_f_Int_Int2_r;
  Pointer_QTree_Int_t lizzieLet44_4Lcall_f_f_Int_Int1_d;
  logic lizzieLet44_4Lcall_f_f_Int_Int1_r;
  Pointer_QTree_Int_t lizzieLet44_4Lcall_f_f_Int_Int0_d;
  logic lizzieLet44_4Lcall_f_f_Int_Int0_r;
  QTree_Int_t lizzieLet44_4Lcall_f_f_Int_Int0_1es_28_1es_29_1_1es_30_2_1QNode_Int_d;
  logic lizzieLet44_4Lcall_f_f_Int_Int0_1es_28_1es_29_1_1es_30_2_1QNode_Int_r;
  QTree_Int_t lizzieLet48_1_argbuf_d;
  logic lizzieLet48_1_argbuf_r;
  CTf_f_Int_Int_t lizzieLet44_4Lcall_f_f_Int_Int1_1es_29_1es_30_1_1sc_0_13_1Lcall_f_f_Int_Int0_d;
  logic lizzieLet44_4Lcall_f_f_Int_Int1_1es_29_1es_30_1_1sc_0_13_1Lcall_f_f_Int_Int0_r;
  CTf_f_Int_Int_t lizzieLet47_1_argbuf_d;
  logic lizzieLet47_1_argbuf_r;
  CTf_f_Int_Int_t lizzieLet44_4Lcall_f_f_Int_Int2_1es_30_1sc_0_12_1q1a8T_2_1t1a8Y_2_1is_z_mapa8E_3_1op_mapa8F_3_1is_z_adda8G_3_1op_adda8H_3_1Lcall_f_f_Int_Int1_d;
  logic lizzieLet44_4Lcall_f_f_Int_Int2_1es_30_1sc_0_12_1q1a8T_2_1t1a8Y_2_1is_z_mapa8E_3_1op_mapa8F_3_1is_z_adda8G_3_1op_adda8H_3_1Lcall_f_f_Int_Int1_r;
  CTf_f_Int_Int_t lizzieLet46_1_argbuf_d;
  logic lizzieLet46_1_argbuf_r;
  CTf_f_Int_Int_t lizzieLet44_4Lcall_f_f_Int_Int3_1sc_0_11_1q1a8T_1_1t1a8Y_1_1is_z_mapa8E_2_1op_mapa8F_2_1is_z_adda8G_2_1op_adda8H_2_1q2a8U_1_1t2a8Z_1_1Lcall_f_f_Int_Int2_d;
  logic lizzieLet44_4Lcall_f_f_Int_Int3_1sc_0_11_1q1a8T_1_1t1a8Y_1_1is_z_mapa8E_2_1op_mapa8F_2_1is_z_adda8G_2_1op_adda8H_2_1q2a8U_1_1t2a8Z_1_1Lcall_f_f_Int_Int2_r;
  CTf_f_Int_Int_t lizzieLet45_1_argbuf_d;
  logic lizzieLet45_1_argbuf_r;
  Pointer_QTree_Int_t lizzieLet44_4Lf_f_Int_Intsbos_1_merge_merge_merge_fork_1_d;
  logic lizzieLet44_4Lf_f_Int_Intsbos_1_merge_merge_merge_fork_1_r;
  Pointer_QTree_Int_t lizzieLet44_4Lf_f_Int_Intsbos_1_merge_merge_merge_fork_2_d;
  logic lizzieLet44_4Lf_f_Int_Intsbos_1_merge_merge_merge_fork_2_r;
  Go_t call_f_f_Int_Int_goConst_d;
  logic call_f_f_Int_Int_goConst_r;
  Pointer_QTree_Int_t f_f_Int_Int_resbuf_d;
  logic f_f_Int_Int_resbuf_r;
  Pointer_QTree_Int_t q1a84_destruct_d;
  logic q1a84_destruct_r;
  Pointer_QTree_Int_t q2a85_destruct_d;
  logic q2a85_destruct_r;
  Pointer_QTree_Int_t q3a86_destruct_d;
  logic q3a86_destruct_r;
  Pointer_QTree_Int_t q4a87_destruct_d;
  logic q4a87_destruct_r;
  QTree_Int_t _8_d;
  logic _8_r;
  assign _8_r = 1'd1;
  QTree_Int_t _7_d;
  logic _7_r;
  assign _7_r = 1'd1;
  QTree_Int_t lizzieLet4_1QNode_Int_d;
  logic lizzieLet4_1QNode_Int_r;
  QTree_Int_t _6_d;
  logic _6_r;
  assign _6_r = 1'd1;
  Go_t lizzieLet4_3QNone_Int_d;
  logic lizzieLet4_3QNone_Int_r;
  Go_t lizzieLet4_3QVal_Int_d;
  logic lizzieLet4_3QVal_Int_r;
  Go_t lizzieLet4_3QNode_Int_d;
  logic lizzieLet4_3QNode_Int_r;
  Go_t lizzieLet4_3QError_Int_d;
  logic lizzieLet4_3QError_Int_r;
  Go_t lizzieLet4_3QError_Int_1_d;
  logic lizzieLet4_3QError_Int_1_r;
  Go_t lizzieLet4_3QError_Int_2_d;
  logic lizzieLet4_3QError_Int_2_r;
  Go_t lizzieLet4_3QError_Int_1_argbuf_d;
  logic lizzieLet4_3QError_Int_1_argbuf_r;
  \Int#_t  lizzieLet4_3QError_Int_1_argbuf_0_d;
  logic lizzieLet4_3QError_Int_1_argbuf_0_r;
  \Int#_t  lizzieLet23_1_1_argbuf_d;
  logic lizzieLet23_1_1_argbuf_r;
  Go_t lizzieLet4_3QError_Int_2_argbuf_d;
  logic lizzieLet4_3QError_Int_2_argbuf_r;
  Go_t lizzieLet4_3QNode_Int_1_argbuf_d;
  logic lizzieLet4_3QNode_Int_1_argbuf_r;
  Go_t lizzieLet4_3QNone_Int_1_d;
  logic lizzieLet4_3QNone_Int_1_r;
  Go_t lizzieLet4_3QNone_Int_2_d;
  logic lizzieLet4_3QNone_Int_2_r;
  Go_t lizzieLet4_3QNone_Int_1_argbuf_d;
  logic lizzieLet4_3QNone_Int_1_argbuf_r;
  \Int#_t  lizzieLet4_3QNone_Int_1_argbuf_0_d;
  logic lizzieLet4_3QNone_Int_1_argbuf_0_r;
  \Int#_t  lizzieLet23_1_argbuf_d;
  logic lizzieLet23_1_argbuf_r;
  Go_t lizzieLet4_3QNone_Int_2_argbuf_d;
  logic lizzieLet4_3QNone_Int_2_argbuf_r;
  C4_t go_15_goMux_choice_d;
  logic go_15_goMux_choice_r;
  Go_t go_15_goMux_data_d;
  logic go_15_goMux_data_r;
  Go_t lizzieLet4_3QVal_Int_1_d;
  logic lizzieLet4_3QVal_Int_1_r;
  Go_t lizzieLet4_3QVal_Int_2_d;
  logic lizzieLet4_3QVal_Int_2_r;
  Go_t lizzieLet4_3QVal_Int_1_argbuf_d;
  logic lizzieLet4_3QVal_Int_1_argbuf_r;
  \Int#_t  lizzieLet4_3QVal_Int_1_argbuf_1_d;
  logic lizzieLet4_3QVal_Int_1_argbuf_1_r;
  \Int#_t  lizzieLet24_1_argbuf_d;
  logic lizzieLet24_1_argbuf_r;
  Go_t lizzieLet4_3QVal_Int_2_argbuf_d;
  logic lizzieLet4_3QVal_Int_2_argbuf_r;
  Pointer_CT$wnnz_t lizzieLet4_4QNone_Int_d;
  logic lizzieLet4_4QNone_Int_r;
  Pointer_CT$wnnz_t lizzieLet4_4QVal_Int_d;
  logic lizzieLet4_4QVal_Int_r;
  Pointer_CT$wnnz_t lizzieLet4_4QNode_Int_d;
  logic lizzieLet4_4QNode_Int_r;
  Pointer_CT$wnnz_t lizzieLet4_4QError_Int_d;
  logic lizzieLet4_4QError_Int_r;
  Pointer_CT$wnnz_t lizzieLet4_4QError_Int_1_argbuf_d;
  logic lizzieLet4_4QError_Int_1_argbuf_r;
  CT$wnnz_t lizzieLet4_4QNode_Int_1q4a87_1q3a86_1q2a85_1Lcall_$wnnz3_d;
  logic lizzieLet4_4QNode_Int_1q4a87_1q3a86_1q2a85_1Lcall_$wnnz3_r;
  CT$wnnz_t lizzieLet5_1_argbuf_d;
  logic lizzieLet5_1_argbuf_r;
  Pointer_CT$wnnz_t lizzieLet4_4QNone_Int_1_argbuf_d;
  logic lizzieLet4_4QNone_Int_1_argbuf_r;
  Pointer_CT$wnnz_t lizzieLet4_4QVal_Int_1_argbuf_d;
  logic lizzieLet4_4QVal_Int_1_argbuf_r;
  Pointer_QTree_Int_t tla8y_destruct_d;
  logic tla8y_destruct_r;
  Pointer_QTree_Int_t tra8z_destruct_d;
  logic tra8z_destruct_r;
  Pointer_QTree_Int_t bla8A_destruct_d;
  logic bla8A_destruct_r;
  Pointer_QTree_Int_t bra8B_destruct_d;
  logic bra8B_destruct_r;
  Int_t va8x_destruct_d;
  logic va8x_destruct_r;
  QTree_Int_t _5_d;
  logic _5_r;
  assign _5_r = 1'd1;
  QTree_Int_t lizzieLet6_1QVal_Int_d;
  logic lizzieLet6_1QVal_Int_r;
  QTree_Int_t lizzieLet6_1QNode_Int_d;
  logic lizzieLet6_1QNode_Int_r;
  QTree_Int_t _4_d;
  logic _4_r;
  assign _4_r = 1'd1;
  Go_t lizzieLet6_3QNone_Int_d;
  logic lizzieLet6_3QNone_Int_r;
  Go_t lizzieLet6_3QVal_Int_d;
  logic lizzieLet6_3QVal_Int_r;
  Go_t lizzieLet6_3QNode_Int_d;
  logic lizzieLet6_3QNode_Int_r;
  Go_t lizzieLet6_3QError_Int_d;
  logic lizzieLet6_3QError_Int_r;
  Go_t lizzieLet6_3QError_Int_1_d;
  logic lizzieLet6_3QError_Int_1_r;
  Go_t lizzieLet6_3QError_Int_2_d;
  logic lizzieLet6_3QError_Int_2_r;
  QTree_Int_t lizzieLet6_3QError_Int_1QError_Int_d;
  logic lizzieLet6_3QError_Int_1QError_Int_r;
  QTree_Int_t lizzieLet11_1_argbuf_d;
  logic lizzieLet11_1_argbuf_r;
  Go_t lizzieLet6_3QError_Int_2_argbuf_d;
  logic lizzieLet6_3QError_Int_2_argbuf_r;
  Go_t lizzieLet6_3QNode_Int_1_argbuf_d;
  logic lizzieLet6_3QNode_Int_1_argbuf_r;
  Go_t lizzieLet6_3QNone_Int_1_d;
  logic lizzieLet6_3QNone_Int_1_r;
  Go_t lizzieLet6_3QNone_Int_2_d;
  logic lizzieLet6_3QNone_Int_2_r;
  QTree_Int_t lizzieLet6_3QNone_Int_1QNone_Int_d;
  logic lizzieLet6_3QNone_Int_1QNone_Int_r;
  QTree_Int_t lizzieLet7_1_argbuf_d;
  logic lizzieLet7_1_argbuf_r;
  Go_t lizzieLet6_3QNone_Int_2_argbuf_d;
  logic lizzieLet6_3QNone_Int_2_argbuf_r;
  C5_t go_16_goMux_choice_d;
  logic go_16_goMux_choice_r;
  Go_t go_16_goMux_data_d;
  logic go_16_goMux_data_r;
  Go_t lizzieLet6_3QVal_Int_1_d;
  logic lizzieLet6_3QVal_Int_1_r;
  Go_t lizzieLet6_3QVal_Int_2_d;
  logic lizzieLet6_3QVal_Int_2_r;
  Go_t lizzieLet6_3QVal_Int_3_d;
  logic lizzieLet6_3QVal_Int_3_r;
  Go_t lizzieLet6_3QVal_Int_1_argbuf_d;
  logic lizzieLet6_3QVal_Int_1_argbuf_r;
  TupGo___MyDTInt_Int___Int_t applyfnInt_Int_5TupGo___MyDTInt_Int___Int3_d;
  logic applyfnInt_Int_5TupGo___MyDTInt_Int___Int3_r;
  Go_t lizzieLet6_3QVal_Int_2_argbuf_d;
  logic lizzieLet6_3QVal_Int_2_argbuf_r;
  TupGo___MyDTInt_Bool___Int_t applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int2_d;
  logic applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int2_r;
  MyDTInt_Bool_t _3_d;
  logic _3_r;
  assign _3_r = 1'd1;
  MyDTInt_Bool_t lizzieLet6_4QVal_Int_d;
  logic lizzieLet6_4QVal_Int_r;
  MyDTInt_Bool_t lizzieLet6_4QNode_Int_d;
  logic lizzieLet6_4QNode_Int_r;
  MyDTInt_Bool_t _2_d;
  logic _2_r;
  assign _2_r = 1'd1;
  MyDTInt_Bool_t lizzieLet6_4QNode_Int_1_d;
  logic lizzieLet6_4QNode_Int_1_r;
  MyDTInt_Bool_t lizzieLet6_4QNode_Int_2_d;
  logic lizzieLet6_4QNode_Int_2_r;
  MyDTInt_Bool_t lizzieLet6_4QNode_Int_2_argbuf_d;
  logic lizzieLet6_4QNode_Int_2_argbuf_r;
  MyDTInt_Bool_t lizzieLet6_4QVal_Int_1_argbuf_d;
  logic lizzieLet6_4QVal_Int_1_argbuf_r;
  MyDTInt_Int_t _1_d;
  logic _1_r;
  assign _1_r = 1'd1;
  MyDTInt_Int_t lizzieLet6_5QVal_Int_d;
  logic lizzieLet6_5QVal_Int_r;
  MyDTInt_Int_t lizzieLet6_5QNode_Int_d;
  logic lizzieLet6_5QNode_Int_r;
  MyDTInt_Int_t _0_d;
  logic _0_r;
  assign _0_r = 1'd1;
  MyDTInt_Int_t lizzieLet6_5QNode_Int_1_d;
  logic lizzieLet6_5QNode_Int_1_r;
  MyDTInt_Int_t lizzieLet6_5QNode_Int_2_d;
  logic lizzieLet6_5QNode_Int_2_r;
  MyDTInt_Int_t lizzieLet6_5QNode_Int_2_argbuf_d;
  logic lizzieLet6_5QNode_Int_2_argbuf_r;
  MyDTInt_Int_t lizzieLet6_5QVal_Int_1_d;
  logic lizzieLet6_5QVal_Int_1_r;
  MyDTInt_Int_t lizzieLet6_5QVal_Int_2_d;
  logic lizzieLet6_5QVal_Int_2_r;
  MyDTInt_Int_t lizzieLet6_5QVal_Int_1_argbuf_d;
  logic lizzieLet6_5QVal_Int_1_argbuf_r;
  \Pointer_CTf''''''''_f''''''''_Int_Int_t  lizzieLet6_6QNone_Int_d;
  logic lizzieLet6_6QNone_Int_r;
  \Pointer_CTf''''''''_f''''''''_Int_Int_t  lizzieLet6_6QVal_Int_d;
  logic lizzieLet6_6QVal_Int_r;
  \Pointer_CTf''''''''_f''''''''_Int_Int_t  lizzieLet6_6QNode_Int_d;
  logic lizzieLet6_6QNode_Int_r;
  \Pointer_CTf''''''''_f''''''''_Int_Int_t  lizzieLet6_6QError_Int_d;
  logic lizzieLet6_6QError_Int_r;
  \Pointer_CTf''''''''_f''''''''_Int_Int_t  lizzieLet6_6QError_Int_1_argbuf_d;
  logic lizzieLet6_6QError_Int_1_argbuf_r;
  \CTf''''''''_f''''''''_Int_Int_t  \lizzieLet6_6QNode_Int_1tla8y_1lizzieLet6_4QNode_Int_1lizzieLet6_5QNode_Int_1tra8z_1bla8A_1Lcall_f''''''''_f''''''''_Int_Int3_d ;
  logic \lizzieLet6_6QNode_Int_1tla8y_1lizzieLet6_4QNode_Int_1lizzieLet6_5QNode_Int_1tra8z_1bla8A_1Lcall_f''''''''_f''''''''_Int_Int3_r ;
  \CTf''''''''_f''''''''_Int_Int_t  lizzieLet10_1_argbuf_d;
  logic lizzieLet10_1_argbuf_r;
  \Pointer_CTf''''''''_f''''''''_Int_Int_t  lizzieLet6_6QNone_Int_1_argbuf_d;
  logic lizzieLet6_6QNone_Int_1_argbuf_r;
  Pointer_QTree_Int_t m1a8C_1_argbuf_d;
  logic m1a8C_1_argbuf_r;
  Pointer_QTree_Int_t m2a8D_1_argbuf_d;
  logic m2a8D_1_argbuf_r;
  MyDTInt_Int_Int_t op_adda8H_2_2_argbuf_d;
  logic op_adda8H_2_2_argbuf_r;
  MyDTInt_Int_Int_t op_adda8H_2_1_d;
  logic op_adda8H_2_1_r;
  MyDTInt_Int_Int_t op_adda8H_2_2_d;
  logic op_adda8H_2_2_r;
  MyDTInt_Int_Int_t op_adda8H_3_2_argbuf_d;
  logic op_adda8H_3_2_argbuf_r;
  MyDTInt_Int_Int_t op_adda8H_3_1_d;
  logic op_adda8H_3_1_r;
  MyDTInt_Int_Int_t op_adda8H_3_2_d;
  logic op_adda8H_3_2_r;
  MyDTInt_Int_Int_t op_adda8H_4_1_argbuf_d;
  logic op_adda8H_4_1_argbuf_r;
  MyDTInt_Int_t op_mapa8F_2_2_argbuf_d;
  logic op_mapa8F_2_2_argbuf_r;
  MyDTInt_Int_t op_mapa8F_2_1_d;
  logic op_mapa8F_2_1_r;
  MyDTInt_Int_t op_mapa8F_2_2_d;
  logic op_mapa8F_2_2_r;
  MyDTInt_Int_t op_mapa8F_3_2_argbuf_d;
  logic op_mapa8F_3_2_argbuf_r;
  MyDTInt_Int_t op_mapa8F_3_1_d;
  logic op_mapa8F_3_1_r;
  MyDTInt_Int_t op_mapa8F_3_2_d;
  logic op_mapa8F_3_2_r;
  MyDTInt_Int_t op_mapa8F_4_1_argbuf_d;
  logic op_mapa8F_4_1_argbuf_r;
  MyDTInt_Int_t op_mapa8w_2_2_argbuf_d;
  logic op_mapa8w_2_2_argbuf_r;
  MyDTInt_Int_t op_mapa8w_2_1_d;
  logic op_mapa8w_2_1_r;
  MyDTInt_Int_t op_mapa8w_2_2_d;
  logic op_mapa8w_2_2_r;
  MyDTInt_Int_t op_mapa8w_3_2_argbuf_d;
  logic op_mapa8w_3_2_argbuf_r;
  MyDTInt_Int_t op_mapa8w_3_1_d;
  logic op_mapa8w_3_1_r;
  MyDTInt_Int_t op_mapa8w_3_2_d;
  logic op_mapa8w_3_2_r;
  MyDTInt_Int_t op_mapa8w_4_1_argbuf_d;
  logic op_mapa8w_4_1_argbuf_r;
  Pointer_QTree_Int_t q1a84_1_argbuf_d;
  logic q1a84_1_argbuf_r;
  Pointer_QTree_Int_t q1a8T_3_1_argbuf_d;
  logic q1a8T_3_1_argbuf_r;
  Pointer_QTree_Int_t q2a85_1_1_argbuf_d;
  logic q2a85_1_1_argbuf_r;
  Pointer_QTree_Int_t q2a8U_2_1_argbuf_d;
  logic q2a8U_2_1_argbuf_r;
  Pointer_QTree_Int_t q3a86_2_1_argbuf_d;
  logic q3a86_2_1_argbuf_r;
  Pointer_QTree_Int_t q3a8V_1_1_argbuf_d;
  logic q3a8V_1_1_argbuf_r;
  Pointer_QTree_Int_t q4a87_3_1_argbuf_d;
  logic q4a87_3_1_argbuf_r;
  Pointer_QTree_Int_t q4a8u_1_argbuf_d;
  logic q4a8u_1_argbuf_r;
  CT$wnnz_t readPointer_CT$wnnzscfarg_0_1_argbuf_rwb_d;
  logic readPointer_CT$wnnzscfarg_0_1_argbuf_rwb_r;
  CT$wnnz_t lizzieLet35_1_d;
  logic lizzieLet35_1_r;
  CT$wnnz_t lizzieLet35_2_d;
  logic lizzieLet35_2_r;
  CT$wnnz_t lizzieLet35_3_d;
  logic lizzieLet35_3_r;
  CT$wnnz_t lizzieLet35_4_d;
  logic lizzieLet35_4_r;
  \CTf''''''''_f''''''''_Int_Int_t  \readPointer_CTf''''''''_f''''''''_Int_Intscfarg_0_1_1_argbuf_rwb_d ;
  logic \readPointer_CTf''''''''_f''''''''_Int_Intscfarg_0_1_1_argbuf_rwb_r ;
  \CTf''''''''_f''''''''_Int_Int_t  lizzieLet39_1_d;
  logic lizzieLet39_1_r;
  \CTf''''''''_f''''''''_Int_Int_t  lizzieLet39_2_d;
  logic lizzieLet39_2_r;
  \CTf''''''''_f''''''''_Int_Int_t  lizzieLet39_3_d;
  logic lizzieLet39_3_r;
  \CTf''''''''_f''''''''_Int_Int_t  lizzieLet39_4_d;
  logic lizzieLet39_4_r;
  CTf_f_Int_Int_t readPointer_CTf_f_Int_Intscfarg_0_2_1_argbuf_rwb_d;
  logic readPointer_CTf_f_Int_Intscfarg_0_2_1_argbuf_rwb_r;
  CTf_f_Int_Int_t lizzieLet44_1_d;
  logic lizzieLet44_1_r;
  CTf_f_Int_Int_t lizzieLet44_2_d;
  logic lizzieLet44_2_r;
  CTf_f_Int_Int_t lizzieLet44_3_d;
  logic lizzieLet44_3_r;
  CTf_f_Int_Int_t lizzieLet44_4_d;
  logic lizzieLet44_4_r;
  QTree_Int_t readPointer_QTree_Intm1a8C_1_argbuf_rwb_d;
  logic readPointer_QTree_Intm1a8C_1_argbuf_rwb_r;
  QTree_Int_t lizzieLet12_1_d;
  logic lizzieLet12_1_r;
  QTree_Int_t lizzieLet12_2_d;
  logic lizzieLet12_2_r;
  QTree_Int_t lizzieLet12_3_d;
  logic lizzieLet12_3_r;
  QTree_Int_t lizzieLet12_4_d;
  logic lizzieLet12_4_r;
  QTree_Int_t lizzieLet12_5_d;
  logic lizzieLet12_5_r;
  QTree_Int_t lizzieLet12_6_d;
  logic lizzieLet12_6_r;
  QTree_Int_t lizzieLet12_7_d;
  logic lizzieLet12_7_r;
  QTree_Int_t lizzieLet12_8_d;
  logic lizzieLet12_8_r;
  QTree_Int_t lizzieLet12_9_d;
  logic lizzieLet12_9_r;
  QTree_Int_t readPointer_QTree_Intm2a8D_1_argbuf_rwb_d;
  logic readPointer_QTree_Intm2a8D_1_argbuf_rwb_r;
  QTree_Int_t readPointer_QTree_Intq4a8u_1_argbuf_rwb_d;
  logic readPointer_QTree_Intq4a8u_1_argbuf_rwb_r;
  QTree_Int_t lizzieLet6_1_d;
  logic lizzieLet6_1_r;
  QTree_Int_t lizzieLet6_2_d;
  logic lizzieLet6_2_r;
  QTree_Int_t lizzieLet6_3_d;
  logic lizzieLet6_3_r;
  QTree_Int_t lizzieLet6_4_d;
  logic lizzieLet6_4_r;
  QTree_Int_t lizzieLet6_5_d;
  logic lizzieLet6_5_r;
  QTree_Int_t lizzieLet6_6_d;
  logic lizzieLet6_6_r;
  QTree_Int_t readPointer_QTree_IntwsiX_1_1_argbuf_rwb_d;
  logic readPointer_QTree_IntwsiX_1_1_argbuf_rwb_r;
  QTree_Int_t lizzieLet4_1_d;
  logic lizzieLet4_1_r;
  QTree_Int_t lizzieLet4_2_d;
  logic lizzieLet4_2_r;
  QTree_Int_t lizzieLet4_3_d;
  logic lizzieLet4_3_r;
  QTree_Int_t lizzieLet4_4_d;
  logic lizzieLet4_4_r;
  \Pointer_CTf''''''''_f''''''''_Int_Int_t  sc_0_10_1_argbuf_d;
  logic sc_0_10_1_argbuf_r;
  Pointer_CTf_f_Int_Int_t sc_0_14_1_argbuf_d;
  logic sc_0_14_1_argbuf_r;
  Pointer_CT$wnnz_t sc_0_6_1_argbuf_d;
  logic sc_0_6_1_argbuf_r;
  \Pointer_CTf''''''''_f''''''''_Int_Int_t  scfarg_0_1_1_argbuf_d;
  logic scfarg_0_1_1_argbuf_r;
  Pointer_CTf_f_Int_Int_t scfarg_0_2_1_argbuf_d;
  logic scfarg_0_2_1_argbuf_r;
  Pointer_CT$wnnz_t scfarg_0_1_argbuf_d;
  logic scfarg_0_1_argbuf_r;
  Pointer_QTree_Int_t t1a8Y_3_1_argbuf_d;
  logic t1a8Y_3_1_argbuf_r;
  Pointer_QTree_Int_t t2a8Z_2_1_argbuf_d;
  logic t2a8Z_2_1_argbuf_r;
  Pointer_QTree_Int_t t3a90_1_1_argbuf_d;
  logic t3a90_1_1_argbuf_r;
  Pointer_QTree_Int_t t4a91_1_argbuf_d;
  logic t4a91_1_argbuf_r;
  Pointer_QTree_Int_t tla8J_1_argbuf_d;
  logic tla8J_1_argbuf_r;
  Pointer_QTree_Int_t tla8y_3_1_argbuf_d;
  logic tla8y_3_1_argbuf_r;
  Pointer_QTree_Int_t tra8K_1_argbuf_d;
  logic tra8K_1_argbuf_r;
  Pointer_QTree_Int_t tra8z_2_1_argbuf_d;
  logic tra8z_2_1_argbuf_r;
  Int_t va8I_1_argbuf_d;
  logic va8I_1_argbuf_r;
  Int_t va8I_1_d;
  logic va8I_1_r;
  Int_t va8I_2_d;
  logic va8I_2_r;
  Int_t va8O_1_argbuf_d;
  logic va8O_1_argbuf_r;
  Int_t va8O_1_d;
  logic va8O_1_r;
  Int_t va8O_2_d;
  logic va8O_2_r;
  Int_t va8x_1_argbuf_d;
  logic va8x_1_argbuf_r;
  Int_t va8x_1_d;
  logic va8x_1_r;
  Int_t va8x_2_d;
  logic va8x_2_r;
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet0_1_argbuf_rwb_d;
  logic writeCT$wnnzlizzieLet0_1_argbuf_rwb_r;
  Pointer_CT$wnnz_t lizzieLet25_1_argbuf_d;
  logic lizzieLet25_1_argbuf_r;
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet36_1_argbuf_rwb_d;
  logic writeCT$wnnzlizzieLet36_1_argbuf_rwb_r;
  Pointer_CT$wnnz_t sca2_1_argbuf_d;
  logic sca2_1_argbuf_r;
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet37_1_argbuf_rwb_d;
  logic writeCT$wnnzlizzieLet37_1_argbuf_rwb_r;
  Pointer_CT$wnnz_t sca1_1_argbuf_d;
  logic sca1_1_argbuf_r;
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet38_1_argbuf_rwb_d;
  logic writeCT$wnnzlizzieLet38_1_argbuf_rwb_r;
  Pointer_CT$wnnz_t sca0_1_argbuf_d;
  logic sca0_1_argbuf_r;
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet5_1_argbuf_rwb_d;
  logic writeCT$wnnzlizzieLet5_1_argbuf_rwb_r;
  Pointer_CT$wnnz_t sca3_1_argbuf_d;
  logic sca3_1_argbuf_r;
  \Pointer_CTf''''''''_f''''''''_Int_Int_t  \writeCTf''''''''_f''''''''_Int_IntlizzieLet10_1_argbuf_rwb_d ;
  logic \writeCTf''''''''_f''''''''_Int_IntlizzieLet10_1_argbuf_rwb_r ;
  \Pointer_CTf''''''''_f''''''''_Int_Int_t  sca3_1_1_argbuf_d;
  logic sca3_1_1_argbuf_r;
  \Pointer_CTf''''''''_f''''''''_Int_Int_t  \writeCTf''''''''_f''''''''_Int_IntlizzieLet33_1_argbuf_rwb_d ;
  logic \writeCTf''''''''_f''''''''_Int_IntlizzieLet33_1_argbuf_rwb_r ;
  \Pointer_CTf''''''''_f''''''''_Int_Int_t  lizzieLet5_1_1_argbuf_d;
  logic lizzieLet5_1_1_argbuf_r;
  \Pointer_CTf''''''''_f''''''''_Int_Int_t  \writeCTf''''''''_f''''''''_Int_IntlizzieLet40_1_argbuf_rwb_d ;
  logic \writeCTf''''''''_f''''''''_Int_IntlizzieLet40_1_argbuf_rwb_r ;
  \Pointer_CTf''''''''_f''''''''_Int_Int_t  sca2_1_1_argbuf_d;
  logic sca2_1_1_argbuf_r;
  \Pointer_CTf''''''''_f''''''''_Int_Int_t  \writeCTf''''''''_f''''''''_Int_IntlizzieLet41_1_argbuf_rwb_d ;
  logic \writeCTf''''''''_f''''''''_Int_IntlizzieLet41_1_argbuf_rwb_r ;
  \Pointer_CTf''''''''_f''''''''_Int_Int_t  sca1_1_1_argbuf_d;
  logic sca1_1_1_argbuf_r;
  \Pointer_CTf''''''''_f''''''''_Int_Int_t  \writeCTf''''''''_f''''''''_Int_IntlizzieLet42_1_argbuf_rwb_d ;
  logic \writeCTf''''''''_f''''''''_Int_IntlizzieLet42_1_argbuf_rwb_r ;
  \Pointer_CTf''''''''_f''''''''_Int_Int_t  sca0_1_1_argbuf_d;
  logic sca0_1_1_argbuf_r;
  Pointer_CTf_f_Int_Int_t writeCTf_f_Int_IntlizzieLet30_1_argbuf_rwb_d;
  logic writeCTf_f_Int_IntlizzieLet30_1_argbuf_rwb_r;
  Pointer_CTf_f_Int_Int_t sca3_2_1_argbuf_d;
  logic sca3_2_1_argbuf_r;
  Pointer_CTf_f_Int_Int_t writeCTf_f_Int_IntlizzieLet34_1_argbuf_rwb_d;
  logic writeCTf_f_Int_IntlizzieLet34_1_argbuf_rwb_r;
  Pointer_CTf_f_Int_Int_t lizzieLet22_1_1_argbuf_d;
  logic lizzieLet22_1_1_argbuf_r;
  Pointer_CTf_f_Int_Int_t writeCTf_f_Int_IntlizzieLet45_1_argbuf_rwb_d;
  logic writeCTf_f_Int_IntlizzieLet45_1_argbuf_rwb_r;
  Pointer_CTf_f_Int_Int_t sca2_2_1_argbuf_d;
  logic sca2_2_1_argbuf_r;
  Pointer_CTf_f_Int_Int_t writeCTf_f_Int_IntlizzieLet46_1_argbuf_rwb_d;
  logic writeCTf_f_Int_IntlizzieLet46_1_argbuf_rwb_r;
  Pointer_CTf_f_Int_Int_t sca1_2_1_argbuf_d;
  logic sca1_2_1_argbuf_r;
  Pointer_CTf_f_Int_Int_t writeCTf_f_Int_IntlizzieLet47_1_argbuf_rwb_d;
  logic writeCTf_f_Int_IntlizzieLet47_1_argbuf_rwb_r;
  Pointer_CTf_f_Int_Int_t sca0_2_1_argbuf_d;
  logic sca0_2_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet11_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet11_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet4_1_1_argbuf_d;
  logic lizzieLet4_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet14_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet14_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet6_1_1_argbuf_d;
  logic lizzieLet6_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet15_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet15_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet7_1_1_argbuf_d;
  logic lizzieLet7_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet16_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet16_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet8_1_1_argbuf_d;
  logic lizzieLet8_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet17_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet17_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet9_1_1_argbuf_d;
  logic lizzieLet9_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet18_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet18_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet10_1_1_argbuf_d;
  logic lizzieLet10_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet20_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet20_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet11_1_1_argbuf_d;
  logic lizzieLet11_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet21_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet21_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet12_1_1_argbuf_d;
  logic lizzieLet12_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet22_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet22_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet13_1_1_argbuf_d;
  logic lizzieLet13_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet23_2_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet23_2_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet14_1_1_argbuf_d;
  logic lizzieLet14_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet24_1_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet24_1_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet15_1_1_argbuf_d;
  logic lizzieLet15_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet25_1_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet25_1_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet16_1_1_argbuf_d;
  logic lizzieLet16_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet26_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet26_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet17_1_1_argbuf_d;
  logic lizzieLet17_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet28_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet28_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet18_1_1_argbuf_d;
  logic lizzieLet18_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet29_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet29_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet19_1_argbuf_d;
  logic lizzieLet19_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet31_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet31_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet20_1_1_argbuf_d;
  logic lizzieLet20_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet32_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet32_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet21_1_1_argbuf_d;
  logic lizzieLet21_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet43_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet43_1_argbuf_rwb_r;
  Pointer_QTree_Int_t contRet_0_1_1_argbuf_d;
  logic contRet_0_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet48_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet48_1_argbuf_rwb_r;
  Pointer_QTree_Int_t contRet_0_2_1_argbuf_d;
  logic contRet_0_2_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet7_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet7_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet1_1_1_argbuf_d;
  logic lizzieLet1_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet8_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet8_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet2_1_1_argbuf_d;
  logic lizzieLet2_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet9_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet9_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet3_1_1_argbuf_d;
  logic lizzieLet3_1_1_argbuf_r;
  Pointer_QTree_Int_t wsiX_1_1_argbuf_d;
  logic wsiX_1_1_argbuf_r;
  CT$wnnz_t lizzieLet37_1_argbuf_d;
  logic lizzieLet37_1_argbuf_r;
  CT$wnnz_t wwsj0_2_1lizzieLet35_4Lcall_$wnnz2_1sc_0_4_1q4a87_2_1Lcall_$wnnz1_d;
  logic wwsj0_2_1lizzieLet35_4Lcall_$wnnz2_1sc_0_4_1q4a87_2_1Lcall_$wnnz1_r;
  CT$wnnz_t lizzieLet38_1_argbuf_d;
  logic lizzieLet38_1_argbuf_r;
  CT$wnnz_t wwsj0_3_1ww1Xju_1_1lizzieLet35_4Lcall_$wnnz1_1sc_0_5_1Lcall_$wnnz0_d;
  logic wwsj0_3_1ww1Xju_1_1lizzieLet35_4Lcall_$wnnz1_1sc_0_5_1Lcall_$wnnz0_r;
  \Int#_t  es_6_2_1ww2Xjx_1_1_Add32_d;
  logic es_6_2_1ww2Xjx_1_1_Add32_r;
  \Int#_t  wwsj0_4_1ww1Xju_2_1_Add32_d;
  logic wwsj0_4_1ww1Xju_2_1_Add32_r;
  Int_t \es_0_1_1I#_d ;
  logic \es_0_1_1I#_r ;
  \Int#_t  x1agS_1lizzieLet0_1_1_Add32_d;
  logic x1agS_1lizzieLet0_1_1_Add32_r;
  
  /* fork (Ty Go) : (sourceGo,Go) > [(go_1,Go),
                                (go_2,Go),
                                (go_3,Go),
                                (go_4,Go),
                                (go_5,Go),
                                (go_6,Go),
                                (go__7,Go),
                                (go__8,Go),
                                (go__9,Go),
                                (go__10,Go),
                                (go__11,Go),
                                (go__12,Go)] */
  logic [11:0] sourceGo_emitted;
  logic [11:0] sourceGo_done;
  assign go_1_d = (sourceGo_d[0] && (! sourceGo_emitted[0]));
  assign go_2_d = (sourceGo_d[0] && (! sourceGo_emitted[1]));
  assign go_3_d = (sourceGo_d[0] && (! sourceGo_emitted[2]));
  assign go_4_d = (sourceGo_d[0] && (! sourceGo_emitted[3]));
  assign go_5_d = (sourceGo_d[0] && (! sourceGo_emitted[4]));
  assign go_6_d = (sourceGo_d[0] && (! sourceGo_emitted[5]));
  assign go__7_d = (sourceGo_d[0] && (! sourceGo_emitted[6]));
  assign go__8_d = (sourceGo_d[0] && (! sourceGo_emitted[7]));
  assign go__9_d = (sourceGo_d[0] && (! sourceGo_emitted[8]));
  assign go__10_d = (sourceGo_d[0] && (! sourceGo_emitted[9]));
  assign go__11_d = (sourceGo_d[0] && (! sourceGo_emitted[10]));
  assign go__12_d = (sourceGo_d[0] && (! sourceGo_emitted[11]));
  assign sourceGo_done = (sourceGo_emitted | ({go__12_d[0],
                                               go__11_d[0],
                                               go__10_d[0],
                                               go__9_d[0],
                                               go__8_d[0],
                                               go__7_d[0],
                                               go_6_d[0],
                                               go_5_d[0],
                                               go_4_d[0],
                                               go_3_d[0],
                                               go_2_d[0],
                                               go_1_d[0]} & {go__12_r,
                                                             go__11_r,
                                                             go__10_r,
                                                             go__9_r,
                                                             go__8_r,
                                                             go__7_r,
                                                             go_6_r,
                                                             go_5_r,
                                                             go_4_r,
                                                             go_3_r,
                                                             go_2_r,
                                                             go_1_r}));
  assign sourceGo_r = (& sourceGo_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) sourceGo_emitted <= 12'd0;
    else
      sourceGo_emitted <= (sourceGo_r ? 12'd0 :
                           sourceGo_done);
  
  /* const (Ty Word16#,Lit 0) : (go__7,Go) > (initHP_CT$wnnz,Word16#) */
  assign initHP_CT$wnnz_d = {16'd0, go__7_d[0]};
  assign go__7_r = initHP_CT$wnnz_r;
  
  /* const (Ty Word16#,
       Lit 1) : (incrHP_CT$wnnz1,Go) > (incrHP_CT$wnnz,Word16#) */
  assign incrHP_CT$wnnz_d = {16'd1, incrHP_CT$wnnz1_d[0]};
  assign incrHP_CT$wnnz1_r = incrHP_CT$wnnz_r;
  
  /* merge (Ty Go) : [(go__8,Go),
                 (incrHP_CT$wnnz2,Go)] > (incrHP_mergeCT$wnnz,Go) */
  logic [1:0] incrHP_mergeCT$wnnz_selected;
  logic [1:0] incrHP_mergeCT$wnnz_select;
  always_comb
    begin
      incrHP_mergeCT$wnnz_selected = 2'd0;
      if ((| incrHP_mergeCT$wnnz_select))
        incrHP_mergeCT$wnnz_selected = incrHP_mergeCT$wnnz_select;
      else
        if (go__8_d[0]) incrHP_mergeCT$wnnz_selected[0] = 1'd1;
        else if (incrHP_CT$wnnz2_d[0])
          incrHP_mergeCT$wnnz_selected[1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeCT$wnnz_select <= 2'd0;
    else
      incrHP_mergeCT$wnnz_select <= (incrHP_mergeCT$wnnz_r ? 2'd0 :
                                     incrHP_mergeCT$wnnz_selected);
  always_comb
    if (incrHP_mergeCT$wnnz_selected[0])
      incrHP_mergeCT$wnnz_d = go__8_d;
    else if (incrHP_mergeCT$wnnz_selected[1])
      incrHP_mergeCT$wnnz_d = incrHP_CT$wnnz2_d;
    else incrHP_mergeCT$wnnz_d = 1'd0;
  assign {incrHP_CT$wnnz2_r,
          go__8_r} = (incrHP_mergeCT$wnnz_r ? incrHP_mergeCT$wnnz_selected :
                      2'd0);
  
  /* fork (Ty Go) : (incrHP_mergeCT$wnnz_buf,Go) > [(incrHP_CT$wnnz1,Go),
                                               (incrHP_CT$wnnz2,Go)] */
  logic [1:0] incrHP_mergeCT$wnnz_buf_emitted;
  logic [1:0] incrHP_mergeCT$wnnz_buf_done;
  assign incrHP_CT$wnnz1_d = (incrHP_mergeCT$wnnz_buf_d[0] && (! incrHP_mergeCT$wnnz_buf_emitted[0]));
  assign incrHP_CT$wnnz2_d = (incrHP_mergeCT$wnnz_buf_d[0] && (! incrHP_mergeCT$wnnz_buf_emitted[1]));
  assign incrHP_mergeCT$wnnz_buf_done = (incrHP_mergeCT$wnnz_buf_emitted | ({incrHP_CT$wnnz2_d[0],
                                                                             incrHP_CT$wnnz1_d[0]} & {incrHP_CT$wnnz2_r,
                                                                                                      incrHP_CT$wnnz1_r}));
  assign incrHP_mergeCT$wnnz_buf_r = (& incrHP_mergeCT$wnnz_buf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeCT$wnnz_buf_emitted <= 2'd0;
    else
      incrHP_mergeCT$wnnz_buf_emitted <= (incrHP_mergeCT$wnnz_buf_r ? 2'd0 :
                                          incrHP_mergeCT$wnnz_buf_done);
  
  /* op_add (Ty Word16#) : (incrHP_CT$wnnz,Word16#) (forkHP1_CT$wnnz,Word16#) > (addHP_CT$wnnz,Word16#) */
  assign addHP_CT$wnnz_d = {(incrHP_CT$wnnz_d[16:1] + forkHP1_CT$wnnz_d[16:1]),
                            (incrHP_CT$wnnz_d[0] && forkHP1_CT$wnnz_d[0])};
  assign {incrHP_CT$wnnz_r,
          forkHP1_CT$wnnz_r} = {2 {(addHP_CT$wnnz_r && addHP_CT$wnnz_d[0])}};
  
  /* merge (Ty Word16#) : [(initHP_CT$wnnz,Word16#),
                      (addHP_CT$wnnz,Word16#)] > (mergeHP_CT$wnnz,Word16#) */
  logic [1:0] mergeHP_CT$wnnz_selected;
  logic [1:0] mergeHP_CT$wnnz_select;
  always_comb
    begin
      mergeHP_CT$wnnz_selected = 2'd0;
      if ((| mergeHP_CT$wnnz_select))
        mergeHP_CT$wnnz_selected = mergeHP_CT$wnnz_select;
      else
        if (initHP_CT$wnnz_d[0]) mergeHP_CT$wnnz_selected[0] = 1'd1;
        else if (addHP_CT$wnnz_d[0]) mergeHP_CT$wnnz_selected[1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_CT$wnnz_select <= 2'd0;
    else
      mergeHP_CT$wnnz_select <= (mergeHP_CT$wnnz_r ? 2'd0 :
                                 mergeHP_CT$wnnz_selected);
  always_comb
    if (mergeHP_CT$wnnz_selected[0])
      mergeHP_CT$wnnz_d = initHP_CT$wnnz_d;
    else if (mergeHP_CT$wnnz_selected[1])
      mergeHP_CT$wnnz_d = addHP_CT$wnnz_d;
    else mergeHP_CT$wnnz_d = {16'd0, 1'd0};
  assign {addHP_CT$wnnz_r,
          initHP_CT$wnnz_r} = (mergeHP_CT$wnnz_r ? mergeHP_CT$wnnz_selected :
                               2'd0);
  
  /* buf (Ty Go) : (incrHP_mergeCT$wnnz,Go) > (incrHP_mergeCT$wnnz_buf,Go) */
  Go_t incrHP_mergeCT$wnnz_bufchan_d;
  logic incrHP_mergeCT$wnnz_bufchan_r;
  assign incrHP_mergeCT$wnnz_r = ((! incrHP_mergeCT$wnnz_bufchan_d[0]) || incrHP_mergeCT$wnnz_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeCT$wnnz_bufchan_d <= 1'd0;
    else
      if (incrHP_mergeCT$wnnz_r)
        incrHP_mergeCT$wnnz_bufchan_d <= incrHP_mergeCT$wnnz_d;
  Go_t incrHP_mergeCT$wnnz_bufchan_buf;
  assign incrHP_mergeCT$wnnz_bufchan_r = (! incrHP_mergeCT$wnnz_bufchan_buf[0]);
  assign incrHP_mergeCT$wnnz_buf_d = (incrHP_mergeCT$wnnz_bufchan_buf[0] ? incrHP_mergeCT$wnnz_bufchan_buf :
                                      incrHP_mergeCT$wnnz_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeCT$wnnz_bufchan_buf <= 1'd0;
    else
      if ((incrHP_mergeCT$wnnz_buf_r && incrHP_mergeCT$wnnz_bufchan_buf[0]))
        incrHP_mergeCT$wnnz_bufchan_buf <= 1'd0;
      else if (((! incrHP_mergeCT$wnnz_buf_r) && (! incrHP_mergeCT$wnnz_bufchan_buf[0])))
        incrHP_mergeCT$wnnz_bufchan_buf <= incrHP_mergeCT$wnnz_bufchan_d;
  
  /* buf (Ty Word16#) : (mergeHP_CT$wnnz,Word16#) > (mergeHP_CT$wnnz_buf,Word16#) */
  \Word16#_t  mergeHP_CT$wnnz_bufchan_d;
  logic mergeHP_CT$wnnz_bufchan_r;
  assign mergeHP_CT$wnnz_r = ((! mergeHP_CT$wnnz_bufchan_d[0]) || mergeHP_CT$wnnz_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_CT$wnnz_bufchan_d <= {16'd0, 1'd0};
    else
      if (mergeHP_CT$wnnz_r)
        mergeHP_CT$wnnz_bufchan_d <= mergeHP_CT$wnnz_d;
  \Word16#_t  mergeHP_CT$wnnz_bufchan_buf;
  assign mergeHP_CT$wnnz_bufchan_r = (! mergeHP_CT$wnnz_bufchan_buf[0]);
  assign mergeHP_CT$wnnz_buf_d = (mergeHP_CT$wnnz_bufchan_buf[0] ? mergeHP_CT$wnnz_bufchan_buf :
                                  mergeHP_CT$wnnz_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_CT$wnnz_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((mergeHP_CT$wnnz_buf_r && mergeHP_CT$wnnz_bufchan_buf[0]))
        mergeHP_CT$wnnz_bufchan_buf <= {16'd0, 1'd0};
      else if (((! mergeHP_CT$wnnz_buf_r) && (! mergeHP_CT$wnnz_bufchan_buf[0])))
        mergeHP_CT$wnnz_bufchan_buf <= mergeHP_CT$wnnz_bufchan_d;
  
  /* fork (Ty Word16#) : (mergeHP_CT$wnnz_buf,Word16#) > [(forkHP1_CT$wnnz,Word16#),
                                                     (forkHP1_CT$wnn2,Word16#),
                                                     (forkHP1_CT$wnn3,Word16#)] */
  logic [2:0] mergeHP_CT$wnnz_buf_emitted;
  logic [2:0] mergeHP_CT$wnnz_buf_done;
  assign forkHP1_CT$wnnz_d = {mergeHP_CT$wnnz_buf_d[16:1],
                              (mergeHP_CT$wnnz_buf_d[0] && (! mergeHP_CT$wnnz_buf_emitted[0]))};
  assign forkHP1_CT$wnn2_d = {mergeHP_CT$wnnz_buf_d[16:1],
                              (mergeHP_CT$wnnz_buf_d[0] && (! mergeHP_CT$wnnz_buf_emitted[1]))};
  assign forkHP1_CT$wnn3_d = {mergeHP_CT$wnnz_buf_d[16:1],
                              (mergeHP_CT$wnnz_buf_d[0] && (! mergeHP_CT$wnnz_buf_emitted[2]))};
  assign mergeHP_CT$wnnz_buf_done = (mergeHP_CT$wnnz_buf_emitted | ({forkHP1_CT$wnn3_d[0],
                                                                     forkHP1_CT$wnn2_d[0],
                                                                     forkHP1_CT$wnnz_d[0]} & {forkHP1_CT$wnn3_r,
                                                                                              forkHP1_CT$wnn2_r,
                                                                                              forkHP1_CT$wnnz_r}));
  assign mergeHP_CT$wnnz_buf_r = (& mergeHP_CT$wnnz_buf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_CT$wnnz_buf_emitted <= 3'd0;
    else
      mergeHP_CT$wnnz_buf_emitted <= (mergeHP_CT$wnnz_buf_r ? 3'd0 :
                                      mergeHP_CT$wnnz_buf_done);
  
  /* mergectrl (Ty C2,
           Ty MemIn_CT$wnnz) : [(dconReadIn_CT$wnnz,MemIn_CT$wnnz),
                                (dconWriteIn_CT$wnnz,MemIn_CT$wnnz)] > (memMergeChoice_CT$wnnz,C2) (memMergeIn_CT$wnnz,MemIn_CT$wnnz) */
  logic [1:0] dconReadIn_CT$wnnz_select_d;
  assign dconReadIn_CT$wnnz_select_d = ((| dconReadIn_CT$wnnz_select_q) ? dconReadIn_CT$wnnz_select_q :
                                        (dconReadIn_CT$wnnz_d[0] ? 2'd1 :
                                         (dconWriteIn_CT$wnnz_d[0] ? 2'd2 :
                                          2'd0)));
  logic [1:0] dconReadIn_CT$wnnz_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) dconReadIn_CT$wnnz_select_q <= 2'd0;
    else
      dconReadIn_CT$wnnz_select_q <= (dconReadIn_CT$wnnz_done ? 2'd0 :
                                      dconReadIn_CT$wnnz_select_d);
  logic [1:0] dconReadIn_CT$wnnz_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) dconReadIn_CT$wnnz_emit_q <= 2'd0;
    else
      dconReadIn_CT$wnnz_emit_q <= (dconReadIn_CT$wnnz_done ? 2'd0 :
                                    dconReadIn_CT$wnnz_emit_d);
  logic [1:0] dconReadIn_CT$wnnz_emit_d;
  assign dconReadIn_CT$wnnz_emit_d = (dconReadIn_CT$wnnz_emit_q | ({memMergeChoice_CT$wnnz_d[0],
                                                                    memMergeIn_CT$wnnz_d[0]} & {memMergeChoice_CT$wnnz_r,
                                                                                                memMergeIn_CT$wnnz_r}));
  logic dconReadIn_CT$wnnz_done;
  assign dconReadIn_CT$wnnz_done = (& dconReadIn_CT$wnnz_emit_d);
  assign {dconWriteIn_CT$wnnz_r,
          dconReadIn_CT$wnnz_r} = (dconReadIn_CT$wnnz_done ? dconReadIn_CT$wnnz_select_d :
                                   2'd0);
  assign memMergeIn_CT$wnnz_d = ((dconReadIn_CT$wnnz_select_d[0] && (! dconReadIn_CT$wnnz_emit_q[0])) ? dconReadIn_CT$wnnz_d :
                                 ((dconReadIn_CT$wnnz_select_d[1] && (! dconReadIn_CT$wnnz_emit_q[0])) ? dconWriteIn_CT$wnnz_d :
                                  {132'd0, 1'd0}));
  assign memMergeChoice_CT$wnnz_d = ((dconReadIn_CT$wnnz_select_d[0] && (! dconReadIn_CT$wnnz_emit_q[1])) ? C1_2_dc(1'd1) :
                                     ((dconReadIn_CT$wnnz_select_d[1] && (! dconReadIn_CT$wnnz_emit_q[1])) ? C2_2_dc(1'd1) :
                                      {1'd0, 1'd0}));
  
  /* bram (Ty MemIn_CT$wnnz,
      Ty MemOut_CT$wnnz) : (memMergeIn_CT$wnnz_dbuf,MemIn_CT$wnnz) > (memOut_CT$wnnz,MemOut_CT$wnnz) */
  logic [114:0] memMergeIn_CT$wnnz_dbuf_mem[65535:0];
  logic [15:0] memMergeIn_CT$wnnz_dbuf_address;
  logic [114:0] memMergeIn_CT$wnnz_dbuf_din;
  logic [114:0] memOut_CT$wnnz_q;
  logic memOut_CT$wnnz_valid;
  logic memMergeIn_CT$wnnz_dbuf_we;
  logic memOut_CT$wnnz_we;
  assign memMergeIn_CT$wnnz_dbuf_din = memMergeIn_CT$wnnz_dbuf_d[132:18];
  assign memMergeIn_CT$wnnz_dbuf_address = memMergeIn_CT$wnnz_dbuf_d[17:2];
  assign memMergeIn_CT$wnnz_dbuf_we = (memMergeIn_CT$wnnz_dbuf_d[1:1] && memMergeIn_CT$wnnz_dbuf_d[0]);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        memOut_CT$wnnz_we <= 1'd0;
        memOut_CT$wnnz_valid <= 1'd0;
      end
    else
      begin
        memOut_CT$wnnz_we <= memMergeIn_CT$wnnz_dbuf_we;
        memOut_CT$wnnz_valid <= memMergeIn_CT$wnnz_dbuf_d[0];
        if (memMergeIn_CT$wnnz_dbuf_we)
          begin
            memMergeIn_CT$wnnz_dbuf_mem[memMergeIn_CT$wnnz_dbuf_address] <= memMergeIn_CT$wnnz_dbuf_din;
            memOut_CT$wnnz_q <= memMergeIn_CT$wnnz_dbuf_din;
          end
        else
          memOut_CT$wnnz_q <= memMergeIn_CT$wnnz_dbuf_mem[memMergeIn_CT$wnnz_dbuf_address];
      end
  assign memOut_CT$wnnz_d = {memOut_CT$wnnz_q,
                             memOut_CT$wnnz_we,
                             memOut_CT$wnnz_valid};
  assign memMergeIn_CT$wnnz_dbuf_r = ((! memOut_CT$wnnz_valid) || memOut_CT$wnnz_r);
  logic [31:0] profiling_MemIn_CT$wnnz_read;
  logic [31:0] profiling_MemIn_CT$wnnz_write;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        profiling_MemIn_CT$wnnz_write <= 0;
        profiling_MemIn_CT$wnnz_read <= 0;
      end
    else
      if ((memMergeIn_CT$wnnz_dbuf_we == 1'd1))
        profiling_MemIn_CT$wnnz_write <= (profiling_MemIn_CT$wnnz_write + 1);
      else
        if ((memOut_CT$wnnz_valid == 1'd1))
          profiling_MemIn_CT$wnnz_read <= (profiling_MemIn_CT$wnnz_read + 1);
  
  /* demux (Ty C2,
       Ty MemOut_CT$wnnz) : (memMergeChoice_CT$wnnz,C2) (memOut_CT$wnnz_dbuf,MemOut_CT$wnnz) > [(memReadOut_CT$wnnz,MemOut_CT$wnnz),
                                                                                                (memWriteOut_CT$wnnz,MemOut_CT$wnnz)] */
  logic [1:0] memOut_CT$wnnz_dbuf_onehotd;
  always_comb
    if ((memMergeChoice_CT$wnnz_d[0] && memOut_CT$wnnz_dbuf_d[0]))
      unique case (memMergeChoice_CT$wnnz_d[1:1])
        1'd0: memOut_CT$wnnz_dbuf_onehotd = 2'd1;
        1'd1: memOut_CT$wnnz_dbuf_onehotd = 2'd2;
        default: memOut_CT$wnnz_dbuf_onehotd = 2'd0;
      endcase
    else memOut_CT$wnnz_dbuf_onehotd = 2'd0;
  assign memReadOut_CT$wnnz_d = {memOut_CT$wnnz_dbuf_d[116:1],
                                 memOut_CT$wnnz_dbuf_onehotd[0]};
  assign memWriteOut_CT$wnnz_d = {memOut_CT$wnnz_dbuf_d[116:1],
                                  memOut_CT$wnnz_dbuf_onehotd[1]};
  assign memOut_CT$wnnz_dbuf_r = (| (memOut_CT$wnnz_dbuf_onehotd & {memWriteOut_CT$wnnz_r,
                                                                    memReadOut_CT$wnnz_r}));
  assign memMergeChoice_CT$wnnz_r = memOut_CT$wnnz_dbuf_r;
  
  /* dbuf (Ty MemIn_CT$wnnz) : (memMergeIn_CT$wnnz_rbuf,MemIn_CT$wnnz) > (memMergeIn_CT$wnnz_dbuf,MemIn_CT$wnnz) */
  assign memMergeIn_CT$wnnz_rbuf_r = ((! memMergeIn_CT$wnnz_dbuf_d[0]) || memMergeIn_CT$wnnz_dbuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memMergeIn_CT$wnnz_dbuf_d <= {132'd0, 1'd0};
    else
      if (memMergeIn_CT$wnnz_rbuf_r)
        memMergeIn_CT$wnnz_dbuf_d <= memMergeIn_CT$wnnz_rbuf_d;
  
  /* rbuf (Ty MemIn_CT$wnnz) : (memMergeIn_CT$wnnz,MemIn_CT$wnnz) > (memMergeIn_CT$wnnz_rbuf,MemIn_CT$wnnz) */
  MemIn_CT$wnnz_t memMergeIn_CT$wnnz_buf;
  assign memMergeIn_CT$wnnz_r = (! memMergeIn_CT$wnnz_buf[0]);
  assign memMergeIn_CT$wnnz_rbuf_d = (memMergeIn_CT$wnnz_buf[0] ? memMergeIn_CT$wnnz_buf :
                                      memMergeIn_CT$wnnz_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memMergeIn_CT$wnnz_buf <= {132'd0, 1'd0};
    else
      if ((memMergeIn_CT$wnnz_rbuf_r && memMergeIn_CT$wnnz_buf[0]))
        memMergeIn_CT$wnnz_buf <= {132'd0, 1'd0};
      else if (((! memMergeIn_CT$wnnz_rbuf_r) && (! memMergeIn_CT$wnnz_buf[0])))
        memMergeIn_CT$wnnz_buf <= memMergeIn_CT$wnnz_d;
  
  /* dbuf (Ty MemOut_CT$wnnz) : (memOut_CT$wnnz_rbuf,MemOut_CT$wnnz) > (memOut_CT$wnnz_dbuf,MemOut_CT$wnnz) */
  assign memOut_CT$wnnz_rbuf_r = ((! memOut_CT$wnnz_dbuf_d[0]) || memOut_CT$wnnz_dbuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memOut_CT$wnnz_dbuf_d <= {116'd0, 1'd0};
    else
      if (memOut_CT$wnnz_rbuf_r)
        memOut_CT$wnnz_dbuf_d <= memOut_CT$wnnz_rbuf_d;
  
  /* rbuf (Ty MemOut_CT$wnnz) : (memOut_CT$wnnz,MemOut_CT$wnnz) > (memOut_CT$wnnz_rbuf,MemOut_CT$wnnz) */
  MemOut_CT$wnnz_t memOut_CT$wnnz_buf;
  assign memOut_CT$wnnz_r = (! memOut_CT$wnnz_buf[0]);
  assign memOut_CT$wnnz_rbuf_d = (memOut_CT$wnnz_buf[0] ? memOut_CT$wnnz_buf :
                                  memOut_CT$wnnz_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memOut_CT$wnnz_buf <= {116'd0, 1'd0};
    else
      if ((memOut_CT$wnnz_rbuf_r && memOut_CT$wnnz_buf[0]))
        memOut_CT$wnnz_buf <= {116'd0, 1'd0};
      else if (((! memOut_CT$wnnz_rbuf_r) && (! memOut_CT$wnnz_buf[0])))
        memOut_CT$wnnz_buf <= memOut_CT$wnnz_d;
  
  /* destruct (Ty Pointer_CT$wnnz,
          Dcon Pointer_CT$wnnz) : (scfarg_0_1_argbuf,Pointer_CT$wnnz) > [(destructReadIn_CT$wnnz,Word16#)] */
  assign destructReadIn_CT$wnnz_d = {scfarg_0_1_argbuf_d[16:1],
                                     scfarg_0_1_argbuf_d[0]};
  assign scfarg_0_1_argbuf_r = destructReadIn_CT$wnnz_r;
  
  /* dcon (Ty MemIn_CT$wnnz,
      Dcon ReadIn_CT$wnnz) : [(destructReadIn_CT$wnnz,Word16#)] > (dconReadIn_CT$wnnz,MemIn_CT$wnnz) */
  assign dconReadIn_CT$wnnz_d = ReadIn_CT$wnnz_dc((& {destructReadIn_CT$wnnz_d[0]}), destructReadIn_CT$wnnz_d);
  assign {destructReadIn_CT$wnnz_r} = {1 {(dconReadIn_CT$wnnz_r && dconReadIn_CT$wnnz_d[0])}};
  
  /* destruct (Ty MemOut_CT$wnnz,
          Dcon ReadOut_CT$wnnz) : (memReadOut_CT$wnnz,MemOut_CT$wnnz) > [(readPointer_CT$wnnzscfarg_0_1_argbuf,CT$wnnz)] */
  assign readPointer_CT$wnnzscfarg_0_1_argbuf_d = {memReadOut_CT$wnnz_d[116:2],
                                                   memReadOut_CT$wnnz_d[0]};
  assign memReadOut_CT$wnnz_r = readPointer_CT$wnnzscfarg_0_1_argbuf_r;
  
  /* mergectrl (Ty C5,Ty CT$wnnz) : [(lizzieLet0_1_argbuf,CT$wnnz),
                                (lizzieLet36_1_argbuf,CT$wnnz),
                                (lizzieLet37_1_argbuf,CT$wnnz),
                                (lizzieLet38_1_argbuf,CT$wnnz),
                                (lizzieLet5_1_argbuf,CT$wnnz)] > (writeMerge_choice_CT$wnnz,C5) (writeMerge_data_CT$wnnz,CT$wnnz) */
  logic [4:0] lizzieLet0_1_argbuf_select_d;
  assign lizzieLet0_1_argbuf_select_d = ((| lizzieLet0_1_argbuf_select_q) ? lizzieLet0_1_argbuf_select_q :
                                         (lizzieLet0_1_argbuf_d[0] ? 5'd1 :
                                          (lizzieLet36_1_argbuf_d[0] ? 5'd2 :
                                           (lizzieLet37_1_argbuf_d[0] ? 5'd4 :
                                            (lizzieLet38_1_argbuf_d[0] ? 5'd8 :
                                             (lizzieLet5_1_argbuf_d[0] ? 5'd16 :
                                              5'd0))))));
  logic [4:0] lizzieLet0_1_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet0_1_argbuf_select_q <= 5'd0;
    else
      lizzieLet0_1_argbuf_select_q <= (lizzieLet0_1_argbuf_done ? 5'd0 :
                                       lizzieLet0_1_argbuf_select_d);
  logic [1:0] lizzieLet0_1_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet0_1_argbuf_emit_q <= 2'd0;
    else
      lizzieLet0_1_argbuf_emit_q <= (lizzieLet0_1_argbuf_done ? 2'd0 :
                                     lizzieLet0_1_argbuf_emit_d);
  logic [1:0] lizzieLet0_1_argbuf_emit_d;
  assign lizzieLet0_1_argbuf_emit_d = (lizzieLet0_1_argbuf_emit_q | ({writeMerge_choice_CT$wnnz_d[0],
                                                                      writeMerge_data_CT$wnnz_d[0]} & {writeMerge_choice_CT$wnnz_r,
                                                                                                       writeMerge_data_CT$wnnz_r}));
  logic lizzieLet0_1_argbuf_done;
  assign lizzieLet0_1_argbuf_done = (& lizzieLet0_1_argbuf_emit_d);
  assign {lizzieLet5_1_argbuf_r,
          lizzieLet38_1_argbuf_r,
          lizzieLet37_1_argbuf_r,
          lizzieLet36_1_argbuf_r,
          lizzieLet0_1_argbuf_r} = (lizzieLet0_1_argbuf_done ? lizzieLet0_1_argbuf_select_d :
                                    5'd0);
  assign writeMerge_data_CT$wnnz_d = ((lizzieLet0_1_argbuf_select_d[0] && (! lizzieLet0_1_argbuf_emit_q[0])) ? lizzieLet0_1_argbuf_d :
                                      ((lizzieLet0_1_argbuf_select_d[1] && (! lizzieLet0_1_argbuf_emit_q[0])) ? lizzieLet36_1_argbuf_d :
                                       ((lizzieLet0_1_argbuf_select_d[2] && (! lizzieLet0_1_argbuf_emit_q[0])) ? lizzieLet37_1_argbuf_d :
                                        ((lizzieLet0_1_argbuf_select_d[3] && (! lizzieLet0_1_argbuf_emit_q[0])) ? lizzieLet38_1_argbuf_d :
                                         ((lizzieLet0_1_argbuf_select_d[4] && (! lizzieLet0_1_argbuf_emit_q[0])) ? lizzieLet5_1_argbuf_d :
                                          {115'd0, 1'd0})))));
  assign writeMerge_choice_CT$wnnz_d = ((lizzieLet0_1_argbuf_select_d[0] && (! lizzieLet0_1_argbuf_emit_q[1])) ? C1_5_dc(1'd1) :
                                        ((lizzieLet0_1_argbuf_select_d[1] && (! lizzieLet0_1_argbuf_emit_q[1])) ? C2_5_dc(1'd1) :
                                         ((lizzieLet0_1_argbuf_select_d[2] && (! lizzieLet0_1_argbuf_emit_q[1])) ? C3_5_dc(1'd1) :
                                          ((lizzieLet0_1_argbuf_select_d[3] && (! lizzieLet0_1_argbuf_emit_q[1])) ? C4_5_dc(1'd1) :
                                           ((lizzieLet0_1_argbuf_select_d[4] && (! lizzieLet0_1_argbuf_emit_q[1])) ? C5_5_dc(1'd1) :
                                            {3'd0, 1'd0})))));
  
  /* demux (Ty C5,
       Ty Pointer_CT$wnnz) : (writeMerge_choice_CT$wnnz,C5) (demuxWriteResult_CT$wnnz,Pointer_CT$wnnz) > [(writeCT$wnnzlizzieLet0_1_argbuf,Pointer_CT$wnnz),
                                                                                                          (writeCT$wnnzlizzieLet36_1_argbuf,Pointer_CT$wnnz),
                                                                                                          (writeCT$wnnzlizzieLet37_1_argbuf,Pointer_CT$wnnz),
                                                                                                          (writeCT$wnnzlizzieLet38_1_argbuf,Pointer_CT$wnnz),
                                                                                                          (writeCT$wnnzlizzieLet5_1_argbuf,Pointer_CT$wnnz)] */
  logic [4:0] demuxWriteResult_CT$wnnz_onehotd;
  always_comb
    if ((writeMerge_choice_CT$wnnz_d[0] && demuxWriteResult_CT$wnnz_d[0]))
      unique case (writeMerge_choice_CT$wnnz_d[3:1])
        3'd0: demuxWriteResult_CT$wnnz_onehotd = 5'd1;
        3'd1: demuxWriteResult_CT$wnnz_onehotd = 5'd2;
        3'd2: demuxWriteResult_CT$wnnz_onehotd = 5'd4;
        3'd3: demuxWriteResult_CT$wnnz_onehotd = 5'd8;
        3'd4: demuxWriteResult_CT$wnnz_onehotd = 5'd16;
        default: demuxWriteResult_CT$wnnz_onehotd = 5'd0;
      endcase
    else demuxWriteResult_CT$wnnz_onehotd = 5'd0;
  assign writeCT$wnnzlizzieLet0_1_argbuf_d = {demuxWriteResult_CT$wnnz_d[16:1],
                                              demuxWriteResult_CT$wnnz_onehotd[0]};
  assign writeCT$wnnzlizzieLet36_1_argbuf_d = {demuxWriteResult_CT$wnnz_d[16:1],
                                               demuxWriteResult_CT$wnnz_onehotd[1]};
  assign writeCT$wnnzlizzieLet37_1_argbuf_d = {demuxWriteResult_CT$wnnz_d[16:1],
                                               demuxWriteResult_CT$wnnz_onehotd[2]};
  assign writeCT$wnnzlizzieLet38_1_argbuf_d = {demuxWriteResult_CT$wnnz_d[16:1],
                                               demuxWriteResult_CT$wnnz_onehotd[3]};
  assign writeCT$wnnzlizzieLet5_1_argbuf_d = {demuxWriteResult_CT$wnnz_d[16:1],
                                              demuxWriteResult_CT$wnnz_onehotd[4]};
  assign demuxWriteResult_CT$wnnz_r = (| (demuxWriteResult_CT$wnnz_onehotd & {writeCT$wnnzlizzieLet5_1_argbuf_r,
                                                                              writeCT$wnnzlizzieLet38_1_argbuf_r,
                                                                              writeCT$wnnzlizzieLet37_1_argbuf_r,
                                                                              writeCT$wnnzlizzieLet36_1_argbuf_r,
                                                                              writeCT$wnnzlizzieLet0_1_argbuf_r}));
  assign writeMerge_choice_CT$wnnz_r = demuxWriteResult_CT$wnnz_r;
  
  /* dcon (Ty MemIn_CT$wnnz,
      Dcon WriteIn_CT$wnnz) : [(forkHP1_CT$wnn2,Word16#),
                               (writeMerge_data_CT$wnnz,CT$wnnz)] > (dconWriteIn_CT$wnnz,MemIn_CT$wnnz) */
  assign dconWriteIn_CT$wnnz_d = WriteIn_CT$wnnz_dc((& {forkHP1_CT$wnn2_d[0],
                                                        writeMerge_data_CT$wnnz_d[0]}), forkHP1_CT$wnn2_d, writeMerge_data_CT$wnnz_d);
  assign {forkHP1_CT$wnn2_r,
          writeMerge_data_CT$wnnz_r} = {2 {(dconWriteIn_CT$wnnz_r && dconWriteIn_CT$wnnz_d[0])}};
  
  /* dcon (Ty Pointer_CT$wnnz,
      Dcon Pointer_CT$wnnz) : [(forkHP1_CT$wnn3,Word16#)] > (dconPtr_CT$wnnz,Pointer_CT$wnnz) */
  assign dconPtr_CT$wnnz_d = Pointer_CT$wnnz_dc((& {forkHP1_CT$wnn3_d[0]}), forkHP1_CT$wnn3_d);
  assign {forkHP1_CT$wnn3_r} = {1 {(dconPtr_CT$wnnz_r && dconPtr_CT$wnnz_d[0])}};
  
  /* demux (Ty MemOut_CT$wnnz,
       Ty Pointer_CT$wnnz) : (memWriteOut_CT$wnnz,MemOut_CT$wnnz) (dconPtr_CT$wnnz,Pointer_CT$wnnz) > [(_84,Pointer_CT$wnnz),
                                                                                                       (demuxWriteResult_CT$wnnz,Pointer_CT$wnnz)] */
  logic [1:0] dconPtr_CT$wnnz_onehotd;
  always_comb
    if ((memWriteOut_CT$wnnz_d[0] && dconPtr_CT$wnnz_d[0]))
      unique case (memWriteOut_CT$wnnz_d[1:1])
        1'd0: dconPtr_CT$wnnz_onehotd = 2'd1;
        1'd1: dconPtr_CT$wnnz_onehotd = 2'd2;
        default: dconPtr_CT$wnnz_onehotd = 2'd0;
      endcase
    else dconPtr_CT$wnnz_onehotd = 2'd0;
  assign _84_d = {dconPtr_CT$wnnz_d[16:1],
                  dconPtr_CT$wnnz_onehotd[0]};
  assign demuxWriteResult_CT$wnnz_d = {dconPtr_CT$wnnz_d[16:1],
                                       dconPtr_CT$wnnz_onehotd[1]};
  assign dconPtr_CT$wnnz_r = (| (dconPtr_CT$wnnz_onehotd & {demuxWriteResult_CT$wnnz_r,
                                                            _84_r}));
  assign memWriteOut_CT$wnnz_r = dconPtr_CT$wnnz_r;
  
  /* const (Ty Word16#,
       Lit 0) : (go__9,Go) > (initHP_CTf''''''''_f''''''''_Int_Int,Word16#) */
  assign \initHP_CTf''''''''_f''''''''_Int_Int_d  = {16'd0,
                                                     go__9_d[0]};
  assign go__9_r = \initHP_CTf''''''''_f''''''''_Int_Int_r ;
  
  /* const (Ty Word16#,
       Lit 1) : (incrHP_CTf''''''''_f''''''''_Int_Int1,Go) > (incrHP_CTf''''''''_f''''''''_Int_Int,Word16#) */
  assign \incrHP_CTf''''''''_f''''''''_Int_Int_d  = {16'd1,
                                                     \incrHP_CTf''''''''_f''''''''_Int_Int1_d [0]};
  assign \incrHP_CTf''''''''_f''''''''_Int_Int1_r  = \incrHP_CTf''''''''_f''''''''_Int_Int_r ;
  
  /* merge (Ty Go) : [(go__10,Go),
                 (incrHP_CTf''''''''_f''''''''_Int_Int2,Go)] > (incrHP_mergeCTf''''''''_f''''''''_Int_Int,Go) */
  logic [1:0] \incrHP_mergeCTf''''''''_f''''''''_Int_Int_selected ;
  logic [1:0] \incrHP_mergeCTf''''''''_f''''''''_Int_Int_select ;
  always_comb
    begin
      \incrHP_mergeCTf''''''''_f''''''''_Int_Int_selected  = 2'd0;
      if ((| \incrHP_mergeCTf''''''''_f''''''''_Int_Int_select ))
        \incrHP_mergeCTf''''''''_f''''''''_Int_Int_selected  = \incrHP_mergeCTf''''''''_f''''''''_Int_Int_select ;
      else
        if (go__10_d[0])
          \incrHP_mergeCTf''''''''_f''''''''_Int_Int_selected [0] = 1'd1;
        else if (\incrHP_CTf''''''''_f''''''''_Int_Int2_d [0])
          \incrHP_mergeCTf''''''''_f''''''''_Int_Int_selected [1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \incrHP_mergeCTf''''''''_f''''''''_Int_Int_select  <= 2'd0;
    else
      \incrHP_mergeCTf''''''''_f''''''''_Int_Int_select  <= (\incrHP_mergeCTf''''''''_f''''''''_Int_Int_r  ? 2'd0 :
                                                             \incrHP_mergeCTf''''''''_f''''''''_Int_Int_selected );
  always_comb
    if (\incrHP_mergeCTf''''''''_f''''''''_Int_Int_selected [0])
      \incrHP_mergeCTf''''''''_f''''''''_Int_Int_d  = go__10_d;
    else if (\incrHP_mergeCTf''''''''_f''''''''_Int_Int_selected [1])
      \incrHP_mergeCTf''''''''_f''''''''_Int_Int_d  = \incrHP_CTf''''''''_f''''''''_Int_Int2_d ;
    else \incrHP_mergeCTf''''''''_f''''''''_Int_Int_d  = 1'd0;
  assign {\incrHP_CTf''''''''_f''''''''_Int_Int2_r ,
          go__10_r} = (\incrHP_mergeCTf''''''''_f''''''''_Int_Int_r  ? \incrHP_mergeCTf''''''''_f''''''''_Int_Int_selected  :
                       2'd0);
  
  /* fork (Ty Go) : (incrHP_mergeCTf''''''''_f''''''''_Int_Int_buf,Go) > [(incrHP_CTf''''''''_f''''''''_Int_Int1,Go),
                                                                     (incrHP_CTf''''''''_f''''''''_Int_Int2,Go)] */
  logic [1:0] \incrHP_mergeCTf''''''''_f''''''''_Int_Int_buf_emitted ;
  logic [1:0] \incrHP_mergeCTf''''''''_f''''''''_Int_Int_buf_done ;
  assign \incrHP_CTf''''''''_f''''''''_Int_Int1_d  = (\incrHP_mergeCTf''''''''_f''''''''_Int_Int_buf_d [0] && (! \incrHP_mergeCTf''''''''_f''''''''_Int_Int_buf_emitted [0]));
  assign \incrHP_CTf''''''''_f''''''''_Int_Int2_d  = (\incrHP_mergeCTf''''''''_f''''''''_Int_Int_buf_d [0] && (! \incrHP_mergeCTf''''''''_f''''''''_Int_Int_buf_emitted [1]));
  assign \incrHP_mergeCTf''''''''_f''''''''_Int_Int_buf_done  = (\incrHP_mergeCTf''''''''_f''''''''_Int_Int_buf_emitted  | ({\incrHP_CTf''''''''_f''''''''_Int_Int2_d [0],
                                                                                                                             \incrHP_CTf''''''''_f''''''''_Int_Int1_d [0]} & {\incrHP_CTf''''''''_f''''''''_Int_Int2_r ,
                                                                                                                                                                              \incrHP_CTf''''''''_f''''''''_Int_Int1_r }));
  assign \incrHP_mergeCTf''''''''_f''''''''_Int_Int_buf_r  = (& \incrHP_mergeCTf''''''''_f''''''''_Int_Int_buf_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \incrHP_mergeCTf''''''''_f''''''''_Int_Int_buf_emitted  <= 2'd0;
    else
      \incrHP_mergeCTf''''''''_f''''''''_Int_Int_buf_emitted  <= (\incrHP_mergeCTf''''''''_f''''''''_Int_Int_buf_r  ? 2'd0 :
                                                                  \incrHP_mergeCTf''''''''_f''''''''_Int_Int_buf_done );
  
  /* op_add (Ty Word16#) : (incrHP_CTf''''''''_f''''''''_Int_Int,Word16#) (forkHP1_CTf''''''''_f''''''''_Int_Int,Word16#) > (addHP_CTf''''''''_f''''''''_Int_Int,Word16#) */
  assign \addHP_CTf''''''''_f''''''''_Int_Int_d  = {(\incrHP_CTf''''''''_f''''''''_Int_Int_d [16:1] + \forkHP1_CTf''''''''_f''''''''_Int_Int_d [16:1]),
                                                    (\incrHP_CTf''''''''_f''''''''_Int_Int_d [0] && \forkHP1_CTf''''''''_f''''''''_Int_Int_d [0])};
  assign {\incrHP_CTf''''''''_f''''''''_Int_Int_r ,
          \forkHP1_CTf''''''''_f''''''''_Int_Int_r } = {2 {(\addHP_CTf''''''''_f''''''''_Int_Int_r  && \addHP_CTf''''''''_f''''''''_Int_Int_d [0])}};
  
  /* merge (Ty Word16#) : [(initHP_CTf''''''''_f''''''''_Int_Int,Word16#),
                      (addHP_CTf''''''''_f''''''''_Int_Int,Word16#)] > (mergeHP_CTf''''''''_f''''''''_Int_Int,Word16#) */
  logic [1:0] \mergeHP_CTf''''''''_f''''''''_Int_Int_selected ;
  logic [1:0] \mergeHP_CTf''''''''_f''''''''_Int_Int_select ;
  always_comb
    begin
      \mergeHP_CTf''''''''_f''''''''_Int_Int_selected  = 2'd0;
      if ((| \mergeHP_CTf''''''''_f''''''''_Int_Int_select ))
        \mergeHP_CTf''''''''_f''''''''_Int_Int_selected  = \mergeHP_CTf''''''''_f''''''''_Int_Int_select ;
      else
        if (\initHP_CTf''''''''_f''''''''_Int_Int_d [0])
          \mergeHP_CTf''''''''_f''''''''_Int_Int_selected [0] = 1'd1;
        else if (\addHP_CTf''''''''_f''''''''_Int_Int_d [0])
          \mergeHP_CTf''''''''_f''''''''_Int_Int_selected [1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \mergeHP_CTf''''''''_f''''''''_Int_Int_select  <= 2'd0;
    else
      \mergeHP_CTf''''''''_f''''''''_Int_Int_select  <= (\mergeHP_CTf''''''''_f''''''''_Int_Int_r  ? 2'd0 :
                                                         \mergeHP_CTf''''''''_f''''''''_Int_Int_selected );
  always_comb
    if (\mergeHP_CTf''''''''_f''''''''_Int_Int_selected [0])
      \mergeHP_CTf''''''''_f''''''''_Int_Int_d  = \initHP_CTf''''''''_f''''''''_Int_Int_d ;
    else if (\mergeHP_CTf''''''''_f''''''''_Int_Int_selected [1])
      \mergeHP_CTf''''''''_f''''''''_Int_Int_d  = \addHP_CTf''''''''_f''''''''_Int_Int_d ;
    else \mergeHP_CTf''''''''_f''''''''_Int_Int_d  = {16'd0, 1'd0};
  assign {\addHP_CTf''''''''_f''''''''_Int_Int_r ,
          \initHP_CTf''''''''_f''''''''_Int_Int_r } = (\mergeHP_CTf''''''''_f''''''''_Int_Int_r  ? \mergeHP_CTf''''''''_f''''''''_Int_Int_selected  :
                                                       2'd0);
  
  /* buf (Ty Go) : (incrHP_mergeCTf''''''''_f''''''''_Int_Int,Go) > (incrHP_mergeCTf''''''''_f''''''''_Int_Int_buf,Go) */
  Go_t \incrHP_mergeCTf''''''''_f''''''''_Int_Int_bufchan_d ;
  logic \incrHP_mergeCTf''''''''_f''''''''_Int_Int_bufchan_r ;
  assign \incrHP_mergeCTf''''''''_f''''''''_Int_Int_r  = ((! \incrHP_mergeCTf''''''''_f''''''''_Int_Int_bufchan_d [0]) || \incrHP_mergeCTf''''''''_f''''''''_Int_Int_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \incrHP_mergeCTf''''''''_f''''''''_Int_Int_bufchan_d  <= 1'd0;
    else
      if (\incrHP_mergeCTf''''''''_f''''''''_Int_Int_r )
        \incrHP_mergeCTf''''''''_f''''''''_Int_Int_bufchan_d  <= \incrHP_mergeCTf''''''''_f''''''''_Int_Int_d ;
  Go_t \incrHP_mergeCTf''''''''_f''''''''_Int_Int_bufchan_buf ;
  assign \incrHP_mergeCTf''''''''_f''''''''_Int_Int_bufchan_r  = (! \incrHP_mergeCTf''''''''_f''''''''_Int_Int_bufchan_buf [0]);
  assign \incrHP_mergeCTf''''''''_f''''''''_Int_Int_buf_d  = (\incrHP_mergeCTf''''''''_f''''''''_Int_Int_bufchan_buf [0] ? \incrHP_mergeCTf''''''''_f''''''''_Int_Int_bufchan_buf  :
                                                              \incrHP_mergeCTf''''''''_f''''''''_Int_Int_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \incrHP_mergeCTf''''''''_f''''''''_Int_Int_bufchan_buf  <= 1'd0;
    else
      if ((\incrHP_mergeCTf''''''''_f''''''''_Int_Int_buf_r  && \incrHP_mergeCTf''''''''_f''''''''_Int_Int_bufchan_buf [0]))
        \incrHP_mergeCTf''''''''_f''''''''_Int_Int_bufchan_buf  <= 1'd0;
      else if (((! \incrHP_mergeCTf''''''''_f''''''''_Int_Int_buf_r ) && (! \incrHP_mergeCTf''''''''_f''''''''_Int_Int_bufchan_buf [0])))
        \incrHP_mergeCTf''''''''_f''''''''_Int_Int_bufchan_buf  <= \incrHP_mergeCTf''''''''_f''''''''_Int_Int_bufchan_d ;
  
  /* buf (Ty Word16#) : (mergeHP_CTf''''''''_f''''''''_Int_Int,Word16#) > (mergeHP_CTf''''''''_f''''''''_Int_Int_buf,Word16#) */
  \Word16#_t  \mergeHP_CTf''''''''_f''''''''_Int_Int_bufchan_d ;
  logic \mergeHP_CTf''''''''_f''''''''_Int_Int_bufchan_r ;
  assign \mergeHP_CTf''''''''_f''''''''_Int_Int_r  = ((! \mergeHP_CTf''''''''_f''''''''_Int_Int_bufchan_d [0]) || \mergeHP_CTf''''''''_f''''''''_Int_Int_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \mergeHP_CTf''''''''_f''''''''_Int_Int_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\mergeHP_CTf''''''''_f''''''''_Int_Int_r )
        \mergeHP_CTf''''''''_f''''''''_Int_Int_bufchan_d  <= \mergeHP_CTf''''''''_f''''''''_Int_Int_d ;
  \Word16#_t  \mergeHP_CTf''''''''_f''''''''_Int_Int_bufchan_buf ;
  assign \mergeHP_CTf''''''''_f''''''''_Int_Int_bufchan_r  = (! \mergeHP_CTf''''''''_f''''''''_Int_Int_bufchan_buf [0]);
  assign \mergeHP_CTf''''''''_f''''''''_Int_Int_buf_d  = (\mergeHP_CTf''''''''_f''''''''_Int_Int_bufchan_buf [0] ? \mergeHP_CTf''''''''_f''''''''_Int_Int_bufchan_buf  :
                                                          \mergeHP_CTf''''''''_f''''''''_Int_Int_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \mergeHP_CTf''''''''_f''''''''_Int_Int_bufchan_buf  <= {16'd0,
                                                              1'd0};
    else
      if ((\mergeHP_CTf''''''''_f''''''''_Int_Int_buf_r  && \mergeHP_CTf''''''''_f''''''''_Int_Int_bufchan_buf [0]))
        \mergeHP_CTf''''''''_f''''''''_Int_Int_bufchan_buf  <= {16'd0,
                                                                1'd0};
      else if (((! \mergeHP_CTf''''''''_f''''''''_Int_Int_buf_r ) && (! \mergeHP_CTf''''''''_f''''''''_Int_Int_bufchan_buf [0])))
        \mergeHP_CTf''''''''_f''''''''_Int_Int_bufchan_buf  <= \mergeHP_CTf''''''''_f''''''''_Int_Int_bufchan_d ;
  
  /* fork (Ty Word16#) : (mergeHP_CTf''''''''_f''''''''_Int_Int_buf,Word16#) > [(forkHP1_CTf''''''''_f''''''''_Int_Int,Word16#),
                                                                           (forkHP1_CTf''''''''_f''''''''_Int_In2,Word16#),
                                                                           (forkHP1_CTf''''''''_f''''''''_Int_In3,Word16#)] */
  logic [2:0] \mergeHP_CTf''''''''_f''''''''_Int_Int_buf_emitted ;
  logic [2:0] \mergeHP_CTf''''''''_f''''''''_Int_Int_buf_done ;
  assign \forkHP1_CTf''''''''_f''''''''_Int_Int_d  = {\mergeHP_CTf''''''''_f''''''''_Int_Int_buf_d [16:1],
                                                      (\mergeHP_CTf''''''''_f''''''''_Int_Int_buf_d [0] && (! \mergeHP_CTf''''''''_f''''''''_Int_Int_buf_emitted [0]))};
  assign \forkHP1_CTf''''''''_f''''''''_Int_In2_d  = {\mergeHP_CTf''''''''_f''''''''_Int_Int_buf_d [16:1],
                                                      (\mergeHP_CTf''''''''_f''''''''_Int_Int_buf_d [0] && (! \mergeHP_CTf''''''''_f''''''''_Int_Int_buf_emitted [1]))};
  assign \forkHP1_CTf''''''''_f''''''''_Int_In3_d  = {\mergeHP_CTf''''''''_f''''''''_Int_Int_buf_d [16:1],
                                                      (\mergeHP_CTf''''''''_f''''''''_Int_Int_buf_d [0] && (! \mergeHP_CTf''''''''_f''''''''_Int_Int_buf_emitted [2]))};
  assign \mergeHP_CTf''''''''_f''''''''_Int_Int_buf_done  = (\mergeHP_CTf''''''''_f''''''''_Int_Int_buf_emitted  | ({\forkHP1_CTf''''''''_f''''''''_Int_In3_d [0],
                                                                                                                     \forkHP1_CTf''''''''_f''''''''_Int_In2_d [0],
                                                                                                                     \forkHP1_CTf''''''''_f''''''''_Int_Int_d [0]} & {\forkHP1_CTf''''''''_f''''''''_Int_In3_r ,
                                                                                                                                                                      \forkHP1_CTf''''''''_f''''''''_Int_In2_r ,
                                                                                                                                                                      \forkHP1_CTf''''''''_f''''''''_Int_Int_r }));
  assign \mergeHP_CTf''''''''_f''''''''_Int_Int_buf_r  = (& \mergeHP_CTf''''''''_f''''''''_Int_Int_buf_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \mergeHP_CTf''''''''_f''''''''_Int_Int_buf_emitted  <= 3'd0;
    else
      \mergeHP_CTf''''''''_f''''''''_Int_Int_buf_emitted  <= (\mergeHP_CTf''''''''_f''''''''_Int_Int_buf_r  ? 3'd0 :
                                                              \mergeHP_CTf''''''''_f''''''''_Int_Int_buf_done );
  
  /* mergectrl (Ty C2,
           Ty MemIn_CTf''''''''_f''''''''_Int_Int) : [(dconReadIn_CTf''''''''_f''''''''_Int_Int,MemIn_CTf''''''''_f''''''''_Int_Int),
                                                      (dconWriteIn_CTf''''''''_f''''''''_Int_Int,MemIn_CTf''''''''_f''''''''_Int_Int)] > (memMergeChoice_CTf''''''''_f''''''''_Int_Int,C2) (memMergeIn_CTf''''''''_f''''''''_Int_Int,MemIn_CTf''''''''_f''''''''_Int_Int) */
  logic [1:0] \dconReadIn_CTf''''''''_f''''''''_Int_Int_select_d ;
  assign \dconReadIn_CTf''''''''_f''''''''_Int_Int_select_d  = ((| \dconReadIn_CTf''''''''_f''''''''_Int_Int_select_q ) ? \dconReadIn_CTf''''''''_f''''''''_Int_Int_select_q  :
                                                                (\dconReadIn_CTf''''''''_f''''''''_Int_Int_d [0] ? 2'd1 :
                                                                 (\dconWriteIn_CTf''''''''_f''''''''_Int_Int_d [0] ? 2'd2 :
                                                                  2'd0)));
  logic [1:0] \dconReadIn_CTf''''''''_f''''''''_Int_Int_select_q ;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \dconReadIn_CTf''''''''_f''''''''_Int_Int_select_q  <= 2'd0;
    else
      \dconReadIn_CTf''''''''_f''''''''_Int_Int_select_q  <= (\dconReadIn_CTf''''''''_f''''''''_Int_Int_done  ? 2'd0 :
                                                              \dconReadIn_CTf''''''''_f''''''''_Int_Int_select_d );
  logic [1:0] \dconReadIn_CTf''''''''_f''''''''_Int_Int_emit_q ;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \dconReadIn_CTf''''''''_f''''''''_Int_Int_emit_q  <= 2'd0;
    else
      \dconReadIn_CTf''''''''_f''''''''_Int_Int_emit_q  <= (\dconReadIn_CTf''''''''_f''''''''_Int_Int_done  ? 2'd0 :
                                                            \dconReadIn_CTf''''''''_f''''''''_Int_Int_emit_d );
  logic [1:0] \dconReadIn_CTf''''''''_f''''''''_Int_Int_emit_d ;
  assign \dconReadIn_CTf''''''''_f''''''''_Int_Int_emit_d  = (\dconReadIn_CTf''''''''_f''''''''_Int_Int_emit_q  | ({\memMergeChoice_CTf''''''''_f''''''''_Int_Int_d [0],
                                                                                                                    \memMergeIn_CTf''''''''_f''''''''_Int_Int_d [0]} & {\memMergeChoice_CTf''''''''_f''''''''_Int_Int_r ,
                                                                                                                                                                        \memMergeIn_CTf''''''''_f''''''''_Int_Int_r }));
  logic \dconReadIn_CTf''''''''_f''''''''_Int_Int_done ;
  assign \dconReadIn_CTf''''''''_f''''''''_Int_Int_done  = (& \dconReadIn_CTf''''''''_f''''''''_Int_Int_emit_d );
  assign {\dconWriteIn_CTf''''''''_f''''''''_Int_Int_r ,
          \dconReadIn_CTf''''''''_f''''''''_Int_Int_r } = (\dconReadIn_CTf''''''''_f''''''''_Int_Int_done  ? \dconReadIn_CTf''''''''_f''''''''_Int_Int_select_d  :
                                                           2'd0);
  assign \memMergeIn_CTf''''''''_f''''''''_Int_Int_d  = ((\dconReadIn_CTf''''''''_f''''''''_Int_Int_select_d [0] && (! \dconReadIn_CTf''''''''_f''''''''_Int_Int_emit_q [0])) ? \dconReadIn_CTf''''''''_f''''''''_Int_Int_d  :
                                                         ((\dconReadIn_CTf''''''''_f''''''''_Int_Int_select_d [1] && (! \dconReadIn_CTf''''''''_f''''''''_Int_Int_emit_q [0])) ? \dconWriteIn_CTf''''''''_f''''''''_Int_Int_d  :
                                                          {84'd0, 1'd0}));
  assign \memMergeChoice_CTf''''''''_f''''''''_Int_Int_d  = ((\dconReadIn_CTf''''''''_f''''''''_Int_Int_select_d [0] && (! \dconReadIn_CTf''''''''_f''''''''_Int_Int_emit_q [1])) ? C1_2_dc(1'd1) :
                                                             ((\dconReadIn_CTf''''''''_f''''''''_Int_Int_select_d [1] && (! \dconReadIn_CTf''''''''_f''''''''_Int_Int_emit_q [1])) ? C2_2_dc(1'd1) :
                                                              {1'd0, 1'd0}));
  
  /* bram (Ty MemIn_CTf''''''''_f''''''''_Int_Int,
      Ty MemOut_CTf''''''''_f''''''''_Int_Int) : (memMergeIn_CTf''''''''_f''''''''_Int_Int_dbuf,MemIn_CTf''''''''_f''''''''_Int_Int) > (memOut_CTf''''''''_f''''''''_Int_Int,MemOut_CTf''''''''_f''''''''_Int_Int) */
  logic [66:0] \memMergeIn_CTf''''''''_f''''''''_Int_Int_dbuf_mem [65535:0];
  logic [15:0] \memMergeIn_CTf''''''''_f''''''''_Int_Int_dbuf_address ;
  logic [66:0] \memMergeIn_CTf''''''''_f''''''''_Int_Int_dbuf_din ;
  logic [66:0] \memOut_CTf''''''''_f''''''''_Int_Int_q ;
  logic \memOut_CTf''''''''_f''''''''_Int_Int_valid ;
  logic \memMergeIn_CTf''''''''_f''''''''_Int_Int_dbuf_we ;
  logic \memOut_CTf''''''''_f''''''''_Int_Int_we ;
  assign \memMergeIn_CTf''''''''_f''''''''_Int_Int_dbuf_din  = \memMergeIn_CTf''''''''_f''''''''_Int_Int_dbuf_d [84:18];
  assign \memMergeIn_CTf''''''''_f''''''''_Int_Int_dbuf_address  = \memMergeIn_CTf''''''''_f''''''''_Int_Int_dbuf_d [17:2];
  assign \memMergeIn_CTf''''''''_f''''''''_Int_Int_dbuf_we  = (\memMergeIn_CTf''''''''_f''''''''_Int_Int_dbuf_d [1:1] && \memMergeIn_CTf''''''''_f''''''''_Int_Int_dbuf_d [0]);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        \memOut_CTf''''''''_f''''''''_Int_Int_we  <= 1'd0;
        \memOut_CTf''''''''_f''''''''_Int_Int_valid  <= 1'd0;
      end
    else
      begin
        \memOut_CTf''''''''_f''''''''_Int_Int_we  <= \memMergeIn_CTf''''''''_f''''''''_Int_Int_dbuf_we ;
        \memOut_CTf''''''''_f''''''''_Int_Int_valid  <= \memMergeIn_CTf''''''''_f''''''''_Int_Int_dbuf_d [0];
        if (\memMergeIn_CTf''''''''_f''''''''_Int_Int_dbuf_we )
          begin
            \memMergeIn_CTf''''''''_f''''''''_Int_Int_dbuf_mem [\memMergeIn_CTf''''''''_f''''''''_Int_Int_dbuf_address ] <= \memMergeIn_CTf''''''''_f''''''''_Int_Int_dbuf_din ;
            \memOut_CTf''''''''_f''''''''_Int_Int_q  <= \memMergeIn_CTf''''''''_f''''''''_Int_Int_dbuf_din ;
          end
        else
          \memOut_CTf''''''''_f''''''''_Int_Int_q  <= \memMergeIn_CTf''''''''_f''''''''_Int_Int_dbuf_mem [\memMergeIn_CTf''''''''_f''''''''_Int_Int_dbuf_address ];
      end
  assign \memOut_CTf''''''''_f''''''''_Int_Int_d  = {\memOut_CTf''''''''_f''''''''_Int_Int_q ,
                                                     \memOut_CTf''''''''_f''''''''_Int_Int_we ,
                                                     \memOut_CTf''''''''_f''''''''_Int_Int_valid };
  assign \memMergeIn_CTf''''''''_f''''''''_Int_Int_dbuf_r  = ((! \memOut_CTf''''''''_f''''''''_Int_Int_valid ) || \memOut_CTf''''''''_f''''''''_Int_Int_r );
  logic [31:0] \profiling_MemIn_CTf''''''''_f''''''''_Int_Int_read ;
  logic [31:0] \profiling_MemIn_CTf''''''''_f''''''''_Int_Int_write ;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        \profiling_MemIn_CTf''''''''_f''''''''_Int_Int_write  <= 0;
        \profiling_MemIn_CTf''''''''_f''''''''_Int_Int_read  <= 0;
      end
    else
      if ((\memMergeIn_CTf''''''''_f''''''''_Int_Int_dbuf_we  == 1'd1))
        \profiling_MemIn_CTf''''''''_f''''''''_Int_Int_write  <= (\profiling_MemIn_CTf''''''''_f''''''''_Int_Int_write  + 1);
      else
        if ((\memOut_CTf''''''''_f''''''''_Int_Int_valid  == 1'd1))
          \profiling_MemIn_CTf''''''''_f''''''''_Int_Int_read  <= (\profiling_MemIn_CTf''''''''_f''''''''_Int_Int_read  + 1);
  
  /* demux (Ty C2,
       Ty MemOut_CTf''''''''_f''''''''_Int_Int) : (memMergeChoice_CTf''''''''_f''''''''_Int_Int,C2) (memOut_CTf''''''''_f''''''''_Int_Int_dbuf,MemOut_CTf''''''''_f''''''''_Int_Int) > [(memReadOut_CTf''''''''_f''''''''_Int_Int,MemOut_CTf''''''''_f''''''''_Int_Int),
                                                                                                                                                                                        (memWriteOut_CTf''''''''_f''''''''_Int_Int,MemOut_CTf''''''''_f''''''''_Int_Int)] */
  logic [1:0] \memOut_CTf''''''''_f''''''''_Int_Int_dbuf_onehotd ;
  always_comb
    if ((\memMergeChoice_CTf''''''''_f''''''''_Int_Int_d [0] && \memOut_CTf''''''''_f''''''''_Int_Int_dbuf_d [0]))
      unique case (\memMergeChoice_CTf''''''''_f''''''''_Int_Int_d [1:1])
        1'd0: \memOut_CTf''''''''_f''''''''_Int_Int_dbuf_onehotd  = 2'd1;
        1'd1: \memOut_CTf''''''''_f''''''''_Int_Int_dbuf_onehotd  = 2'd2;
        default:
          \memOut_CTf''''''''_f''''''''_Int_Int_dbuf_onehotd  = 2'd0;
      endcase
    else \memOut_CTf''''''''_f''''''''_Int_Int_dbuf_onehotd  = 2'd0;
  assign \memReadOut_CTf''''''''_f''''''''_Int_Int_d  = {\memOut_CTf''''''''_f''''''''_Int_Int_dbuf_d [68:1],
                                                         \memOut_CTf''''''''_f''''''''_Int_Int_dbuf_onehotd [0]};
  assign \memWriteOut_CTf''''''''_f''''''''_Int_Int_d  = {\memOut_CTf''''''''_f''''''''_Int_Int_dbuf_d [68:1],
                                                          \memOut_CTf''''''''_f''''''''_Int_Int_dbuf_onehotd [1]};
  assign \memOut_CTf''''''''_f''''''''_Int_Int_dbuf_r  = (| (\memOut_CTf''''''''_f''''''''_Int_Int_dbuf_onehotd  & {\memWriteOut_CTf''''''''_f''''''''_Int_Int_r ,
                                                                                                                    \memReadOut_CTf''''''''_f''''''''_Int_Int_r }));
  assign \memMergeChoice_CTf''''''''_f''''''''_Int_Int_r  = \memOut_CTf''''''''_f''''''''_Int_Int_dbuf_r ;
  
  /* dbuf (Ty MemIn_CTf''''''''_f''''''''_Int_Int) : (memMergeIn_CTf''''''''_f''''''''_Int_Int_rbuf,MemIn_CTf''''''''_f''''''''_Int_Int) > (memMergeIn_CTf''''''''_f''''''''_Int_Int_dbuf,MemIn_CTf''''''''_f''''''''_Int_Int) */
  assign \memMergeIn_CTf''''''''_f''''''''_Int_Int_rbuf_r  = ((! \memMergeIn_CTf''''''''_f''''''''_Int_Int_dbuf_d [0]) || \memMergeIn_CTf''''''''_f''''''''_Int_Int_dbuf_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \memMergeIn_CTf''''''''_f''''''''_Int_Int_dbuf_d  <= {84'd0, 1'd0};
    else
      if (\memMergeIn_CTf''''''''_f''''''''_Int_Int_rbuf_r )
        \memMergeIn_CTf''''''''_f''''''''_Int_Int_dbuf_d  <= \memMergeIn_CTf''''''''_f''''''''_Int_Int_rbuf_d ;
  
  /* rbuf (Ty MemIn_CTf''''''''_f''''''''_Int_Int) : (memMergeIn_CTf''''''''_f''''''''_Int_Int,MemIn_CTf''''''''_f''''''''_Int_Int) > (memMergeIn_CTf''''''''_f''''''''_Int_Int_rbuf,MemIn_CTf''''''''_f''''''''_Int_Int) */
  \MemIn_CTf''''''''_f''''''''_Int_Int_t  \memMergeIn_CTf''''''''_f''''''''_Int_Int_buf ;
  assign \memMergeIn_CTf''''''''_f''''''''_Int_Int_r  = (! \memMergeIn_CTf''''''''_f''''''''_Int_Int_buf [0]);
  assign \memMergeIn_CTf''''''''_f''''''''_Int_Int_rbuf_d  = (\memMergeIn_CTf''''''''_f''''''''_Int_Int_buf [0] ? \memMergeIn_CTf''''''''_f''''''''_Int_Int_buf  :
                                                              \memMergeIn_CTf''''''''_f''''''''_Int_Int_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \memMergeIn_CTf''''''''_f''''''''_Int_Int_buf  <= {84'd0, 1'd0};
    else
      if ((\memMergeIn_CTf''''''''_f''''''''_Int_Int_rbuf_r  && \memMergeIn_CTf''''''''_f''''''''_Int_Int_buf [0]))
        \memMergeIn_CTf''''''''_f''''''''_Int_Int_buf  <= {84'd0, 1'd0};
      else if (((! \memMergeIn_CTf''''''''_f''''''''_Int_Int_rbuf_r ) && (! \memMergeIn_CTf''''''''_f''''''''_Int_Int_buf [0])))
        \memMergeIn_CTf''''''''_f''''''''_Int_Int_buf  <= \memMergeIn_CTf''''''''_f''''''''_Int_Int_d ;
  
  /* dbuf (Ty MemOut_CTf''''''''_f''''''''_Int_Int) : (memOut_CTf''''''''_f''''''''_Int_Int_rbuf,MemOut_CTf''''''''_f''''''''_Int_Int) > (memOut_CTf''''''''_f''''''''_Int_Int_dbuf,MemOut_CTf''''''''_f''''''''_Int_Int) */
  assign \memOut_CTf''''''''_f''''''''_Int_Int_rbuf_r  = ((! \memOut_CTf''''''''_f''''''''_Int_Int_dbuf_d [0]) || \memOut_CTf''''''''_f''''''''_Int_Int_dbuf_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \memOut_CTf''''''''_f''''''''_Int_Int_dbuf_d  <= {68'd0, 1'd0};
    else
      if (\memOut_CTf''''''''_f''''''''_Int_Int_rbuf_r )
        \memOut_CTf''''''''_f''''''''_Int_Int_dbuf_d  <= \memOut_CTf''''''''_f''''''''_Int_Int_rbuf_d ;
  
  /* rbuf (Ty MemOut_CTf''''''''_f''''''''_Int_Int) : (memOut_CTf''''''''_f''''''''_Int_Int,MemOut_CTf''''''''_f''''''''_Int_Int) > (memOut_CTf''''''''_f''''''''_Int_Int_rbuf,MemOut_CTf''''''''_f''''''''_Int_Int) */
  \MemOut_CTf''''''''_f''''''''_Int_Int_t  \memOut_CTf''''''''_f''''''''_Int_Int_buf ;
  assign \memOut_CTf''''''''_f''''''''_Int_Int_r  = (! \memOut_CTf''''''''_f''''''''_Int_Int_buf [0]);
  assign \memOut_CTf''''''''_f''''''''_Int_Int_rbuf_d  = (\memOut_CTf''''''''_f''''''''_Int_Int_buf [0] ? \memOut_CTf''''''''_f''''''''_Int_Int_buf  :
                                                          \memOut_CTf''''''''_f''''''''_Int_Int_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \memOut_CTf''''''''_f''''''''_Int_Int_buf  <= {68'd0, 1'd0};
    else
      if ((\memOut_CTf''''''''_f''''''''_Int_Int_rbuf_r  && \memOut_CTf''''''''_f''''''''_Int_Int_buf [0]))
        \memOut_CTf''''''''_f''''''''_Int_Int_buf  <= {68'd0, 1'd0};
      else if (((! \memOut_CTf''''''''_f''''''''_Int_Int_rbuf_r ) && (! \memOut_CTf''''''''_f''''''''_Int_Int_buf [0])))
        \memOut_CTf''''''''_f''''''''_Int_Int_buf  <= \memOut_CTf''''''''_f''''''''_Int_Int_d ;
  
  /* destruct (Ty Pointer_CTf''''''''_f''''''''_Int_Int,
          Dcon Pointer_CTf''''''''_f''''''''_Int_Int) : (scfarg_0_1_1_argbuf,Pointer_CTf''''''''_f''''''''_Int_Int) > [(destructReadIn_CTf''''''''_f''''''''_Int_Int,Word16#)] */
  assign \destructReadIn_CTf''''''''_f''''''''_Int_Int_d  = {scfarg_0_1_1_argbuf_d[16:1],
                                                             scfarg_0_1_1_argbuf_d[0]};
  assign scfarg_0_1_1_argbuf_r = \destructReadIn_CTf''''''''_f''''''''_Int_Int_r ;
  
  /* dcon (Ty MemIn_CTf''''''''_f''''''''_Int_Int,
      Dcon ReadIn_CTf''''''''_f''''''''_Int_Int) : [(destructReadIn_CTf''''''''_f''''''''_Int_Int,Word16#)] > (dconReadIn_CTf''''''''_f''''''''_Int_Int,MemIn_CTf''''''''_f''''''''_Int_Int) */
  assign \dconReadIn_CTf''''''''_f''''''''_Int_Int_d  = \ReadIn_CTf''''''''_f''''''''_Int_Int_dc ((& {\destructReadIn_CTf''''''''_f''''''''_Int_Int_d [0]}), \destructReadIn_CTf''''''''_f''''''''_Int_Int_d );
  assign {\destructReadIn_CTf''''''''_f''''''''_Int_Int_r } = {1 {(\dconReadIn_CTf''''''''_f''''''''_Int_Int_r  && \dconReadIn_CTf''''''''_f''''''''_Int_Int_d [0])}};
  
  /* destruct (Ty MemOut_CTf''''''''_f''''''''_Int_Int,
          Dcon ReadOut_CTf''''''''_f''''''''_Int_Int) : (memReadOut_CTf''''''''_f''''''''_Int_Int,MemOut_CTf''''''''_f''''''''_Int_Int) > [(readPointer_CTf''''''''_f''''''''_Int_Intscfarg_0_1_1_argbuf,CTf''''''''_f''''''''_Int_Int)] */
  assign \readPointer_CTf''''''''_f''''''''_Int_Intscfarg_0_1_1_argbuf_d  = {\memReadOut_CTf''''''''_f''''''''_Int_Int_d [68:2],
                                                                             \memReadOut_CTf''''''''_f''''''''_Int_Int_d [0]};
  assign \memReadOut_CTf''''''''_f''''''''_Int_Int_r  = \readPointer_CTf''''''''_f''''''''_Int_Intscfarg_0_1_1_argbuf_r ;
  
  /* mergectrl (Ty C5,
           Ty CTf''''''''_f''''''''_Int_Int) : [(lizzieLet10_1_argbuf,CTf''''''''_f''''''''_Int_Int),
                                                (lizzieLet33_1_argbuf,CTf''''''''_f''''''''_Int_Int),
                                                (lizzieLet40_1_argbuf,CTf''''''''_f''''''''_Int_Int),
                                                (lizzieLet41_1_argbuf,CTf''''''''_f''''''''_Int_Int),
                                                (lizzieLet42_1_argbuf,CTf''''''''_f''''''''_Int_Int)] > (writeMerge_choice_CTf''''''''_f''''''''_Int_Int,C5) (writeMerge_data_CTf''''''''_f''''''''_Int_Int,CTf''''''''_f''''''''_Int_Int) */
  logic [4:0] lizzieLet10_1_argbuf_select_d;
  assign lizzieLet10_1_argbuf_select_d = ((| lizzieLet10_1_argbuf_select_q) ? lizzieLet10_1_argbuf_select_q :
                                          (lizzieLet10_1_argbuf_d[0] ? 5'd1 :
                                           (lizzieLet33_1_argbuf_d[0] ? 5'd2 :
                                            (lizzieLet40_1_argbuf_d[0] ? 5'd4 :
                                             (lizzieLet41_1_argbuf_d[0] ? 5'd8 :
                                              (lizzieLet42_1_argbuf_d[0] ? 5'd16 :
                                               5'd0))))));
  logic [4:0] lizzieLet10_1_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet10_1_argbuf_select_q <= 5'd0;
    else
      lizzieLet10_1_argbuf_select_q <= (lizzieLet10_1_argbuf_done ? 5'd0 :
                                        lizzieLet10_1_argbuf_select_d);
  logic [1:0] lizzieLet10_1_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet10_1_argbuf_emit_q <= 2'd0;
    else
      lizzieLet10_1_argbuf_emit_q <= (lizzieLet10_1_argbuf_done ? 2'd0 :
                                      lizzieLet10_1_argbuf_emit_d);
  logic [1:0] lizzieLet10_1_argbuf_emit_d;
  assign lizzieLet10_1_argbuf_emit_d = (lizzieLet10_1_argbuf_emit_q | ({\writeMerge_choice_CTf''''''''_f''''''''_Int_Int_d [0],
                                                                        \writeMerge_data_CTf''''''''_f''''''''_Int_Int_d [0]} & {\writeMerge_choice_CTf''''''''_f''''''''_Int_Int_r ,
                                                                                                                                 \writeMerge_data_CTf''''''''_f''''''''_Int_Int_r }));
  logic lizzieLet10_1_argbuf_done;
  assign lizzieLet10_1_argbuf_done = (& lizzieLet10_1_argbuf_emit_d);
  assign {lizzieLet42_1_argbuf_r,
          lizzieLet41_1_argbuf_r,
          lizzieLet40_1_argbuf_r,
          lizzieLet33_1_argbuf_r,
          lizzieLet10_1_argbuf_r} = (lizzieLet10_1_argbuf_done ? lizzieLet10_1_argbuf_select_d :
                                     5'd0);
  assign \writeMerge_data_CTf''''''''_f''''''''_Int_Int_d  = ((lizzieLet10_1_argbuf_select_d[0] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet10_1_argbuf_d :
                                                              ((lizzieLet10_1_argbuf_select_d[1] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet33_1_argbuf_d :
                                                               ((lizzieLet10_1_argbuf_select_d[2] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet40_1_argbuf_d :
                                                                ((lizzieLet10_1_argbuf_select_d[3] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet41_1_argbuf_d :
                                                                 ((lizzieLet10_1_argbuf_select_d[4] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet42_1_argbuf_d :
                                                                  {67'd0, 1'd0})))));
  assign \writeMerge_choice_CTf''''''''_f''''''''_Int_Int_d  = ((lizzieLet10_1_argbuf_select_d[0] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C1_5_dc(1'd1) :
                                                                ((lizzieLet10_1_argbuf_select_d[1] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C2_5_dc(1'd1) :
                                                                 ((lizzieLet10_1_argbuf_select_d[2] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C3_5_dc(1'd1) :
                                                                  ((lizzieLet10_1_argbuf_select_d[3] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C4_5_dc(1'd1) :
                                                                   ((lizzieLet10_1_argbuf_select_d[4] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C5_5_dc(1'd1) :
                                                                    {3'd0, 1'd0})))));
  
  /* demux (Ty C5,
       Ty Pointer_CTf''''''''_f''''''''_Int_Int) : (writeMerge_choice_CTf''''''''_f''''''''_Int_Int,C5) (demuxWriteResult_CTf''''''''_f''''''''_Int_Int,Pointer_CTf''''''''_f''''''''_Int_Int) > [(writeCTf''''''''_f''''''''_Int_IntlizzieLet10_1_argbuf,Pointer_CTf''''''''_f''''''''_Int_Int),
                                                                                                                                                                                                  (writeCTf''''''''_f''''''''_Int_IntlizzieLet33_1_argbuf,Pointer_CTf''''''''_f''''''''_Int_Int),
                                                                                                                                                                                                  (writeCTf''''''''_f''''''''_Int_IntlizzieLet40_1_argbuf,Pointer_CTf''''''''_f''''''''_Int_Int),
                                                                                                                                                                                                  (writeCTf''''''''_f''''''''_Int_IntlizzieLet41_1_argbuf,Pointer_CTf''''''''_f''''''''_Int_Int),
                                                                                                                                                                                                  (writeCTf''''''''_f''''''''_Int_IntlizzieLet42_1_argbuf,Pointer_CTf''''''''_f''''''''_Int_Int)] */
  logic [4:0] \demuxWriteResult_CTf''''''''_f''''''''_Int_Int_onehotd ;
  always_comb
    if ((\writeMerge_choice_CTf''''''''_f''''''''_Int_Int_d [0] && \demuxWriteResult_CTf''''''''_f''''''''_Int_Int_d [0]))
      unique case (\writeMerge_choice_CTf''''''''_f''''''''_Int_Int_d [3:1])
        3'd0:
          \demuxWriteResult_CTf''''''''_f''''''''_Int_Int_onehotd  = 5'd1;
        3'd1:
          \demuxWriteResult_CTf''''''''_f''''''''_Int_Int_onehotd  = 5'd2;
        3'd2:
          \demuxWriteResult_CTf''''''''_f''''''''_Int_Int_onehotd  = 5'd4;
        3'd3:
          \demuxWriteResult_CTf''''''''_f''''''''_Int_Int_onehotd  = 5'd8;
        3'd4:
          \demuxWriteResult_CTf''''''''_f''''''''_Int_Int_onehotd  = 5'd16;
        default:
          \demuxWriteResult_CTf''''''''_f''''''''_Int_Int_onehotd  = 5'd0;
      endcase
    else
      \demuxWriteResult_CTf''''''''_f''''''''_Int_Int_onehotd  = 5'd0;
  assign \writeCTf''''''''_f''''''''_Int_IntlizzieLet10_1_argbuf_d  = {\demuxWriteResult_CTf''''''''_f''''''''_Int_Int_d [16:1],
                                                                       \demuxWriteResult_CTf''''''''_f''''''''_Int_Int_onehotd [0]};
  assign \writeCTf''''''''_f''''''''_Int_IntlizzieLet33_1_argbuf_d  = {\demuxWriteResult_CTf''''''''_f''''''''_Int_Int_d [16:1],
                                                                       \demuxWriteResult_CTf''''''''_f''''''''_Int_Int_onehotd [1]};
  assign \writeCTf''''''''_f''''''''_Int_IntlizzieLet40_1_argbuf_d  = {\demuxWriteResult_CTf''''''''_f''''''''_Int_Int_d [16:1],
                                                                       \demuxWriteResult_CTf''''''''_f''''''''_Int_Int_onehotd [2]};
  assign \writeCTf''''''''_f''''''''_Int_IntlizzieLet41_1_argbuf_d  = {\demuxWriteResult_CTf''''''''_f''''''''_Int_Int_d [16:1],
                                                                       \demuxWriteResult_CTf''''''''_f''''''''_Int_Int_onehotd [3]};
  assign \writeCTf''''''''_f''''''''_Int_IntlizzieLet42_1_argbuf_d  = {\demuxWriteResult_CTf''''''''_f''''''''_Int_Int_d [16:1],
                                                                       \demuxWriteResult_CTf''''''''_f''''''''_Int_Int_onehotd [4]};
  assign \demuxWriteResult_CTf''''''''_f''''''''_Int_Int_r  = (| (\demuxWriteResult_CTf''''''''_f''''''''_Int_Int_onehotd  & {\writeCTf''''''''_f''''''''_Int_IntlizzieLet42_1_argbuf_r ,
                                                                                                                              \writeCTf''''''''_f''''''''_Int_IntlizzieLet41_1_argbuf_r ,
                                                                                                                              \writeCTf''''''''_f''''''''_Int_IntlizzieLet40_1_argbuf_r ,
                                                                                                                              \writeCTf''''''''_f''''''''_Int_IntlizzieLet33_1_argbuf_r ,
                                                                                                                              \writeCTf''''''''_f''''''''_Int_IntlizzieLet10_1_argbuf_r }));
  assign \writeMerge_choice_CTf''''''''_f''''''''_Int_Int_r  = \demuxWriteResult_CTf''''''''_f''''''''_Int_Int_r ;
  
  /* dcon (Ty MemIn_CTf''''''''_f''''''''_Int_Int,
      Dcon WriteIn_CTf''''''''_f''''''''_Int_Int) : [(forkHP1_CTf''''''''_f''''''''_Int_In2,Word16#),
                                                     (writeMerge_data_CTf''''''''_f''''''''_Int_Int,CTf''''''''_f''''''''_Int_Int)] > (dconWriteIn_CTf''''''''_f''''''''_Int_Int,MemIn_CTf''''''''_f''''''''_Int_Int) */
  assign \dconWriteIn_CTf''''''''_f''''''''_Int_Int_d  = \WriteIn_CTf''''''''_f''''''''_Int_Int_dc ((& {\forkHP1_CTf''''''''_f''''''''_Int_In2_d [0],
                                                                                                        \writeMerge_data_CTf''''''''_f''''''''_Int_Int_d [0]}), \forkHP1_CTf''''''''_f''''''''_Int_In2_d , \writeMerge_data_CTf''''''''_f''''''''_Int_Int_d );
  assign {\forkHP1_CTf''''''''_f''''''''_Int_In2_r ,
          \writeMerge_data_CTf''''''''_f''''''''_Int_Int_r } = {2 {(\dconWriteIn_CTf''''''''_f''''''''_Int_Int_r  && \dconWriteIn_CTf''''''''_f''''''''_Int_Int_d [0])}};
  
  /* dcon (Ty Pointer_CTf''''''''_f''''''''_Int_Int,
      Dcon Pointer_CTf''''''''_f''''''''_Int_Int) : [(forkHP1_CTf''''''''_f''''''''_Int_In3,Word16#)] > (dconPtr_CTf''''''''_f''''''''_Int_Int,Pointer_CTf''''''''_f''''''''_Int_Int) */
  assign \dconPtr_CTf''''''''_f''''''''_Int_Int_d  = \Pointer_CTf''''''''_f''''''''_Int_Int_dc ((& {\forkHP1_CTf''''''''_f''''''''_Int_In3_d [0]}), \forkHP1_CTf''''''''_f''''''''_Int_In3_d );
  assign {\forkHP1_CTf''''''''_f''''''''_Int_In3_r } = {1 {(\dconPtr_CTf''''''''_f''''''''_Int_Int_r  && \dconPtr_CTf''''''''_f''''''''_Int_Int_d [0])}};
  
  /* demux (Ty MemOut_CTf''''''''_f''''''''_Int_Int,
       Ty Pointer_CTf''''''''_f''''''''_Int_Int) : (memWriteOut_CTf''''''''_f''''''''_Int_Int,MemOut_CTf''''''''_f''''''''_Int_Int) (dconPtr_CTf''''''''_f''''''''_Int_Int,Pointer_CTf''''''''_f''''''''_Int_Int) > [(_83,Pointer_CTf''''''''_f''''''''_Int_Int),
                                                                                                                                                                                                                     (demuxWriteResult_CTf''''''''_f''''''''_Int_Int,Pointer_CTf''''''''_f''''''''_Int_Int)] */
  logic [1:0] \dconPtr_CTf''''''''_f''''''''_Int_Int_onehotd ;
  always_comb
    if ((\memWriteOut_CTf''''''''_f''''''''_Int_Int_d [0] && \dconPtr_CTf''''''''_f''''''''_Int_Int_d [0]))
      unique case (\memWriteOut_CTf''''''''_f''''''''_Int_Int_d [1:1])
        1'd0: \dconPtr_CTf''''''''_f''''''''_Int_Int_onehotd  = 2'd1;
        1'd1: \dconPtr_CTf''''''''_f''''''''_Int_Int_onehotd  = 2'd2;
        default: \dconPtr_CTf''''''''_f''''''''_Int_Int_onehotd  = 2'd0;
      endcase
    else \dconPtr_CTf''''''''_f''''''''_Int_Int_onehotd  = 2'd0;
  assign _83_d = {\dconPtr_CTf''''''''_f''''''''_Int_Int_d [16:1],
                  \dconPtr_CTf''''''''_f''''''''_Int_Int_onehotd [0]};
  assign \demuxWriteResult_CTf''''''''_f''''''''_Int_Int_d  = {\dconPtr_CTf''''''''_f''''''''_Int_Int_d [16:1],
                                                               \dconPtr_CTf''''''''_f''''''''_Int_Int_onehotd [1]};
  assign \dconPtr_CTf''''''''_f''''''''_Int_Int_r  = (| (\dconPtr_CTf''''''''_f''''''''_Int_Int_onehotd  & {\demuxWriteResult_CTf''''''''_f''''''''_Int_Int_r ,
                                                                                                            _83_r}));
  assign \memWriteOut_CTf''''''''_f''''''''_Int_Int_r  = \dconPtr_CTf''''''''_f''''''''_Int_Int_r ;
  
  /* const (Ty Word16#,
       Lit 0) : (go_1_dummy_write_QTree_Int,Go) > (initHP_QTree_Int,Word16#) */
  assign initHP_QTree_Int_d = {16'd0,
                               go_1_dummy_write_QTree_Int_d[0]};
  assign go_1_dummy_write_QTree_Int_r = initHP_QTree_Int_r;
  
  /* const (Ty Word16#,
       Lit 1) : (incrHP_QTree_Int1,Go) > (incrHP_QTree_Int,Word16#) */
  assign incrHP_QTree_Int_d = {16'd1, incrHP_QTree_Int1_d[0]};
  assign incrHP_QTree_Int1_r = incrHP_QTree_Int_r;
  
  /* merge (Ty Go) : [(go_2_dummy_write_QTree_Int,Go),
                 (incrHP_QTree_Int2,Go)] > (incrHP_mergeQTree_Int,Go) */
  logic [1:0] incrHP_mergeQTree_Int_selected;
  logic [1:0] incrHP_mergeQTree_Int_select;
  always_comb
    begin
      incrHP_mergeQTree_Int_selected = 2'd0;
      if ((| incrHP_mergeQTree_Int_select))
        incrHP_mergeQTree_Int_selected = incrHP_mergeQTree_Int_select;
      else
        if (go_2_dummy_write_QTree_Int_d[0])
          incrHP_mergeQTree_Int_selected[0] = 1'd1;
        else if (incrHP_QTree_Int2_d[0])
          incrHP_mergeQTree_Int_selected[1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeQTree_Int_select <= 2'd0;
    else
      incrHP_mergeQTree_Int_select <= (incrHP_mergeQTree_Int_r ? 2'd0 :
                                       incrHP_mergeQTree_Int_selected);
  always_comb
    if (incrHP_mergeQTree_Int_selected[0])
      incrHP_mergeQTree_Int_d = go_2_dummy_write_QTree_Int_d;
    else if (incrHP_mergeQTree_Int_selected[1])
      incrHP_mergeQTree_Int_d = incrHP_QTree_Int2_d;
    else incrHP_mergeQTree_Int_d = 1'd0;
  assign {incrHP_QTree_Int2_r,
          go_2_dummy_write_QTree_Int_r} = (incrHP_mergeQTree_Int_r ? incrHP_mergeQTree_Int_selected :
                                           2'd0);
  
  /* fork (Ty Go) : (incrHP_mergeQTree_Int_buf,Go) > [(incrHP_QTree_Int1,Go),
                                                 (incrHP_QTree_Int2,Go)] */
  logic [1:0] incrHP_mergeQTree_Int_buf_emitted;
  logic [1:0] incrHP_mergeQTree_Int_buf_done;
  assign incrHP_QTree_Int1_d = (incrHP_mergeQTree_Int_buf_d[0] && (! incrHP_mergeQTree_Int_buf_emitted[0]));
  assign incrHP_QTree_Int2_d = (incrHP_mergeQTree_Int_buf_d[0] && (! incrHP_mergeQTree_Int_buf_emitted[1]));
  assign incrHP_mergeQTree_Int_buf_done = (incrHP_mergeQTree_Int_buf_emitted | ({incrHP_QTree_Int2_d[0],
                                                                                 incrHP_QTree_Int1_d[0]} & {incrHP_QTree_Int2_r,
                                                                                                            incrHP_QTree_Int1_r}));
  assign incrHP_mergeQTree_Int_buf_r = (& incrHP_mergeQTree_Int_buf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeQTree_Int_buf_emitted <= 2'd0;
    else
      incrHP_mergeQTree_Int_buf_emitted <= (incrHP_mergeQTree_Int_buf_r ? 2'd0 :
                                            incrHP_mergeQTree_Int_buf_done);
  
  /* op_add (Ty Word16#) : (incrHP_QTree_Int,Word16#) (forkHP1_QTree_Int,Word16#) > (addHP_QTree_Int,Word16#) */
  assign addHP_QTree_Int_d = {(incrHP_QTree_Int_d[16:1] + forkHP1_QTree_Int_d[16:1]),
                              (incrHP_QTree_Int_d[0] && forkHP1_QTree_Int_d[0])};
  assign {incrHP_QTree_Int_r,
          forkHP1_QTree_Int_r} = {2 {(addHP_QTree_Int_r && addHP_QTree_Int_d[0])}};
  
  /* merge (Ty Word16#) : [(initHP_QTree_Int,Word16#),
                      (addHP_QTree_Int,Word16#)] > (mergeHP_QTree_Int,Word16#) */
  logic [1:0] mergeHP_QTree_Int_selected;
  logic [1:0] mergeHP_QTree_Int_select;
  always_comb
    begin
      mergeHP_QTree_Int_selected = 2'd0;
      if ((| mergeHP_QTree_Int_select))
        mergeHP_QTree_Int_selected = mergeHP_QTree_Int_select;
      else
        if (initHP_QTree_Int_d[0]) mergeHP_QTree_Int_selected[0] = 1'd1;
        else if (addHP_QTree_Int_d[0])
          mergeHP_QTree_Int_selected[1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_QTree_Int_select <= 2'd0;
    else
      mergeHP_QTree_Int_select <= (mergeHP_QTree_Int_r ? 2'd0 :
                                   mergeHP_QTree_Int_selected);
  always_comb
    if (mergeHP_QTree_Int_selected[0])
      mergeHP_QTree_Int_d = initHP_QTree_Int_d;
    else if (mergeHP_QTree_Int_selected[1])
      mergeHP_QTree_Int_d = addHP_QTree_Int_d;
    else mergeHP_QTree_Int_d = {16'd0, 1'd0};
  assign {addHP_QTree_Int_r,
          initHP_QTree_Int_r} = (mergeHP_QTree_Int_r ? mergeHP_QTree_Int_selected :
                                 2'd0);
  
  /* buf (Ty Go) : (incrHP_mergeQTree_Int,Go) > (incrHP_mergeQTree_Int_buf,Go) */
  Go_t incrHP_mergeQTree_Int_bufchan_d;
  logic incrHP_mergeQTree_Int_bufchan_r;
  assign incrHP_mergeQTree_Int_r = ((! incrHP_mergeQTree_Int_bufchan_d[0]) || incrHP_mergeQTree_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeQTree_Int_bufchan_d <= 1'd0;
    else
      if (incrHP_mergeQTree_Int_r)
        incrHP_mergeQTree_Int_bufchan_d <= incrHP_mergeQTree_Int_d;
  Go_t incrHP_mergeQTree_Int_bufchan_buf;
  assign incrHP_mergeQTree_Int_bufchan_r = (! incrHP_mergeQTree_Int_bufchan_buf[0]);
  assign incrHP_mergeQTree_Int_buf_d = (incrHP_mergeQTree_Int_bufchan_buf[0] ? incrHP_mergeQTree_Int_bufchan_buf :
                                        incrHP_mergeQTree_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeQTree_Int_bufchan_buf <= 1'd0;
    else
      if ((incrHP_mergeQTree_Int_buf_r && incrHP_mergeQTree_Int_bufchan_buf[0]))
        incrHP_mergeQTree_Int_bufchan_buf <= 1'd0;
      else if (((! incrHP_mergeQTree_Int_buf_r) && (! incrHP_mergeQTree_Int_bufchan_buf[0])))
        incrHP_mergeQTree_Int_bufchan_buf <= incrHP_mergeQTree_Int_bufchan_d;
  
  /* buf (Ty Word16#) : (mergeHP_QTree_Int,Word16#) > (mergeHP_QTree_Int_buf,Word16#) */
  \Word16#_t  mergeHP_QTree_Int_bufchan_d;
  logic mergeHP_QTree_Int_bufchan_r;
  assign mergeHP_QTree_Int_r = ((! mergeHP_QTree_Int_bufchan_d[0]) || mergeHP_QTree_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_QTree_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (mergeHP_QTree_Int_r)
        mergeHP_QTree_Int_bufchan_d <= mergeHP_QTree_Int_d;
  \Word16#_t  mergeHP_QTree_Int_bufchan_buf;
  assign mergeHP_QTree_Int_bufchan_r = (! mergeHP_QTree_Int_bufchan_buf[0]);
  assign mergeHP_QTree_Int_buf_d = (mergeHP_QTree_Int_bufchan_buf[0] ? mergeHP_QTree_Int_bufchan_buf :
                                    mergeHP_QTree_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      mergeHP_QTree_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((mergeHP_QTree_Int_buf_r && mergeHP_QTree_Int_bufchan_buf[0]))
        mergeHP_QTree_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! mergeHP_QTree_Int_buf_r) && (! mergeHP_QTree_Int_bufchan_buf[0])))
        mergeHP_QTree_Int_bufchan_buf <= mergeHP_QTree_Int_bufchan_d;
  
  /* sink (Ty Word16#) : (forkHP1_QTree_Int_snk,Word16#) > */
  assign {forkHP1_QTree_Int_snk_r,
          forkHP1_QTree_Int_snk_dout} = {forkHP1_QTree_Int_snk_rout,
                                         forkHP1_QTree_Int_snk_d};
  
  /* source (Ty Go) : > (\QTree_Int_src,Go) */
  
  /* fork (Ty Go) : (\QTree_Int_src,Go) > [(go_1_dummy_write_QTree_Int,Go),
                                      (go_2_dummy_write_QTree_Int,Go)] */
  logic [1:0] \\QTree_Int_src_emitted ;
  logic [1:0] \\QTree_Int_src_done ;
  assign go_1_dummy_write_QTree_Int_d = (\\QTree_Int_src_d [0] && (! \\QTree_Int_src_emitted [0]));
  assign go_2_dummy_write_QTree_Int_d = (\\QTree_Int_src_d [0] && (! \\QTree_Int_src_emitted [1]));
  assign \\QTree_Int_src_done  = (\\QTree_Int_src_emitted  | ({go_2_dummy_write_QTree_Int_d[0],
                                                               go_1_dummy_write_QTree_Int_d[0]} & {go_2_dummy_write_QTree_Int_r,
                                                                                                   go_1_dummy_write_QTree_Int_r}));
  assign \\QTree_Int_src_r  = (& \\QTree_Int_src_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \\QTree_Int_src_emitted  <= 2'd0;
    else
      \\QTree_Int_src_emitted  <= (\\QTree_Int_src_r  ? 2'd0 :
                                   \\QTree_Int_src_done );
  
  /* source (Ty QTree_Int) : > (dummy_write_QTree_Int,QTree_Int) */
  
  /* sink (Ty Pointer_QTree_Int) : (dummy_write_QTree_Int_sink,Pointer_QTree_Int) > */
  assign {dummy_write_QTree_Int_sink_r,
          dummy_write_QTree_Int_sink_dout} = {dummy_write_QTree_Int_sink_rout,
                                              dummy_write_QTree_Int_sink_d};
  
  /* fork (Ty Word16#) : (mergeHP_QTree_Int_buf,Word16#) > [(forkHP1_QTree_Int,Word16#),
                                                       (forkHP1_QTree_Int_snk,Word16#),
                                                       (forkHP1_QTree_In3,Word16#),
                                                       (forkHP1_QTree_In4,Word16#)] */
  logic [3:0] mergeHP_QTree_Int_buf_emitted;
  logic [3:0] mergeHP_QTree_Int_buf_done;
  assign forkHP1_QTree_Int_d = {mergeHP_QTree_Int_buf_d[16:1],
                                (mergeHP_QTree_Int_buf_d[0] && (! mergeHP_QTree_Int_buf_emitted[0]))};
  assign forkHP1_QTree_Int_snk_d = {mergeHP_QTree_Int_buf_d[16:1],
                                    (mergeHP_QTree_Int_buf_d[0] && (! mergeHP_QTree_Int_buf_emitted[1]))};
  assign forkHP1_QTree_In3_d = {mergeHP_QTree_Int_buf_d[16:1],
                                (mergeHP_QTree_Int_buf_d[0] && (! mergeHP_QTree_Int_buf_emitted[2]))};
  assign forkHP1_QTree_In4_d = {mergeHP_QTree_Int_buf_d[16:1],
                                (mergeHP_QTree_Int_buf_d[0] && (! mergeHP_QTree_Int_buf_emitted[3]))};
  assign mergeHP_QTree_Int_buf_done = (mergeHP_QTree_Int_buf_emitted | ({forkHP1_QTree_In4_d[0],
                                                                         forkHP1_QTree_In3_d[0],
                                                                         forkHP1_QTree_Int_snk_d[0],
                                                                         forkHP1_QTree_Int_d[0]} & {forkHP1_QTree_In4_r,
                                                                                                    forkHP1_QTree_In3_r,
                                                                                                    forkHP1_QTree_Int_snk_r,
                                                                                                    forkHP1_QTree_Int_r}));
  assign mergeHP_QTree_Int_buf_r = (& mergeHP_QTree_Int_buf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_QTree_Int_buf_emitted <= 4'd0;
    else
      mergeHP_QTree_Int_buf_emitted <= (mergeHP_QTree_Int_buf_r ? 4'd0 :
                                        mergeHP_QTree_Int_buf_done);
  
  /* mergectrl (Ty C2,
           Ty MemIn_QTree_Int) : [(dconReadIn_QTree_Int,MemIn_QTree_Int),
                                  (dconWriteIn_QTree_Int,MemIn_QTree_Int)] > (memMergeChoice_QTree_Int,C2) (memMergeIn_QTree_Int,MemIn_QTree_Int) */
  logic [1:0] dconReadIn_QTree_Int_select_d;
  assign dconReadIn_QTree_Int_select_d = ((| dconReadIn_QTree_Int_select_q) ? dconReadIn_QTree_Int_select_q :
                                          (dconReadIn_QTree_Int_d[0] ? 2'd1 :
                                           (dconWriteIn_QTree_Int_d[0] ? 2'd2 :
                                            2'd0)));
  logic [1:0] dconReadIn_QTree_Int_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) dconReadIn_QTree_Int_select_q <= 2'd0;
    else
      dconReadIn_QTree_Int_select_q <= (dconReadIn_QTree_Int_done ? 2'd0 :
                                        dconReadIn_QTree_Int_select_d);
  logic [1:0] dconReadIn_QTree_Int_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) dconReadIn_QTree_Int_emit_q <= 2'd0;
    else
      dconReadIn_QTree_Int_emit_q <= (dconReadIn_QTree_Int_done ? 2'd0 :
                                      dconReadIn_QTree_Int_emit_d);
  logic [1:0] dconReadIn_QTree_Int_emit_d;
  assign dconReadIn_QTree_Int_emit_d = (dconReadIn_QTree_Int_emit_q | ({memMergeChoice_QTree_Int_d[0],
                                                                        memMergeIn_QTree_Int_d[0]} & {memMergeChoice_QTree_Int_r,
                                                                                                      memMergeIn_QTree_Int_r}));
  logic dconReadIn_QTree_Int_done;
  assign dconReadIn_QTree_Int_done = (& dconReadIn_QTree_Int_emit_d);
  assign {dconWriteIn_QTree_Int_r,
          dconReadIn_QTree_Int_r} = (dconReadIn_QTree_Int_done ? dconReadIn_QTree_Int_select_d :
                                     2'd0);
  assign memMergeIn_QTree_Int_d = ((dconReadIn_QTree_Int_select_d[0] && (! dconReadIn_QTree_Int_emit_q[0])) ? dconReadIn_QTree_Int_d :
                                   ((dconReadIn_QTree_Int_select_d[1] && (! dconReadIn_QTree_Int_emit_q[0])) ? dconWriteIn_QTree_Int_d :
                                    {83'd0, 1'd0}));
  assign memMergeChoice_QTree_Int_d = ((dconReadIn_QTree_Int_select_d[0] && (! dconReadIn_QTree_Int_emit_q[1])) ? C1_2_dc(1'd1) :
                                       ((dconReadIn_QTree_Int_select_d[1] && (! dconReadIn_QTree_Int_emit_q[1])) ? C2_2_dc(1'd1) :
                                        {1'd0, 1'd0}));
  
  /* bram (Ty MemIn_QTree_Int,
      Ty MemOut_QTree_Int) : (memMergeIn_QTree_Int_dbuf,MemIn_QTree_Int) > (memOut_QTree_Int,MemOut_QTree_Int) */
  logic [65:0] memMergeIn_QTree_Int_dbuf_mem[65535:0];
  logic [15:0] memMergeIn_QTree_Int_dbuf_address;
  logic [65:0] memMergeIn_QTree_Int_dbuf_din;
  logic [65:0] memOut_QTree_Int_q;
  logic memOut_QTree_Int_valid;
  logic memMergeIn_QTree_Int_dbuf_we;
  logic memOut_QTree_Int_we;
  assign memMergeIn_QTree_Int_dbuf_din = memMergeIn_QTree_Int_dbuf_d[83:18];
  assign memMergeIn_QTree_Int_dbuf_address = memMergeIn_QTree_Int_dbuf_d[17:2];
  assign memMergeIn_QTree_Int_dbuf_we = (memMergeIn_QTree_Int_dbuf_d[1:1] && memMergeIn_QTree_Int_dbuf_d[0]);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        memOut_QTree_Int_we <= 1'd0;
        memOut_QTree_Int_valid <= 1'd0;
      end
    else
      begin
        memOut_QTree_Int_we <= memMergeIn_QTree_Int_dbuf_we;
        memOut_QTree_Int_valid <= memMergeIn_QTree_Int_dbuf_d[0];
        if (memMergeIn_QTree_Int_dbuf_we)
          begin
            memMergeIn_QTree_Int_dbuf_mem[memMergeIn_QTree_Int_dbuf_address] <= memMergeIn_QTree_Int_dbuf_din;
            memOut_QTree_Int_q <= memMergeIn_QTree_Int_dbuf_din;
          end
        else
          memOut_QTree_Int_q <= memMergeIn_QTree_Int_dbuf_mem[memMergeIn_QTree_Int_dbuf_address];
      end
  assign memOut_QTree_Int_d = {memOut_QTree_Int_q,
                               memOut_QTree_Int_we,
                               memOut_QTree_Int_valid};
  assign memMergeIn_QTree_Int_dbuf_r = ((! memOut_QTree_Int_valid) || memOut_QTree_Int_r);
  logic [31:0] profiling_MemIn_QTree_Int_read;
  logic [31:0] profiling_MemIn_QTree_Int_write;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        profiling_MemIn_QTree_Int_write <= 0;
        profiling_MemIn_QTree_Int_read <= 0;
      end
    else
      if ((memMergeIn_QTree_Int_dbuf_we == 1'd1))
        profiling_MemIn_QTree_Int_write <= (profiling_MemIn_QTree_Int_write + 1);
      else
        if ((memOut_QTree_Int_valid == 1'd1))
          profiling_MemIn_QTree_Int_read <= (profiling_MemIn_QTree_Int_read + 1);
  
  /* demux (Ty C2,
       Ty MemOut_QTree_Int) : (memMergeChoice_QTree_Int,C2) (memOut_QTree_Int_dbuf,MemOut_QTree_Int) > [(memReadOut_QTree_Int,MemOut_QTree_Int),
                                                                                                        (memWriteOut_QTree_Int,MemOut_QTree_Int)] */
  logic [1:0] memOut_QTree_Int_dbuf_onehotd;
  always_comb
    if ((memMergeChoice_QTree_Int_d[0] && memOut_QTree_Int_dbuf_d[0]))
      unique case (memMergeChoice_QTree_Int_d[1:1])
        1'd0: memOut_QTree_Int_dbuf_onehotd = 2'd1;
        1'd1: memOut_QTree_Int_dbuf_onehotd = 2'd2;
        default: memOut_QTree_Int_dbuf_onehotd = 2'd0;
      endcase
    else memOut_QTree_Int_dbuf_onehotd = 2'd0;
  assign memReadOut_QTree_Int_d = {memOut_QTree_Int_dbuf_d[67:1],
                                   memOut_QTree_Int_dbuf_onehotd[0]};
  assign memWriteOut_QTree_Int_d = {memOut_QTree_Int_dbuf_d[67:1],
                                    memOut_QTree_Int_dbuf_onehotd[1]};
  assign memOut_QTree_Int_dbuf_r = (| (memOut_QTree_Int_dbuf_onehotd & {memWriteOut_QTree_Int_r,
                                                                        memReadOut_QTree_Int_r}));
  assign memMergeChoice_QTree_Int_r = memOut_QTree_Int_dbuf_r;
  
  /* dbuf (Ty MemIn_QTree_Int) : (memMergeIn_QTree_Int_rbuf,MemIn_QTree_Int) > (memMergeIn_QTree_Int_dbuf,MemIn_QTree_Int) */
  assign memMergeIn_QTree_Int_rbuf_r = ((! memMergeIn_QTree_Int_dbuf_d[0]) || memMergeIn_QTree_Int_dbuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memMergeIn_QTree_Int_dbuf_d <= {83'd0, 1'd0};
    else
      if (memMergeIn_QTree_Int_rbuf_r)
        memMergeIn_QTree_Int_dbuf_d <= memMergeIn_QTree_Int_rbuf_d;
  
  /* rbuf (Ty MemIn_QTree_Int) : (memMergeIn_QTree_Int,MemIn_QTree_Int) > (memMergeIn_QTree_Int_rbuf,MemIn_QTree_Int) */
  MemIn_QTree_Int_t memMergeIn_QTree_Int_buf;
  assign memMergeIn_QTree_Int_r = (! memMergeIn_QTree_Int_buf[0]);
  assign memMergeIn_QTree_Int_rbuf_d = (memMergeIn_QTree_Int_buf[0] ? memMergeIn_QTree_Int_buf :
                                        memMergeIn_QTree_Int_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memMergeIn_QTree_Int_buf <= {83'd0, 1'd0};
    else
      if ((memMergeIn_QTree_Int_rbuf_r && memMergeIn_QTree_Int_buf[0]))
        memMergeIn_QTree_Int_buf <= {83'd0, 1'd0};
      else if (((! memMergeIn_QTree_Int_rbuf_r) && (! memMergeIn_QTree_Int_buf[0])))
        memMergeIn_QTree_Int_buf <= memMergeIn_QTree_Int_d;
  
  /* dbuf (Ty MemOut_QTree_Int) : (memOut_QTree_Int_rbuf,MemOut_QTree_Int) > (memOut_QTree_Int_dbuf,MemOut_QTree_Int) */
  assign memOut_QTree_Int_rbuf_r = ((! memOut_QTree_Int_dbuf_d[0]) || memOut_QTree_Int_dbuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memOut_QTree_Int_dbuf_d <= {67'd0, 1'd0};
    else
      if (memOut_QTree_Int_rbuf_r)
        memOut_QTree_Int_dbuf_d <= memOut_QTree_Int_rbuf_d;
  
  /* rbuf (Ty MemOut_QTree_Int) : (memOut_QTree_Int,MemOut_QTree_Int) > (memOut_QTree_Int_rbuf,MemOut_QTree_Int) */
  MemOut_QTree_Int_t memOut_QTree_Int_buf;
  assign memOut_QTree_Int_r = (! memOut_QTree_Int_buf[0]);
  assign memOut_QTree_Int_rbuf_d = (memOut_QTree_Int_buf[0] ? memOut_QTree_Int_buf :
                                    memOut_QTree_Int_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memOut_QTree_Int_buf <= {67'd0, 1'd0};
    else
      if ((memOut_QTree_Int_rbuf_r && memOut_QTree_Int_buf[0]))
        memOut_QTree_Int_buf <= {67'd0, 1'd0};
      else if (((! memOut_QTree_Int_rbuf_r) && (! memOut_QTree_Int_buf[0])))
        memOut_QTree_Int_buf <= memOut_QTree_Int_d;
  
  /* mergectrl (Ty C4,
           Ty Pointer_QTree_Int) : [(m1a8C_1_argbuf,Pointer_QTree_Int),
                                    (m2a8D_1_argbuf,Pointer_QTree_Int),
                                    (q4a8u_1_argbuf,Pointer_QTree_Int),
                                    (wsiX_1_1_argbuf,Pointer_QTree_Int)] > (readMerge_choice_QTree_Int,C4) (readMerge_data_QTree_Int,Pointer_QTree_Int) */
  logic [3:0] m1a8C_1_argbuf_select_d;
  assign m1a8C_1_argbuf_select_d = ((| m1a8C_1_argbuf_select_q) ? m1a8C_1_argbuf_select_q :
                                    (m1a8C_1_argbuf_d[0] ? 4'd1 :
                                     (m2a8D_1_argbuf_d[0] ? 4'd2 :
                                      (q4a8u_1_argbuf_d[0] ? 4'd4 :
                                       (wsiX_1_1_argbuf_d[0] ? 4'd8 :
                                        4'd0)))));
  logic [3:0] m1a8C_1_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m1a8C_1_argbuf_select_q <= 4'd0;
    else
      m1a8C_1_argbuf_select_q <= (m1a8C_1_argbuf_done ? 4'd0 :
                                  m1a8C_1_argbuf_select_d);
  logic [1:0] m1a8C_1_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m1a8C_1_argbuf_emit_q <= 2'd0;
    else
      m1a8C_1_argbuf_emit_q <= (m1a8C_1_argbuf_done ? 2'd0 :
                                m1a8C_1_argbuf_emit_d);
  logic [1:0] m1a8C_1_argbuf_emit_d;
  assign m1a8C_1_argbuf_emit_d = (m1a8C_1_argbuf_emit_q | ({readMerge_choice_QTree_Int_d[0],
                                                            readMerge_data_QTree_Int_d[0]} & {readMerge_choice_QTree_Int_r,
                                                                                              readMerge_data_QTree_Int_r}));
  logic m1a8C_1_argbuf_done;
  assign m1a8C_1_argbuf_done = (& m1a8C_1_argbuf_emit_d);
  assign {wsiX_1_1_argbuf_r,
          q4a8u_1_argbuf_r,
          m2a8D_1_argbuf_r,
          m1a8C_1_argbuf_r} = (m1a8C_1_argbuf_done ? m1a8C_1_argbuf_select_d :
                               4'd0);
  assign readMerge_data_QTree_Int_d = ((m1a8C_1_argbuf_select_d[0] && (! m1a8C_1_argbuf_emit_q[0])) ? m1a8C_1_argbuf_d :
                                       ((m1a8C_1_argbuf_select_d[1] && (! m1a8C_1_argbuf_emit_q[0])) ? m2a8D_1_argbuf_d :
                                        ((m1a8C_1_argbuf_select_d[2] && (! m1a8C_1_argbuf_emit_q[0])) ? q4a8u_1_argbuf_d :
                                         ((m1a8C_1_argbuf_select_d[3] && (! m1a8C_1_argbuf_emit_q[0])) ? wsiX_1_1_argbuf_d :
                                          {16'd0, 1'd0}))));
  assign readMerge_choice_QTree_Int_d = ((m1a8C_1_argbuf_select_d[0] && (! m1a8C_1_argbuf_emit_q[1])) ? C1_4_dc(1'd1) :
                                         ((m1a8C_1_argbuf_select_d[1] && (! m1a8C_1_argbuf_emit_q[1])) ? C2_4_dc(1'd1) :
                                          ((m1a8C_1_argbuf_select_d[2] && (! m1a8C_1_argbuf_emit_q[1])) ? C3_4_dc(1'd1) :
                                           ((m1a8C_1_argbuf_select_d[3] && (! m1a8C_1_argbuf_emit_q[1])) ? C4_4_dc(1'd1) :
                                            {2'd0, 1'd0}))));
  
  /* demux (Ty C4,
       Ty QTree_Int) : (readMerge_choice_QTree_Int,C4) (destructReadOut_QTree_Int,QTree_Int) > [(readPointer_QTree_Intm1a8C_1_argbuf,QTree_Int),
                                                                                                (readPointer_QTree_Intm2a8D_1_argbuf,QTree_Int),
                                                                                                (readPointer_QTree_Intq4a8u_1_argbuf,QTree_Int),
                                                                                                (readPointer_QTree_IntwsiX_1_1_argbuf,QTree_Int)] */
  logic [3:0] destructReadOut_QTree_Int_onehotd;
  always_comb
    if ((readMerge_choice_QTree_Int_d[0] && destructReadOut_QTree_Int_d[0]))
      unique case (readMerge_choice_QTree_Int_d[2:1])
        2'd0: destructReadOut_QTree_Int_onehotd = 4'd1;
        2'd1: destructReadOut_QTree_Int_onehotd = 4'd2;
        2'd2: destructReadOut_QTree_Int_onehotd = 4'd4;
        2'd3: destructReadOut_QTree_Int_onehotd = 4'd8;
        default: destructReadOut_QTree_Int_onehotd = 4'd0;
      endcase
    else destructReadOut_QTree_Int_onehotd = 4'd0;
  assign readPointer_QTree_Intm1a8C_1_argbuf_d = {destructReadOut_QTree_Int_d[66:1],
                                                  destructReadOut_QTree_Int_onehotd[0]};
  assign readPointer_QTree_Intm2a8D_1_argbuf_d = {destructReadOut_QTree_Int_d[66:1],
                                                  destructReadOut_QTree_Int_onehotd[1]};
  assign readPointer_QTree_Intq4a8u_1_argbuf_d = {destructReadOut_QTree_Int_d[66:1],
                                                  destructReadOut_QTree_Int_onehotd[2]};
  assign readPointer_QTree_IntwsiX_1_1_argbuf_d = {destructReadOut_QTree_Int_d[66:1],
                                                   destructReadOut_QTree_Int_onehotd[3]};
  assign destructReadOut_QTree_Int_r = (| (destructReadOut_QTree_Int_onehotd & {readPointer_QTree_IntwsiX_1_1_argbuf_r,
                                                                                readPointer_QTree_Intq4a8u_1_argbuf_r,
                                                                                readPointer_QTree_Intm2a8D_1_argbuf_r,
                                                                                readPointer_QTree_Intm1a8C_1_argbuf_r}));
  assign readMerge_choice_QTree_Int_r = destructReadOut_QTree_Int_r;
  
  /* destruct (Ty Pointer_QTree_Int,
          Dcon Pointer_QTree_Int) : (readMerge_data_QTree_Int,Pointer_QTree_Int) > [(destructReadIn_QTree_Int,Word16#)] */
  assign destructReadIn_QTree_Int_d = {readMerge_data_QTree_Int_d[16:1],
                                       readMerge_data_QTree_Int_d[0]};
  assign readMerge_data_QTree_Int_r = destructReadIn_QTree_Int_r;
  
  /* dcon (Ty MemIn_QTree_Int,
      Dcon ReadIn_QTree_Int) : [(destructReadIn_QTree_Int,Word16#)] > (dconReadIn_QTree_Int,MemIn_QTree_Int) */
  assign dconReadIn_QTree_Int_d = ReadIn_QTree_Int_dc((& {destructReadIn_QTree_Int_d[0]}), destructReadIn_QTree_Int_d);
  assign {destructReadIn_QTree_Int_r} = {1 {(dconReadIn_QTree_Int_r && dconReadIn_QTree_Int_d[0])}};
  
  /* destruct (Ty MemOut_QTree_Int,
          Dcon ReadOut_QTree_Int) : (memReadOut_QTree_Int,MemOut_QTree_Int) > [(destructReadOut_QTree_Int,QTree_Int)] */
  assign destructReadOut_QTree_Int_d = {memReadOut_QTree_Int_d[67:2],
                                        memReadOut_QTree_Int_d[0]};
  assign memReadOut_QTree_Int_r = destructReadOut_QTree_Int_r;
  
  /* mergectrl (Ty C23,
           Ty QTree_Int) : [(lizzieLet11_1_argbuf,QTree_Int),
                            (lizzieLet14_1_argbuf,QTree_Int),
                            (lizzieLet15_1_argbuf,QTree_Int),
                            (lizzieLet16_1_argbuf,QTree_Int),
                            (lizzieLet17_1_argbuf,QTree_Int),
                            (lizzieLet18_1_argbuf,QTree_Int),
                            (lizzieLet20_1_argbuf,QTree_Int),
                            (lizzieLet21_1_argbuf,QTree_Int),
                            (lizzieLet22_1_argbuf,QTree_Int),
                            (lizzieLet23_2_1_argbuf,QTree_Int),
                            (lizzieLet24_1_1_argbuf,QTree_Int),
                            (lizzieLet25_1_1_argbuf,QTree_Int),
                            (lizzieLet26_1_argbuf,QTree_Int),
                            (lizzieLet28_1_argbuf,QTree_Int),
                            (lizzieLet29_1_argbuf,QTree_Int),
                            (lizzieLet31_1_argbuf,QTree_Int),
                            (lizzieLet32_1_argbuf,QTree_Int),
                            (lizzieLet43_1_argbuf,QTree_Int),
                            (lizzieLet48_1_argbuf,QTree_Int),
                            (lizzieLet7_1_argbuf,QTree_Int),
                            (lizzieLet8_1_argbuf,QTree_Int),
                            (lizzieLet9_1_argbuf,QTree_Int),
                            (dummy_write_QTree_Int,QTree_Int)] > (writeMerge_choice_QTree_Int,C23) (writeMerge_data_QTree_Int,QTree_Int) */
  logic [22:0] lizzieLet11_1_argbuf_select_d;
  assign lizzieLet11_1_argbuf_select_d = ((| lizzieLet11_1_argbuf_select_q) ? lizzieLet11_1_argbuf_select_q :
                                          (lizzieLet11_1_argbuf_d[0] ? 23'd1 :
                                           (lizzieLet14_1_argbuf_d[0] ? 23'd2 :
                                            (lizzieLet15_1_argbuf_d[0] ? 23'd4 :
                                             (lizzieLet16_1_argbuf_d[0] ? 23'd8 :
                                              (lizzieLet17_1_argbuf_d[0] ? 23'd16 :
                                               (lizzieLet18_1_argbuf_d[0] ? 23'd32 :
                                                (lizzieLet20_1_argbuf_d[0] ? 23'd64 :
                                                 (lizzieLet21_1_argbuf_d[0] ? 23'd128 :
                                                  (lizzieLet22_1_argbuf_d[0] ? 23'd256 :
                                                   (lizzieLet23_2_1_argbuf_d[0] ? 23'd512 :
                                                    (lizzieLet24_1_1_argbuf_d[0] ? 23'd1024 :
                                                     (lizzieLet25_1_1_argbuf_d[0] ? 23'd2048 :
                                                      (lizzieLet26_1_argbuf_d[0] ? 23'd4096 :
                                                       (lizzieLet28_1_argbuf_d[0] ? 23'd8192 :
                                                        (lizzieLet29_1_argbuf_d[0] ? 23'd16384 :
                                                         (lizzieLet31_1_argbuf_d[0] ? 23'd32768 :
                                                          (lizzieLet32_1_argbuf_d[0] ? 23'd65536 :
                                                           (lizzieLet43_1_argbuf_d[0] ? 23'd131072 :
                                                            (lizzieLet48_1_argbuf_d[0] ? 23'd262144 :
                                                             (lizzieLet7_1_argbuf_d[0] ? 23'd524288 :
                                                              (lizzieLet8_1_argbuf_d[0] ? 23'd1048576 :
                                                               (lizzieLet9_1_argbuf_d[0] ? 23'd2097152 :
                                                                (dummy_write_QTree_Int_d[0] ? 23'd4194304 :
                                                                 23'd0))))))))))))))))))))))));
  logic [22:0] lizzieLet11_1_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet11_1_argbuf_select_q <= 23'd0;
    else
      lizzieLet11_1_argbuf_select_q <= (lizzieLet11_1_argbuf_done ? 23'd0 :
                                        lizzieLet11_1_argbuf_select_d);
  logic [1:0] lizzieLet11_1_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet11_1_argbuf_emit_q <= 2'd0;
    else
      lizzieLet11_1_argbuf_emit_q <= (lizzieLet11_1_argbuf_done ? 2'd0 :
                                      lizzieLet11_1_argbuf_emit_d);
  logic [1:0] lizzieLet11_1_argbuf_emit_d;
  assign lizzieLet11_1_argbuf_emit_d = (lizzieLet11_1_argbuf_emit_q | ({writeMerge_choice_QTree_Int_d[0],
                                                                        writeMerge_data_QTree_Int_d[0]} & {writeMerge_choice_QTree_Int_r,
                                                                                                           writeMerge_data_QTree_Int_r}));
  logic lizzieLet11_1_argbuf_done;
  assign lizzieLet11_1_argbuf_done = (& lizzieLet11_1_argbuf_emit_d);
  assign {dummy_write_QTree_Int_r,
          lizzieLet9_1_argbuf_r,
          lizzieLet8_1_argbuf_r,
          lizzieLet7_1_argbuf_r,
          lizzieLet48_1_argbuf_r,
          lizzieLet43_1_argbuf_r,
          lizzieLet32_1_argbuf_r,
          lizzieLet31_1_argbuf_r,
          lizzieLet29_1_argbuf_r,
          lizzieLet28_1_argbuf_r,
          lizzieLet26_1_argbuf_r,
          lizzieLet25_1_1_argbuf_r,
          lizzieLet24_1_1_argbuf_r,
          lizzieLet23_2_1_argbuf_r,
          lizzieLet22_1_argbuf_r,
          lizzieLet21_1_argbuf_r,
          lizzieLet20_1_argbuf_r,
          lizzieLet18_1_argbuf_r,
          lizzieLet17_1_argbuf_r,
          lizzieLet16_1_argbuf_r,
          lizzieLet15_1_argbuf_r,
          lizzieLet14_1_argbuf_r,
          lizzieLet11_1_argbuf_r} = (lizzieLet11_1_argbuf_done ? lizzieLet11_1_argbuf_select_d :
                                     23'd0);
  assign writeMerge_data_QTree_Int_d = ((lizzieLet11_1_argbuf_select_d[0] && (! lizzieLet11_1_argbuf_emit_q[0])) ? lizzieLet11_1_argbuf_d :
                                        ((lizzieLet11_1_argbuf_select_d[1] && (! lizzieLet11_1_argbuf_emit_q[0])) ? lizzieLet14_1_argbuf_d :
                                         ((lizzieLet11_1_argbuf_select_d[2] && (! lizzieLet11_1_argbuf_emit_q[0])) ? lizzieLet15_1_argbuf_d :
                                          ((lizzieLet11_1_argbuf_select_d[3] && (! lizzieLet11_1_argbuf_emit_q[0])) ? lizzieLet16_1_argbuf_d :
                                           ((lizzieLet11_1_argbuf_select_d[4] && (! lizzieLet11_1_argbuf_emit_q[0])) ? lizzieLet17_1_argbuf_d :
                                            ((lizzieLet11_1_argbuf_select_d[5] && (! lizzieLet11_1_argbuf_emit_q[0])) ? lizzieLet18_1_argbuf_d :
                                             ((lizzieLet11_1_argbuf_select_d[6] && (! lizzieLet11_1_argbuf_emit_q[0])) ? lizzieLet20_1_argbuf_d :
                                              ((lizzieLet11_1_argbuf_select_d[7] && (! lizzieLet11_1_argbuf_emit_q[0])) ? lizzieLet21_1_argbuf_d :
                                               ((lizzieLet11_1_argbuf_select_d[8] && (! lizzieLet11_1_argbuf_emit_q[0])) ? lizzieLet22_1_argbuf_d :
                                                ((lizzieLet11_1_argbuf_select_d[9] && (! lizzieLet11_1_argbuf_emit_q[0])) ? lizzieLet23_2_1_argbuf_d :
                                                 ((lizzieLet11_1_argbuf_select_d[10] && (! lizzieLet11_1_argbuf_emit_q[0])) ? lizzieLet24_1_1_argbuf_d :
                                                  ((lizzieLet11_1_argbuf_select_d[11] && (! lizzieLet11_1_argbuf_emit_q[0])) ? lizzieLet25_1_1_argbuf_d :
                                                   ((lizzieLet11_1_argbuf_select_d[12] && (! lizzieLet11_1_argbuf_emit_q[0])) ? lizzieLet26_1_argbuf_d :
                                                    ((lizzieLet11_1_argbuf_select_d[13] && (! lizzieLet11_1_argbuf_emit_q[0])) ? lizzieLet28_1_argbuf_d :
                                                     ((lizzieLet11_1_argbuf_select_d[14] && (! lizzieLet11_1_argbuf_emit_q[0])) ? lizzieLet29_1_argbuf_d :
                                                      ((lizzieLet11_1_argbuf_select_d[15] && (! lizzieLet11_1_argbuf_emit_q[0])) ? lizzieLet31_1_argbuf_d :
                                                       ((lizzieLet11_1_argbuf_select_d[16] && (! lizzieLet11_1_argbuf_emit_q[0])) ? lizzieLet32_1_argbuf_d :
                                                        ((lizzieLet11_1_argbuf_select_d[17] && (! lizzieLet11_1_argbuf_emit_q[0])) ? lizzieLet43_1_argbuf_d :
                                                         ((lizzieLet11_1_argbuf_select_d[18] && (! lizzieLet11_1_argbuf_emit_q[0])) ? lizzieLet48_1_argbuf_d :
                                                          ((lizzieLet11_1_argbuf_select_d[19] && (! lizzieLet11_1_argbuf_emit_q[0])) ? lizzieLet7_1_argbuf_d :
                                                           ((lizzieLet11_1_argbuf_select_d[20] && (! lizzieLet11_1_argbuf_emit_q[0])) ? lizzieLet8_1_argbuf_d :
                                                            ((lizzieLet11_1_argbuf_select_d[21] && (! lizzieLet11_1_argbuf_emit_q[0])) ? lizzieLet9_1_argbuf_d :
                                                             ((lizzieLet11_1_argbuf_select_d[22] && (! lizzieLet11_1_argbuf_emit_q[0])) ? dummy_write_QTree_Int_d :
                                                              {66'd0, 1'd0})))))))))))))))))))))));
  assign writeMerge_choice_QTree_Int_d = ((lizzieLet11_1_argbuf_select_d[0] && (! lizzieLet11_1_argbuf_emit_q[1])) ? C1_23_dc(1'd1) :
                                          ((lizzieLet11_1_argbuf_select_d[1] && (! lizzieLet11_1_argbuf_emit_q[1])) ? C2_23_dc(1'd1) :
                                           ((lizzieLet11_1_argbuf_select_d[2] && (! lizzieLet11_1_argbuf_emit_q[1])) ? C3_23_dc(1'd1) :
                                            ((lizzieLet11_1_argbuf_select_d[3] && (! lizzieLet11_1_argbuf_emit_q[1])) ? C4_23_dc(1'd1) :
                                             ((lizzieLet11_1_argbuf_select_d[4] && (! lizzieLet11_1_argbuf_emit_q[1])) ? C5_23_dc(1'd1) :
                                              ((lizzieLet11_1_argbuf_select_d[5] && (! lizzieLet11_1_argbuf_emit_q[1])) ? C6_23_dc(1'd1) :
                                               ((lizzieLet11_1_argbuf_select_d[6] && (! lizzieLet11_1_argbuf_emit_q[1])) ? C7_23_dc(1'd1) :
                                                ((lizzieLet11_1_argbuf_select_d[7] && (! lizzieLet11_1_argbuf_emit_q[1])) ? C8_23_dc(1'd1) :
                                                 ((lizzieLet11_1_argbuf_select_d[8] && (! lizzieLet11_1_argbuf_emit_q[1])) ? C9_23_dc(1'd1) :
                                                  ((lizzieLet11_1_argbuf_select_d[9] && (! lizzieLet11_1_argbuf_emit_q[1])) ? C10_23_dc(1'd1) :
                                                   ((lizzieLet11_1_argbuf_select_d[10] && (! lizzieLet11_1_argbuf_emit_q[1])) ? C11_23_dc(1'd1) :
                                                    ((lizzieLet11_1_argbuf_select_d[11] && (! lizzieLet11_1_argbuf_emit_q[1])) ? C12_23_dc(1'd1) :
                                                     ((lizzieLet11_1_argbuf_select_d[12] && (! lizzieLet11_1_argbuf_emit_q[1])) ? C13_23_dc(1'd1) :
                                                      ((lizzieLet11_1_argbuf_select_d[13] && (! lizzieLet11_1_argbuf_emit_q[1])) ? C14_23_dc(1'd1) :
                                                       ((lizzieLet11_1_argbuf_select_d[14] && (! lizzieLet11_1_argbuf_emit_q[1])) ? C15_23_dc(1'd1) :
                                                        ((lizzieLet11_1_argbuf_select_d[15] && (! lizzieLet11_1_argbuf_emit_q[1])) ? C16_23_dc(1'd1) :
                                                         ((lizzieLet11_1_argbuf_select_d[16] && (! lizzieLet11_1_argbuf_emit_q[1])) ? C17_23_dc(1'd1) :
                                                          ((lizzieLet11_1_argbuf_select_d[17] && (! lizzieLet11_1_argbuf_emit_q[1])) ? C18_23_dc(1'd1) :
                                                           ((lizzieLet11_1_argbuf_select_d[18] && (! lizzieLet11_1_argbuf_emit_q[1])) ? C19_23_dc(1'd1) :
                                                            ((lizzieLet11_1_argbuf_select_d[19] && (! lizzieLet11_1_argbuf_emit_q[1])) ? C20_23_dc(1'd1) :
                                                             ((lizzieLet11_1_argbuf_select_d[20] && (! lizzieLet11_1_argbuf_emit_q[1])) ? C21_23_dc(1'd1) :
                                                              ((lizzieLet11_1_argbuf_select_d[21] && (! lizzieLet11_1_argbuf_emit_q[1])) ? C22_23_dc(1'd1) :
                                                               ((lizzieLet11_1_argbuf_select_d[22] && (! lizzieLet11_1_argbuf_emit_q[1])) ? C23_23_dc(1'd1) :
                                                                {5'd0, 1'd0})))))))))))))))))))))));
  
  /* demux (Ty C23,
       Ty Pointer_QTree_Int) : (writeMerge_choice_QTree_Int,C23) (demuxWriteResult_QTree_Int,Pointer_QTree_Int) > [(writeQTree_IntlizzieLet11_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet14_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet15_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet16_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet17_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet18_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet20_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet21_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet22_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet23_2_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet24_1_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet25_1_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet26_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet28_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet29_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet31_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet32_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet43_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet48_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet7_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet8_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet9_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (dummy_write_QTree_Int_sink,Pointer_QTree_Int)] */
  logic [22:0] demuxWriteResult_QTree_Int_onehotd;
  always_comb
    if ((writeMerge_choice_QTree_Int_d[0] && demuxWriteResult_QTree_Int_d[0]))
      unique case (writeMerge_choice_QTree_Int_d[5:1])
        5'd0: demuxWriteResult_QTree_Int_onehotd = 23'd1;
        5'd1: demuxWriteResult_QTree_Int_onehotd = 23'd2;
        5'd2: demuxWriteResult_QTree_Int_onehotd = 23'd4;
        5'd3: demuxWriteResult_QTree_Int_onehotd = 23'd8;
        5'd4: demuxWriteResult_QTree_Int_onehotd = 23'd16;
        5'd5: demuxWriteResult_QTree_Int_onehotd = 23'd32;
        5'd6: demuxWriteResult_QTree_Int_onehotd = 23'd64;
        5'd7: demuxWriteResult_QTree_Int_onehotd = 23'd128;
        5'd8: demuxWriteResult_QTree_Int_onehotd = 23'd256;
        5'd9: demuxWriteResult_QTree_Int_onehotd = 23'd512;
        5'd10: demuxWriteResult_QTree_Int_onehotd = 23'd1024;
        5'd11: demuxWriteResult_QTree_Int_onehotd = 23'd2048;
        5'd12: demuxWriteResult_QTree_Int_onehotd = 23'd4096;
        5'd13: demuxWriteResult_QTree_Int_onehotd = 23'd8192;
        5'd14: demuxWriteResult_QTree_Int_onehotd = 23'd16384;
        5'd15: demuxWriteResult_QTree_Int_onehotd = 23'd32768;
        5'd16: demuxWriteResult_QTree_Int_onehotd = 23'd65536;
        5'd17: demuxWriteResult_QTree_Int_onehotd = 23'd131072;
        5'd18: demuxWriteResult_QTree_Int_onehotd = 23'd262144;
        5'd19: demuxWriteResult_QTree_Int_onehotd = 23'd524288;
        5'd20: demuxWriteResult_QTree_Int_onehotd = 23'd1048576;
        5'd21: demuxWriteResult_QTree_Int_onehotd = 23'd2097152;
        5'd22: demuxWriteResult_QTree_Int_onehotd = 23'd4194304;
        default: demuxWriteResult_QTree_Int_onehotd = 23'd0;
      endcase
    else demuxWriteResult_QTree_Int_onehotd = 23'd0;
  assign writeQTree_IntlizzieLet11_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                 demuxWriteResult_QTree_Int_onehotd[0]};
  assign writeQTree_IntlizzieLet14_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                 demuxWriteResult_QTree_Int_onehotd[1]};
  assign writeQTree_IntlizzieLet15_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                 demuxWriteResult_QTree_Int_onehotd[2]};
  assign writeQTree_IntlizzieLet16_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                 demuxWriteResult_QTree_Int_onehotd[3]};
  assign writeQTree_IntlizzieLet17_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                 demuxWriteResult_QTree_Int_onehotd[4]};
  assign writeQTree_IntlizzieLet18_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                 demuxWriteResult_QTree_Int_onehotd[5]};
  assign writeQTree_IntlizzieLet20_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                 demuxWriteResult_QTree_Int_onehotd[6]};
  assign writeQTree_IntlizzieLet21_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                 demuxWriteResult_QTree_Int_onehotd[7]};
  assign writeQTree_IntlizzieLet22_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                 demuxWriteResult_QTree_Int_onehotd[8]};
  assign writeQTree_IntlizzieLet23_2_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                   demuxWriteResult_QTree_Int_onehotd[9]};
  assign writeQTree_IntlizzieLet24_1_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                   demuxWriteResult_QTree_Int_onehotd[10]};
  assign writeQTree_IntlizzieLet25_1_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                   demuxWriteResult_QTree_Int_onehotd[11]};
  assign writeQTree_IntlizzieLet26_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                 demuxWriteResult_QTree_Int_onehotd[12]};
  assign writeQTree_IntlizzieLet28_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                 demuxWriteResult_QTree_Int_onehotd[13]};
  assign writeQTree_IntlizzieLet29_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                 demuxWriteResult_QTree_Int_onehotd[14]};
  assign writeQTree_IntlizzieLet31_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                 demuxWriteResult_QTree_Int_onehotd[15]};
  assign writeQTree_IntlizzieLet32_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                 demuxWriteResult_QTree_Int_onehotd[16]};
  assign writeQTree_IntlizzieLet43_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                 demuxWriteResult_QTree_Int_onehotd[17]};
  assign writeQTree_IntlizzieLet48_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                 demuxWriteResult_QTree_Int_onehotd[18]};
  assign writeQTree_IntlizzieLet7_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                demuxWriteResult_QTree_Int_onehotd[19]};
  assign writeQTree_IntlizzieLet8_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                demuxWriteResult_QTree_Int_onehotd[20]};
  assign writeQTree_IntlizzieLet9_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                demuxWriteResult_QTree_Int_onehotd[21]};
  assign dummy_write_QTree_Int_sink_d = {demuxWriteResult_QTree_Int_d[16:1],
                                         demuxWriteResult_QTree_Int_onehotd[22]};
  assign demuxWriteResult_QTree_Int_r = (| (demuxWriteResult_QTree_Int_onehotd & {dummy_write_QTree_Int_sink_r,
                                                                                  writeQTree_IntlizzieLet9_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet8_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet7_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet48_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet43_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet32_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet31_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet29_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet28_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet26_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet25_1_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet24_1_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet23_2_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet22_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet21_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet20_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet18_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet17_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet16_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet15_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet14_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet11_1_argbuf_r}));
  assign writeMerge_choice_QTree_Int_r = demuxWriteResult_QTree_Int_r;
  
  /* dcon (Ty MemIn_QTree_Int,
      Dcon WriteIn_QTree_Int) : [(forkHP1_QTree_In3,Word16#),
                                 (writeMerge_data_QTree_Int,QTree_Int)] > (dconWriteIn_QTree_Int,MemIn_QTree_Int) */
  assign dconWriteIn_QTree_Int_d = WriteIn_QTree_Int_dc((& {forkHP1_QTree_In3_d[0],
                                                            writeMerge_data_QTree_Int_d[0]}), forkHP1_QTree_In3_d, writeMerge_data_QTree_Int_d);
  assign {forkHP1_QTree_In3_r,
          writeMerge_data_QTree_Int_r} = {2 {(dconWriteIn_QTree_Int_r && dconWriteIn_QTree_Int_d[0])}};
  
  /* dcon (Ty Pointer_QTree_Int,
      Dcon Pointer_QTree_Int) : [(forkHP1_QTree_In4,Word16#)] > (dconPtr_QTree_Int,Pointer_QTree_Int) */
  assign dconPtr_QTree_Int_d = Pointer_QTree_Int_dc((& {forkHP1_QTree_In4_d[0]}), forkHP1_QTree_In4_d);
  assign {forkHP1_QTree_In4_r} = {1 {(dconPtr_QTree_Int_r && dconPtr_QTree_Int_d[0])}};
  
  /* demux (Ty MemOut_QTree_Int,
       Ty Pointer_QTree_Int) : (memWriteOut_QTree_Int,MemOut_QTree_Int) (dconPtr_QTree_Int,Pointer_QTree_Int) > [(_82,Pointer_QTree_Int),
                                                                                                                 (demuxWriteResult_QTree_Int,Pointer_QTree_Int)] */
  logic [1:0] dconPtr_QTree_Int_onehotd;
  always_comb
    if ((memWriteOut_QTree_Int_d[0] && dconPtr_QTree_Int_d[0]))
      unique case (memWriteOut_QTree_Int_d[1:1])
        1'd0: dconPtr_QTree_Int_onehotd = 2'd1;
        1'd1: dconPtr_QTree_Int_onehotd = 2'd2;
        default: dconPtr_QTree_Int_onehotd = 2'd0;
      endcase
    else dconPtr_QTree_Int_onehotd = 2'd0;
  assign _82_d = {dconPtr_QTree_Int_d[16:1],
                  dconPtr_QTree_Int_onehotd[0]};
  assign demuxWriteResult_QTree_Int_d = {dconPtr_QTree_Int_d[16:1],
                                         dconPtr_QTree_Int_onehotd[1]};
  assign dconPtr_QTree_Int_r = (| (dconPtr_QTree_Int_onehotd & {demuxWriteResult_QTree_Int_r,
                                                                _82_r}));
  assign memWriteOut_QTree_Int_r = dconPtr_QTree_Int_r;
  
  /* const (Ty Word16#,
       Lit 0) : (go__11,Go) > (initHP_CTf_f_Int_Int,Word16#) */
  assign initHP_CTf_f_Int_Int_d = {16'd0, go__11_d[0]};
  assign go__11_r = initHP_CTf_f_Int_Int_r;
  
  /* const (Ty Word16#,
       Lit 1) : (incrHP_CTf_f_Int_Int1,Go) > (incrHP_CTf_f_Int_Int,Word16#) */
  assign incrHP_CTf_f_Int_Int_d = {16'd1,
                                   incrHP_CTf_f_Int_Int1_d[0]};
  assign incrHP_CTf_f_Int_Int1_r = incrHP_CTf_f_Int_Int_r;
  
  /* merge (Ty Go) : [(go__12,Go),
                 (incrHP_CTf_f_Int_Int2,Go)] > (incrHP_mergeCTf_f_Int_Int,Go) */
  logic [1:0] incrHP_mergeCTf_f_Int_Int_selected;
  logic [1:0] incrHP_mergeCTf_f_Int_Int_select;
  always_comb
    begin
      incrHP_mergeCTf_f_Int_Int_selected = 2'd0;
      if ((| incrHP_mergeCTf_f_Int_Int_select))
        incrHP_mergeCTf_f_Int_Int_selected = incrHP_mergeCTf_f_Int_Int_select;
      else
        if (go__12_d[0]) incrHP_mergeCTf_f_Int_Int_selected[0] = 1'd1;
        else if (incrHP_CTf_f_Int_Int2_d[0])
          incrHP_mergeCTf_f_Int_Int_selected[1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeCTf_f_Int_Int_select <= 2'd0;
    else
      incrHP_mergeCTf_f_Int_Int_select <= (incrHP_mergeCTf_f_Int_Int_r ? 2'd0 :
                                           incrHP_mergeCTf_f_Int_Int_selected);
  always_comb
    if (incrHP_mergeCTf_f_Int_Int_selected[0])
      incrHP_mergeCTf_f_Int_Int_d = go__12_d;
    else if (incrHP_mergeCTf_f_Int_Int_selected[1])
      incrHP_mergeCTf_f_Int_Int_d = incrHP_CTf_f_Int_Int2_d;
    else incrHP_mergeCTf_f_Int_Int_d = 1'd0;
  assign {incrHP_CTf_f_Int_Int2_r,
          go__12_r} = (incrHP_mergeCTf_f_Int_Int_r ? incrHP_mergeCTf_f_Int_Int_selected :
                       2'd0);
  
  /* fork (Ty Go) : (incrHP_mergeCTf_f_Int_Int_buf,Go) > [(incrHP_CTf_f_Int_Int1,Go),
                                                     (incrHP_CTf_f_Int_Int2,Go)] */
  logic [1:0] incrHP_mergeCTf_f_Int_Int_buf_emitted;
  logic [1:0] incrHP_mergeCTf_f_Int_Int_buf_done;
  assign incrHP_CTf_f_Int_Int1_d = (incrHP_mergeCTf_f_Int_Int_buf_d[0] && (! incrHP_mergeCTf_f_Int_Int_buf_emitted[0]));
  assign incrHP_CTf_f_Int_Int2_d = (incrHP_mergeCTf_f_Int_Int_buf_d[0] && (! incrHP_mergeCTf_f_Int_Int_buf_emitted[1]));
  assign incrHP_mergeCTf_f_Int_Int_buf_done = (incrHP_mergeCTf_f_Int_Int_buf_emitted | ({incrHP_CTf_f_Int_Int2_d[0],
                                                                                         incrHP_CTf_f_Int_Int1_d[0]} & {incrHP_CTf_f_Int_Int2_r,
                                                                                                                        incrHP_CTf_f_Int_Int1_r}));
  assign incrHP_mergeCTf_f_Int_Int_buf_r = (& incrHP_mergeCTf_f_Int_Int_buf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeCTf_f_Int_Int_buf_emitted <= 2'd0;
    else
      incrHP_mergeCTf_f_Int_Int_buf_emitted <= (incrHP_mergeCTf_f_Int_Int_buf_r ? 2'd0 :
                                                incrHP_mergeCTf_f_Int_Int_buf_done);
  
  /* op_add (Ty Word16#) : (incrHP_CTf_f_Int_Int,Word16#) (forkHP1_CTf_f_Int_Int,Word16#) > (addHP_CTf_f_Int_Int,Word16#) */
  assign addHP_CTf_f_Int_Int_d = {(incrHP_CTf_f_Int_Int_d[16:1] + forkHP1_CTf_f_Int_Int_d[16:1]),
                                  (incrHP_CTf_f_Int_Int_d[0] && forkHP1_CTf_f_Int_Int_d[0])};
  assign {incrHP_CTf_f_Int_Int_r,
          forkHP1_CTf_f_Int_Int_r} = {2 {(addHP_CTf_f_Int_Int_r && addHP_CTf_f_Int_Int_d[0])}};
  
  /* merge (Ty Word16#) : [(initHP_CTf_f_Int_Int,Word16#),
                      (addHP_CTf_f_Int_Int,Word16#)] > (mergeHP_CTf_f_Int_Int,Word16#) */
  logic [1:0] mergeHP_CTf_f_Int_Int_selected;
  logic [1:0] mergeHP_CTf_f_Int_Int_select;
  always_comb
    begin
      mergeHP_CTf_f_Int_Int_selected = 2'd0;
      if ((| mergeHP_CTf_f_Int_Int_select))
        mergeHP_CTf_f_Int_Int_selected = mergeHP_CTf_f_Int_Int_select;
      else
        if (initHP_CTf_f_Int_Int_d[0])
          mergeHP_CTf_f_Int_Int_selected[0] = 1'd1;
        else if (addHP_CTf_f_Int_Int_d[0])
          mergeHP_CTf_f_Int_Int_selected[1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_CTf_f_Int_Int_select <= 2'd0;
    else
      mergeHP_CTf_f_Int_Int_select <= (mergeHP_CTf_f_Int_Int_r ? 2'd0 :
                                       mergeHP_CTf_f_Int_Int_selected);
  always_comb
    if (mergeHP_CTf_f_Int_Int_selected[0])
      mergeHP_CTf_f_Int_Int_d = initHP_CTf_f_Int_Int_d;
    else if (mergeHP_CTf_f_Int_Int_selected[1])
      mergeHP_CTf_f_Int_Int_d = addHP_CTf_f_Int_Int_d;
    else mergeHP_CTf_f_Int_Int_d = {16'd0, 1'd0};
  assign {addHP_CTf_f_Int_Int_r,
          initHP_CTf_f_Int_Int_r} = (mergeHP_CTf_f_Int_Int_r ? mergeHP_CTf_f_Int_Int_selected :
                                     2'd0);
  
  /* buf (Ty Go) : (incrHP_mergeCTf_f_Int_Int,Go) > (incrHP_mergeCTf_f_Int_Int_buf,Go) */
  Go_t incrHP_mergeCTf_f_Int_Int_bufchan_d;
  logic incrHP_mergeCTf_f_Int_Int_bufchan_r;
  assign incrHP_mergeCTf_f_Int_Int_r = ((! incrHP_mergeCTf_f_Int_Int_bufchan_d[0]) || incrHP_mergeCTf_f_Int_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeCTf_f_Int_Int_bufchan_d <= 1'd0;
    else
      if (incrHP_mergeCTf_f_Int_Int_r)
        incrHP_mergeCTf_f_Int_Int_bufchan_d <= incrHP_mergeCTf_f_Int_Int_d;
  Go_t incrHP_mergeCTf_f_Int_Int_bufchan_buf;
  assign incrHP_mergeCTf_f_Int_Int_bufchan_r = (! incrHP_mergeCTf_f_Int_Int_bufchan_buf[0]);
  assign incrHP_mergeCTf_f_Int_Int_buf_d = (incrHP_mergeCTf_f_Int_Int_bufchan_buf[0] ? incrHP_mergeCTf_f_Int_Int_bufchan_buf :
                                            incrHP_mergeCTf_f_Int_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeCTf_f_Int_Int_bufchan_buf <= 1'd0;
    else
      if ((incrHP_mergeCTf_f_Int_Int_buf_r && incrHP_mergeCTf_f_Int_Int_bufchan_buf[0]))
        incrHP_mergeCTf_f_Int_Int_bufchan_buf <= 1'd0;
      else if (((! incrHP_mergeCTf_f_Int_Int_buf_r) && (! incrHP_mergeCTf_f_Int_Int_bufchan_buf[0])))
        incrHP_mergeCTf_f_Int_Int_bufchan_buf <= incrHP_mergeCTf_f_Int_Int_bufchan_d;
  
  /* buf (Ty Word16#) : (mergeHP_CTf_f_Int_Int,Word16#) > (mergeHP_CTf_f_Int_Int_buf,Word16#) */
  \Word16#_t  mergeHP_CTf_f_Int_Int_bufchan_d;
  logic mergeHP_CTf_f_Int_Int_bufchan_r;
  assign mergeHP_CTf_f_Int_Int_r = ((! mergeHP_CTf_f_Int_Int_bufchan_d[0]) || mergeHP_CTf_f_Int_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      mergeHP_CTf_f_Int_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (mergeHP_CTf_f_Int_Int_r)
        mergeHP_CTf_f_Int_Int_bufchan_d <= mergeHP_CTf_f_Int_Int_d;
  \Word16#_t  mergeHP_CTf_f_Int_Int_bufchan_buf;
  assign mergeHP_CTf_f_Int_Int_bufchan_r = (! mergeHP_CTf_f_Int_Int_bufchan_buf[0]);
  assign mergeHP_CTf_f_Int_Int_buf_d = (mergeHP_CTf_f_Int_Int_bufchan_buf[0] ? mergeHP_CTf_f_Int_Int_bufchan_buf :
                                        mergeHP_CTf_f_Int_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      mergeHP_CTf_f_Int_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((mergeHP_CTf_f_Int_Int_buf_r && mergeHP_CTf_f_Int_Int_bufchan_buf[0]))
        mergeHP_CTf_f_Int_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! mergeHP_CTf_f_Int_Int_buf_r) && (! mergeHP_CTf_f_Int_Int_bufchan_buf[0])))
        mergeHP_CTf_f_Int_Int_bufchan_buf <= mergeHP_CTf_f_Int_Int_bufchan_d;
  
  /* fork (Ty Word16#) : (mergeHP_CTf_f_Int_Int_buf,Word16#) > [(forkHP1_CTf_f_Int_Int,Word16#),
                                                           (forkHP1_CTf_f_Int_In2,Word16#),
                                                           (forkHP1_CTf_f_Int_In3,Word16#)] */
  logic [2:0] mergeHP_CTf_f_Int_Int_buf_emitted;
  logic [2:0] mergeHP_CTf_f_Int_Int_buf_done;
  assign forkHP1_CTf_f_Int_Int_d = {mergeHP_CTf_f_Int_Int_buf_d[16:1],
                                    (mergeHP_CTf_f_Int_Int_buf_d[0] && (! mergeHP_CTf_f_Int_Int_buf_emitted[0]))};
  assign forkHP1_CTf_f_Int_In2_d = {mergeHP_CTf_f_Int_Int_buf_d[16:1],
                                    (mergeHP_CTf_f_Int_Int_buf_d[0] && (! mergeHP_CTf_f_Int_Int_buf_emitted[1]))};
  assign forkHP1_CTf_f_Int_In3_d = {mergeHP_CTf_f_Int_Int_buf_d[16:1],
                                    (mergeHP_CTf_f_Int_Int_buf_d[0] && (! mergeHP_CTf_f_Int_Int_buf_emitted[2]))};
  assign mergeHP_CTf_f_Int_Int_buf_done = (mergeHP_CTf_f_Int_Int_buf_emitted | ({forkHP1_CTf_f_Int_In3_d[0],
                                                                                 forkHP1_CTf_f_Int_In2_d[0],
                                                                                 forkHP1_CTf_f_Int_Int_d[0]} & {forkHP1_CTf_f_Int_In3_r,
                                                                                                                forkHP1_CTf_f_Int_In2_r,
                                                                                                                forkHP1_CTf_f_Int_Int_r}));
  assign mergeHP_CTf_f_Int_Int_buf_r = (& mergeHP_CTf_f_Int_Int_buf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_CTf_f_Int_Int_buf_emitted <= 3'd0;
    else
      mergeHP_CTf_f_Int_Int_buf_emitted <= (mergeHP_CTf_f_Int_Int_buf_r ? 3'd0 :
                                            mergeHP_CTf_f_Int_Int_buf_done);
  
  /* mergectrl (Ty C2,
           Ty MemIn_CTf_f_Int_Int) : [(dconReadIn_CTf_f_Int_Int,MemIn_CTf_f_Int_Int),
                                      (dconWriteIn_CTf_f_Int_Int,MemIn_CTf_f_Int_Int)] > (memMergeChoice_CTf_f_Int_Int,C2) (memMergeIn_CTf_f_Int_Int,MemIn_CTf_f_Int_Int) */
  logic [1:0] dconReadIn_CTf_f_Int_Int_select_d;
  assign dconReadIn_CTf_f_Int_Int_select_d = ((| dconReadIn_CTf_f_Int_Int_select_q) ? dconReadIn_CTf_f_Int_Int_select_q :
                                              (dconReadIn_CTf_f_Int_Int_d[0] ? 2'd1 :
                                               (dconWriteIn_CTf_f_Int_Int_d[0] ? 2'd2 :
                                                2'd0)));
  logic [1:0] dconReadIn_CTf_f_Int_Int_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) dconReadIn_CTf_f_Int_Int_select_q <= 2'd0;
    else
      dconReadIn_CTf_f_Int_Int_select_q <= (dconReadIn_CTf_f_Int_Int_done ? 2'd0 :
                                            dconReadIn_CTf_f_Int_Int_select_d);
  logic [1:0] dconReadIn_CTf_f_Int_Int_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) dconReadIn_CTf_f_Int_Int_emit_q <= 2'd0;
    else
      dconReadIn_CTf_f_Int_Int_emit_q <= (dconReadIn_CTf_f_Int_Int_done ? 2'd0 :
                                          dconReadIn_CTf_f_Int_Int_emit_d);
  logic [1:0] dconReadIn_CTf_f_Int_Int_emit_d;
  assign dconReadIn_CTf_f_Int_Int_emit_d = (dconReadIn_CTf_f_Int_Int_emit_q | ({memMergeChoice_CTf_f_Int_Int_d[0],
                                                                                memMergeIn_CTf_f_Int_Int_d[0]} & {memMergeChoice_CTf_f_Int_Int_r,
                                                                                                                  memMergeIn_CTf_f_Int_Int_r}));
  logic dconReadIn_CTf_f_Int_Int_done;
  assign dconReadIn_CTf_f_Int_Int_done = (& dconReadIn_CTf_f_Int_Int_emit_d);
  assign {dconWriteIn_CTf_f_Int_Int_r,
          dconReadIn_CTf_f_Int_Int_r} = (dconReadIn_CTf_f_Int_Int_done ? dconReadIn_CTf_f_Int_Int_select_d :
                                         2'd0);
  assign memMergeIn_CTf_f_Int_Int_d = ((dconReadIn_CTf_f_Int_Int_select_d[0] && (! dconReadIn_CTf_f_Int_Int_emit_q[0])) ? dconReadIn_CTf_f_Int_Int_d :
                                       ((dconReadIn_CTf_f_Int_Int_select_d[1] && (! dconReadIn_CTf_f_Int_Int_emit_q[0])) ? dconWriteIn_CTf_f_Int_Int_d :
                                        {132'd0, 1'd0}));
  assign memMergeChoice_CTf_f_Int_Int_d = ((dconReadIn_CTf_f_Int_Int_select_d[0] && (! dconReadIn_CTf_f_Int_Int_emit_q[1])) ? C1_2_dc(1'd1) :
                                           ((dconReadIn_CTf_f_Int_Int_select_d[1] && (! dconReadIn_CTf_f_Int_Int_emit_q[1])) ? C2_2_dc(1'd1) :
                                            {1'd0, 1'd0}));
  
  /* bram (Ty MemIn_CTf_f_Int_Int,
      Ty MemOut_CTf_f_Int_Int) : (memMergeIn_CTf_f_Int_Int_dbuf,MemIn_CTf_f_Int_Int) > (memOut_CTf_f_Int_Int,MemOut_CTf_f_Int_Int) */
  logic [114:0] memMergeIn_CTf_f_Int_Int_dbuf_mem[65535:0];
  logic [15:0] memMergeIn_CTf_f_Int_Int_dbuf_address;
  logic [114:0] memMergeIn_CTf_f_Int_Int_dbuf_din;
  logic [114:0] memOut_CTf_f_Int_Int_q;
  logic memOut_CTf_f_Int_Int_valid;
  logic memMergeIn_CTf_f_Int_Int_dbuf_we;
  logic memOut_CTf_f_Int_Int_we;
  assign memMergeIn_CTf_f_Int_Int_dbuf_din = memMergeIn_CTf_f_Int_Int_dbuf_d[132:18];
  assign memMergeIn_CTf_f_Int_Int_dbuf_address = memMergeIn_CTf_f_Int_Int_dbuf_d[17:2];
  assign memMergeIn_CTf_f_Int_Int_dbuf_we = (memMergeIn_CTf_f_Int_Int_dbuf_d[1:1] && memMergeIn_CTf_f_Int_Int_dbuf_d[0]);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        memOut_CTf_f_Int_Int_we <= 1'd0;
        memOut_CTf_f_Int_Int_valid <= 1'd0;
      end
    else
      begin
        memOut_CTf_f_Int_Int_we <= memMergeIn_CTf_f_Int_Int_dbuf_we;
        memOut_CTf_f_Int_Int_valid <= memMergeIn_CTf_f_Int_Int_dbuf_d[0];
        if (memMergeIn_CTf_f_Int_Int_dbuf_we)
          begin
            memMergeIn_CTf_f_Int_Int_dbuf_mem[memMergeIn_CTf_f_Int_Int_dbuf_address] <= memMergeIn_CTf_f_Int_Int_dbuf_din;
            memOut_CTf_f_Int_Int_q <= memMergeIn_CTf_f_Int_Int_dbuf_din;
          end
        else
          memOut_CTf_f_Int_Int_q <= memMergeIn_CTf_f_Int_Int_dbuf_mem[memMergeIn_CTf_f_Int_Int_dbuf_address];
      end
  assign memOut_CTf_f_Int_Int_d = {memOut_CTf_f_Int_Int_q,
                                   memOut_CTf_f_Int_Int_we,
                                   memOut_CTf_f_Int_Int_valid};
  assign memMergeIn_CTf_f_Int_Int_dbuf_r = ((! memOut_CTf_f_Int_Int_valid) || memOut_CTf_f_Int_Int_r);
  logic [31:0] profiling_MemIn_CTf_f_Int_Int_read;
  logic [31:0] profiling_MemIn_CTf_f_Int_Int_write;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        profiling_MemIn_CTf_f_Int_Int_write <= 0;
        profiling_MemIn_CTf_f_Int_Int_read <= 0;
      end
    else
      if ((memMergeIn_CTf_f_Int_Int_dbuf_we == 1'd1))
        profiling_MemIn_CTf_f_Int_Int_write <= (profiling_MemIn_CTf_f_Int_Int_write + 1);
      else
        if ((memOut_CTf_f_Int_Int_valid == 1'd1))
          profiling_MemIn_CTf_f_Int_Int_read <= (profiling_MemIn_CTf_f_Int_Int_read + 1);
  
  /* demux (Ty C2,
       Ty MemOut_CTf_f_Int_Int) : (memMergeChoice_CTf_f_Int_Int,C2) (memOut_CTf_f_Int_Int_dbuf,MemOut_CTf_f_Int_Int) > [(memReadOut_CTf_f_Int_Int,MemOut_CTf_f_Int_Int),
                                                                                                                        (memWriteOut_CTf_f_Int_Int,MemOut_CTf_f_Int_Int)] */
  logic [1:0] memOut_CTf_f_Int_Int_dbuf_onehotd;
  always_comb
    if ((memMergeChoice_CTf_f_Int_Int_d[0] && memOut_CTf_f_Int_Int_dbuf_d[0]))
      unique case (memMergeChoice_CTf_f_Int_Int_d[1:1])
        1'd0: memOut_CTf_f_Int_Int_dbuf_onehotd = 2'd1;
        1'd1: memOut_CTf_f_Int_Int_dbuf_onehotd = 2'd2;
        default: memOut_CTf_f_Int_Int_dbuf_onehotd = 2'd0;
      endcase
    else memOut_CTf_f_Int_Int_dbuf_onehotd = 2'd0;
  assign memReadOut_CTf_f_Int_Int_d = {memOut_CTf_f_Int_Int_dbuf_d[116:1],
                                       memOut_CTf_f_Int_Int_dbuf_onehotd[0]};
  assign memWriteOut_CTf_f_Int_Int_d = {memOut_CTf_f_Int_Int_dbuf_d[116:1],
                                        memOut_CTf_f_Int_Int_dbuf_onehotd[1]};
  assign memOut_CTf_f_Int_Int_dbuf_r = (| (memOut_CTf_f_Int_Int_dbuf_onehotd & {memWriteOut_CTf_f_Int_Int_r,
                                                                                memReadOut_CTf_f_Int_Int_r}));
  assign memMergeChoice_CTf_f_Int_Int_r = memOut_CTf_f_Int_Int_dbuf_r;
  
  /* dbuf (Ty MemIn_CTf_f_Int_Int) : (memMergeIn_CTf_f_Int_Int_rbuf,MemIn_CTf_f_Int_Int) > (memMergeIn_CTf_f_Int_Int_dbuf,MemIn_CTf_f_Int_Int) */
  assign memMergeIn_CTf_f_Int_Int_rbuf_r = ((! memMergeIn_CTf_f_Int_Int_dbuf_d[0]) || memMergeIn_CTf_f_Int_Int_dbuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      memMergeIn_CTf_f_Int_Int_dbuf_d <= {132'd0, 1'd0};
    else
      if (memMergeIn_CTf_f_Int_Int_rbuf_r)
        memMergeIn_CTf_f_Int_Int_dbuf_d <= memMergeIn_CTf_f_Int_Int_rbuf_d;
  
  /* rbuf (Ty MemIn_CTf_f_Int_Int) : (memMergeIn_CTf_f_Int_Int,MemIn_CTf_f_Int_Int) > (memMergeIn_CTf_f_Int_Int_rbuf,MemIn_CTf_f_Int_Int) */
  MemIn_CTf_f_Int_Int_t memMergeIn_CTf_f_Int_Int_buf;
  assign memMergeIn_CTf_f_Int_Int_r = (! memMergeIn_CTf_f_Int_Int_buf[0]);
  assign memMergeIn_CTf_f_Int_Int_rbuf_d = (memMergeIn_CTf_f_Int_Int_buf[0] ? memMergeIn_CTf_f_Int_Int_buf :
                                            memMergeIn_CTf_f_Int_Int_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      memMergeIn_CTf_f_Int_Int_buf <= {132'd0, 1'd0};
    else
      if ((memMergeIn_CTf_f_Int_Int_rbuf_r && memMergeIn_CTf_f_Int_Int_buf[0]))
        memMergeIn_CTf_f_Int_Int_buf <= {132'd0, 1'd0};
      else if (((! memMergeIn_CTf_f_Int_Int_rbuf_r) && (! memMergeIn_CTf_f_Int_Int_buf[0])))
        memMergeIn_CTf_f_Int_Int_buf <= memMergeIn_CTf_f_Int_Int_d;
  
  /* dbuf (Ty MemOut_CTf_f_Int_Int) : (memOut_CTf_f_Int_Int_rbuf,MemOut_CTf_f_Int_Int) > (memOut_CTf_f_Int_Int_dbuf,MemOut_CTf_f_Int_Int) */
  assign memOut_CTf_f_Int_Int_rbuf_r = ((! memOut_CTf_f_Int_Int_dbuf_d[0]) || memOut_CTf_f_Int_Int_dbuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memOut_CTf_f_Int_Int_dbuf_d <= {116'd0, 1'd0};
    else
      if (memOut_CTf_f_Int_Int_rbuf_r)
        memOut_CTf_f_Int_Int_dbuf_d <= memOut_CTf_f_Int_Int_rbuf_d;
  
  /* rbuf (Ty MemOut_CTf_f_Int_Int) : (memOut_CTf_f_Int_Int,MemOut_CTf_f_Int_Int) > (memOut_CTf_f_Int_Int_rbuf,MemOut_CTf_f_Int_Int) */
  MemOut_CTf_f_Int_Int_t memOut_CTf_f_Int_Int_buf;
  assign memOut_CTf_f_Int_Int_r = (! memOut_CTf_f_Int_Int_buf[0]);
  assign memOut_CTf_f_Int_Int_rbuf_d = (memOut_CTf_f_Int_Int_buf[0] ? memOut_CTf_f_Int_Int_buf :
                                        memOut_CTf_f_Int_Int_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memOut_CTf_f_Int_Int_buf <= {116'd0, 1'd0};
    else
      if ((memOut_CTf_f_Int_Int_rbuf_r && memOut_CTf_f_Int_Int_buf[0]))
        memOut_CTf_f_Int_Int_buf <= {116'd0, 1'd0};
      else if (((! memOut_CTf_f_Int_Int_rbuf_r) && (! memOut_CTf_f_Int_Int_buf[0])))
        memOut_CTf_f_Int_Int_buf <= memOut_CTf_f_Int_Int_d;
  
  /* destruct (Ty Pointer_CTf_f_Int_Int,
          Dcon Pointer_CTf_f_Int_Int) : (scfarg_0_2_1_argbuf,Pointer_CTf_f_Int_Int) > [(destructReadIn_CTf_f_Int_Int,Word16#)] */
  assign destructReadIn_CTf_f_Int_Int_d = {scfarg_0_2_1_argbuf_d[16:1],
                                           scfarg_0_2_1_argbuf_d[0]};
  assign scfarg_0_2_1_argbuf_r = destructReadIn_CTf_f_Int_Int_r;
  
  /* dcon (Ty MemIn_CTf_f_Int_Int,
      Dcon ReadIn_CTf_f_Int_Int) : [(destructReadIn_CTf_f_Int_Int,Word16#)] > (dconReadIn_CTf_f_Int_Int,MemIn_CTf_f_Int_Int) */
  assign dconReadIn_CTf_f_Int_Int_d = ReadIn_CTf_f_Int_Int_dc((& {destructReadIn_CTf_f_Int_Int_d[0]}), destructReadIn_CTf_f_Int_Int_d);
  assign {destructReadIn_CTf_f_Int_Int_r} = {1 {(dconReadIn_CTf_f_Int_Int_r && dconReadIn_CTf_f_Int_Int_d[0])}};
  
  /* destruct (Ty MemOut_CTf_f_Int_Int,
          Dcon ReadOut_CTf_f_Int_Int) : (memReadOut_CTf_f_Int_Int,MemOut_CTf_f_Int_Int) > [(readPointer_CTf_f_Int_Intscfarg_0_2_1_argbuf,CTf_f_Int_Int)] */
  assign readPointer_CTf_f_Int_Intscfarg_0_2_1_argbuf_d = {memReadOut_CTf_f_Int_Int_d[116:2],
                                                           memReadOut_CTf_f_Int_Int_d[0]};
  assign memReadOut_CTf_f_Int_Int_r = readPointer_CTf_f_Int_Intscfarg_0_2_1_argbuf_r;
  
  /* mergectrl (Ty C5,
           Ty CTf_f_Int_Int) : [(lizzieLet30_1_argbuf,CTf_f_Int_Int),
                                (lizzieLet34_1_argbuf,CTf_f_Int_Int),
                                (lizzieLet45_1_argbuf,CTf_f_Int_Int),
                                (lizzieLet46_1_argbuf,CTf_f_Int_Int),
                                (lizzieLet47_1_argbuf,CTf_f_Int_Int)] > (writeMerge_choice_CTf_f_Int_Int,C5) (writeMerge_data_CTf_f_Int_Int,CTf_f_Int_Int) */
  logic [4:0] lizzieLet30_1_argbuf_select_d;
  assign lizzieLet30_1_argbuf_select_d = ((| lizzieLet30_1_argbuf_select_q) ? lizzieLet30_1_argbuf_select_q :
                                          (lizzieLet30_1_argbuf_d[0] ? 5'd1 :
                                           (lizzieLet34_1_argbuf_d[0] ? 5'd2 :
                                            (lizzieLet45_1_argbuf_d[0] ? 5'd4 :
                                             (lizzieLet46_1_argbuf_d[0] ? 5'd8 :
                                              (lizzieLet47_1_argbuf_d[0] ? 5'd16 :
                                               5'd0))))));
  logic [4:0] lizzieLet30_1_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet30_1_argbuf_select_q <= 5'd0;
    else
      lizzieLet30_1_argbuf_select_q <= (lizzieLet30_1_argbuf_done ? 5'd0 :
                                        lizzieLet30_1_argbuf_select_d);
  logic [1:0] lizzieLet30_1_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet30_1_argbuf_emit_q <= 2'd0;
    else
      lizzieLet30_1_argbuf_emit_q <= (lizzieLet30_1_argbuf_done ? 2'd0 :
                                      lizzieLet30_1_argbuf_emit_d);
  logic [1:0] lizzieLet30_1_argbuf_emit_d;
  assign lizzieLet30_1_argbuf_emit_d = (lizzieLet30_1_argbuf_emit_q | ({writeMerge_choice_CTf_f_Int_Int_d[0],
                                                                        writeMerge_data_CTf_f_Int_Int_d[0]} & {writeMerge_choice_CTf_f_Int_Int_r,
                                                                                                               writeMerge_data_CTf_f_Int_Int_r}));
  logic lizzieLet30_1_argbuf_done;
  assign lizzieLet30_1_argbuf_done = (& lizzieLet30_1_argbuf_emit_d);
  assign {lizzieLet47_1_argbuf_r,
          lizzieLet46_1_argbuf_r,
          lizzieLet45_1_argbuf_r,
          lizzieLet34_1_argbuf_r,
          lizzieLet30_1_argbuf_r} = (lizzieLet30_1_argbuf_done ? lizzieLet30_1_argbuf_select_d :
                                     5'd0);
  assign writeMerge_data_CTf_f_Int_Int_d = ((lizzieLet30_1_argbuf_select_d[0] && (! lizzieLet30_1_argbuf_emit_q[0])) ? lizzieLet30_1_argbuf_d :
                                            ((lizzieLet30_1_argbuf_select_d[1] && (! lizzieLet30_1_argbuf_emit_q[0])) ? lizzieLet34_1_argbuf_d :
                                             ((lizzieLet30_1_argbuf_select_d[2] && (! lizzieLet30_1_argbuf_emit_q[0])) ? lizzieLet45_1_argbuf_d :
                                              ((lizzieLet30_1_argbuf_select_d[3] && (! lizzieLet30_1_argbuf_emit_q[0])) ? lizzieLet46_1_argbuf_d :
                                               ((lizzieLet30_1_argbuf_select_d[4] && (! lizzieLet30_1_argbuf_emit_q[0])) ? lizzieLet47_1_argbuf_d :
                                                {115'd0, 1'd0})))));
  assign writeMerge_choice_CTf_f_Int_Int_d = ((lizzieLet30_1_argbuf_select_d[0] && (! lizzieLet30_1_argbuf_emit_q[1])) ? C1_5_dc(1'd1) :
                                              ((lizzieLet30_1_argbuf_select_d[1] && (! lizzieLet30_1_argbuf_emit_q[1])) ? C2_5_dc(1'd1) :
                                               ((lizzieLet30_1_argbuf_select_d[2] && (! lizzieLet30_1_argbuf_emit_q[1])) ? C3_5_dc(1'd1) :
                                                ((lizzieLet30_1_argbuf_select_d[3] && (! lizzieLet30_1_argbuf_emit_q[1])) ? C4_5_dc(1'd1) :
                                                 ((lizzieLet30_1_argbuf_select_d[4] && (! lizzieLet30_1_argbuf_emit_q[1])) ? C5_5_dc(1'd1) :
                                                  {3'd0, 1'd0})))));
  
  /* demux (Ty C5,
       Ty Pointer_CTf_f_Int_Int) : (writeMerge_choice_CTf_f_Int_Int,C5) (demuxWriteResult_CTf_f_Int_Int,Pointer_CTf_f_Int_Int) > [(writeCTf_f_Int_IntlizzieLet30_1_argbuf,Pointer_CTf_f_Int_Int),
                                                                                                                                  (writeCTf_f_Int_IntlizzieLet34_1_argbuf,Pointer_CTf_f_Int_Int),
                                                                                                                                  (writeCTf_f_Int_IntlizzieLet45_1_argbuf,Pointer_CTf_f_Int_Int),
                                                                                                                                  (writeCTf_f_Int_IntlizzieLet46_1_argbuf,Pointer_CTf_f_Int_Int),
                                                                                                                                  (writeCTf_f_Int_IntlizzieLet47_1_argbuf,Pointer_CTf_f_Int_Int)] */
  logic [4:0] demuxWriteResult_CTf_f_Int_Int_onehotd;
  always_comb
    if ((writeMerge_choice_CTf_f_Int_Int_d[0] && demuxWriteResult_CTf_f_Int_Int_d[0]))
      unique case (writeMerge_choice_CTf_f_Int_Int_d[3:1])
        3'd0: demuxWriteResult_CTf_f_Int_Int_onehotd = 5'd1;
        3'd1: demuxWriteResult_CTf_f_Int_Int_onehotd = 5'd2;
        3'd2: demuxWriteResult_CTf_f_Int_Int_onehotd = 5'd4;
        3'd3: demuxWriteResult_CTf_f_Int_Int_onehotd = 5'd8;
        3'd4: demuxWriteResult_CTf_f_Int_Int_onehotd = 5'd16;
        default: demuxWriteResult_CTf_f_Int_Int_onehotd = 5'd0;
      endcase
    else demuxWriteResult_CTf_f_Int_Int_onehotd = 5'd0;
  assign writeCTf_f_Int_IntlizzieLet30_1_argbuf_d = {demuxWriteResult_CTf_f_Int_Int_d[16:1],
                                                     demuxWriteResult_CTf_f_Int_Int_onehotd[0]};
  assign writeCTf_f_Int_IntlizzieLet34_1_argbuf_d = {demuxWriteResult_CTf_f_Int_Int_d[16:1],
                                                     demuxWriteResult_CTf_f_Int_Int_onehotd[1]};
  assign writeCTf_f_Int_IntlizzieLet45_1_argbuf_d = {demuxWriteResult_CTf_f_Int_Int_d[16:1],
                                                     demuxWriteResult_CTf_f_Int_Int_onehotd[2]};
  assign writeCTf_f_Int_IntlizzieLet46_1_argbuf_d = {demuxWriteResult_CTf_f_Int_Int_d[16:1],
                                                     demuxWriteResult_CTf_f_Int_Int_onehotd[3]};
  assign writeCTf_f_Int_IntlizzieLet47_1_argbuf_d = {demuxWriteResult_CTf_f_Int_Int_d[16:1],
                                                     demuxWriteResult_CTf_f_Int_Int_onehotd[4]};
  assign demuxWriteResult_CTf_f_Int_Int_r = (| (demuxWriteResult_CTf_f_Int_Int_onehotd & {writeCTf_f_Int_IntlizzieLet47_1_argbuf_r,
                                                                                          writeCTf_f_Int_IntlizzieLet46_1_argbuf_r,
                                                                                          writeCTf_f_Int_IntlizzieLet45_1_argbuf_r,
                                                                                          writeCTf_f_Int_IntlizzieLet34_1_argbuf_r,
                                                                                          writeCTf_f_Int_IntlizzieLet30_1_argbuf_r}));
  assign writeMerge_choice_CTf_f_Int_Int_r = demuxWriteResult_CTf_f_Int_Int_r;
  
  /* dcon (Ty MemIn_CTf_f_Int_Int,
      Dcon WriteIn_CTf_f_Int_Int) : [(forkHP1_CTf_f_Int_In2,Word16#),
                                     (writeMerge_data_CTf_f_Int_Int,CTf_f_Int_Int)] > (dconWriteIn_CTf_f_Int_Int,MemIn_CTf_f_Int_Int) */
  assign dconWriteIn_CTf_f_Int_Int_d = WriteIn_CTf_f_Int_Int_dc((& {forkHP1_CTf_f_Int_In2_d[0],
                                                                    writeMerge_data_CTf_f_Int_Int_d[0]}), forkHP1_CTf_f_Int_In2_d, writeMerge_data_CTf_f_Int_Int_d);
  assign {forkHP1_CTf_f_Int_In2_r,
          writeMerge_data_CTf_f_Int_Int_r} = {2 {(dconWriteIn_CTf_f_Int_Int_r && dconWriteIn_CTf_f_Int_Int_d[0])}};
  
  /* dcon (Ty Pointer_CTf_f_Int_Int,
      Dcon Pointer_CTf_f_Int_Int) : [(forkHP1_CTf_f_Int_In3,Word16#)] > (dconPtr_CTf_f_Int_Int,Pointer_CTf_f_Int_Int) */
  assign dconPtr_CTf_f_Int_Int_d = Pointer_CTf_f_Int_Int_dc((& {forkHP1_CTf_f_Int_In3_d[0]}), forkHP1_CTf_f_Int_In3_d);
  assign {forkHP1_CTf_f_Int_In3_r} = {1 {(dconPtr_CTf_f_Int_Int_r && dconPtr_CTf_f_Int_Int_d[0])}};
  
  /* demux (Ty MemOut_CTf_f_Int_Int,
       Ty Pointer_CTf_f_Int_Int) : (memWriteOut_CTf_f_Int_Int,MemOut_CTf_f_Int_Int) (dconPtr_CTf_f_Int_Int,Pointer_CTf_f_Int_Int) > [(_81,Pointer_CTf_f_Int_Int),
                                                                                                                                     (demuxWriteResult_CTf_f_Int_Int,Pointer_CTf_f_Int_Int)] */
  logic [1:0] dconPtr_CTf_f_Int_Int_onehotd;
  always_comb
    if ((memWriteOut_CTf_f_Int_Int_d[0] && dconPtr_CTf_f_Int_Int_d[0]))
      unique case (memWriteOut_CTf_f_Int_Int_d[1:1])
        1'd0: dconPtr_CTf_f_Int_Int_onehotd = 2'd1;
        1'd1: dconPtr_CTf_f_Int_Int_onehotd = 2'd2;
        default: dconPtr_CTf_f_Int_Int_onehotd = 2'd0;
      endcase
    else dconPtr_CTf_f_Int_Int_onehotd = 2'd0;
  assign _81_d = {dconPtr_CTf_f_Int_Int_d[16:1],
                  dconPtr_CTf_f_Int_Int_onehotd[0]};
  assign demuxWriteResult_CTf_f_Int_Int_d = {dconPtr_CTf_f_Int_Int_d[16:1],
                                             dconPtr_CTf_f_Int_Int_onehotd[1]};
  assign dconPtr_CTf_f_Int_Int_r = (| (dconPtr_CTf_f_Int_Int_onehotd & {demuxWriteResult_CTf_f_Int_Int_r,
                                                                        _81_r}));
  assign memWriteOut_CTf_f_Int_Int_r = dconPtr_CTf_f_Int_Int_r;
  
  /* source (Ty Go) : > (sourceGo,Go) */
  
  /* source (Ty Pointer_QTree_Int) : > (m1aey_0,Pointer_QTree_Int) */
  
  /* source (Ty Pointer_QTree_Int) : > (m2aez_1,Pointer_QTree_Int) */
  
  /* destruct (Ty TupGo___Pointer_QTree_Int,
          Dcon TupGo___Pointer_QTree_Int) : ($wnnzTupGo___Pointer_QTree_Int_1,TupGo___Pointer_QTree_Int) > [($wnnzTupGo___Pointer_QTree_Intgo_7,Go),
                                                                                                            ($wnnzTupGo___Pointer_QTree_IntwsiX,Pointer_QTree_Int)] */
  logic [1:0] \$wnnzTupGo___Pointer_QTree_Int_1_emitted ;
  logic [1:0] \$wnnzTupGo___Pointer_QTree_Int_1_done ;
  assign \$wnnzTupGo___Pointer_QTree_Intgo_7_d  = (\$wnnzTupGo___Pointer_QTree_Int_1_d [0] && (! \$wnnzTupGo___Pointer_QTree_Int_1_emitted [0]));
  assign \$wnnzTupGo___Pointer_QTree_IntwsiX_d  = {\$wnnzTupGo___Pointer_QTree_Int_1_d [16:1],
                                                   (\$wnnzTupGo___Pointer_QTree_Int_1_d [0] && (! \$wnnzTupGo___Pointer_QTree_Int_1_emitted [1]))};
  assign \$wnnzTupGo___Pointer_QTree_Int_1_done  = (\$wnnzTupGo___Pointer_QTree_Int_1_emitted  | ({\$wnnzTupGo___Pointer_QTree_IntwsiX_d [0],
                                                                                                   \$wnnzTupGo___Pointer_QTree_Intgo_7_d [0]} & {\$wnnzTupGo___Pointer_QTree_IntwsiX_r ,
                                                                                                                                                 \$wnnzTupGo___Pointer_QTree_Intgo_7_r }));
  assign \$wnnzTupGo___Pointer_QTree_Int_1_r  = (& \$wnnzTupGo___Pointer_QTree_Int_1_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \$wnnzTupGo___Pointer_QTree_Int_1_emitted  <= 2'd0;
    else
      \$wnnzTupGo___Pointer_QTree_Int_1_emitted  <= (\$wnnzTupGo___Pointer_QTree_Int_1_r  ? 2'd0 :
                                                     \$wnnzTupGo___Pointer_QTree_Int_1_done );
  
  /* fork (Ty Go) : ($wnnzTupGo___Pointer_QTree_Intgo_7,Go) > [(go_7_1,Go),
                                                          (go_7_2,Go)] */
  logic [1:0] \$wnnzTupGo___Pointer_QTree_Intgo_7_emitted ;
  logic [1:0] \$wnnzTupGo___Pointer_QTree_Intgo_7_done ;
  assign go_7_1_d = (\$wnnzTupGo___Pointer_QTree_Intgo_7_d [0] && (! \$wnnzTupGo___Pointer_QTree_Intgo_7_emitted [0]));
  assign go_7_2_d = (\$wnnzTupGo___Pointer_QTree_Intgo_7_d [0] && (! \$wnnzTupGo___Pointer_QTree_Intgo_7_emitted [1]));
  assign \$wnnzTupGo___Pointer_QTree_Intgo_7_done  = (\$wnnzTupGo___Pointer_QTree_Intgo_7_emitted  | ({go_7_2_d[0],
                                                                                                       go_7_1_d[0]} & {go_7_2_r,
                                                                                                                       go_7_1_r}));
  assign \$wnnzTupGo___Pointer_QTree_Intgo_7_r  = (& \$wnnzTupGo___Pointer_QTree_Intgo_7_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \$wnnzTupGo___Pointer_QTree_Intgo_7_emitted  <= 2'd0;
    else
      \$wnnzTupGo___Pointer_QTree_Intgo_7_emitted  <= (\$wnnzTupGo___Pointer_QTree_Intgo_7_r  ? 2'd0 :
                                                       \$wnnzTupGo___Pointer_QTree_Intgo_7_done );
  
  /* buf (Ty Pointer_QTree_Int) : ($wnnzTupGo___Pointer_QTree_IntwsiX,Pointer_QTree_Int) > (wsiX_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t \$wnnzTupGo___Pointer_QTree_IntwsiX_bufchan_d ;
  logic \$wnnzTupGo___Pointer_QTree_IntwsiX_bufchan_r ;
  assign \$wnnzTupGo___Pointer_QTree_IntwsiX_r  = ((! \$wnnzTupGo___Pointer_QTree_IntwsiX_bufchan_d [0]) || \$wnnzTupGo___Pointer_QTree_IntwsiX_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \$wnnzTupGo___Pointer_QTree_IntwsiX_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\$wnnzTupGo___Pointer_QTree_IntwsiX_r )
        \$wnnzTupGo___Pointer_QTree_IntwsiX_bufchan_d  <= \$wnnzTupGo___Pointer_QTree_IntwsiX_d ;
  Pointer_QTree_Int_t \$wnnzTupGo___Pointer_QTree_IntwsiX_bufchan_buf ;
  assign \$wnnzTupGo___Pointer_QTree_IntwsiX_bufchan_r  = (! \$wnnzTupGo___Pointer_QTree_IntwsiX_bufchan_buf [0]);
  assign wsiX_1_argbuf_d = (\$wnnzTupGo___Pointer_QTree_IntwsiX_bufchan_buf [0] ? \$wnnzTupGo___Pointer_QTree_IntwsiX_bufchan_buf  :
                            \$wnnzTupGo___Pointer_QTree_IntwsiX_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \$wnnzTupGo___Pointer_QTree_IntwsiX_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((wsiX_1_argbuf_r && \$wnnzTupGo___Pointer_QTree_IntwsiX_bufchan_buf [0]))
        \$wnnzTupGo___Pointer_QTree_IntwsiX_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! wsiX_1_argbuf_r) && (! \$wnnzTupGo___Pointer_QTree_IntwsiX_bufchan_buf [0])))
        \$wnnzTupGo___Pointer_QTree_IntwsiX_bufchan_buf  <= \$wnnzTupGo___Pointer_QTree_IntwsiX_bufchan_d ;
  
  /* dcon (Ty Int,Dcon I#) : [($wnnz_resbuf,Int#)] > (es_7_1I#,Int) */
  assign \es_7_1I#_d  = \I#_dc ((& {\$wnnz_resbuf_d [0]}), \$wnnz_resbuf_d );
  assign {\$wnnz_resbuf_r } = {1 {(\es_7_1I#_r  && \es_7_1I#_d [0])}};
  
  /* mergectrl (Ty C5,
           Ty TupGo___MyDTInt_Bool___Int) : [(applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1,TupGo___MyDTInt_Bool___Int),
                                             (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int2,TupGo___MyDTInt_Bool___Int),
                                             (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int3,TupGo___MyDTInt_Bool___Int),
                                             (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int4,TupGo___MyDTInt_Bool___Int),
                                             (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int5,TupGo___MyDTInt_Bool___Int)] > (applyfnInt_Bool_5_choice,C5) (applyfnInt_Bool_5_data,TupGo___MyDTInt_Bool___Int) */
  logic [4:0] applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_select_d;
  assign applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_select_d = ((| applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_select_q) ? applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_select_q :
                                                                   (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_d[0] ? 5'd1 :
                                                                    (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int2_d[0] ? 5'd2 :
                                                                     (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int3_d[0] ? 5'd4 :
                                                                      (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int4_d[0] ? 5'd8 :
                                                                       (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int5_d[0] ? 5'd16 :
                                                                        5'd0))))));
  logic [4:0] applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_select_q <= 5'd0;
    else
      applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_select_q <= (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_done ? 5'd0 :
                                                                 applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_select_d);
  logic [1:0] applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_emit_q <= 2'd0;
    else
      applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_emit_q <= (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_done ? 2'd0 :
                                                               applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_emit_d);
  logic [1:0] applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_emit_d;
  assign applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_emit_d = (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_emit_q | ({applyfnInt_Bool_5_choice_d[0],
                                                                                                                          applyfnInt_Bool_5_data_d[0]} & {applyfnInt_Bool_5_choice_r,
                                                                                                                                                          applyfnInt_Bool_5_data_r}));
  logic applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_done;
  assign applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_done = (& applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_emit_d);
  assign {applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int5_r,
          applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int4_r,
          applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int3_r,
          applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int2_r,
          applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_r} = (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_done ? applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_select_d :
                                                              5'd0);
  assign applyfnInt_Bool_5_data_d = ((applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_select_d[0] && (! applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_emit_q[0])) ? applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_d :
                                     ((applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_select_d[1] && (! applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_emit_q[0])) ? applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int2_d :
                                      ((applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_select_d[2] && (! applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_emit_q[0])) ? applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int3_d :
                                       ((applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_select_d[3] && (! applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_emit_q[0])) ? applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int4_d :
                                        ((applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_select_d[4] && (! applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_emit_q[0])) ? applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int5_d :
                                         {32'd0, 1'd0})))));
  assign applyfnInt_Bool_5_choice_d = ((applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_select_d[0] && (! applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_emit_q[1])) ? C1_5_dc(1'd1) :
                                       ((applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_select_d[1] && (! applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_emit_q[1])) ? C2_5_dc(1'd1) :
                                        ((applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_select_d[2] && (! applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_emit_q[1])) ? C3_5_dc(1'd1) :
                                         ((applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_select_d[3] && (! applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_emit_q[1])) ? C4_5_dc(1'd1) :
                                          ((applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_select_d[4] && (! applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_emit_q[1])) ? C5_5_dc(1'd1) :
                                           {3'd0, 1'd0})))));
  
  /* fork (Ty MyDTInt_Bool) : (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0,MyDTInt_Bool) > [(arg0_1,MyDTInt_Bool),
                                                                                           (arg0_2,MyDTInt_Bool),
                                                                                           (arg0_3,MyDTInt_Bool)] */
  logic [2:0] applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_emitted;
  logic [2:0] applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_done;
  assign arg0_1_d = (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_d[0] && (! applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_emitted[0]));
  assign arg0_2_d = (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_d[0] && (! applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_emitted[1]));
  assign arg0_3_d = (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_d[0] && (! applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_emitted[2]));
  assign applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_done = (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_emitted | ({arg0_3_d[0],
                                                                                                                             arg0_2_d[0],
                                                                                                                             arg0_1_d[0]} & {arg0_3_r,
                                                                                                                                             arg0_2_r,
                                                                                                                                             arg0_1_r}));
  assign applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_r = (& applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_emitted <= 3'd0;
    else
      applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_emitted <= (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_r ? 3'd0 :
                                                                  applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_done);
  
  /* buf (Ty MyBool) : (applyfnInt_Bool_5_1,MyBool) > (applyfnInt_Bool_5_resbuf,MyBool) */
  MyBool_t applyfnInt_Bool_5_1_bufchan_d;
  logic applyfnInt_Bool_5_1_bufchan_r;
  assign applyfnInt_Bool_5_1_r = ((! applyfnInt_Bool_5_1_bufchan_d[0]) || applyfnInt_Bool_5_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) applyfnInt_Bool_5_1_bufchan_d <= {1'd0, 1'd0};
    else
      if (applyfnInt_Bool_5_1_r)
        applyfnInt_Bool_5_1_bufchan_d <= applyfnInt_Bool_5_1_d;
  MyBool_t applyfnInt_Bool_5_1_bufchan_buf;
  assign applyfnInt_Bool_5_1_bufchan_r = (! applyfnInt_Bool_5_1_bufchan_buf[0]);
  assign applyfnInt_Bool_5_resbuf_d = (applyfnInt_Bool_5_1_bufchan_buf[0] ? applyfnInt_Bool_5_1_bufchan_buf :
                                       applyfnInt_Bool_5_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Bool_5_1_bufchan_buf <= {1'd0, 1'd0};
    else
      if ((applyfnInt_Bool_5_resbuf_r && applyfnInt_Bool_5_1_bufchan_buf[0]))
        applyfnInt_Bool_5_1_bufchan_buf <= {1'd0, 1'd0};
      else if (((! applyfnInt_Bool_5_resbuf_r) && (! applyfnInt_Bool_5_1_bufchan_buf[0])))
        applyfnInt_Bool_5_1_bufchan_buf <= applyfnInt_Bool_5_1_bufchan_d;
  
  /* buf (Ty MyBool) : (applyfnInt_Bool_5_2,MyBool) > (applyfnInt_Bool_5_2_argbuf,MyBool) */
  MyBool_t applyfnInt_Bool_5_2_bufchan_d;
  logic applyfnInt_Bool_5_2_bufchan_r;
  assign applyfnInt_Bool_5_2_r = ((! applyfnInt_Bool_5_2_bufchan_d[0]) || applyfnInt_Bool_5_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) applyfnInt_Bool_5_2_bufchan_d <= {1'd0, 1'd0};
    else
      if (applyfnInt_Bool_5_2_r)
        applyfnInt_Bool_5_2_bufchan_d <= applyfnInt_Bool_5_2_d;
  MyBool_t applyfnInt_Bool_5_2_bufchan_buf;
  assign applyfnInt_Bool_5_2_bufchan_r = (! applyfnInt_Bool_5_2_bufchan_buf[0]);
  assign applyfnInt_Bool_5_2_argbuf_d = (applyfnInt_Bool_5_2_bufchan_buf[0] ? applyfnInt_Bool_5_2_bufchan_buf :
                                         applyfnInt_Bool_5_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Bool_5_2_bufchan_buf <= {1'd0, 1'd0};
    else
      if ((applyfnInt_Bool_5_2_argbuf_r && applyfnInt_Bool_5_2_bufchan_buf[0]))
        applyfnInt_Bool_5_2_bufchan_buf <= {1'd0, 1'd0};
      else if (((! applyfnInt_Bool_5_2_argbuf_r) && (! applyfnInt_Bool_5_2_bufchan_buf[0])))
        applyfnInt_Bool_5_2_bufchan_buf <= applyfnInt_Bool_5_2_bufchan_d;
  
  /* fork (Ty MyBool) : (applyfnInt_Bool_5_2_argbuf,MyBool) > [(es_2_1,MyBool),
                                                          (es_2_2,MyBool),
                                                          (es_2_3,MyBool),
                                                          (es_2_4,MyBool)] */
  logic [3:0] applyfnInt_Bool_5_2_argbuf_emitted;
  logic [3:0] applyfnInt_Bool_5_2_argbuf_done;
  assign es_2_1_d = {applyfnInt_Bool_5_2_argbuf_d[1:1],
                     (applyfnInt_Bool_5_2_argbuf_d[0] && (! applyfnInt_Bool_5_2_argbuf_emitted[0]))};
  assign es_2_2_d = {applyfnInt_Bool_5_2_argbuf_d[1:1],
                     (applyfnInt_Bool_5_2_argbuf_d[0] && (! applyfnInt_Bool_5_2_argbuf_emitted[1]))};
  assign es_2_3_d = {applyfnInt_Bool_5_2_argbuf_d[1:1],
                     (applyfnInt_Bool_5_2_argbuf_d[0] && (! applyfnInt_Bool_5_2_argbuf_emitted[2]))};
  assign es_2_4_d = {applyfnInt_Bool_5_2_argbuf_d[1:1],
                     (applyfnInt_Bool_5_2_argbuf_d[0] && (! applyfnInt_Bool_5_2_argbuf_emitted[3]))};
  assign applyfnInt_Bool_5_2_argbuf_done = (applyfnInt_Bool_5_2_argbuf_emitted | ({es_2_4_d[0],
                                                                                   es_2_3_d[0],
                                                                                   es_2_2_d[0],
                                                                                   es_2_1_d[0]} & {es_2_4_r,
                                                                                                   es_2_3_r,
                                                                                                   es_2_2_r,
                                                                                                   es_2_1_r}));
  assign applyfnInt_Bool_5_2_argbuf_r = (& applyfnInt_Bool_5_2_argbuf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) applyfnInt_Bool_5_2_argbuf_emitted <= 4'd0;
    else
      applyfnInt_Bool_5_2_argbuf_emitted <= (applyfnInt_Bool_5_2_argbuf_r ? 4'd0 :
                                             applyfnInt_Bool_5_2_argbuf_done);
  
  /* buf (Ty MyBool) : (applyfnInt_Bool_5_3,MyBool) > (applyfnInt_Bool_5_3_argbuf,MyBool) */
  MyBool_t applyfnInt_Bool_5_3_bufchan_d;
  logic applyfnInt_Bool_5_3_bufchan_r;
  assign applyfnInt_Bool_5_3_r = ((! applyfnInt_Bool_5_3_bufchan_d[0]) || applyfnInt_Bool_5_3_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) applyfnInt_Bool_5_3_bufchan_d <= {1'd0, 1'd0};
    else
      if (applyfnInt_Bool_5_3_r)
        applyfnInt_Bool_5_3_bufchan_d <= applyfnInt_Bool_5_3_d;
  MyBool_t applyfnInt_Bool_5_3_bufchan_buf;
  assign applyfnInt_Bool_5_3_bufchan_r = (! applyfnInt_Bool_5_3_bufchan_buf[0]);
  assign applyfnInt_Bool_5_3_argbuf_d = (applyfnInt_Bool_5_3_bufchan_buf[0] ? applyfnInt_Bool_5_3_bufchan_buf :
                                         applyfnInt_Bool_5_3_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Bool_5_3_bufchan_buf <= {1'd0, 1'd0};
    else
      if ((applyfnInt_Bool_5_3_argbuf_r && applyfnInt_Bool_5_3_bufchan_buf[0]))
        applyfnInt_Bool_5_3_bufchan_buf <= {1'd0, 1'd0};
      else if (((! applyfnInt_Bool_5_3_argbuf_r) && (! applyfnInt_Bool_5_3_bufchan_buf[0])))
        applyfnInt_Bool_5_3_bufchan_buf <= applyfnInt_Bool_5_3_bufchan_d;
  
  /* fork (Ty MyBool) : (applyfnInt_Bool_5_3_argbuf,MyBool) > [(es_10_1,MyBool),
                                                          (es_10_2,MyBool),
                                                          (es_10_3,MyBool),
                                                          (es_10_4,MyBool)] */
  logic [3:0] applyfnInt_Bool_5_3_argbuf_emitted;
  logic [3:0] applyfnInt_Bool_5_3_argbuf_done;
  assign es_10_1_d = {applyfnInt_Bool_5_3_argbuf_d[1:1],
                      (applyfnInt_Bool_5_3_argbuf_d[0] && (! applyfnInt_Bool_5_3_argbuf_emitted[0]))};
  assign es_10_2_d = {applyfnInt_Bool_5_3_argbuf_d[1:1],
                      (applyfnInt_Bool_5_3_argbuf_d[0] && (! applyfnInt_Bool_5_3_argbuf_emitted[1]))};
  assign es_10_3_d = {applyfnInt_Bool_5_3_argbuf_d[1:1],
                      (applyfnInt_Bool_5_3_argbuf_d[0] && (! applyfnInt_Bool_5_3_argbuf_emitted[2]))};
  assign es_10_4_d = {applyfnInt_Bool_5_3_argbuf_d[1:1],
                      (applyfnInt_Bool_5_3_argbuf_d[0] && (! applyfnInt_Bool_5_3_argbuf_emitted[3]))};
  assign applyfnInt_Bool_5_3_argbuf_done = (applyfnInt_Bool_5_3_argbuf_emitted | ({es_10_4_d[0],
                                                                                   es_10_3_d[0],
                                                                                   es_10_2_d[0],
                                                                                   es_10_1_d[0]} & {es_10_4_r,
                                                                                                    es_10_3_r,
                                                                                                    es_10_2_r,
                                                                                                    es_10_1_r}));
  assign applyfnInt_Bool_5_3_argbuf_r = (& applyfnInt_Bool_5_3_argbuf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) applyfnInt_Bool_5_3_argbuf_emitted <= 4'd0;
    else
      applyfnInt_Bool_5_3_argbuf_emitted <= (applyfnInt_Bool_5_3_argbuf_r ? 4'd0 :
                                             applyfnInt_Bool_5_3_argbuf_done);
  
  /* buf (Ty MyBool) : (applyfnInt_Bool_5_4,MyBool) > (applyfnInt_Bool_5_4_argbuf,MyBool) */
  MyBool_t applyfnInt_Bool_5_4_bufchan_d;
  logic applyfnInt_Bool_5_4_bufchan_r;
  assign applyfnInt_Bool_5_4_r = ((! applyfnInt_Bool_5_4_bufchan_d[0]) || applyfnInt_Bool_5_4_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) applyfnInt_Bool_5_4_bufchan_d <= {1'd0, 1'd0};
    else
      if (applyfnInt_Bool_5_4_r)
        applyfnInt_Bool_5_4_bufchan_d <= applyfnInt_Bool_5_4_d;
  MyBool_t applyfnInt_Bool_5_4_bufchan_buf;
  assign applyfnInt_Bool_5_4_bufchan_r = (! applyfnInt_Bool_5_4_bufchan_buf[0]);
  assign applyfnInt_Bool_5_4_argbuf_d = (applyfnInt_Bool_5_4_bufchan_buf[0] ? applyfnInt_Bool_5_4_bufchan_buf :
                                         applyfnInt_Bool_5_4_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Bool_5_4_bufchan_buf <= {1'd0, 1'd0};
    else
      if ((applyfnInt_Bool_5_4_argbuf_r && applyfnInt_Bool_5_4_bufchan_buf[0]))
        applyfnInt_Bool_5_4_bufchan_buf <= {1'd0, 1'd0};
      else if (((! applyfnInt_Bool_5_4_argbuf_r) && (! applyfnInt_Bool_5_4_bufchan_buf[0])))
        applyfnInt_Bool_5_4_bufchan_buf <= applyfnInt_Bool_5_4_bufchan_d;
  
  /* fork (Ty MyBool) : (applyfnInt_Bool_5_4_argbuf,MyBool) > [(es_14_1,MyBool),
                                                          (es_14_2,MyBool),
                                                          (es_14_3,MyBool),
                                                          (es_14_4,MyBool),
                                                          (es_14_5,MyBool),
                                                          (es_14_6,MyBool),
                                                          (es_14_7,MyBool)] */
  logic [6:0] applyfnInt_Bool_5_4_argbuf_emitted;
  logic [6:0] applyfnInt_Bool_5_4_argbuf_done;
  assign es_14_1_d = {applyfnInt_Bool_5_4_argbuf_d[1:1],
                      (applyfnInt_Bool_5_4_argbuf_d[0] && (! applyfnInt_Bool_5_4_argbuf_emitted[0]))};
  assign es_14_2_d = {applyfnInt_Bool_5_4_argbuf_d[1:1],
                      (applyfnInt_Bool_5_4_argbuf_d[0] && (! applyfnInt_Bool_5_4_argbuf_emitted[1]))};
  assign es_14_3_d = {applyfnInt_Bool_5_4_argbuf_d[1:1],
                      (applyfnInt_Bool_5_4_argbuf_d[0] && (! applyfnInt_Bool_5_4_argbuf_emitted[2]))};
  assign es_14_4_d = {applyfnInt_Bool_5_4_argbuf_d[1:1],
                      (applyfnInt_Bool_5_4_argbuf_d[0] && (! applyfnInt_Bool_5_4_argbuf_emitted[3]))};
  assign es_14_5_d = {applyfnInt_Bool_5_4_argbuf_d[1:1],
                      (applyfnInt_Bool_5_4_argbuf_d[0] && (! applyfnInt_Bool_5_4_argbuf_emitted[4]))};
  assign es_14_6_d = {applyfnInt_Bool_5_4_argbuf_d[1:1],
                      (applyfnInt_Bool_5_4_argbuf_d[0] && (! applyfnInt_Bool_5_4_argbuf_emitted[5]))};
  assign es_14_7_d = {applyfnInt_Bool_5_4_argbuf_d[1:1],
                      (applyfnInt_Bool_5_4_argbuf_d[0] && (! applyfnInt_Bool_5_4_argbuf_emitted[6]))};
  assign applyfnInt_Bool_5_4_argbuf_done = (applyfnInt_Bool_5_4_argbuf_emitted | ({es_14_7_d[0],
                                                                                   es_14_6_d[0],
                                                                                   es_14_5_d[0],
                                                                                   es_14_4_d[0],
                                                                                   es_14_3_d[0],
                                                                                   es_14_2_d[0],
                                                                                   es_14_1_d[0]} & {es_14_7_r,
                                                                                                    es_14_6_r,
                                                                                                    es_14_5_r,
                                                                                                    es_14_4_r,
                                                                                                    es_14_3_r,
                                                                                                    es_14_2_r,
                                                                                                    es_14_1_r}));
  assign applyfnInt_Bool_5_4_argbuf_r = (& applyfnInt_Bool_5_4_argbuf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) applyfnInt_Bool_5_4_argbuf_emitted <= 7'd0;
    else
      applyfnInt_Bool_5_4_argbuf_emitted <= (applyfnInt_Bool_5_4_argbuf_r ? 7'd0 :
                                             applyfnInt_Bool_5_4_argbuf_done);
  
  /* buf (Ty MyBool) : (applyfnInt_Bool_5_5,MyBool) > (applyfnInt_Bool_5_5_argbuf,MyBool) */
  MyBool_t applyfnInt_Bool_5_5_bufchan_d;
  logic applyfnInt_Bool_5_5_bufchan_r;
  assign applyfnInt_Bool_5_5_r = ((! applyfnInt_Bool_5_5_bufchan_d[0]) || applyfnInt_Bool_5_5_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) applyfnInt_Bool_5_5_bufchan_d <= {1'd0, 1'd0};
    else
      if (applyfnInt_Bool_5_5_r)
        applyfnInt_Bool_5_5_bufchan_d <= applyfnInt_Bool_5_5_d;
  MyBool_t applyfnInt_Bool_5_5_bufchan_buf;
  assign applyfnInt_Bool_5_5_bufchan_r = (! applyfnInt_Bool_5_5_bufchan_buf[0]);
  assign applyfnInt_Bool_5_5_argbuf_d = (applyfnInt_Bool_5_5_bufchan_buf[0] ? applyfnInt_Bool_5_5_bufchan_buf :
                                         applyfnInt_Bool_5_5_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Bool_5_5_bufchan_buf <= {1'd0, 1'd0};
    else
      if ((applyfnInt_Bool_5_5_argbuf_r && applyfnInt_Bool_5_5_bufchan_buf[0]))
        applyfnInt_Bool_5_5_bufchan_buf <= {1'd0, 1'd0};
      else if (((! applyfnInt_Bool_5_5_argbuf_r) && (! applyfnInt_Bool_5_5_bufchan_buf[0])))
        applyfnInt_Bool_5_5_bufchan_buf <= applyfnInt_Bool_5_5_bufchan_d;
  
  /* fork (Ty MyBool) : (applyfnInt_Bool_5_5_argbuf,MyBool) > [(es_19_1,MyBool),
                                                          (es_19_2,MyBool),
                                                          (es_19_3,MyBool),
                                                          (es_19_4,MyBool),
                                                          (es_19_5,MyBool),
                                                          (es_19_6,MyBool)] */
  logic [5:0] applyfnInt_Bool_5_5_argbuf_emitted;
  logic [5:0] applyfnInt_Bool_5_5_argbuf_done;
  assign es_19_1_d = {applyfnInt_Bool_5_5_argbuf_d[1:1],
                      (applyfnInt_Bool_5_5_argbuf_d[0] && (! applyfnInt_Bool_5_5_argbuf_emitted[0]))};
  assign es_19_2_d = {applyfnInt_Bool_5_5_argbuf_d[1:1],
                      (applyfnInt_Bool_5_5_argbuf_d[0] && (! applyfnInt_Bool_5_5_argbuf_emitted[1]))};
  assign es_19_3_d = {applyfnInt_Bool_5_5_argbuf_d[1:1],
                      (applyfnInt_Bool_5_5_argbuf_d[0] && (! applyfnInt_Bool_5_5_argbuf_emitted[2]))};
  assign es_19_4_d = {applyfnInt_Bool_5_5_argbuf_d[1:1],
                      (applyfnInt_Bool_5_5_argbuf_d[0] && (! applyfnInt_Bool_5_5_argbuf_emitted[3]))};
  assign es_19_5_d = {applyfnInt_Bool_5_5_argbuf_d[1:1],
                      (applyfnInt_Bool_5_5_argbuf_d[0] && (! applyfnInt_Bool_5_5_argbuf_emitted[4]))};
  assign es_19_6_d = {applyfnInt_Bool_5_5_argbuf_d[1:1],
                      (applyfnInt_Bool_5_5_argbuf_d[0] && (! applyfnInt_Bool_5_5_argbuf_emitted[5]))};
  assign applyfnInt_Bool_5_5_argbuf_done = (applyfnInt_Bool_5_5_argbuf_emitted | ({es_19_6_d[0],
                                                                                   es_19_5_d[0],
                                                                                   es_19_4_d[0],
                                                                                   es_19_3_d[0],
                                                                                   es_19_2_d[0],
                                                                                   es_19_1_d[0]} & {es_19_6_r,
                                                                                                    es_19_5_r,
                                                                                                    es_19_4_r,
                                                                                                    es_19_3_r,
                                                                                                    es_19_2_r,
                                                                                                    es_19_1_r}));
  assign applyfnInt_Bool_5_5_argbuf_r = (& applyfnInt_Bool_5_5_argbuf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) applyfnInt_Bool_5_5_argbuf_emitted <= 6'd0;
    else
      applyfnInt_Bool_5_5_argbuf_emitted <= (applyfnInt_Bool_5_5_argbuf_r ? 6'd0 :
                                             applyfnInt_Bool_5_5_argbuf_done);
  
  /* demux (Ty C5,
       Ty MyBool) : (applyfnInt_Bool_5_choice,C5) (lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux,MyBool) > [(applyfnInt_Bool_5_1,MyBool),
                                                                                                                                 (applyfnInt_Bool_5_2,MyBool),
                                                                                                                                 (applyfnInt_Bool_5_3,MyBool),
                                                                                                                                 (applyfnInt_Bool_5_4,MyBool),
                                                                                                                                 (applyfnInt_Bool_5_5,MyBool)] */
  logic [4:0] lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_onehotd;
  always_comb
    if ((applyfnInt_Bool_5_choice_d[0] && lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_d[0]))
      unique case (applyfnInt_Bool_5_choice_d[3:1])
        3'd0:
          lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_onehotd = 5'd1;
        3'd1:
          lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_onehotd = 5'd2;
        3'd2:
          lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_onehotd = 5'd4;
        3'd3:
          lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_onehotd = 5'd8;
        3'd4:
          lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_onehotd = 5'd16;
        default:
          lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_onehotd = 5'd0;
      endcase
    else
      lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_onehotd = 5'd0;
  assign applyfnInt_Bool_5_1_d = {lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_d[1:1],
                                  lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_onehotd[0]};
  assign applyfnInt_Bool_5_2_d = {lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_d[1:1],
                                  lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_onehotd[1]};
  assign applyfnInt_Bool_5_3_d = {lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_d[1:1],
                                  lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_onehotd[2]};
  assign applyfnInt_Bool_5_4_d = {lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_d[1:1],
                                  lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_onehotd[3]};
  assign applyfnInt_Bool_5_5_d = {lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_d[1:1],
                                  lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_onehotd[4]};
  assign lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_r = (| (lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_onehotd & {applyfnInt_Bool_5_5_r,
                                                                                                                                                                  applyfnInt_Bool_5_4_r,
                                                                                                                                                                  applyfnInt_Bool_5_3_r,
                                                                                                                                                                  applyfnInt_Bool_5_2_r,
                                                                                                                                                                  applyfnInt_Bool_5_1_r}));
  assign applyfnInt_Bool_5_choice_r = lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_r;
  
  /* destruct (Ty TupGo___MyDTInt_Bool___Int,
          Dcon TupGo___MyDTInt_Bool___Int) : (applyfnInt_Bool_5_data,TupGo___MyDTInt_Bool___Int) > [(applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intgo_8,Go),
                                                                                                    (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0,MyDTInt_Bool),
                                                                                                    (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg1,Int)] */
  logic [2:0] applyfnInt_Bool_5_data_emitted;
  logic [2:0] applyfnInt_Bool_5_data_done;
  assign applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intgo_8_d = (applyfnInt_Bool_5_data_d[0] && (! applyfnInt_Bool_5_data_emitted[0]));
  assign applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_d = (applyfnInt_Bool_5_data_d[0] && (! applyfnInt_Bool_5_data_emitted[1]));
  assign applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg1_d = {applyfnInt_Bool_5_data_d[32:1],
                                                              (applyfnInt_Bool_5_data_d[0] && (! applyfnInt_Bool_5_data_emitted[2]))};
  assign applyfnInt_Bool_5_data_done = (applyfnInt_Bool_5_data_emitted | ({applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg1_d[0],
                                                                           applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_d[0],
                                                                           applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intgo_8_d[0]} & {applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg1_r,
                                                                                                                                    applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_r,
                                                                                                                                    applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intgo_8_r}));
  assign applyfnInt_Bool_5_data_r = (& applyfnInt_Bool_5_data_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) applyfnInt_Bool_5_data_emitted <= 3'd0;
    else
      applyfnInt_Bool_5_data_emitted <= (applyfnInt_Bool_5_data_r ? 3'd0 :
                                         applyfnInt_Bool_5_data_done);
  
  /* fork (Ty MyBool) : (applyfnInt_Bool_5_resbuf,MyBool) > [(es_2_1_1,MyBool),
                                                        (es_2_1_2,MyBool),
                                                        (es_2_1_3,MyBool),
                                                        (es_2_1_4,MyBool)] */
  logic [3:0] applyfnInt_Bool_5_resbuf_emitted;
  logic [3:0] applyfnInt_Bool_5_resbuf_done;
  assign es_2_1_1_d = {applyfnInt_Bool_5_resbuf_d[1:1],
                       (applyfnInt_Bool_5_resbuf_d[0] && (! applyfnInt_Bool_5_resbuf_emitted[0]))};
  assign es_2_1_2_d = {applyfnInt_Bool_5_resbuf_d[1:1],
                       (applyfnInt_Bool_5_resbuf_d[0] && (! applyfnInt_Bool_5_resbuf_emitted[1]))};
  assign es_2_1_3_d = {applyfnInt_Bool_5_resbuf_d[1:1],
                       (applyfnInt_Bool_5_resbuf_d[0] && (! applyfnInt_Bool_5_resbuf_emitted[2]))};
  assign es_2_1_4_d = {applyfnInt_Bool_5_resbuf_d[1:1],
                       (applyfnInt_Bool_5_resbuf_d[0] && (! applyfnInt_Bool_5_resbuf_emitted[3]))};
  assign applyfnInt_Bool_5_resbuf_done = (applyfnInt_Bool_5_resbuf_emitted | ({es_2_1_4_d[0],
                                                                               es_2_1_3_d[0],
                                                                               es_2_1_2_d[0],
                                                                               es_2_1_1_d[0]} & {es_2_1_4_r,
                                                                                                 es_2_1_3_r,
                                                                                                 es_2_1_2_r,
                                                                                                 es_2_1_1_r}));
  assign applyfnInt_Bool_5_resbuf_r = (& applyfnInt_Bool_5_resbuf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) applyfnInt_Bool_5_resbuf_emitted <= 4'd0;
    else
      applyfnInt_Bool_5_resbuf_emitted <= (applyfnInt_Bool_5_resbuf_r ? 4'd0 :
                                           applyfnInt_Bool_5_resbuf_done);
  
  /* mergectrl (Ty C8,
           Ty TupGo___MyDTInt_Int___Int) : [(applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1,TupGo___MyDTInt_Int___Int),
                                            (applyfnInt_Int_5TupGo___MyDTInt_Int___Int2,TupGo___MyDTInt_Int___Int),
                                            (applyfnInt_Int_5TupGo___MyDTInt_Int___Int3,TupGo___MyDTInt_Int___Int),
                                            (applyfnInt_Int_5TupGo___MyDTInt_Int___Int4,TupGo___MyDTInt_Int___Int),
                                            (applyfnInt_Int_5TupGo___MyDTInt_Int___Int5,TupGo___MyDTInt_Int___Int),
                                            (applyfnInt_Int_5TupGo___MyDTInt_Int___Int6,TupGo___MyDTInt_Int___Int),
                                            (applyfnInt_Int_5TupGo___MyDTInt_Int___Int7,TupGo___MyDTInt_Int___Int),
                                            (applyfnInt_Int_5TupGo___MyDTInt_Int___Int8,TupGo___MyDTInt_Int___Int)] > (applyfnInt_Int_5_choice,C8) (applyfnInt_Int_5_data,TupGo___MyDTInt_Int___Int) */
  logic [7:0] applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_select_d;
  assign applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_select_d = ((| applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_select_q) ? applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_select_q :
                                                                 (applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_d[0] ? 8'd1 :
                                                                  (applyfnInt_Int_5TupGo___MyDTInt_Int___Int2_d[0] ? 8'd2 :
                                                                   (applyfnInt_Int_5TupGo___MyDTInt_Int___Int3_d[0] ? 8'd4 :
                                                                    (applyfnInt_Int_5TupGo___MyDTInt_Int___Int4_d[0] ? 8'd8 :
                                                                     (applyfnInt_Int_5TupGo___MyDTInt_Int___Int5_d[0] ? 8'd16 :
                                                                      (applyfnInt_Int_5TupGo___MyDTInt_Int___Int6_d[0] ? 8'd32 :
                                                                       (applyfnInt_Int_5TupGo___MyDTInt_Int___Int7_d[0] ? 8'd64 :
                                                                        (applyfnInt_Int_5TupGo___MyDTInt_Int___Int8_d[0] ? 8'd128 :
                                                                         8'd0)))))))));
  logic [7:0] applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_select_q <= 8'd0;
    else
      applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_select_q <= (applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_done ? 8'd0 :
                                                               applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_select_d);
  logic [1:0] applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_emit_q <= 2'd0;
    else
      applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_emit_q <= (applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_done ? 2'd0 :
                                                             applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_emit_d);
  logic [1:0] applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_emit_d;
  assign applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_emit_d = (applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_emit_q | ({applyfnInt_Int_5_choice_d[0],
                                                                                                                      applyfnInt_Int_5_data_d[0]} & {applyfnInt_Int_5_choice_r,
                                                                                                                                                     applyfnInt_Int_5_data_r}));
  logic applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_done;
  assign applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_done = (& applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_emit_d);
  assign {applyfnInt_Int_5TupGo___MyDTInt_Int___Int8_r,
          applyfnInt_Int_5TupGo___MyDTInt_Int___Int7_r,
          applyfnInt_Int_5TupGo___MyDTInt_Int___Int6_r,
          applyfnInt_Int_5TupGo___MyDTInt_Int___Int5_r,
          applyfnInt_Int_5TupGo___MyDTInt_Int___Int4_r,
          applyfnInt_Int_5TupGo___MyDTInt_Int___Int3_r,
          applyfnInt_Int_5TupGo___MyDTInt_Int___Int2_r,
          applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_r} = (applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_done ? applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_select_d :
                                                            8'd0);
  assign applyfnInt_Int_5_data_d = ((applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_select_d[0] && (! applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_emit_q[0])) ? applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_d :
                                    ((applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_select_d[1] && (! applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_emit_q[0])) ? applyfnInt_Int_5TupGo___MyDTInt_Int___Int2_d :
                                     ((applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_select_d[2] && (! applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_emit_q[0])) ? applyfnInt_Int_5TupGo___MyDTInt_Int___Int3_d :
                                      ((applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_select_d[3] && (! applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_emit_q[0])) ? applyfnInt_Int_5TupGo___MyDTInt_Int___Int4_d :
                                       ((applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_select_d[4] && (! applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_emit_q[0])) ? applyfnInt_Int_5TupGo___MyDTInt_Int___Int5_d :
                                        ((applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_select_d[5] && (! applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_emit_q[0])) ? applyfnInt_Int_5TupGo___MyDTInt_Int___Int6_d :
                                         ((applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_select_d[6] && (! applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_emit_q[0])) ? applyfnInt_Int_5TupGo___MyDTInt_Int___Int7_d :
                                          ((applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_select_d[7] && (! applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_emit_q[0])) ? applyfnInt_Int_5TupGo___MyDTInt_Int___Int8_d :
                                           {32'd0, 1'd0}))))))));
  assign applyfnInt_Int_5_choice_d = ((applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_select_d[0] && (! applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_emit_q[1])) ? C1_8_dc(1'd1) :
                                      ((applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_select_d[1] && (! applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_emit_q[1])) ? C2_8_dc(1'd1) :
                                       ((applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_select_d[2] && (! applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_emit_q[1])) ? C3_8_dc(1'd1) :
                                        ((applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_select_d[3] && (! applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_emit_q[1])) ? C4_8_dc(1'd1) :
                                         ((applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_select_d[4] && (! applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_emit_q[1])) ? C5_8_dc(1'd1) :
                                          ((applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_select_d[5] && (! applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_emit_q[1])) ? C6_8_dc(1'd1) :
                                           ((applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_select_d[6] && (! applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_emit_q[1])) ? C7_8_dc(1'd1) :
                                            ((applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_select_d[7] && (! applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_emit_q[1])) ? C8_8_dc(1'd1) :
                                             {3'd0, 1'd0}))))))));
  
  /* fork (Ty MyDTInt_Int) : (applyfnInt_Int_5TupGo___MyDTInt_Int___Intarg0_2,MyDTInt_Int) > [(arg0_2_1,MyDTInt_Int),
                                                                                         (arg0_2_2,MyDTInt_Int),
                                                                                         (arg0_2_3,MyDTInt_Int)] */
  logic [2:0] applyfnInt_Int_5TupGo___MyDTInt_Int___Intarg0_2_emitted;
  logic [2:0] applyfnInt_Int_5TupGo___MyDTInt_Int___Intarg0_2_done;
  assign arg0_2_1_d = (applyfnInt_Int_5TupGo___MyDTInt_Int___Intarg0_2_d[0] && (! applyfnInt_Int_5TupGo___MyDTInt_Int___Intarg0_2_emitted[0]));
  assign arg0_2_2_d = (applyfnInt_Int_5TupGo___MyDTInt_Int___Intarg0_2_d[0] && (! applyfnInt_Int_5TupGo___MyDTInt_Int___Intarg0_2_emitted[1]));
  assign arg0_2_3_d = (applyfnInt_Int_5TupGo___MyDTInt_Int___Intarg0_2_d[0] && (! applyfnInt_Int_5TupGo___MyDTInt_Int___Intarg0_2_emitted[2]));
  assign applyfnInt_Int_5TupGo___MyDTInt_Int___Intarg0_2_done = (applyfnInt_Int_5TupGo___MyDTInt_Int___Intarg0_2_emitted | ({arg0_2_3_d[0],
                                                                                                                             arg0_2_2_d[0],
                                                                                                                             arg0_2_1_d[0]} & {arg0_2_3_r,
                                                                                                                                               arg0_2_2_r,
                                                                                                                                               arg0_2_1_r}));
  assign applyfnInt_Int_5TupGo___MyDTInt_Int___Intarg0_2_r = (& applyfnInt_Int_5TupGo___MyDTInt_Int___Intarg0_2_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_5TupGo___MyDTInt_Int___Intarg0_2_emitted <= 3'd0;
    else
      applyfnInt_Int_5TupGo___MyDTInt_Int___Intarg0_2_emitted <= (applyfnInt_Int_5TupGo___MyDTInt_Int___Intarg0_2_r ? 3'd0 :
                                                                  applyfnInt_Int_5TupGo___MyDTInt_Int___Intarg0_2_done);
  
  /* buf (Ty Int) : (applyfnInt_Int_5_1,Int) > (applyfnInt_Int_5_resbuf,Int) */
  Int_t applyfnInt_Int_5_1_bufchan_d;
  logic applyfnInt_Int_5_1_bufchan_r;
  assign applyfnInt_Int_5_1_r = ((! applyfnInt_Int_5_1_bufchan_d[0]) || applyfnInt_Int_5_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) applyfnInt_Int_5_1_bufchan_d <= {32'd0, 1'd0};
    else
      if (applyfnInt_Int_5_1_r)
        applyfnInt_Int_5_1_bufchan_d <= applyfnInt_Int_5_1_d;
  Int_t applyfnInt_Int_5_1_bufchan_buf;
  assign applyfnInt_Int_5_1_bufchan_r = (! applyfnInt_Int_5_1_bufchan_buf[0]);
  assign applyfnInt_Int_5_resbuf_d = (applyfnInt_Int_5_1_bufchan_buf[0] ? applyfnInt_Int_5_1_bufchan_buf :
                                      applyfnInt_Int_5_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_5_1_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((applyfnInt_Int_5_resbuf_r && applyfnInt_Int_5_1_bufchan_buf[0]))
        applyfnInt_Int_5_1_bufchan_buf <= {32'd0, 1'd0};
      else if (((! applyfnInt_Int_5_resbuf_r) && (! applyfnInt_Int_5_1_bufchan_buf[0])))
        applyfnInt_Int_5_1_bufchan_buf <= applyfnInt_Int_5_1_bufchan_d;
  
  /* buf (Ty Int) : (applyfnInt_Int_5_2,Int) > (applyfnInt_Int_5_2_argbuf,Int) */
  Int_t applyfnInt_Int_5_2_bufchan_d;
  logic applyfnInt_Int_5_2_bufchan_r;
  assign applyfnInt_Int_5_2_r = ((! applyfnInt_Int_5_2_bufchan_d[0]) || applyfnInt_Int_5_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) applyfnInt_Int_5_2_bufchan_d <= {32'd0, 1'd0};
    else
      if (applyfnInt_Int_5_2_r)
        applyfnInt_Int_5_2_bufchan_d <= applyfnInt_Int_5_2_d;
  Int_t applyfnInt_Int_5_2_bufchan_buf;
  assign applyfnInt_Int_5_2_bufchan_r = (! applyfnInt_Int_5_2_bufchan_buf[0]);
  assign applyfnInt_Int_5_2_argbuf_d = (applyfnInt_Int_5_2_bufchan_buf[0] ? applyfnInt_Int_5_2_bufchan_buf :
                                        applyfnInt_Int_5_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_5_2_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((applyfnInt_Int_5_2_argbuf_r && applyfnInt_Int_5_2_bufchan_buf[0]))
        applyfnInt_Int_5_2_bufchan_buf <= {32'd0, 1'd0};
      else if (((! applyfnInt_Int_5_2_argbuf_r) && (! applyfnInt_Int_5_2_bufchan_buf[0])))
        applyfnInt_Int_5_2_bufchan_buf <= applyfnInt_Int_5_2_bufchan_d;
  
  /* dcon (Ty QTree_Int,
      Dcon QVal_Int) : [(applyfnInt_Int_5_2_argbuf,Int)] > (es_3_2_1QVal_Int,QTree_Int) */
  assign es_3_2_1QVal_Int_d = QVal_Int_dc((& {applyfnInt_Int_5_2_argbuf_d[0]}), applyfnInt_Int_5_2_argbuf_d);
  assign {applyfnInt_Int_5_2_argbuf_r} = {1 {(es_3_2_1QVal_Int_r && es_3_2_1QVal_Int_d[0])}};
  
  /* buf (Ty Int) : (applyfnInt_Int_5_3,Int) > (applyfnInt_Int_5_3_argbuf,Int) */
  Int_t applyfnInt_Int_5_3_bufchan_d;
  logic applyfnInt_Int_5_3_bufchan_r;
  assign applyfnInt_Int_5_3_r = ((! applyfnInt_Int_5_3_bufchan_d[0]) || applyfnInt_Int_5_3_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) applyfnInt_Int_5_3_bufchan_d <= {32'd0, 1'd0};
    else
      if (applyfnInt_Int_5_3_r)
        applyfnInt_Int_5_3_bufchan_d <= applyfnInt_Int_5_3_d;
  Int_t applyfnInt_Int_5_3_bufchan_buf;
  assign applyfnInt_Int_5_3_bufchan_r = (! applyfnInt_Int_5_3_bufchan_buf[0]);
  assign applyfnInt_Int_5_3_argbuf_d = (applyfnInt_Int_5_3_bufchan_buf[0] ? applyfnInt_Int_5_3_bufchan_buf :
                                        applyfnInt_Int_5_3_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_5_3_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((applyfnInt_Int_5_3_argbuf_r && applyfnInt_Int_5_3_bufchan_buf[0]))
        applyfnInt_Int_5_3_bufchan_buf <= {32'd0, 1'd0};
      else if (((! applyfnInt_Int_5_3_argbuf_r) && (! applyfnInt_Int_5_3_bufchan_buf[0])))
        applyfnInt_Int_5_3_bufchan_buf <= applyfnInt_Int_5_3_bufchan_d;
  
  /* buf (Ty Int) : (applyfnInt_Int_5_3_argbuf,Int) > (es_1_1_argbuf,Int) */
  Int_t applyfnInt_Int_5_3_argbuf_bufchan_d;
  logic applyfnInt_Int_5_3_argbuf_bufchan_r;
  assign applyfnInt_Int_5_3_argbuf_r = ((! applyfnInt_Int_5_3_argbuf_bufchan_d[0]) || applyfnInt_Int_5_3_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_5_3_argbuf_bufchan_d <= {32'd0, 1'd0};
    else
      if (applyfnInt_Int_5_3_argbuf_r)
        applyfnInt_Int_5_3_argbuf_bufchan_d <= applyfnInt_Int_5_3_argbuf_d;
  Int_t applyfnInt_Int_5_3_argbuf_bufchan_buf;
  assign applyfnInt_Int_5_3_argbuf_bufchan_r = (! applyfnInt_Int_5_3_argbuf_bufchan_buf[0]);
  assign es_1_1_argbuf_d = (applyfnInt_Int_5_3_argbuf_bufchan_buf[0] ? applyfnInt_Int_5_3_argbuf_bufchan_buf :
                            applyfnInt_Int_5_3_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_5_3_argbuf_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((es_1_1_argbuf_r && applyfnInt_Int_5_3_argbuf_bufchan_buf[0]))
        applyfnInt_Int_5_3_argbuf_bufchan_buf <= {32'd0, 1'd0};
      else if (((! es_1_1_argbuf_r) && (! applyfnInt_Int_5_3_argbuf_bufchan_buf[0])))
        applyfnInt_Int_5_3_argbuf_bufchan_buf <= applyfnInt_Int_5_3_argbuf_bufchan_d;
  
  /* buf (Ty Int) : (applyfnInt_Int_5_4,Int) > (applyfnInt_Int_5_4_argbuf,Int) */
  Int_t applyfnInt_Int_5_4_bufchan_d;
  logic applyfnInt_Int_5_4_bufchan_r;
  assign applyfnInt_Int_5_4_r = ((! applyfnInt_Int_5_4_bufchan_d[0]) || applyfnInt_Int_5_4_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) applyfnInt_Int_5_4_bufchan_d <= {32'd0, 1'd0};
    else
      if (applyfnInt_Int_5_4_r)
        applyfnInt_Int_5_4_bufchan_d <= applyfnInt_Int_5_4_d;
  Int_t applyfnInt_Int_5_4_bufchan_buf;
  assign applyfnInt_Int_5_4_bufchan_r = (! applyfnInt_Int_5_4_bufchan_buf[0]);
  assign applyfnInt_Int_5_4_argbuf_d = (applyfnInt_Int_5_4_bufchan_buf[0] ? applyfnInt_Int_5_4_bufchan_buf :
                                        applyfnInt_Int_5_4_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_5_4_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((applyfnInt_Int_5_4_argbuf_r && applyfnInt_Int_5_4_bufchan_buf[0]))
        applyfnInt_Int_5_4_bufchan_buf <= {32'd0, 1'd0};
      else if (((! applyfnInt_Int_5_4_argbuf_r) && (! applyfnInt_Int_5_4_bufchan_buf[0])))
        applyfnInt_Int_5_4_bufchan_buf <= applyfnInt_Int_5_4_bufchan_d;
  
  /* dcon (Ty QTree_Int,
      Dcon QVal_Int) : [(applyfnInt_Int_5_4_argbuf,Int)] > (es_3_1_1QVal_Int,QTree_Int) */
  assign es_3_1_1QVal_Int_d = QVal_Int_dc((& {applyfnInt_Int_5_4_argbuf_d[0]}), applyfnInt_Int_5_4_argbuf_d);
  assign {applyfnInt_Int_5_4_argbuf_r} = {1 {(es_3_1_1QVal_Int_r && es_3_1_1QVal_Int_d[0])}};
  
  /* buf (Ty Int) : (applyfnInt_Int_5_5,Int) > (applyfnInt_Int_5_5_argbuf,Int) */
  Int_t applyfnInt_Int_5_5_bufchan_d;
  logic applyfnInt_Int_5_5_bufchan_r;
  assign applyfnInt_Int_5_5_r = ((! applyfnInt_Int_5_5_bufchan_d[0]) || applyfnInt_Int_5_5_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) applyfnInt_Int_5_5_bufchan_d <= {32'd0, 1'd0};
    else
      if (applyfnInt_Int_5_5_r)
        applyfnInt_Int_5_5_bufchan_d <= applyfnInt_Int_5_5_d;
  Int_t applyfnInt_Int_5_5_bufchan_buf;
  assign applyfnInt_Int_5_5_bufchan_r = (! applyfnInt_Int_5_5_bufchan_buf[0]);
  assign applyfnInt_Int_5_5_argbuf_d = (applyfnInt_Int_5_5_bufchan_buf[0] ? applyfnInt_Int_5_5_bufchan_buf :
                                        applyfnInt_Int_5_5_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_5_5_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((applyfnInt_Int_5_5_argbuf_r && applyfnInt_Int_5_5_bufchan_buf[0]))
        applyfnInt_Int_5_5_bufchan_buf <= {32'd0, 1'd0};
      else if (((! applyfnInt_Int_5_5_argbuf_r) && (! applyfnInt_Int_5_5_bufchan_buf[0])))
        applyfnInt_Int_5_5_bufchan_buf <= applyfnInt_Int_5_5_bufchan_d;
  
  /* buf (Ty Int) : (applyfnInt_Int_5_5_argbuf,Int) > (es_9_1_argbuf,Int) */
  Int_t applyfnInt_Int_5_5_argbuf_bufchan_d;
  logic applyfnInt_Int_5_5_argbuf_bufchan_r;
  assign applyfnInt_Int_5_5_argbuf_r = ((! applyfnInt_Int_5_5_argbuf_bufchan_d[0]) || applyfnInt_Int_5_5_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_5_5_argbuf_bufchan_d <= {32'd0, 1'd0};
    else
      if (applyfnInt_Int_5_5_argbuf_r)
        applyfnInt_Int_5_5_argbuf_bufchan_d <= applyfnInt_Int_5_5_argbuf_d;
  Int_t applyfnInt_Int_5_5_argbuf_bufchan_buf;
  assign applyfnInt_Int_5_5_argbuf_bufchan_r = (! applyfnInt_Int_5_5_argbuf_bufchan_buf[0]);
  assign es_9_1_argbuf_d = (applyfnInt_Int_5_5_argbuf_bufchan_buf[0] ? applyfnInt_Int_5_5_argbuf_bufchan_buf :
                            applyfnInt_Int_5_5_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_5_5_argbuf_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((es_9_1_argbuf_r && applyfnInt_Int_5_5_argbuf_bufchan_buf[0]))
        applyfnInt_Int_5_5_argbuf_bufchan_buf <= {32'd0, 1'd0};
      else if (((! es_9_1_argbuf_r) && (! applyfnInt_Int_5_5_argbuf_bufchan_buf[0])))
        applyfnInt_Int_5_5_argbuf_bufchan_buf <= applyfnInt_Int_5_5_argbuf_bufchan_d;
  
  /* buf (Ty Int) : (applyfnInt_Int_5_6,Int) > (applyfnInt_Int_5_6_argbuf,Int) */
  Int_t applyfnInt_Int_5_6_bufchan_d;
  logic applyfnInt_Int_5_6_bufchan_r;
  assign applyfnInt_Int_5_6_r = ((! applyfnInt_Int_5_6_bufchan_d[0]) || applyfnInt_Int_5_6_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) applyfnInt_Int_5_6_bufchan_d <= {32'd0, 1'd0};
    else
      if (applyfnInt_Int_5_6_r)
        applyfnInt_Int_5_6_bufchan_d <= applyfnInt_Int_5_6_d;
  Int_t applyfnInt_Int_5_6_bufchan_buf;
  assign applyfnInt_Int_5_6_bufchan_r = (! applyfnInt_Int_5_6_bufchan_buf[0]);
  assign applyfnInt_Int_5_6_argbuf_d = (applyfnInt_Int_5_6_bufchan_buf[0] ? applyfnInt_Int_5_6_bufchan_buf :
                                        applyfnInt_Int_5_6_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_5_6_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((applyfnInt_Int_5_6_argbuf_r && applyfnInt_Int_5_6_bufchan_buf[0]))
        applyfnInt_Int_5_6_bufchan_buf <= {32'd0, 1'd0};
      else if (((! applyfnInt_Int_5_6_argbuf_r) && (! applyfnInt_Int_5_6_bufchan_buf[0])))
        applyfnInt_Int_5_6_bufchan_buf <= applyfnInt_Int_5_6_bufchan_d;
  
  /* dcon (Ty QTree_Int,
      Dcon QVal_Int) : [(applyfnInt_Int_5_6_argbuf,Int)] > (es_11_1QVal_Int,QTree_Int) */
  assign es_11_1QVal_Int_d = QVal_Int_dc((& {applyfnInt_Int_5_6_argbuf_d[0]}), applyfnInt_Int_5_6_argbuf_d);
  assign {applyfnInt_Int_5_6_argbuf_r} = {1 {(es_11_1QVal_Int_r && es_11_1QVal_Int_d[0])}};
  
  /* buf (Ty Int) : (applyfnInt_Int_5_7,Int) > (applyfnInt_Int_5_7_argbuf,Int) */
  Int_t applyfnInt_Int_5_7_bufchan_d;
  logic applyfnInt_Int_5_7_bufchan_r;
  assign applyfnInt_Int_5_7_r = ((! applyfnInt_Int_5_7_bufchan_d[0]) || applyfnInt_Int_5_7_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) applyfnInt_Int_5_7_bufchan_d <= {32'd0, 1'd0};
    else
      if (applyfnInt_Int_5_7_r)
        applyfnInt_Int_5_7_bufchan_d <= applyfnInt_Int_5_7_d;
  Int_t applyfnInt_Int_5_7_bufchan_buf;
  assign applyfnInt_Int_5_7_bufchan_r = (! applyfnInt_Int_5_7_bufchan_buf[0]);
  assign applyfnInt_Int_5_7_argbuf_d = (applyfnInt_Int_5_7_bufchan_buf[0] ? applyfnInt_Int_5_7_bufchan_buf :
                                        applyfnInt_Int_5_7_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_5_7_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((applyfnInt_Int_5_7_argbuf_r && applyfnInt_Int_5_7_bufchan_buf[0]))
        applyfnInt_Int_5_7_bufchan_buf <= {32'd0, 1'd0};
      else if (((! applyfnInt_Int_5_7_argbuf_r) && (! applyfnInt_Int_5_7_bufchan_buf[0])))
        applyfnInt_Int_5_7_bufchan_buf <= applyfnInt_Int_5_7_bufchan_d;
  
  /* buf (Ty Int) : (applyfnInt_Int_5_7_argbuf,Int) > (es_16_1_argbuf,Int) */
  Int_t applyfnInt_Int_5_7_argbuf_bufchan_d;
  logic applyfnInt_Int_5_7_argbuf_bufchan_r;
  assign applyfnInt_Int_5_7_argbuf_r = ((! applyfnInt_Int_5_7_argbuf_bufchan_d[0]) || applyfnInt_Int_5_7_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_5_7_argbuf_bufchan_d <= {32'd0, 1'd0};
    else
      if (applyfnInt_Int_5_7_argbuf_r)
        applyfnInt_Int_5_7_argbuf_bufchan_d <= applyfnInt_Int_5_7_argbuf_d;
  Int_t applyfnInt_Int_5_7_argbuf_bufchan_buf;
  assign applyfnInt_Int_5_7_argbuf_bufchan_r = (! applyfnInt_Int_5_7_argbuf_bufchan_buf[0]);
  assign es_16_1_argbuf_d = (applyfnInt_Int_5_7_argbuf_bufchan_buf[0] ? applyfnInt_Int_5_7_argbuf_bufchan_buf :
                             applyfnInt_Int_5_7_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_5_7_argbuf_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((es_16_1_argbuf_r && applyfnInt_Int_5_7_argbuf_bufchan_buf[0]))
        applyfnInt_Int_5_7_argbuf_bufchan_buf <= {32'd0, 1'd0};
      else if (((! es_16_1_argbuf_r) && (! applyfnInt_Int_5_7_argbuf_bufchan_buf[0])))
        applyfnInt_Int_5_7_argbuf_bufchan_buf <= applyfnInt_Int_5_7_argbuf_bufchan_d;
  
  /* buf (Ty Int) : (applyfnInt_Int_5_8,Int) > (applyfnInt_Int_5_8_argbuf,Int) */
  Int_t applyfnInt_Int_5_8_bufchan_d;
  logic applyfnInt_Int_5_8_bufchan_r;
  assign applyfnInt_Int_5_8_r = ((! applyfnInt_Int_5_8_bufchan_d[0]) || applyfnInt_Int_5_8_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) applyfnInt_Int_5_8_bufchan_d <= {32'd0, 1'd0};
    else
      if (applyfnInt_Int_5_8_r)
        applyfnInt_Int_5_8_bufchan_d <= applyfnInt_Int_5_8_d;
  Int_t applyfnInt_Int_5_8_bufchan_buf;
  assign applyfnInt_Int_5_8_bufchan_r = (! applyfnInt_Int_5_8_bufchan_buf[0]);
  assign applyfnInt_Int_5_8_argbuf_d = (applyfnInt_Int_5_8_bufchan_buf[0] ? applyfnInt_Int_5_8_bufchan_buf :
                                        applyfnInt_Int_5_8_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_5_8_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((applyfnInt_Int_5_8_argbuf_r && applyfnInt_Int_5_8_bufchan_buf[0]))
        applyfnInt_Int_5_8_bufchan_buf <= {32'd0, 1'd0};
      else if (((! applyfnInt_Int_5_8_argbuf_r) && (! applyfnInt_Int_5_8_bufchan_buf[0])))
        applyfnInt_Int_5_8_bufchan_buf <= applyfnInt_Int_5_8_bufchan_d;
  
  /* dcon (Ty QTree_Int,
      Dcon QVal_Int) : [(applyfnInt_Int_5_8_argbuf,Int)] > (es_20_1QVal_Int,QTree_Int) */
  assign es_20_1QVal_Int_d = QVal_Int_dc((& {applyfnInt_Int_5_8_argbuf_d[0]}), applyfnInt_Int_5_8_argbuf_d);
  assign {applyfnInt_Int_5_8_argbuf_r} = {1 {(es_20_1QVal_Int_r && es_20_1QVal_Int_d[0])}};
  
  /* demux (Ty C8,
       Ty Int) : (applyfnInt_Int_5_choice,C8) (es_0_1_1I#_mux_mux,Int) > [(applyfnInt_Int_5_1,Int),
                                                                          (applyfnInt_Int_5_2,Int),
                                                                          (applyfnInt_Int_5_3,Int),
                                                                          (applyfnInt_Int_5_4,Int),
                                                                          (applyfnInt_Int_5_5,Int),
                                                                          (applyfnInt_Int_5_6,Int),
                                                                          (applyfnInt_Int_5_7,Int),
                                                                          (applyfnInt_Int_5_8,Int)] */
  logic [7:0] \es_0_1_1I#_mux_mux_onehotd ;
  always_comb
    if ((applyfnInt_Int_5_choice_d[0] && \es_0_1_1I#_mux_mux_d [0]))
      unique case (applyfnInt_Int_5_choice_d[3:1])
        3'd0: \es_0_1_1I#_mux_mux_onehotd  = 8'd1;
        3'd1: \es_0_1_1I#_mux_mux_onehotd  = 8'd2;
        3'd2: \es_0_1_1I#_mux_mux_onehotd  = 8'd4;
        3'd3: \es_0_1_1I#_mux_mux_onehotd  = 8'd8;
        3'd4: \es_0_1_1I#_mux_mux_onehotd  = 8'd16;
        3'd5: \es_0_1_1I#_mux_mux_onehotd  = 8'd32;
        3'd6: \es_0_1_1I#_mux_mux_onehotd  = 8'd64;
        3'd7: \es_0_1_1I#_mux_mux_onehotd  = 8'd128;
        default: \es_0_1_1I#_mux_mux_onehotd  = 8'd0;
      endcase
    else \es_0_1_1I#_mux_mux_onehotd  = 8'd0;
  assign applyfnInt_Int_5_1_d = {\es_0_1_1I#_mux_mux_d [32:1],
                                 \es_0_1_1I#_mux_mux_onehotd [0]};
  assign applyfnInt_Int_5_2_d = {\es_0_1_1I#_mux_mux_d [32:1],
                                 \es_0_1_1I#_mux_mux_onehotd [1]};
  assign applyfnInt_Int_5_3_d = {\es_0_1_1I#_mux_mux_d [32:1],
                                 \es_0_1_1I#_mux_mux_onehotd [2]};
  assign applyfnInt_Int_5_4_d = {\es_0_1_1I#_mux_mux_d [32:1],
                                 \es_0_1_1I#_mux_mux_onehotd [3]};
  assign applyfnInt_Int_5_5_d = {\es_0_1_1I#_mux_mux_d [32:1],
                                 \es_0_1_1I#_mux_mux_onehotd [4]};
  assign applyfnInt_Int_5_6_d = {\es_0_1_1I#_mux_mux_d [32:1],
                                 \es_0_1_1I#_mux_mux_onehotd [5]};
  assign applyfnInt_Int_5_7_d = {\es_0_1_1I#_mux_mux_d [32:1],
                                 \es_0_1_1I#_mux_mux_onehotd [6]};
  assign applyfnInt_Int_5_8_d = {\es_0_1_1I#_mux_mux_d [32:1],
                                 \es_0_1_1I#_mux_mux_onehotd [7]};
  assign \es_0_1_1I#_mux_mux_r  = (| (\es_0_1_1I#_mux_mux_onehotd  & {applyfnInt_Int_5_8_r,
                                                                      applyfnInt_Int_5_7_r,
                                                                      applyfnInt_Int_5_6_r,
                                                                      applyfnInt_Int_5_5_r,
                                                                      applyfnInt_Int_5_4_r,
                                                                      applyfnInt_Int_5_3_r,
                                                                      applyfnInt_Int_5_2_r,
                                                                      applyfnInt_Int_5_1_r}));
  assign applyfnInt_Int_5_choice_r = \es_0_1_1I#_mux_mux_r ;
  
  /* destruct (Ty TupGo___MyDTInt_Int___Int,
          Dcon TupGo___MyDTInt_Int___Int) : (applyfnInt_Int_5_data,TupGo___MyDTInt_Int___Int) > [(applyfnInt_Int_5TupGo___MyDTInt_Int___Intgo_9,Go),
                                                                                                 (applyfnInt_Int_5TupGo___MyDTInt_Int___Intarg0_2,MyDTInt_Int),
                                                                                                 (applyfnInt_Int_5TupGo___MyDTInt_Int___Intarg1_1,Int)] */
  logic [2:0] applyfnInt_Int_5_data_emitted;
  logic [2:0] applyfnInt_Int_5_data_done;
  assign applyfnInt_Int_5TupGo___MyDTInt_Int___Intgo_9_d = (applyfnInt_Int_5_data_d[0] && (! applyfnInt_Int_5_data_emitted[0]));
  assign applyfnInt_Int_5TupGo___MyDTInt_Int___Intarg0_2_d = (applyfnInt_Int_5_data_d[0] && (! applyfnInt_Int_5_data_emitted[1]));
  assign applyfnInt_Int_5TupGo___MyDTInt_Int___Intarg1_1_d = {applyfnInt_Int_5_data_d[32:1],
                                                              (applyfnInt_Int_5_data_d[0] && (! applyfnInt_Int_5_data_emitted[2]))};
  assign applyfnInt_Int_5_data_done = (applyfnInt_Int_5_data_emitted | ({applyfnInt_Int_5TupGo___MyDTInt_Int___Intarg1_1_d[0],
                                                                         applyfnInt_Int_5TupGo___MyDTInt_Int___Intarg0_2_d[0],
                                                                         applyfnInt_Int_5TupGo___MyDTInt_Int___Intgo_9_d[0]} & {applyfnInt_Int_5TupGo___MyDTInt_Int___Intarg1_1_r,
                                                                                                                                applyfnInt_Int_5TupGo___MyDTInt_Int___Intarg0_2_r,
                                                                                                                                applyfnInt_Int_5TupGo___MyDTInt_Int___Intgo_9_r}));
  assign applyfnInt_Int_5_data_r = (& applyfnInt_Int_5_data_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) applyfnInt_Int_5_data_emitted <= 3'd0;
    else
      applyfnInt_Int_5_data_emitted <= (applyfnInt_Int_5_data_r ? 3'd0 :
                                        applyfnInt_Int_5_data_done);
  
  /* buf (Ty Int) : (applyfnInt_Int_5_resbuf,Int) > (es_1_1_1_argbuf,Int) */
  Int_t applyfnInt_Int_5_resbuf_bufchan_d;
  logic applyfnInt_Int_5_resbuf_bufchan_r;
  assign applyfnInt_Int_5_resbuf_r = ((! applyfnInt_Int_5_resbuf_bufchan_d[0]) || applyfnInt_Int_5_resbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_5_resbuf_bufchan_d <= {32'd0, 1'd0};
    else
      if (applyfnInt_Int_5_resbuf_r)
        applyfnInt_Int_5_resbuf_bufchan_d <= applyfnInt_Int_5_resbuf_d;
  Int_t applyfnInt_Int_5_resbuf_bufchan_buf;
  assign applyfnInt_Int_5_resbuf_bufchan_r = (! applyfnInt_Int_5_resbuf_bufchan_buf[0]);
  assign es_1_1_1_argbuf_d = (applyfnInt_Int_5_resbuf_bufchan_buf[0] ? applyfnInt_Int_5_resbuf_bufchan_buf :
                              applyfnInt_Int_5_resbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_5_resbuf_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((es_1_1_1_argbuf_r && applyfnInt_Int_5_resbuf_bufchan_buf[0]))
        applyfnInt_Int_5_resbuf_bufchan_buf <= {32'd0, 1'd0};
      else if (((! es_1_1_1_argbuf_r) && (! applyfnInt_Int_5_resbuf_bufchan_buf[0])))
        applyfnInt_Int_5_resbuf_bufchan_buf <= applyfnInt_Int_5_resbuf_bufchan_d;
  
  /* mergectrl (Ty C3,
           Ty TupMyDTInt_Int_Int___Int___Int) : [(applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1,TupMyDTInt_Int_Int___Int___Int),
                                                 (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int2,TupMyDTInt_Int_Int___Int___Int),
                                                 (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int3,TupMyDTInt_Int_Int___Int___Int)] > (applyfnInt_Int_Int_5_choice,C3) (applyfnInt_Int_Int_5_data,TupMyDTInt_Int_Int___Int___Int) */
  logic [2:0] applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_select_d;
  assign applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_select_d = ((| applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_select_q) ? applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_select_q :
                                                                          (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_d[0] ? 3'd1 :
                                                                           (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int2_d[0] ? 3'd2 :
                                                                            (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int3_d[0] ? 3'd4 :
                                                                             3'd0))));
  logic [2:0] applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_select_q <= 3'd0;
    else
      applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_select_q <= (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_done ? 3'd0 :
                                                                        applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_select_d);
  logic [1:0] applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_emit_q <= 2'd0;
    else
      applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_emit_q <= (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_done ? 2'd0 :
                                                                      applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_emit_d);
  logic [1:0] applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_emit_d;
  assign applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_emit_d = (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_emit_q | ({applyfnInt_Int_Int_5_choice_d[0],
                                                                                                                                        applyfnInt_Int_Int_5_data_d[0]} & {applyfnInt_Int_Int_5_choice_r,
                                                                                                                                                                           applyfnInt_Int_Int_5_data_r}));
  logic applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_done;
  assign applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_done = (& applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_emit_d);
  assign {applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int3_r,
          applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int2_r,
          applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_r} = (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_done ? applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_select_d :
                                                                     3'd0);
  assign applyfnInt_Int_Int_5_data_d = ((applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_select_d[0] && (! applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_emit_q[0])) ? applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_d :
                                        ((applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_select_d[1] && (! applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_emit_q[0])) ? applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int2_d :
                                         ((applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_select_d[2] && (! applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_emit_q[0])) ? applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int3_d :
                                          {64'd0, 1'd0})));
  assign applyfnInt_Int_Int_5_choice_d = ((applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_select_d[0] && (! applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_emit_q[1])) ? C1_3_dc(1'd1) :
                                          ((applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_select_d[1] && (! applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_emit_q[1])) ? C2_3_dc(1'd1) :
                                           ((applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_select_d[2] && (! applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_emit_q[1])) ? C3_3_dc(1'd1) :
                                            {2'd0, 1'd0})));
  
  /* fork (Ty MyDTInt_Int_Int) : (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_4,MyDTInt_Int_Int) > [(arg0_4_1,MyDTInt_Int_Int),
                                                                                                          (arg0_4_2,MyDTInt_Int_Int),
                                                                                                          (arg0_4_3,MyDTInt_Int_Int)] */
  logic [2:0] applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_4_emitted;
  logic [2:0] applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_4_done;
  assign arg0_4_1_d = (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_4_d[0] && (! applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_4_emitted[0]));
  assign arg0_4_2_d = (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_4_d[0] && (! applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_4_emitted[1]));
  assign arg0_4_3_d = (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_4_d[0] && (! applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_4_emitted[2]));
  assign applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_4_done = (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_4_emitted | ({arg0_4_3_d[0],
                                                                                                                                               arg0_4_2_d[0],
                                                                                                                                               arg0_4_1_d[0]} & {arg0_4_3_r,
                                                                                                                                                                 arg0_4_2_r,
                                                                                                                                                                 arg0_4_1_r}));
  assign applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_4_r = (& applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_4_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_4_emitted <= 3'd0;
    else
      applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_4_emitted <= (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_4_r ? 3'd0 :
                                                                           applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_4_done);
  
  /* buf (Ty Int) : (applyfnInt_Int_Int_5_1,Int) > (applyfnInt_Int_Int_5_resbuf,Int) */
  Int_t applyfnInt_Int_Int_5_1_bufchan_d;
  logic applyfnInt_Int_Int_5_1_bufchan_r;
  assign applyfnInt_Int_Int_5_1_r = ((! applyfnInt_Int_Int_5_1_bufchan_d[0]) || applyfnInt_Int_Int_5_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_Int_5_1_bufchan_d <= {32'd0, 1'd0};
    else
      if (applyfnInt_Int_Int_5_1_r)
        applyfnInt_Int_Int_5_1_bufchan_d <= applyfnInt_Int_Int_5_1_d;
  Int_t applyfnInt_Int_Int_5_1_bufchan_buf;
  assign applyfnInt_Int_Int_5_1_bufchan_r = (! applyfnInt_Int_Int_5_1_bufchan_buf[0]);
  assign applyfnInt_Int_Int_5_resbuf_d = (applyfnInt_Int_Int_5_1_bufchan_buf[0] ? applyfnInt_Int_Int_5_1_bufchan_buf :
                                          applyfnInt_Int_Int_5_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_Int_5_1_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((applyfnInt_Int_Int_5_resbuf_r && applyfnInt_Int_Int_5_1_bufchan_buf[0]))
        applyfnInt_Int_Int_5_1_bufchan_buf <= {32'd0, 1'd0};
      else if (((! applyfnInt_Int_Int_5_resbuf_r) && (! applyfnInt_Int_Int_5_1_bufchan_buf[0])))
        applyfnInt_Int_Int_5_1_bufchan_buf <= applyfnInt_Int_Int_5_1_bufchan_d;
  
  /* buf (Ty Int) : (applyfnInt_Int_Int_5_2,Int) > (applyfnInt_Int_Int_5_2_argbuf,Int) */
  Int_t applyfnInt_Int_Int_5_2_bufchan_d;
  logic applyfnInt_Int_Int_5_2_bufchan_r;
  assign applyfnInt_Int_Int_5_2_r = ((! applyfnInt_Int_Int_5_2_bufchan_d[0]) || applyfnInt_Int_Int_5_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_Int_5_2_bufchan_d <= {32'd0, 1'd0};
    else
      if (applyfnInt_Int_Int_5_2_r)
        applyfnInt_Int_Int_5_2_bufchan_d <= applyfnInt_Int_Int_5_2_d;
  Int_t applyfnInt_Int_Int_5_2_bufchan_buf;
  assign applyfnInt_Int_Int_5_2_bufchan_r = (! applyfnInt_Int_Int_5_2_bufchan_buf[0]);
  assign applyfnInt_Int_Int_5_2_argbuf_d = (applyfnInt_Int_Int_5_2_bufchan_buf[0] ? applyfnInt_Int_Int_5_2_bufchan_buf :
                                            applyfnInt_Int_Int_5_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_Int_5_2_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((applyfnInt_Int_Int_5_2_argbuf_r && applyfnInt_Int_Int_5_2_bufchan_buf[0]))
        applyfnInt_Int_Int_5_2_bufchan_buf <= {32'd0, 1'd0};
      else if (((! applyfnInt_Int_Int_5_2_argbuf_r) && (! applyfnInt_Int_Int_5_2_bufchan_buf[0])))
        applyfnInt_Int_Int_5_2_bufchan_buf <= applyfnInt_Int_Int_5_2_bufchan_d;
  
  /* buf (Ty Int) : (applyfnInt_Int_Int_5_2_argbuf,Int) > (es_18_1_argbuf,Int) */
  Int_t applyfnInt_Int_Int_5_2_argbuf_bufchan_d;
  logic applyfnInt_Int_Int_5_2_argbuf_bufchan_r;
  assign applyfnInt_Int_Int_5_2_argbuf_r = ((! applyfnInt_Int_Int_5_2_argbuf_bufchan_d[0]) || applyfnInt_Int_Int_5_2_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_Int_5_2_argbuf_bufchan_d <= {32'd0, 1'd0};
    else
      if (applyfnInt_Int_Int_5_2_argbuf_r)
        applyfnInt_Int_Int_5_2_argbuf_bufchan_d <= applyfnInt_Int_Int_5_2_argbuf_d;
  Int_t applyfnInt_Int_Int_5_2_argbuf_bufchan_buf;
  assign applyfnInt_Int_Int_5_2_argbuf_bufchan_r = (! applyfnInt_Int_Int_5_2_argbuf_bufchan_buf[0]);
  assign es_18_1_argbuf_d = (applyfnInt_Int_Int_5_2_argbuf_bufchan_buf[0] ? applyfnInt_Int_Int_5_2_argbuf_bufchan_buf :
                             applyfnInt_Int_Int_5_2_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_Int_5_2_argbuf_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((es_18_1_argbuf_r && applyfnInt_Int_Int_5_2_argbuf_bufchan_buf[0]))
        applyfnInt_Int_Int_5_2_argbuf_bufchan_buf <= {32'd0, 1'd0};
      else if (((! es_18_1_argbuf_r) && (! applyfnInt_Int_Int_5_2_argbuf_bufchan_buf[0])))
        applyfnInt_Int_Int_5_2_argbuf_bufchan_buf <= applyfnInt_Int_Int_5_2_argbuf_bufchan_d;
  
  /* buf (Ty Int) : (applyfnInt_Int_Int_5_3,Int) > (applyfnInt_Int_Int_5_3_argbuf,Int) */
  Int_t applyfnInt_Int_Int_5_3_bufchan_d;
  logic applyfnInt_Int_Int_5_3_bufchan_r;
  assign applyfnInt_Int_Int_5_3_r = ((! applyfnInt_Int_Int_5_3_bufchan_d[0]) || applyfnInt_Int_Int_5_3_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_Int_5_3_bufchan_d <= {32'd0, 1'd0};
    else
      if (applyfnInt_Int_Int_5_3_r)
        applyfnInt_Int_Int_5_3_bufchan_d <= applyfnInt_Int_Int_5_3_d;
  Int_t applyfnInt_Int_Int_5_3_bufchan_buf;
  assign applyfnInt_Int_Int_5_3_bufchan_r = (! applyfnInt_Int_Int_5_3_bufchan_buf[0]);
  assign applyfnInt_Int_Int_5_3_argbuf_d = (applyfnInt_Int_Int_5_3_bufchan_buf[0] ? applyfnInt_Int_Int_5_3_bufchan_buf :
                                            applyfnInt_Int_Int_5_3_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_Int_5_3_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((applyfnInt_Int_Int_5_3_argbuf_r && applyfnInt_Int_Int_5_3_bufchan_buf[0]))
        applyfnInt_Int_Int_5_3_bufchan_buf <= {32'd0, 1'd0};
      else if (((! applyfnInt_Int_Int_5_3_argbuf_r) && (! applyfnInt_Int_Int_5_3_bufchan_buf[0])))
        applyfnInt_Int_Int_5_3_bufchan_buf <= applyfnInt_Int_Int_5_3_bufchan_d;
  
  /* buf (Ty Int) : (applyfnInt_Int_Int_5_3_argbuf,Int) > (es_22_1_argbuf,Int) */
  Int_t applyfnInt_Int_Int_5_3_argbuf_bufchan_d;
  logic applyfnInt_Int_Int_5_3_argbuf_bufchan_r;
  assign applyfnInt_Int_Int_5_3_argbuf_r = ((! applyfnInt_Int_Int_5_3_argbuf_bufchan_d[0]) || applyfnInt_Int_Int_5_3_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_Int_5_3_argbuf_bufchan_d <= {32'd0, 1'd0};
    else
      if (applyfnInt_Int_Int_5_3_argbuf_r)
        applyfnInt_Int_Int_5_3_argbuf_bufchan_d <= applyfnInt_Int_Int_5_3_argbuf_d;
  Int_t applyfnInt_Int_Int_5_3_argbuf_bufchan_buf;
  assign applyfnInt_Int_Int_5_3_argbuf_bufchan_r = (! applyfnInt_Int_Int_5_3_argbuf_bufchan_buf[0]);
  assign es_22_1_argbuf_d = (applyfnInt_Int_Int_5_3_argbuf_bufchan_buf[0] ? applyfnInt_Int_Int_5_3_argbuf_bufchan_buf :
                             applyfnInt_Int_Int_5_3_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_Int_5_3_argbuf_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((es_22_1_argbuf_r && applyfnInt_Int_Int_5_3_argbuf_bufchan_buf[0]))
        applyfnInt_Int_Int_5_3_argbuf_bufchan_buf <= {32'd0, 1'd0};
      else if (((! es_22_1_argbuf_r) && (! applyfnInt_Int_Int_5_3_argbuf_bufchan_buf[0])))
        applyfnInt_Int_Int_5_3_argbuf_bufchan_buf <= applyfnInt_Int_Int_5_3_argbuf_bufchan_d;
  
  /* demux (Ty C3,
       Ty Int) : (applyfnInt_Int_Int_5_choice,C3) (es_0_2_1I#_mux_mux_mux,Int) > [(applyfnInt_Int_Int_5_1,Int),
                                                                                  (applyfnInt_Int_Int_5_2,Int),
                                                                                  (applyfnInt_Int_Int_5_3,Int)] */
  logic [2:0] \es_0_2_1I#_mux_mux_mux_onehotd ;
  always_comb
    if ((applyfnInt_Int_Int_5_choice_d[0] && \es_0_2_1I#_mux_mux_mux_d [0]))
      unique case (applyfnInt_Int_Int_5_choice_d[2:1])
        2'd0: \es_0_2_1I#_mux_mux_mux_onehotd  = 3'd1;
        2'd1: \es_0_2_1I#_mux_mux_mux_onehotd  = 3'd2;
        2'd2: \es_0_2_1I#_mux_mux_mux_onehotd  = 3'd4;
        default: \es_0_2_1I#_mux_mux_mux_onehotd  = 3'd0;
      endcase
    else \es_0_2_1I#_mux_mux_mux_onehotd  = 3'd0;
  assign applyfnInt_Int_Int_5_1_d = {\es_0_2_1I#_mux_mux_mux_d [32:1],
                                     \es_0_2_1I#_mux_mux_mux_onehotd [0]};
  assign applyfnInt_Int_Int_5_2_d = {\es_0_2_1I#_mux_mux_mux_d [32:1],
                                     \es_0_2_1I#_mux_mux_mux_onehotd [1]};
  assign applyfnInt_Int_Int_5_3_d = {\es_0_2_1I#_mux_mux_mux_d [32:1],
                                     \es_0_2_1I#_mux_mux_mux_onehotd [2]};
  assign \es_0_2_1I#_mux_mux_mux_r  = (| (\es_0_2_1I#_mux_mux_mux_onehotd  & {applyfnInt_Int_Int_5_3_r,
                                                                              applyfnInt_Int_Int_5_2_r,
                                                                              applyfnInt_Int_Int_5_1_r}));
  assign applyfnInt_Int_Int_5_choice_r = \es_0_2_1I#_mux_mux_mux_r ;
  
  /* destruct (Ty TupMyDTInt_Int_Int___Int___Int,
          Dcon TupMyDTInt_Int_Int___Int___Int) : (applyfnInt_Int_Int_5_data,TupMyDTInt_Int_Int___Int___Int) > [(applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_4,MyDTInt_Int_Int),
                                                                                                               (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg2,Int),
                                                                                                               (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg1_2,Int)] */
  logic [2:0] applyfnInt_Int_Int_5_data_emitted;
  logic [2:0] applyfnInt_Int_Int_5_data_done;
  assign applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_4_d = (applyfnInt_Int_Int_5_data_d[0] && (! applyfnInt_Int_Int_5_data_emitted[0]));
  assign applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg2_d = {applyfnInt_Int_Int_5_data_d[32:1],
                                                                     (applyfnInt_Int_Int_5_data_d[0] && (! applyfnInt_Int_Int_5_data_emitted[1]))};
  assign applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg1_2_d = {applyfnInt_Int_Int_5_data_d[64:33],
                                                                       (applyfnInt_Int_Int_5_data_d[0] && (! applyfnInt_Int_Int_5_data_emitted[2]))};
  assign applyfnInt_Int_Int_5_data_done = (applyfnInt_Int_Int_5_data_emitted | ({applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg1_2_d[0],
                                                                                 applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg2_d[0],
                                                                                 applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_4_d[0]} & {applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg1_2_r,
                                                                                                                                                   applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg2_r,
                                                                                                                                                   applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_4_r}));
  assign applyfnInt_Int_Int_5_data_r = (& applyfnInt_Int_Int_5_data_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) applyfnInt_Int_Int_5_data_emitted <= 3'd0;
    else
      applyfnInt_Int_Int_5_data_emitted <= (applyfnInt_Int_Int_5_data_r ? 3'd0 :
                                            applyfnInt_Int_Int_5_data_done);
  
  /* buf (Ty Int) : (applyfnInt_Int_Int_5_resbuf,Int) > (es_13_1_argbuf,Int) */
  Int_t applyfnInt_Int_Int_5_resbuf_bufchan_d;
  logic applyfnInt_Int_Int_5_resbuf_bufchan_r;
  assign applyfnInt_Int_Int_5_resbuf_r = ((! applyfnInt_Int_Int_5_resbuf_bufchan_d[0]) || applyfnInt_Int_Int_5_resbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_Int_5_resbuf_bufchan_d <= {32'd0, 1'd0};
    else
      if (applyfnInt_Int_Int_5_resbuf_r)
        applyfnInt_Int_Int_5_resbuf_bufchan_d <= applyfnInt_Int_Int_5_resbuf_d;
  Int_t applyfnInt_Int_Int_5_resbuf_bufchan_buf;
  assign applyfnInt_Int_Int_5_resbuf_bufchan_r = (! applyfnInt_Int_Int_5_resbuf_bufchan_buf[0]);
  assign es_13_1_argbuf_d = (applyfnInt_Int_Int_5_resbuf_bufchan_buf[0] ? applyfnInt_Int_Int_5_resbuf_bufchan_buf :
                             applyfnInt_Int_Int_5_resbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_Int_5_resbuf_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((es_13_1_argbuf_r && applyfnInt_Int_Int_5_resbuf_bufchan_buf[0]))
        applyfnInt_Int_Int_5_resbuf_bufchan_buf <= {32'd0, 1'd0};
      else if (((! es_13_1_argbuf_r) && (! applyfnInt_Int_Int_5_resbuf_bufchan_buf[0])))
        applyfnInt_Int_Int_5_resbuf_bufchan_buf <= applyfnInt_Int_Int_5_resbuf_bufchan_d;
  
  /* demux (Ty MyDTInt_Bool,
       Ty Int) : (arg0_1,MyDTInt_Bool) (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg1,Int) > [(arg0_1Dcon_is_z_1,Int)] */
  assign arg0_1Dcon_is_z_1_d = {applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg1_d[32:1],
                                (arg0_1_d[0] && applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg1_d[0])};
  assign applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg1_r = (arg0_1Dcon_is_z_1_r && (arg0_1_d[0] && applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg1_d[0]));
  assign arg0_1_r = (arg0_1Dcon_is_z_1_r && (arg0_1_d[0] && applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg1_d[0]));
  
  /* fork (Ty Int) : (arg0_1Dcon_is_z_1,Int) > [(arg0_1Dcon_is_z_1_1,Int),
                                           (arg0_1Dcon_is_z_1_2,Int),
                                           (arg0_1Dcon_is_z_1_3,Int),
                                           (arg0_1Dcon_is_z_1_4,Int)] */
  logic [3:0] arg0_1Dcon_is_z_1_emitted;
  logic [3:0] arg0_1Dcon_is_z_1_done;
  assign arg0_1Dcon_is_z_1_1_d = {arg0_1Dcon_is_z_1_d[32:1],
                                  (arg0_1Dcon_is_z_1_d[0] && (! arg0_1Dcon_is_z_1_emitted[0]))};
  assign arg0_1Dcon_is_z_1_2_d = {arg0_1Dcon_is_z_1_d[32:1],
                                  (arg0_1Dcon_is_z_1_d[0] && (! arg0_1Dcon_is_z_1_emitted[1]))};
  assign arg0_1Dcon_is_z_1_3_d = {arg0_1Dcon_is_z_1_d[32:1],
                                  (arg0_1Dcon_is_z_1_d[0] && (! arg0_1Dcon_is_z_1_emitted[2]))};
  assign arg0_1Dcon_is_z_1_4_d = {arg0_1Dcon_is_z_1_d[32:1],
                                  (arg0_1Dcon_is_z_1_d[0] && (! arg0_1Dcon_is_z_1_emitted[3]))};
  assign arg0_1Dcon_is_z_1_done = (arg0_1Dcon_is_z_1_emitted | ({arg0_1Dcon_is_z_1_4_d[0],
                                                                 arg0_1Dcon_is_z_1_3_d[0],
                                                                 arg0_1Dcon_is_z_1_2_d[0],
                                                                 arg0_1Dcon_is_z_1_1_d[0]} & {arg0_1Dcon_is_z_1_4_r,
                                                                                              arg0_1Dcon_is_z_1_3_r,
                                                                                              arg0_1Dcon_is_z_1_2_r,
                                                                                              arg0_1Dcon_is_z_1_1_r}));
  assign arg0_1Dcon_is_z_1_r = (& arg0_1Dcon_is_z_1_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) arg0_1Dcon_is_z_1_emitted <= 4'd0;
    else
      arg0_1Dcon_is_z_1_emitted <= (arg0_1Dcon_is_z_1_r ? 4'd0 :
                                    arg0_1Dcon_is_z_1_done);
  
  /* destruct (Ty Int,
          Dcon I#) : (arg0_1Dcon_is_z_1_1I#,Int) > [(x1ah2_destruct,Int#)] */
  assign x1ah2_destruct_d = {\arg0_1Dcon_is_z_1_1I#_d [32:1],
                             \arg0_1Dcon_is_z_1_1I#_d [0]};
  assign \arg0_1Dcon_is_z_1_1I#_r  = x1ah2_destruct_r;
  
  /* demux (Ty Int,
       Ty Int) : (arg0_1Dcon_is_z_1_2,Int) (arg0_1Dcon_is_z_1_1,Int) > [(arg0_1Dcon_is_z_1_1I#,Int)] */
  assign \arg0_1Dcon_is_z_1_1I#_d  = {arg0_1Dcon_is_z_1_1_d[32:1],
                                      (arg0_1Dcon_is_z_1_2_d[0] && arg0_1Dcon_is_z_1_1_d[0])};
  assign arg0_1Dcon_is_z_1_1_r = (\arg0_1Dcon_is_z_1_1I#_r  && (arg0_1Dcon_is_z_1_2_d[0] && arg0_1Dcon_is_z_1_1_d[0]));
  assign arg0_1Dcon_is_z_1_2_r = (\arg0_1Dcon_is_z_1_1I#_r  && (arg0_1Dcon_is_z_1_2_d[0] && arg0_1Dcon_is_z_1_1_d[0]));
  
  /* demux (Ty Int,
       Ty Go) : (arg0_1Dcon_is_z_1_3,Int) (arg0_2Dcon_is_z_1,Go) > [(arg0_1Dcon_is_z_1_3I#,Go)] */
  assign \arg0_1Dcon_is_z_1_3I#_d  = (arg0_1Dcon_is_z_1_3_d[0] && arg0_2Dcon_is_z_1_d[0]);
  assign arg0_2Dcon_is_z_1_r = (\arg0_1Dcon_is_z_1_3I#_r  && (arg0_1Dcon_is_z_1_3_d[0] && arg0_2Dcon_is_z_1_d[0]));
  assign arg0_1Dcon_is_z_1_3_r = (\arg0_1Dcon_is_z_1_3I#_r  && (arg0_1Dcon_is_z_1_3_d[0] && arg0_2Dcon_is_z_1_d[0]));
  
  /* fork (Ty Go) : (arg0_1Dcon_is_z_1_3I#,Go) > [(arg0_1Dcon_is_z_1_3I#_1,Go),
                                             (arg0_1Dcon_is_z_1_3I#_2,Go),
                                             (arg0_1Dcon_is_z_1_3I#_3,Go)] */
  logic [2:0] \arg0_1Dcon_is_z_1_3I#_emitted ;
  logic [2:0] \arg0_1Dcon_is_z_1_3I#_done ;
  assign \arg0_1Dcon_is_z_1_3I#_1_d  = (\arg0_1Dcon_is_z_1_3I#_d [0] && (! \arg0_1Dcon_is_z_1_3I#_emitted [0]));
  assign \arg0_1Dcon_is_z_1_3I#_2_d  = (\arg0_1Dcon_is_z_1_3I#_d [0] && (! \arg0_1Dcon_is_z_1_3I#_emitted [1]));
  assign \arg0_1Dcon_is_z_1_3I#_3_d  = (\arg0_1Dcon_is_z_1_3I#_d [0] && (! \arg0_1Dcon_is_z_1_3I#_emitted [2]));
  assign \arg0_1Dcon_is_z_1_3I#_done  = (\arg0_1Dcon_is_z_1_3I#_emitted  | ({\arg0_1Dcon_is_z_1_3I#_3_d [0],
                                                                             \arg0_1Dcon_is_z_1_3I#_2_d [0],
                                                                             \arg0_1Dcon_is_z_1_3I#_1_d [0]} & {\arg0_1Dcon_is_z_1_3I#_3_r ,
                                                                                                                \arg0_1Dcon_is_z_1_3I#_2_r ,
                                                                                                                \arg0_1Dcon_is_z_1_3I#_1_r }));
  assign \arg0_1Dcon_is_z_1_3I#_r  = (& \arg0_1Dcon_is_z_1_3I#_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \arg0_1Dcon_is_z_1_3I#_emitted  <= 3'd0;
    else
      \arg0_1Dcon_is_z_1_3I#_emitted  <= (\arg0_1Dcon_is_z_1_3I#_r  ? 3'd0 :
                                          \arg0_1Dcon_is_z_1_3I#_done );
  
  /* buf (Ty Go) : (arg0_1Dcon_is_z_1_3I#_1,Go) > (arg0_1Dcon_is_z_1_3I#_1_argbuf,Go) */
  Go_t \arg0_1Dcon_is_z_1_3I#_1_bufchan_d ;
  logic \arg0_1Dcon_is_z_1_3I#_1_bufchan_r ;
  assign \arg0_1Dcon_is_z_1_3I#_1_r  = ((! \arg0_1Dcon_is_z_1_3I#_1_bufchan_d [0]) || \arg0_1Dcon_is_z_1_3I#_1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \arg0_1Dcon_is_z_1_3I#_1_bufchan_d  <= 1'd0;
    else
      if (\arg0_1Dcon_is_z_1_3I#_1_r )
        \arg0_1Dcon_is_z_1_3I#_1_bufchan_d  <= \arg0_1Dcon_is_z_1_3I#_1_d ;
  Go_t \arg0_1Dcon_is_z_1_3I#_1_bufchan_buf ;
  assign \arg0_1Dcon_is_z_1_3I#_1_bufchan_r  = (! \arg0_1Dcon_is_z_1_3I#_1_bufchan_buf [0]);
  assign \arg0_1Dcon_is_z_1_3I#_1_argbuf_d  = (\arg0_1Dcon_is_z_1_3I#_1_bufchan_buf [0] ? \arg0_1Dcon_is_z_1_3I#_1_bufchan_buf  :
                                               \arg0_1Dcon_is_z_1_3I#_1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \arg0_1Dcon_is_z_1_3I#_1_bufchan_buf  <= 1'd0;
    else
      if ((\arg0_1Dcon_is_z_1_3I#_1_argbuf_r  && \arg0_1Dcon_is_z_1_3I#_1_bufchan_buf [0]))
        \arg0_1Dcon_is_z_1_3I#_1_bufchan_buf  <= 1'd0;
      else if (((! \arg0_1Dcon_is_z_1_3I#_1_argbuf_r ) && (! \arg0_1Dcon_is_z_1_3I#_1_bufchan_buf [0])))
        \arg0_1Dcon_is_z_1_3I#_1_bufchan_buf  <= \arg0_1Dcon_is_z_1_3I#_1_bufchan_d ;
  
  /* const (Ty Int#,
       Lit 0) : (arg0_1Dcon_is_z_1_3I#_1_argbuf,Go) > (arg0_1Dcon_is_z_1_3I#_1_argbuf_0,Int#) */
  assign \arg0_1Dcon_is_z_1_3I#_1_argbuf_0_d  = {32'd0,
                                                 \arg0_1Dcon_is_z_1_3I#_1_argbuf_d [0]};
  assign \arg0_1Dcon_is_z_1_3I#_1_argbuf_r  = \arg0_1Dcon_is_z_1_3I#_1_argbuf_0_r ;
  
  /* op_eq (Ty Int#) : (arg0_1Dcon_is_z_1_3I#_1_argbuf_0,Int#) (x1ah2_destruct,Int#) > (lizzieLet1_1wild1Xr_1_Eq,Bool) */
  assign lizzieLet1_1wild1Xr_1_Eq_d = {(\arg0_1Dcon_is_z_1_3I#_1_argbuf_0_d [32:1] == x1ah2_destruct_d[32:1]),
                                       (\arg0_1Dcon_is_z_1_3I#_1_argbuf_0_d [0] && x1ah2_destruct_d[0])};
  assign {\arg0_1Dcon_is_z_1_3I#_1_argbuf_0_r ,
          x1ah2_destruct_r} = {2 {(lizzieLet1_1wild1Xr_1_Eq_r && lizzieLet1_1wild1Xr_1_Eq_d[0])}};
  
  /* buf (Ty Go) : (arg0_1Dcon_is_z_1_3I#_2,Go) > (arg0_1Dcon_is_z_1_3I#_2_argbuf,Go) */
  Go_t \arg0_1Dcon_is_z_1_3I#_2_bufchan_d ;
  logic \arg0_1Dcon_is_z_1_3I#_2_bufchan_r ;
  assign \arg0_1Dcon_is_z_1_3I#_2_r  = ((! \arg0_1Dcon_is_z_1_3I#_2_bufchan_d [0]) || \arg0_1Dcon_is_z_1_3I#_2_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \arg0_1Dcon_is_z_1_3I#_2_bufchan_d  <= 1'd0;
    else
      if (\arg0_1Dcon_is_z_1_3I#_2_r )
        \arg0_1Dcon_is_z_1_3I#_2_bufchan_d  <= \arg0_1Dcon_is_z_1_3I#_2_d ;
  Go_t \arg0_1Dcon_is_z_1_3I#_2_bufchan_buf ;
  assign \arg0_1Dcon_is_z_1_3I#_2_bufchan_r  = (! \arg0_1Dcon_is_z_1_3I#_2_bufchan_buf [0]);
  assign \arg0_1Dcon_is_z_1_3I#_2_argbuf_d  = (\arg0_1Dcon_is_z_1_3I#_2_bufchan_buf [0] ? \arg0_1Dcon_is_z_1_3I#_2_bufchan_buf  :
                                               \arg0_1Dcon_is_z_1_3I#_2_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \arg0_1Dcon_is_z_1_3I#_2_bufchan_buf  <= 1'd0;
    else
      if ((\arg0_1Dcon_is_z_1_3I#_2_argbuf_r  && \arg0_1Dcon_is_z_1_3I#_2_bufchan_buf [0]))
        \arg0_1Dcon_is_z_1_3I#_2_bufchan_buf  <= 1'd0;
      else if (((! \arg0_1Dcon_is_z_1_3I#_2_argbuf_r ) && (! \arg0_1Dcon_is_z_1_3I#_2_bufchan_buf [0])))
        \arg0_1Dcon_is_z_1_3I#_2_bufchan_buf  <= \arg0_1Dcon_is_z_1_3I#_2_bufchan_d ;
  
  /* dcon (Ty TupGo___Bool,
      Dcon TupGo___Bool) : [(arg0_1Dcon_is_z_1_3I#_2_argbuf,Go),
                            (lizzieLet2_1_argbuf,Bool)] > (boolConvert_1TupGo___Bool_1,TupGo___Bool) */
  assign boolConvert_1TupGo___Bool_1_d = TupGo___Bool_dc((& {\arg0_1Dcon_is_z_1_3I#_2_argbuf_d [0],
                                                             lizzieLet2_1_argbuf_d[0]}), \arg0_1Dcon_is_z_1_3I#_2_argbuf_d , lizzieLet2_1_argbuf_d);
  assign {\arg0_1Dcon_is_z_1_3I#_2_argbuf_r ,
          lizzieLet2_1_argbuf_r} = {2 {(boolConvert_1TupGo___Bool_1_r && boolConvert_1TupGo___Bool_1_d[0])}};
  
  /* mux (Ty Int,
     Ty MyBool) : (arg0_1Dcon_is_z_1_4,Int) [(lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux,MyBool)] > (lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux,MyBool) */
  assign lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_d = {lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_d[1:1],
                                                                             (arg0_1Dcon_is_z_1_4_d[0] && lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_d[0])};
  assign lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_r = (lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_r && (arg0_1Dcon_is_z_1_4_d[0] && lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_d[0]));
  assign arg0_1Dcon_is_z_1_4_r = (lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_r && (arg0_1Dcon_is_z_1_4_d[0] && lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_d[0]));
  
  /* demux (Ty MyDTInt_Bool,
       Ty Go) : (arg0_2,MyDTInt_Bool) (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intgo_8,Go) > [(arg0_2Dcon_is_z_1,Go)] */
  assign arg0_2Dcon_is_z_1_d = (arg0_2_d[0] && applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intgo_8_d[0]);
  assign applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intgo_8_r = (arg0_2Dcon_is_z_1_r && (arg0_2_d[0] && applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intgo_8_d[0]));
  assign arg0_2_r = (arg0_2Dcon_is_z_1_r && (arg0_2_d[0] && applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intgo_8_d[0]));
  
  /* demux (Ty MyDTInt_Int,
       Ty Int) : (arg0_2_1,MyDTInt_Int) (applyfnInt_Int_5TupGo___MyDTInt_Int___Intarg1_1,Int) > [(arg0_2_1Dcon_main1,Int)] */
  assign arg0_2_1Dcon_main1_d = {applyfnInt_Int_5TupGo___MyDTInt_Int___Intarg1_1_d[32:1],
                                 (arg0_2_1_d[0] && applyfnInt_Int_5TupGo___MyDTInt_Int___Intarg1_1_d[0])};
  assign applyfnInt_Int_5TupGo___MyDTInt_Int___Intarg1_1_r = (arg0_2_1Dcon_main1_r && (arg0_2_1_d[0] && applyfnInt_Int_5TupGo___MyDTInt_Int___Intarg1_1_d[0]));
  assign arg0_2_1_r = (arg0_2_1Dcon_main1_r && (arg0_2_1_d[0] && applyfnInt_Int_5TupGo___MyDTInt_Int___Intarg1_1_d[0]));
  
  /* fork (Ty Int) : (arg0_2_1Dcon_main1,Int) > [(arg0_2_1Dcon_main1_1,Int),
                                            (arg0_2_1Dcon_main1_2,Int),
                                            (arg0_2_1Dcon_main1_3,Int),
                                            (arg0_2_1Dcon_main1_4,Int)] */
  logic [3:0] arg0_2_1Dcon_main1_emitted;
  logic [3:0] arg0_2_1Dcon_main1_done;
  assign arg0_2_1Dcon_main1_1_d = {arg0_2_1Dcon_main1_d[32:1],
                                   (arg0_2_1Dcon_main1_d[0] && (! arg0_2_1Dcon_main1_emitted[0]))};
  assign arg0_2_1Dcon_main1_2_d = {arg0_2_1Dcon_main1_d[32:1],
                                   (arg0_2_1Dcon_main1_d[0] && (! arg0_2_1Dcon_main1_emitted[1]))};
  assign arg0_2_1Dcon_main1_3_d = {arg0_2_1Dcon_main1_d[32:1],
                                   (arg0_2_1Dcon_main1_d[0] && (! arg0_2_1Dcon_main1_emitted[2]))};
  assign arg0_2_1Dcon_main1_4_d = {arg0_2_1Dcon_main1_d[32:1],
                                   (arg0_2_1Dcon_main1_d[0] && (! arg0_2_1Dcon_main1_emitted[3]))};
  assign arg0_2_1Dcon_main1_done = (arg0_2_1Dcon_main1_emitted | ({arg0_2_1Dcon_main1_4_d[0],
                                                                   arg0_2_1Dcon_main1_3_d[0],
                                                                   arg0_2_1Dcon_main1_2_d[0],
                                                                   arg0_2_1Dcon_main1_1_d[0]} & {arg0_2_1Dcon_main1_4_r,
                                                                                                 arg0_2_1Dcon_main1_3_r,
                                                                                                 arg0_2_1Dcon_main1_2_r,
                                                                                                 arg0_2_1Dcon_main1_1_r}));
  assign arg0_2_1Dcon_main1_r = (& arg0_2_1Dcon_main1_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) arg0_2_1Dcon_main1_emitted <= 4'd0;
    else
      arg0_2_1Dcon_main1_emitted <= (arg0_2_1Dcon_main1_r ? 4'd0 :
                                     arg0_2_1Dcon_main1_done);
  
  /* destruct (Ty Int,
          Dcon I#) : (arg0_2_1Dcon_main1_1I#,Int) > [(x1agS_destruct,Int#)] */
  assign x1agS_destruct_d = {\arg0_2_1Dcon_main1_1I#_d [32:1],
                             \arg0_2_1Dcon_main1_1I#_d [0]};
  assign \arg0_2_1Dcon_main1_1I#_r  = x1agS_destruct_r;
  
  /* demux (Ty Int,
       Ty Int) : (arg0_2_1Dcon_main1_2,Int) (arg0_2_1Dcon_main1_1,Int) > [(arg0_2_1Dcon_main1_1I#,Int)] */
  assign \arg0_2_1Dcon_main1_1I#_d  = {arg0_2_1Dcon_main1_1_d[32:1],
                                       (arg0_2_1Dcon_main1_2_d[0] && arg0_2_1Dcon_main1_1_d[0])};
  assign arg0_2_1Dcon_main1_1_r = (\arg0_2_1Dcon_main1_1I#_r  && (arg0_2_1Dcon_main1_2_d[0] && arg0_2_1Dcon_main1_1_d[0]));
  assign arg0_2_1Dcon_main1_2_r = (\arg0_2_1Dcon_main1_1I#_r  && (arg0_2_1Dcon_main1_2_d[0] && arg0_2_1Dcon_main1_1_d[0]));
  
  /* demux (Ty Int,
       Ty Go) : (arg0_2_1Dcon_main1_3,Int) (arg0_2_2Dcon_main1,Go) > [(arg0_2_1Dcon_main1_3I#,Go)] */
  assign \arg0_2_1Dcon_main1_3I#_d  = (arg0_2_1Dcon_main1_3_d[0] && arg0_2_2Dcon_main1_d[0]);
  assign arg0_2_2Dcon_main1_r = (\arg0_2_1Dcon_main1_3I#_r  && (arg0_2_1Dcon_main1_3_d[0] && arg0_2_2Dcon_main1_d[0]));
  assign arg0_2_1Dcon_main1_3_r = (\arg0_2_1Dcon_main1_3I#_r  && (arg0_2_1Dcon_main1_3_d[0] && arg0_2_2Dcon_main1_d[0]));
  
  /* buf (Ty Go) : (arg0_2_1Dcon_main1_3I#,Go) > (arg0_2_1Dcon_main1_3I#_1_argbuf,Go) */
  Go_t \arg0_2_1Dcon_main1_3I#_bufchan_d ;
  logic \arg0_2_1Dcon_main1_3I#_bufchan_r ;
  assign \arg0_2_1Dcon_main1_3I#_r  = ((! \arg0_2_1Dcon_main1_3I#_bufchan_d [0]) || \arg0_2_1Dcon_main1_3I#_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \arg0_2_1Dcon_main1_3I#_bufchan_d  <= 1'd0;
    else
      if (\arg0_2_1Dcon_main1_3I#_r )
        \arg0_2_1Dcon_main1_3I#_bufchan_d  <= \arg0_2_1Dcon_main1_3I#_d ;
  Go_t \arg0_2_1Dcon_main1_3I#_bufchan_buf ;
  assign \arg0_2_1Dcon_main1_3I#_bufchan_r  = (! \arg0_2_1Dcon_main1_3I#_bufchan_buf [0]);
  assign \arg0_2_1Dcon_main1_3I#_1_argbuf_d  = (\arg0_2_1Dcon_main1_3I#_bufchan_buf [0] ? \arg0_2_1Dcon_main1_3I#_bufchan_buf  :
                                                \arg0_2_1Dcon_main1_3I#_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \arg0_2_1Dcon_main1_3I#_bufchan_buf  <= 1'd0;
    else
      if ((\arg0_2_1Dcon_main1_3I#_1_argbuf_r  && \arg0_2_1Dcon_main1_3I#_bufchan_buf [0]))
        \arg0_2_1Dcon_main1_3I#_bufchan_buf  <= 1'd0;
      else if (((! \arg0_2_1Dcon_main1_3I#_1_argbuf_r ) && (! \arg0_2_1Dcon_main1_3I#_bufchan_buf [0])))
        \arg0_2_1Dcon_main1_3I#_bufchan_buf  <= \arg0_2_1Dcon_main1_3I#_bufchan_d ;
  
  /* const (Ty Int#,
       Lit 2) : (arg0_2_1Dcon_main1_3I#_1_argbuf,Go) > (arg0_2_1Dcon_main1_3I#_1_argbuf_2,Int#) */
  assign \arg0_2_1Dcon_main1_3I#_1_argbuf_2_d  = {32'd2,
                                                  \arg0_2_1Dcon_main1_3I#_1_argbuf_d [0]};
  assign \arg0_2_1Dcon_main1_3I#_1_argbuf_r  = \arg0_2_1Dcon_main1_3I#_1_argbuf_2_r ;
  
  /* mux (Ty Int,
     Ty Int) : (arg0_2_1Dcon_main1_4,Int) [(es_0_1_1I#,Int)] > (es_0_1_1I#_mux,Int) */
  assign \es_0_1_1I#_mux_d  = {\es_0_1_1I#_d [32:1],
                               (arg0_2_1Dcon_main1_4_d[0] && \es_0_1_1I#_d [0])};
  assign \es_0_1_1I#_r  = (\es_0_1_1I#_mux_r  && (arg0_2_1Dcon_main1_4_d[0] && \es_0_1_1I#_d [0]));
  assign arg0_2_1Dcon_main1_4_r = (\es_0_1_1I#_mux_r  && (arg0_2_1Dcon_main1_4_d[0] && \es_0_1_1I#_d [0]));
  
  /* demux (Ty MyDTInt_Int,
       Ty Go) : (arg0_2_2,MyDTInt_Int) (applyfnInt_Int_5TupGo___MyDTInt_Int___Intgo_9,Go) > [(arg0_2_2Dcon_main1,Go)] */
  assign arg0_2_2Dcon_main1_d = (arg0_2_2_d[0] && applyfnInt_Int_5TupGo___MyDTInt_Int___Intgo_9_d[0]);
  assign applyfnInt_Int_5TupGo___MyDTInt_Int___Intgo_9_r = (arg0_2_2Dcon_main1_r && (arg0_2_2_d[0] && applyfnInt_Int_5TupGo___MyDTInt_Int___Intgo_9_d[0]));
  assign arg0_2_2_r = (arg0_2_2Dcon_main1_r && (arg0_2_2_d[0] && applyfnInt_Int_5TupGo___MyDTInt_Int___Intgo_9_d[0]));
  
  /* mux (Ty MyDTInt_Int,
     Ty Int) : (arg0_2_3,MyDTInt_Int) [(es_0_1_1I#_mux,Int)] > (es_0_1_1I#_mux_mux,Int) */
  assign \es_0_1_1I#_mux_mux_d  = {\es_0_1_1I#_mux_d [32:1],
                                   (arg0_2_3_d[0] && \es_0_1_1I#_mux_d [0])};
  assign \es_0_1_1I#_mux_r  = (\es_0_1_1I#_mux_mux_r  && (arg0_2_3_d[0] && \es_0_1_1I#_mux_d [0]));
  assign arg0_2_3_r = (\es_0_1_1I#_mux_mux_r  && (arg0_2_3_d[0] && \es_0_1_1I#_mux_d [0]));
  
  /* mux (Ty MyDTInt_Bool,
     Ty MyBool) : (arg0_3,MyDTInt_Bool) [(lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux,MyBool)] > (lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux,MyBool) */
  assign lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_d = {lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_d[1:1],
                                                                                 (arg0_3_d[0] && lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_d[0])};
  assign lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_r = (lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_r && (arg0_3_d[0] && lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_d[0]));
  assign arg0_3_r = (lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_r && (arg0_3_d[0] && lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_d[0]));
  
  /* demux (Ty MyDTInt_Int_Int,
       Ty Int) : (arg0_4_1,MyDTInt_Int_Int) (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg1_2,Int) > [(arg0_4_1Dcon_$fNumInt_$c+,Int)] */
  assign \arg0_4_1Dcon_$fNumInt_$c+_d  = {applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg1_2_d[32:1],
                                          (arg0_4_1_d[0] && applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg1_2_d[0])};
  assign applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg1_2_r = (\arg0_4_1Dcon_$fNumInt_$c+_r  && (arg0_4_1_d[0] && applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg1_2_d[0]));
  assign arg0_4_1_r = (\arg0_4_1Dcon_$fNumInt_$c+_r  && (arg0_4_1_d[0] && applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg1_2_d[0]));
  
  /* demux (Ty MyDTInt_Int_Int,
       Ty Int) : (arg0_4_2,MyDTInt_Int_Int) (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg2,Int) > [(arg0_4_2Dcon_$fNumInt_$c+,Int)] */
  assign \arg0_4_2Dcon_$fNumInt_$c+_d  = {applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg2_d[32:1],
                                          (arg0_4_2_d[0] && applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg2_d[0])};
  assign applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg2_r = (\arg0_4_2Dcon_$fNumInt_$c+_r  && (arg0_4_2_d[0] && applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg2_d[0]));
  assign arg0_4_2_r = (\arg0_4_2Dcon_$fNumInt_$c+_r  && (arg0_4_2_d[0] && applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg2_d[0]));
  
  /* fork (Ty Int) : (arg0_4_2Dcon_$fNumInt_$c+,Int) > [(arg0_4_2Dcon_$fNumInt_$c+_1,Int),
                                                   (arg0_4_2Dcon_$fNumInt_$c+_2,Int),
                                                   (arg0_4_2Dcon_$fNumInt_$c+_3,Int),
                                                   (arg0_4_2Dcon_$fNumInt_$c+_4,Int)] */
  logic [3:0] \arg0_4_2Dcon_$fNumInt_$c+_emitted ;
  logic [3:0] \arg0_4_2Dcon_$fNumInt_$c+_done ;
  assign \arg0_4_2Dcon_$fNumInt_$c+_1_d  = {\arg0_4_2Dcon_$fNumInt_$c+_d [32:1],
                                            (\arg0_4_2Dcon_$fNumInt_$c+_d [0] && (! \arg0_4_2Dcon_$fNumInt_$c+_emitted [0]))};
  assign \arg0_4_2Dcon_$fNumInt_$c+_2_d  = {\arg0_4_2Dcon_$fNumInt_$c+_d [32:1],
                                            (\arg0_4_2Dcon_$fNumInt_$c+_d [0] && (! \arg0_4_2Dcon_$fNumInt_$c+_emitted [1]))};
  assign \arg0_4_2Dcon_$fNumInt_$c+_3_d  = {\arg0_4_2Dcon_$fNumInt_$c+_d [32:1],
                                            (\arg0_4_2Dcon_$fNumInt_$c+_d [0] && (! \arg0_4_2Dcon_$fNumInt_$c+_emitted [2]))};
  assign \arg0_4_2Dcon_$fNumInt_$c+_4_d  = {\arg0_4_2Dcon_$fNumInt_$c+_d [32:1],
                                            (\arg0_4_2Dcon_$fNumInt_$c+_d [0] && (! \arg0_4_2Dcon_$fNumInt_$c+_emitted [3]))};
  assign \arg0_4_2Dcon_$fNumInt_$c+_done  = (\arg0_4_2Dcon_$fNumInt_$c+_emitted  | ({\arg0_4_2Dcon_$fNumInt_$c+_4_d [0],
                                                                                     \arg0_4_2Dcon_$fNumInt_$c+_3_d [0],
                                                                                     \arg0_4_2Dcon_$fNumInt_$c+_2_d [0],
                                                                                     \arg0_4_2Dcon_$fNumInt_$c+_1_d [0]} & {\arg0_4_2Dcon_$fNumInt_$c+_4_r ,
                                                                                                                            \arg0_4_2Dcon_$fNumInt_$c+_3_r ,
                                                                                                                            \arg0_4_2Dcon_$fNumInt_$c+_2_r ,
                                                                                                                            \arg0_4_2Dcon_$fNumInt_$c+_1_r }));
  assign \arg0_4_2Dcon_$fNumInt_$c+_r  = (& \arg0_4_2Dcon_$fNumInt_$c+_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \arg0_4_2Dcon_$fNumInt_$c+_emitted  <= 4'd0;
    else
      \arg0_4_2Dcon_$fNumInt_$c+_emitted  <= (\arg0_4_2Dcon_$fNumInt_$c+_r  ? 4'd0 :
                                              \arg0_4_2Dcon_$fNumInt_$c+_done );
  
  /* destruct (Ty Int,
          Dcon I#) : (arg0_4_2Dcon_$fNumInt_$c+_1I#,Int) > [(xa1lV_destruct,Int#)] */
  assign xa1lV_destruct_d = {\arg0_4_2Dcon_$fNumInt_$c+_1I#_d [32:1],
                             \arg0_4_2Dcon_$fNumInt_$c+_1I#_d [0]};
  assign \arg0_4_2Dcon_$fNumInt_$c+_1I#_r  = xa1lV_destruct_r;
  
  /* demux (Ty Int,
       Ty Int) : (arg0_4_2Dcon_$fNumInt_$c+_2,Int) (arg0_4_2Dcon_$fNumInt_$c+_1,Int) > [(arg0_4_2Dcon_$fNumInt_$c+_1I#,Int)] */
  assign \arg0_4_2Dcon_$fNumInt_$c+_1I#_d  = {\arg0_4_2Dcon_$fNumInt_$c+_1_d [32:1],
                                              (\arg0_4_2Dcon_$fNumInt_$c+_2_d [0] && \arg0_4_2Dcon_$fNumInt_$c+_1_d [0])};
  assign \arg0_4_2Dcon_$fNumInt_$c+_1_r  = (\arg0_4_2Dcon_$fNumInt_$c+_1I#_r  && (\arg0_4_2Dcon_$fNumInt_$c+_2_d [0] && \arg0_4_2Dcon_$fNumInt_$c+_1_d [0]));
  assign \arg0_4_2Dcon_$fNumInt_$c+_2_r  = (\arg0_4_2Dcon_$fNumInt_$c+_1I#_r  && (\arg0_4_2Dcon_$fNumInt_$c+_2_d [0] && \arg0_4_2Dcon_$fNumInt_$c+_1_d [0]));
  
  /* demux (Ty Int,
       Ty Int) : (arg0_4_2Dcon_$fNumInt_$c+_3,Int) (arg0_4_1Dcon_$fNumInt_$c+,Int) > [(arg0_4_2Dcon_$fNumInt_$c+_3I#,Int)] */
  assign \arg0_4_2Dcon_$fNumInt_$c+_3I#_d  = {\arg0_4_1Dcon_$fNumInt_$c+_d [32:1],
                                              (\arg0_4_2Dcon_$fNumInt_$c+_3_d [0] && \arg0_4_1Dcon_$fNumInt_$c+_d [0])};
  assign \arg0_4_1Dcon_$fNumInt_$c+_r  = (\arg0_4_2Dcon_$fNumInt_$c+_3I#_r  && (\arg0_4_2Dcon_$fNumInt_$c+_3_d [0] && \arg0_4_1Dcon_$fNumInt_$c+_d [0]));
  assign \arg0_4_2Dcon_$fNumInt_$c+_3_r  = (\arg0_4_2Dcon_$fNumInt_$c+_3I#_r  && (\arg0_4_2Dcon_$fNumInt_$c+_3_d [0] && \arg0_4_1Dcon_$fNumInt_$c+_d [0]));
  
  /* fork (Ty Int) : (arg0_4_2Dcon_$fNumInt_$c+_3I#,Int) > [(arg0_4_2Dcon_$fNumInt_$c+_3I#_1,Int),
                                                       (arg0_4_2Dcon_$fNumInt_$c+_3I#_2,Int),
                                                       (arg0_4_2Dcon_$fNumInt_$c+_3I#_3,Int),
                                                       (arg0_4_2Dcon_$fNumInt_$c+_3I#_4,Int)] */
  logic [3:0] \arg0_4_2Dcon_$fNumInt_$c+_3I#_emitted ;
  logic [3:0] \arg0_4_2Dcon_$fNumInt_$c+_3I#_done ;
  assign \arg0_4_2Dcon_$fNumInt_$c+_3I#_1_d  = {\arg0_4_2Dcon_$fNumInt_$c+_3I#_d [32:1],
                                                (\arg0_4_2Dcon_$fNumInt_$c+_3I#_d [0] && (! \arg0_4_2Dcon_$fNumInt_$c+_3I#_emitted [0]))};
  assign \arg0_4_2Dcon_$fNumInt_$c+_3I#_2_d  = {\arg0_4_2Dcon_$fNumInt_$c+_3I#_d [32:1],
                                                (\arg0_4_2Dcon_$fNumInt_$c+_3I#_d [0] && (! \arg0_4_2Dcon_$fNumInt_$c+_3I#_emitted [1]))};
  assign \arg0_4_2Dcon_$fNumInt_$c+_3I#_3_d  = {\arg0_4_2Dcon_$fNumInt_$c+_3I#_d [32:1],
                                                (\arg0_4_2Dcon_$fNumInt_$c+_3I#_d [0] && (! \arg0_4_2Dcon_$fNumInt_$c+_3I#_emitted [2]))};
  assign \arg0_4_2Dcon_$fNumInt_$c+_3I#_4_d  = {\arg0_4_2Dcon_$fNumInt_$c+_3I#_d [32:1],
                                                (\arg0_4_2Dcon_$fNumInt_$c+_3I#_d [0] && (! \arg0_4_2Dcon_$fNumInt_$c+_3I#_emitted [3]))};
  assign \arg0_4_2Dcon_$fNumInt_$c+_3I#_done  = (\arg0_4_2Dcon_$fNumInt_$c+_3I#_emitted  | ({\arg0_4_2Dcon_$fNumInt_$c+_3I#_4_d [0],
                                                                                             \arg0_4_2Dcon_$fNumInt_$c+_3I#_3_d [0],
                                                                                             \arg0_4_2Dcon_$fNumInt_$c+_3I#_2_d [0],
                                                                                             \arg0_4_2Dcon_$fNumInt_$c+_3I#_1_d [0]} & {\arg0_4_2Dcon_$fNumInt_$c+_3I#_4_r ,
                                                                                                                                        \arg0_4_2Dcon_$fNumInt_$c+_3I#_3_r ,
                                                                                                                                        \arg0_4_2Dcon_$fNumInt_$c+_3I#_2_r ,
                                                                                                                                        \arg0_4_2Dcon_$fNumInt_$c+_3I#_1_r }));
  assign \arg0_4_2Dcon_$fNumInt_$c+_3I#_r  = (& \arg0_4_2Dcon_$fNumInt_$c+_3I#_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \arg0_4_2Dcon_$fNumInt_$c+_3I#_emitted  <= 4'd0;
    else
      \arg0_4_2Dcon_$fNumInt_$c+_3I#_emitted  <= (\arg0_4_2Dcon_$fNumInt_$c+_3I#_r  ? 4'd0 :
                                                  \arg0_4_2Dcon_$fNumInt_$c+_3I#_done );
  
  /* destruct (Ty Int,
          Dcon I#) : (arg0_4_2Dcon_$fNumInt_$c+_3I#_1I#,Int) > [(ya1lW_destruct,Int#)] */
  assign ya1lW_destruct_d = {\arg0_4_2Dcon_$fNumInt_$c+_3I#_1I#_d [32:1],
                             \arg0_4_2Dcon_$fNumInt_$c+_3I#_1I#_d [0]};
  assign \arg0_4_2Dcon_$fNumInt_$c+_3I#_1I#_r  = ya1lW_destruct_r;
  
  /* demux (Ty Int,
       Ty Int) : (arg0_4_2Dcon_$fNumInt_$c+_3I#_2,Int) (arg0_4_2Dcon_$fNumInt_$c+_3I#_1,Int) > [(arg0_4_2Dcon_$fNumInt_$c+_3I#_1I#,Int)] */
  assign \arg0_4_2Dcon_$fNumInt_$c+_3I#_1I#_d  = {\arg0_4_2Dcon_$fNumInt_$c+_3I#_1_d [32:1],
                                                  (\arg0_4_2Dcon_$fNumInt_$c+_3I#_2_d [0] && \arg0_4_2Dcon_$fNumInt_$c+_3I#_1_d [0])};
  assign \arg0_4_2Dcon_$fNumInt_$c+_3I#_1_r  = (\arg0_4_2Dcon_$fNumInt_$c+_3I#_1I#_r  && (\arg0_4_2Dcon_$fNumInt_$c+_3I#_2_d [0] && \arg0_4_2Dcon_$fNumInt_$c+_3I#_1_d [0]));
  assign \arg0_4_2Dcon_$fNumInt_$c+_3I#_2_r  = (\arg0_4_2Dcon_$fNumInt_$c+_3I#_1I#_r  && (\arg0_4_2Dcon_$fNumInt_$c+_3I#_2_d [0] && \arg0_4_2Dcon_$fNumInt_$c+_3I#_1_d [0]));
  
  /* demux (Ty Int,
       Ty Int#) : (arg0_4_2Dcon_$fNumInt_$c+_3I#_3,Int) (xa1lV_destruct,Int#) > [(arg0_4_2Dcon_$fNumInt_$c+_3I#_3I#,Int#)] */
  assign \arg0_4_2Dcon_$fNumInt_$c+_3I#_3I#_d  = {xa1lV_destruct_d[32:1],
                                                  (\arg0_4_2Dcon_$fNumInt_$c+_3I#_3_d [0] && xa1lV_destruct_d[0])};
  assign xa1lV_destruct_r = (\arg0_4_2Dcon_$fNumInt_$c+_3I#_3I#_r  && (\arg0_4_2Dcon_$fNumInt_$c+_3I#_3_d [0] && xa1lV_destruct_d[0]));
  assign \arg0_4_2Dcon_$fNumInt_$c+_3I#_3_r  = (\arg0_4_2Dcon_$fNumInt_$c+_3I#_3I#_r  && (\arg0_4_2Dcon_$fNumInt_$c+_3I#_3_d [0] && xa1lV_destruct_d[0]));
  
  /* op_add (Ty Int#) : (arg0_4_2Dcon_$fNumInt_$c+_3I#_3I#,Int#) (ya1lW_destruct,Int#) > (arg0_4_2Dcon_$fNumInt_$c+_3I#_3I#_1ya1lW_1_Add32,Int#) */
  assign \arg0_4_2Dcon_$fNumInt_$c+_3I#_3I#_1ya1lW_1_Add32_d  = {(\arg0_4_2Dcon_$fNumInt_$c+_3I#_3I#_d [32:1] + ya1lW_destruct_d[32:1]),
                                                                 (\arg0_4_2Dcon_$fNumInt_$c+_3I#_3I#_d [0] && ya1lW_destruct_d[0])};
  assign {\arg0_4_2Dcon_$fNumInt_$c+_3I#_3I#_r ,
          ya1lW_destruct_r} = {2 {(\arg0_4_2Dcon_$fNumInt_$c+_3I#_3I#_1ya1lW_1_Add32_r  && \arg0_4_2Dcon_$fNumInt_$c+_3I#_3I#_1ya1lW_1_Add32_d [0])}};
  
  /* dcon (Ty Int,
      Dcon I#) : [(arg0_4_2Dcon_$fNumInt_$c+_3I#_3I#_1ya1lW_1_Add32,Int#)] > (es_0_2_1I#,Int) */
  assign \es_0_2_1I#_d  = \I#_dc ((& {\arg0_4_2Dcon_$fNumInt_$c+_3I#_3I#_1ya1lW_1_Add32_d [0]}), \arg0_4_2Dcon_$fNumInt_$c+_3I#_3I#_1ya1lW_1_Add32_d );
  assign {\arg0_4_2Dcon_$fNumInt_$c+_3I#_3I#_1ya1lW_1_Add32_r } = {1 {(\es_0_2_1I#_r  && \es_0_2_1I#_d [0])}};
  
  /* mux (Ty Int,
     Ty Int) : (arg0_4_2Dcon_$fNumInt_$c+_3I#_4,Int) [(es_0_2_1I#,Int)] > (es_0_2_1I#_mux,Int) */
  assign \es_0_2_1I#_mux_d  = {\es_0_2_1I#_d [32:1],
                               (\arg0_4_2Dcon_$fNumInt_$c+_3I#_4_d [0] && \es_0_2_1I#_d [0])};
  assign \es_0_2_1I#_r  = (\es_0_2_1I#_mux_r  && (\arg0_4_2Dcon_$fNumInt_$c+_3I#_4_d [0] && \es_0_2_1I#_d [0]));
  assign \arg0_4_2Dcon_$fNumInt_$c+_3I#_4_r  = (\es_0_2_1I#_mux_r  && (\arg0_4_2Dcon_$fNumInt_$c+_3I#_4_d [0] && \es_0_2_1I#_d [0]));
  
  /* mux (Ty Int,
     Ty Int) : (arg0_4_2Dcon_$fNumInt_$c+_4,Int) [(es_0_2_1I#_mux,Int)] > (es_0_2_1I#_mux_mux,Int) */
  assign \es_0_2_1I#_mux_mux_d  = {\es_0_2_1I#_mux_d [32:1],
                                   (\arg0_4_2Dcon_$fNumInt_$c+_4_d [0] && \es_0_2_1I#_mux_d [0])};
  assign \es_0_2_1I#_mux_r  = (\es_0_2_1I#_mux_mux_r  && (\arg0_4_2Dcon_$fNumInt_$c+_4_d [0] && \es_0_2_1I#_mux_d [0]));
  assign \arg0_4_2Dcon_$fNumInt_$c+_4_r  = (\es_0_2_1I#_mux_mux_r  && (\arg0_4_2Dcon_$fNumInt_$c+_4_d [0] && \es_0_2_1I#_mux_d [0]));
  
  /* mux (Ty MyDTInt_Int_Int,
     Ty Int) : (arg0_4_3,MyDTInt_Int_Int) [(es_0_2_1I#_mux_mux,Int)] > (es_0_2_1I#_mux_mux_mux,Int) */
  assign \es_0_2_1I#_mux_mux_mux_d  = {\es_0_2_1I#_mux_mux_d [32:1],
                                       (arg0_4_3_d[0] && \es_0_2_1I#_mux_mux_d [0])};
  assign \es_0_2_1I#_mux_mux_r  = (\es_0_2_1I#_mux_mux_mux_r  && (arg0_4_3_d[0] && \es_0_2_1I#_mux_mux_d [0]));
  assign arg0_4_3_r = (\es_0_2_1I#_mux_mux_mux_r  && (arg0_4_3_d[0] && \es_0_2_1I#_mux_mux_d [0]));
  
  /* buf (Ty Pointer_QTree_Int) : (bla8A_1_destruct,Pointer_QTree_Int) > (bla8A_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t bla8A_1_destruct_bufchan_d;
  logic bla8A_1_destruct_bufchan_r;
  assign bla8A_1_destruct_r = ((! bla8A_1_destruct_bufchan_d[0]) || bla8A_1_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) bla8A_1_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (bla8A_1_destruct_r)
        bla8A_1_destruct_bufchan_d <= bla8A_1_destruct_d;
  Pointer_QTree_Int_t bla8A_1_destruct_bufchan_buf;
  assign bla8A_1_destruct_bufchan_r = (! bla8A_1_destruct_bufchan_buf[0]);
  assign bla8A_1_1_argbuf_d = (bla8A_1_destruct_bufchan_buf[0] ? bla8A_1_destruct_bufchan_buf :
                               bla8A_1_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) bla8A_1_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((bla8A_1_1_argbuf_r && bla8A_1_destruct_bufchan_buf[0]))
        bla8A_1_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! bla8A_1_1_argbuf_r) && (! bla8A_1_destruct_bufchan_buf[0])))
        bla8A_1_destruct_bufchan_buf <= bla8A_1_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (bla8L_destruct,Pointer_QTree_Int) > (bla8L_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t bla8L_destruct_bufchan_d;
  logic bla8L_destruct_bufchan_r;
  assign bla8L_destruct_r = ((! bla8L_destruct_bufchan_d[0]) || bla8L_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) bla8L_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (bla8L_destruct_r) bla8L_destruct_bufchan_d <= bla8L_destruct_d;
  Pointer_QTree_Int_t bla8L_destruct_bufchan_buf;
  assign bla8L_destruct_bufchan_r = (! bla8L_destruct_bufchan_buf[0]);
  assign bla8L_1_argbuf_d = (bla8L_destruct_bufchan_buf[0] ? bla8L_destruct_bufchan_buf :
                             bla8L_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) bla8L_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((bla8L_1_argbuf_r && bla8L_destruct_bufchan_buf[0]))
        bla8L_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! bla8L_1_argbuf_r) && (! bla8L_destruct_bufchan_buf[0])))
        bla8L_destruct_bufchan_buf <= bla8L_destruct_bufchan_d;
  
  /* destruct (Ty TupGo___Bool,
          Dcon TupGo___Bool) : (boolConvert_1TupGo___Bool_1,TupGo___Bool) > [(boolConvert_1TupGo___Boolgo_1,Go),
                                                                             (boolConvert_1TupGo___Boolbool,Bool)] */
  logic [1:0] boolConvert_1TupGo___Bool_1_emitted;
  logic [1:0] boolConvert_1TupGo___Bool_1_done;
  assign boolConvert_1TupGo___Boolgo_1_d = (boolConvert_1TupGo___Bool_1_d[0] && (! boolConvert_1TupGo___Bool_1_emitted[0]));
  assign boolConvert_1TupGo___Boolbool_d = {boolConvert_1TupGo___Bool_1_d[1:1],
                                            (boolConvert_1TupGo___Bool_1_d[0] && (! boolConvert_1TupGo___Bool_1_emitted[1]))};
  assign boolConvert_1TupGo___Bool_1_done = (boolConvert_1TupGo___Bool_1_emitted | ({boolConvert_1TupGo___Boolbool_d[0],
                                                                                     boolConvert_1TupGo___Boolgo_1_d[0]} & {boolConvert_1TupGo___Boolbool_r,
                                                                                                                            boolConvert_1TupGo___Boolgo_1_r}));
  assign boolConvert_1TupGo___Bool_1_r = (& boolConvert_1TupGo___Bool_1_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) boolConvert_1TupGo___Bool_1_emitted <= 2'd0;
    else
      boolConvert_1TupGo___Bool_1_emitted <= (boolConvert_1TupGo___Bool_1_r ? 2'd0 :
                                              boolConvert_1TupGo___Bool_1_done);
  
  /* fork (Ty Bool) : (boolConvert_1TupGo___Boolbool,Bool) > [(bool_1,Bool),
                                                         (bool_2,Bool)] */
  logic [1:0] boolConvert_1TupGo___Boolbool_emitted;
  logic [1:0] boolConvert_1TupGo___Boolbool_done;
  assign bool_1_d = {boolConvert_1TupGo___Boolbool_d[1:1],
                     (boolConvert_1TupGo___Boolbool_d[0] && (! boolConvert_1TupGo___Boolbool_emitted[0]))};
  assign bool_2_d = {boolConvert_1TupGo___Boolbool_d[1:1],
                     (boolConvert_1TupGo___Boolbool_d[0] && (! boolConvert_1TupGo___Boolbool_emitted[1]))};
  assign boolConvert_1TupGo___Boolbool_done = (boolConvert_1TupGo___Boolbool_emitted | ({bool_2_d[0],
                                                                                         bool_1_d[0]} & {bool_2_r,
                                                                                                         bool_1_r}));
  assign boolConvert_1TupGo___Boolbool_r = (& boolConvert_1TupGo___Boolbool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) boolConvert_1TupGo___Boolbool_emitted <= 2'd0;
    else
      boolConvert_1TupGo___Boolbool_emitted <= (boolConvert_1TupGo___Boolbool_r ? 2'd0 :
                                                boolConvert_1TupGo___Boolbool_done);
  
  /* fork (Ty MyBool) : (boolConvert_1_resbuf,MyBool) > [(lizzieLet3_1,MyBool),
                                                    (lizzieLet3_2,MyBool)] */
  logic [1:0] boolConvert_1_resbuf_emitted;
  logic [1:0] boolConvert_1_resbuf_done;
  assign lizzieLet3_1_d = {boolConvert_1_resbuf_d[1:1],
                           (boolConvert_1_resbuf_d[0] && (! boolConvert_1_resbuf_emitted[0]))};
  assign lizzieLet3_2_d = {boolConvert_1_resbuf_d[1:1],
                           (boolConvert_1_resbuf_d[0] && (! boolConvert_1_resbuf_emitted[1]))};
  assign boolConvert_1_resbuf_done = (boolConvert_1_resbuf_emitted | ({lizzieLet3_2_d[0],
                                                                       lizzieLet3_1_d[0]} & {lizzieLet3_2_r,
                                                                                             lizzieLet3_1_r}));
  assign boolConvert_1_resbuf_r = (& boolConvert_1_resbuf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) boolConvert_1_resbuf_emitted <= 2'd0;
    else
      boolConvert_1_resbuf_emitted <= (boolConvert_1_resbuf_r ? 2'd0 :
                                       boolConvert_1_resbuf_done);
  
  /* demux (Ty Bool,
       Ty Go) : (bool_1,Bool) (boolConvert_1TupGo___Boolgo_1,Go) > [(bool_1False,Go),
                                                                    (bool_1True,Go)] */
  logic [1:0] boolConvert_1TupGo___Boolgo_1_onehotd;
  always_comb
    if ((bool_1_d[0] && boolConvert_1TupGo___Boolgo_1_d[0]))
      unique case (bool_1_d[1:1])
        1'd0: boolConvert_1TupGo___Boolgo_1_onehotd = 2'd1;
        1'd1: boolConvert_1TupGo___Boolgo_1_onehotd = 2'd2;
        default: boolConvert_1TupGo___Boolgo_1_onehotd = 2'd0;
      endcase
    else boolConvert_1TupGo___Boolgo_1_onehotd = 2'd0;
  assign bool_1False_d = boolConvert_1TupGo___Boolgo_1_onehotd[0];
  assign bool_1True_d = boolConvert_1TupGo___Boolgo_1_onehotd[1];
  assign boolConvert_1TupGo___Boolgo_1_r = (| (boolConvert_1TupGo___Boolgo_1_onehotd & {bool_1True_r,
                                                                                        bool_1False_r}));
  assign bool_1_r = boolConvert_1TupGo___Boolgo_1_r;
  
  /* dcon (Ty MyBool,
      Dcon MyFalse) : [(bool_1False,Go)] > (bool_1False_1MyFalse,MyBool) */
  assign bool_1False_1MyFalse_d = MyFalse_dc((& {bool_1False_d[0]}), bool_1False_d);
  assign {bool_1False_r} = {1 {(bool_1False_1MyFalse_r && bool_1False_1MyFalse_d[0])}};
  
  /* buf (Ty MyBool) : (bool_1False_1MyFalsebool_1True_1MyTrue_mux,MyBool) > (boolConvert_1_resbuf,MyBool) */
  MyBool_t bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_d;
  logic bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_r;
  assign bool_1False_1MyFalsebool_1True_1MyTrue_mux_r = ((! bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_d[0]) || bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_d <= {1'd0,
                                                               1'd0};
    else
      if (bool_1False_1MyFalsebool_1True_1MyTrue_mux_r)
        bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_d <= bool_1False_1MyFalsebool_1True_1MyTrue_mux_d;
  MyBool_t bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_buf;
  assign bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_r = (! bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_buf[0]);
  assign boolConvert_1_resbuf_d = (bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_buf[0] ? bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_buf :
                                   bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_buf <= {1'd0,
                                                                 1'd0};
    else
      if ((boolConvert_1_resbuf_r && bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_buf[0]))
        bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_buf <= {1'd0,
                                                                   1'd0};
      else if (((! boolConvert_1_resbuf_r) && (! bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_buf[0])))
        bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_buf <= bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_d;
  
  /* dcon (Ty MyBool,
      Dcon MyTrue) : [(bool_1True,Go)] > (bool_1True_1MyTrue,MyBool) */
  assign bool_1True_1MyTrue_d = MyTrue_dc((& {bool_1True_d[0]}), bool_1True_d);
  assign {bool_1True_r} = {1 {(bool_1True_1MyTrue_r && bool_1True_1MyTrue_d[0])}};
  
  /* mux (Ty Bool,
     Ty MyBool) : (bool_2,Bool) [(bool_1False_1MyFalse,MyBool),
                                 (bool_1True_1MyTrue,MyBool)] > (bool_1False_1MyFalsebool_1True_1MyTrue_mux,MyBool) */
  logic [1:0] bool_1False_1MyFalsebool_1True_1MyTrue_mux_mux;
  logic [1:0] bool_1False_1MyFalsebool_1True_1MyTrue_mux_onehot;
  always_comb
    unique case (bool_2_d[1:1])
      1'd0:
        {bool_1False_1MyFalsebool_1True_1MyTrue_mux_onehot,
         bool_1False_1MyFalsebool_1True_1MyTrue_mux_mux} = {2'd1,
                                                            bool_1False_1MyFalse_d};
      1'd1:
        {bool_1False_1MyFalsebool_1True_1MyTrue_mux_onehot,
         bool_1False_1MyFalsebool_1True_1MyTrue_mux_mux} = {2'd2,
                                                            bool_1True_1MyTrue_d};
      default:
        {bool_1False_1MyFalsebool_1True_1MyTrue_mux_onehot,
         bool_1False_1MyFalsebool_1True_1MyTrue_mux_mux} = {2'd0,
                                                            {1'd0, 1'd0}};
    endcase
  assign bool_1False_1MyFalsebool_1True_1MyTrue_mux_d = {bool_1False_1MyFalsebool_1True_1MyTrue_mux_mux[1:1],
                                                         (bool_1False_1MyFalsebool_1True_1MyTrue_mux_mux[0] && bool_2_d[0])};
  assign bool_2_r = (bool_1False_1MyFalsebool_1True_1MyTrue_mux_d[0] && bool_1False_1MyFalsebool_1True_1MyTrue_mux_r);
  assign {bool_1True_1MyTrue_r,
          bool_1False_1MyFalse_r} = (bool_2_r ? bool_1False_1MyFalsebool_1True_1MyTrue_mux_onehot :
                                     2'd0);
  
  /* buf (Ty Pointer_QTree_Int) : (bra8B_destruct,Pointer_QTree_Int) > (bra8B_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t bra8B_destruct_bufchan_d;
  logic bra8B_destruct_bufchan_r;
  assign bra8B_destruct_r = ((! bra8B_destruct_bufchan_d[0]) || bra8B_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) bra8B_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (bra8B_destruct_r) bra8B_destruct_bufchan_d <= bra8B_destruct_d;
  Pointer_QTree_Int_t bra8B_destruct_bufchan_buf;
  assign bra8B_destruct_bufchan_r = (! bra8B_destruct_bufchan_buf[0]);
  assign bra8B_1_argbuf_d = (bra8B_destruct_bufchan_buf[0] ? bra8B_destruct_bufchan_buf :
                             bra8B_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) bra8B_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((bra8B_1_argbuf_r && bra8B_destruct_bufchan_buf[0]))
        bra8B_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! bra8B_1_argbuf_r) && (! bra8B_destruct_bufchan_buf[0])))
        bra8B_destruct_bufchan_buf <= bra8B_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (bra8M_destruct,Pointer_QTree_Int) > (bra8M_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t bra8M_destruct_bufchan_d;
  logic bra8M_destruct_bufchan_r;
  assign bra8M_destruct_r = ((! bra8M_destruct_bufchan_d[0]) || bra8M_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) bra8M_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (bra8M_destruct_r) bra8M_destruct_bufchan_d <= bra8M_destruct_d;
  Pointer_QTree_Int_t bra8M_destruct_bufchan_buf;
  assign bra8M_destruct_bufchan_r = (! bra8M_destruct_bufchan_buf[0]);
  assign bra8M_1_argbuf_d = (bra8M_destruct_bufchan_buf[0] ? bra8M_destruct_bufchan_buf :
                             bra8M_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) bra8M_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((bra8M_1_argbuf_r && bra8M_destruct_bufchan_buf[0]))
        bra8M_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! bra8M_1_argbuf_r) && (! bra8M_destruct_bufchan_buf[0])))
        bra8M_destruct_bufchan_buf <= bra8M_destruct_bufchan_d;
  
  /* destruct (Ty TupGo___Pointer_QTree_Int___Pointer_CT$wnnz,
          Dcon TupGo___Pointer_QTree_Int___Pointer_CT$wnnz) : (call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_1,TupGo___Pointer_QTree_Int___Pointer_CT$wnnz) > [(call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnzgo_10,Go),
                                                                                                                                                                       (call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnzwsiX_1,Pointer_QTree_Int),
                                                                                                                                                                       (call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnzsc_0,Pointer_CT$wnnz)] */
  logic [2:0] call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_1_emitted;
  logic [2:0] call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_1_done;
  assign call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnzgo_10_d = (call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_1_d[0] && (! call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_1_emitted[0]));
  assign call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnzwsiX_1_d = {call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_1_d[16:1],
                                                                          (call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_1_d[0] && (! call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_1_emitted[1]))};
  assign call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnzsc_0_d = {call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_1_d[32:17],
                                                                        (call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_1_d[0] && (! call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_1_emitted[2]))};
  assign call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_1_done = (call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_1_emitted | ({call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnzsc_0_d[0],
                                                                                                                                             call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnzwsiX_1_d[0],
                                                                                                                                             call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnzgo_10_d[0]} & {call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnzsc_0_r,
                                                                                                                                                                                                                 call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnzwsiX_1_r,
                                                                                                                                                                                                                 call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnzgo_10_r}));
  assign call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_1_r = (& call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_1_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_1_emitted <= 3'd0;
    else
      call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_1_emitted <= (call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_1_r ? 3'd0 :
                                                                          call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_1_done);
  
  /* rbuf (Ty Go) : (call_$wnnz_goConst,Go) > (call_$wnnz_initBufi,Go) */
  Go_t call_$wnnz_goConst_buf;
  assign call_$wnnz_goConst_r = (! call_$wnnz_goConst_buf[0]);
  assign call_$wnnz_initBufi_d = (call_$wnnz_goConst_buf[0] ? call_$wnnz_goConst_buf :
                                  call_$wnnz_goConst_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_$wnnz_goConst_buf <= 1'd0;
    else
      if ((call_$wnnz_initBufi_r && call_$wnnz_goConst_buf[0]))
        call_$wnnz_goConst_buf <= 1'd0;
      else if (((! call_$wnnz_initBufi_r) && (! call_$wnnz_goConst_buf[0])))
        call_$wnnz_goConst_buf <= call_$wnnz_goConst_d;
  
  /* mergectrl (Ty C5,Ty Go) : [(call_$wnnz_goMux1,Go),
                           (lizzieLet35_3Lcall_$wnnz3_1_argbuf,Go),
                           (lizzieLet35_3Lcall_$wnnz2_1_argbuf,Go),
                           (lizzieLet35_3Lcall_$wnnz1_1_argbuf,Go),
                           (lizzieLet4_3QNode_Int_1_argbuf,Go)] > (go_10_goMux_choice,C5) (go_10_goMux_data,Go) */
  logic [4:0] call_$wnnz_goMux1_select_d;
  assign call_$wnnz_goMux1_select_d = ((| call_$wnnz_goMux1_select_q) ? call_$wnnz_goMux1_select_q :
                                       (call_$wnnz_goMux1_d[0] ? 5'd1 :
                                        (lizzieLet35_3Lcall_$wnnz3_1_argbuf_d[0] ? 5'd2 :
                                         (lizzieLet35_3Lcall_$wnnz2_1_argbuf_d[0] ? 5'd4 :
                                          (lizzieLet35_3Lcall_$wnnz1_1_argbuf_d[0] ? 5'd8 :
                                           (lizzieLet4_3QNode_Int_1_argbuf_d[0] ? 5'd16 :
                                            5'd0))))));
  logic [4:0] call_$wnnz_goMux1_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_$wnnz_goMux1_select_q <= 5'd0;
    else
      call_$wnnz_goMux1_select_q <= (call_$wnnz_goMux1_done ? 5'd0 :
                                     call_$wnnz_goMux1_select_d);
  logic [1:0] call_$wnnz_goMux1_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_$wnnz_goMux1_emit_q <= 2'd0;
    else
      call_$wnnz_goMux1_emit_q <= (call_$wnnz_goMux1_done ? 2'd0 :
                                   call_$wnnz_goMux1_emit_d);
  logic [1:0] call_$wnnz_goMux1_emit_d;
  assign call_$wnnz_goMux1_emit_d = (call_$wnnz_goMux1_emit_q | ({go_10_goMux_choice_d[0],
                                                                  go_10_goMux_data_d[0]} & {go_10_goMux_choice_r,
                                                                                            go_10_goMux_data_r}));
  logic call_$wnnz_goMux1_done;
  assign call_$wnnz_goMux1_done = (& call_$wnnz_goMux1_emit_d);
  assign {lizzieLet4_3QNode_Int_1_argbuf_r,
          lizzieLet35_3Lcall_$wnnz1_1_argbuf_r,
          lizzieLet35_3Lcall_$wnnz2_1_argbuf_r,
          lizzieLet35_3Lcall_$wnnz3_1_argbuf_r,
          call_$wnnz_goMux1_r} = (call_$wnnz_goMux1_done ? call_$wnnz_goMux1_select_d :
                                  5'd0);
  assign go_10_goMux_data_d = ((call_$wnnz_goMux1_select_d[0] && (! call_$wnnz_goMux1_emit_q[0])) ? call_$wnnz_goMux1_d :
                               ((call_$wnnz_goMux1_select_d[1] && (! call_$wnnz_goMux1_emit_q[0])) ? lizzieLet35_3Lcall_$wnnz3_1_argbuf_d :
                                ((call_$wnnz_goMux1_select_d[2] && (! call_$wnnz_goMux1_emit_q[0])) ? lizzieLet35_3Lcall_$wnnz2_1_argbuf_d :
                                 ((call_$wnnz_goMux1_select_d[3] && (! call_$wnnz_goMux1_emit_q[0])) ? lizzieLet35_3Lcall_$wnnz1_1_argbuf_d :
                                  ((call_$wnnz_goMux1_select_d[4] && (! call_$wnnz_goMux1_emit_q[0])) ? lizzieLet4_3QNode_Int_1_argbuf_d :
                                   1'd0)))));
  assign go_10_goMux_choice_d = ((call_$wnnz_goMux1_select_d[0] && (! call_$wnnz_goMux1_emit_q[1])) ? C1_5_dc(1'd1) :
                                 ((call_$wnnz_goMux1_select_d[1] && (! call_$wnnz_goMux1_emit_q[1])) ? C2_5_dc(1'd1) :
                                  ((call_$wnnz_goMux1_select_d[2] && (! call_$wnnz_goMux1_emit_q[1])) ? C3_5_dc(1'd1) :
                                   ((call_$wnnz_goMux1_select_d[3] && (! call_$wnnz_goMux1_emit_q[1])) ? C4_5_dc(1'd1) :
                                    ((call_$wnnz_goMux1_select_d[4] && (! call_$wnnz_goMux1_emit_q[1])) ? C5_5_dc(1'd1) :
                                     {3'd0, 1'd0})))));
  
  /* fork (Ty Go) : (call_$wnnz_initBuf,Go) > [(call_$wnnz_unlockFork1,Go),
                                          (call_$wnnz_unlockFork2,Go),
                                          (call_$wnnz_unlockFork3,Go)] */
  logic [2:0] call_$wnnz_initBuf_emitted;
  logic [2:0] call_$wnnz_initBuf_done;
  assign call_$wnnz_unlockFork1_d = (call_$wnnz_initBuf_d[0] && (! call_$wnnz_initBuf_emitted[0]));
  assign call_$wnnz_unlockFork2_d = (call_$wnnz_initBuf_d[0] && (! call_$wnnz_initBuf_emitted[1]));
  assign call_$wnnz_unlockFork3_d = (call_$wnnz_initBuf_d[0] && (! call_$wnnz_initBuf_emitted[2]));
  assign call_$wnnz_initBuf_done = (call_$wnnz_initBuf_emitted | ({call_$wnnz_unlockFork3_d[0],
                                                                   call_$wnnz_unlockFork2_d[0],
                                                                   call_$wnnz_unlockFork1_d[0]} & {call_$wnnz_unlockFork3_r,
                                                                                                   call_$wnnz_unlockFork2_r,
                                                                                                   call_$wnnz_unlockFork1_r}));
  assign call_$wnnz_initBuf_r = (& call_$wnnz_initBuf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_$wnnz_initBuf_emitted <= 3'd0;
    else
      call_$wnnz_initBuf_emitted <= (call_$wnnz_initBuf_r ? 3'd0 :
                                     call_$wnnz_initBuf_done);
  
  /* initbuf (Ty Go,
         Dcon Go) : (call_$wnnz_initBufi,Go) > (call_$wnnz_initBuf,Go) */
  assign call_$wnnz_initBufi_r = ((! call_$wnnz_initBuf_d[0]) || call_$wnnz_initBuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_$wnnz_initBuf_d <= Go_dc(1'd1);
    else
      if (call_$wnnz_initBufi_r)
        call_$wnnz_initBuf_d <= call_$wnnz_initBufi_d;
  
  /* mux (Ty Go,
     Ty Go) : (call_$wnnz_unlockFork1,Go) [(call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnzgo_10,Go)] > (call_$wnnz_goMux1,Go) */
  assign call_$wnnz_goMux1_d = (call_$wnnz_unlockFork1_d[0] && call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnzgo_10_d[0]);
  assign call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnzgo_10_r = (call_$wnnz_goMux1_r && (call_$wnnz_unlockFork1_d[0] && call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnzgo_10_d[0]));
  assign call_$wnnz_unlockFork1_r = (call_$wnnz_goMux1_r && (call_$wnnz_unlockFork1_d[0] && call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnzgo_10_d[0]));
  
  /* mux (Ty Go,
     Ty Pointer_QTree_Int) : (call_$wnnz_unlockFork2,Go) [(call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnzwsiX_1,Pointer_QTree_Int)] > (call_$wnnz_goMux2,Pointer_QTree_Int) */
  assign call_$wnnz_goMux2_d = {call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnzwsiX_1_d[16:1],
                                (call_$wnnz_unlockFork2_d[0] && call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnzwsiX_1_d[0])};
  assign call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnzwsiX_1_r = (call_$wnnz_goMux2_r && (call_$wnnz_unlockFork2_d[0] && call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnzwsiX_1_d[0]));
  assign call_$wnnz_unlockFork2_r = (call_$wnnz_goMux2_r && (call_$wnnz_unlockFork2_d[0] && call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnzwsiX_1_d[0]));
  
  /* mux (Ty Go,
     Ty Pointer_CT$wnnz) : (call_$wnnz_unlockFork3,Go) [(call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnzsc_0,Pointer_CT$wnnz)] > (call_$wnnz_goMux3,Pointer_CT$wnnz) */
  assign call_$wnnz_goMux3_d = {call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnzsc_0_d[16:1],
                                (call_$wnnz_unlockFork3_d[0] && call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnzsc_0_d[0])};
  assign call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnzsc_0_r = (call_$wnnz_goMux3_r && (call_$wnnz_unlockFork3_d[0] && call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnzsc_0_d[0]));
  assign call_$wnnz_unlockFork3_r = (call_$wnnz_goMux3_r && (call_$wnnz_unlockFork3_d[0] && call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnzsc_0_d[0]));
  
  /* destruct (Ty TupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf''''''''_f''''''''_Int_Int,
          Dcon TupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf''''''''_f''''''''_Int_Int) : (call_f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf''''''''_f''''''''_Int_Int_1,TupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf''''''''_f''''''''_Int_Int) > [(call_f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf''''''''_f''''''''_Int_Intgo_11,Go),
                                                                                                                                                                                                                                                                                                                                                      (call_f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf''''''''_f''''''''_Int_Intq4a8u,Pointer_QTree_Int),
                                                                                                                                                                                                                                                                                                                                                      (call_f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf''''''''_f''''''''_Int_Intis_z_mapa8v,MyDTInt_Bool),
                                                                                                                                                                                                                                                                                                                                                      (call_f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf''''''''_f''''''''_Int_Intop_mapa8w,MyDTInt_Int),
                                                                                                                                                                                                                                                                                                                                                      (call_f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf''''''''_f''''''''_Int_Intsc_0_1,Pointer_CTf''''''''_f''''''''_Int_Int)] */
  logic [4:0] \call_f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf''''''''_f''''''''_Int_Int_1_emitted ;
  logic [4:0] \call_f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf''''''''_f''''''''_Int_Int_1_done ;
  assign \call_f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf''''''''_f''''''''_Int_Intgo_11_d  = (\call_f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf''''''''_f''''''''_Int_Int_1_d [0] && (! \call_f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf''''''''_f''''''''_Int_Int_1_emitted [0]));
  assign \call_f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf''''''''_f''''''''_Int_Intq4a8u_d  = {\call_f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf''''''''_f''''''''_Int_Int_1_d [16:1],
                                                                                                                                                    (\call_f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf''''''''_f''''''''_Int_Int_1_d [0] && (! \call_f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf''''''''_f''''''''_Int_Int_1_emitted [1]))};
  assign \call_f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf''''''''_f''''''''_Int_Intis_z_mapa8v_d  = (\call_f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf''''''''_f''''''''_Int_Int_1_d [0] && (! \call_f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf''''''''_f''''''''_Int_Int_1_emitted [2]));
  assign \call_f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf''''''''_f''''''''_Int_Intop_mapa8w_d  = (\call_f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf''''''''_f''''''''_Int_Int_1_d [0] && (! \call_f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf''''''''_f''''''''_Int_Int_1_emitted [3]));
  assign \call_f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf''''''''_f''''''''_Int_Intsc_0_1_d  = {\call_f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf''''''''_f''''''''_Int_Int_1_d [32:17],
                                                                                                                                                     (\call_f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf''''''''_f''''''''_Int_Int_1_d [0] && (! \call_f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf''''''''_f''''''''_Int_Int_1_emitted [4]))};
  assign \call_f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf''''''''_f''''''''_Int_Int_1_done  = (\call_f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf''''''''_f''''''''_Int_Int_1_emitted  | ({\call_f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf''''''''_f''''''''_Int_Intsc_0_1_d [0],
                                                                                                                                                                                                                                                                                                   \call_f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf''''''''_f''''''''_Int_Intop_mapa8w_d [0],
                                                                                                                                                                                                                                                                                                   \call_f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf''''''''_f''''''''_Int_Intis_z_mapa8v_d [0],
                                                                                                                                                                                                                                                                                                   \call_f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf''''''''_f''''''''_Int_Intq4a8u_d [0],
                                                                                                                                                                                                                                                                                                   \call_f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf''''''''_f''''''''_Int_Intgo_11_d [0]} & {\call_f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf''''''''_f''''''''_Int_Intsc_0_1_r ,
                                                                                                                                                                                                                                                                                                                                                                                                                                                  \call_f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf''''''''_f''''''''_Int_Intop_mapa8w_r ,
                                                                                                                                                                                                                                                                                                                                                                                                                                                  \call_f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf''''''''_f''''''''_Int_Intis_z_mapa8v_r ,
                                                                                                                                                                                                                                                                                                                                                                                                                                                  \call_f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf''''''''_f''''''''_Int_Intq4a8u_r ,
                                                                                                                                                                                                                                                                                                                                                                                                                                                  \call_f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf''''''''_f''''''''_Int_Intgo_11_r }));
  assign \call_f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf''''''''_f''''''''_Int_Int_1_r  = (& \call_f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf''''''''_f''''''''_Int_Int_1_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \call_f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf''''''''_f''''''''_Int_Int_1_emitted  <= 5'd0;
    else
      \call_f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf''''''''_f''''''''_Int_Int_1_emitted  <= (\call_f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf''''''''_f''''''''_Int_Int_1_r  ? 5'd0 :
                                                                                                                                                     \call_f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf''''''''_f''''''''_Int_Int_1_done );
  
  /* rbuf (Ty Go) : (call_f''''''''_f''''''''_Int_Int_goConst,Go) > (call_f''''''''_f''''''''_Int_Int_initBufi,Go) */
  Go_t \call_f''''''''_f''''''''_Int_Int_goConst_buf ;
  assign \call_f''''''''_f''''''''_Int_Int_goConst_r  = (! \call_f''''''''_f''''''''_Int_Int_goConst_buf [0]);
  assign \call_f''''''''_f''''''''_Int_Int_initBufi_d  = (\call_f''''''''_f''''''''_Int_Int_goConst_buf [0] ? \call_f''''''''_f''''''''_Int_Int_goConst_buf  :
                                                          \call_f''''''''_f''''''''_Int_Int_goConst_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \call_f''''''''_f''''''''_Int_Int_goConst_buf  <= 1'd0;
    else
      if ((\call_f''''''''_f''''''''_Int_Int_initBufi_r  && \call_f''''''''_f''''''''_Int_Int_goConst_buf [0]))
        \call_f''''''''_f''''''''_Int_Int_goConst_buf  <= 1'd0;
      else if (((! \call_f''''''''_f''''''''_Int_Int_initBufi_r ) && (! \call_f''''''''_f''''''''_Int_Int_goConst_buf [0])))
        \call_f''''''''_f''''''''_Int_Int_goConst_buf  <= \call_f''''''''_f''''''''_Int_Int_goConst_d ;
  
  /* mergectrl (Ty C5,
           Ty Go) : [(call_f''''''''_f''''''''_Int_Int_goMux1,Go),
                     (lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int3_1_argbuf,Go),
                     (lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int2_1_argbuf,Go),
                     (lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int1_1_argbuf,Go),
                     (lizzieLet6_3QNode_Int_1_argbuf,Go)] > (go_11_goMux_choice,C5) (go_11_goMux_data,Go) */
  logic [4:0] \call_f''''''''_f''''''''_Int_Int_goMux1_select_d ;
  assign \call_f''''''''_f''''''''_Int_Int_goMux1_select_d  = ((| \call_f''''''''_f''''''''_Int_Int_goMux1_select_q ) ? \call_f''''''''_f''''''''_Int_Int_goMux1_select_q  :
                                                               (\call_f''''''''_f''''''''_Int_Int_goMux1_d [0] ? 5'd1 :
                                                                (\lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int3_1_argbuf_d [0] ? 5'd2 :
                                                                 (\lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int2_1_argbuf_d [0] ? 5'd4 :
                                                                  (\lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int1_1_argbuf_d [0] ? 5'd8 :
                                                                   (lizzieLet6_3QNode_Int_1_argbuf_d[0] ? 5'd16 :
                                                                    5'd0))))));
  logic [4:0] \call_f''''''''_f''''''''_Int_Int_goMux1_select_q ;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \call_f''''''''_f''''''''_Int_Int_goMux1_select_q  <= 5'd0;
    else
      \call_f''''''''_f''''''''_Int_Int_goMux1_select_q  <= (\call_f''''''''_f''''''''_Int_Int_goMux1_done  ? 5'd0 :
                                                             \call_f''''''''_f''''''''_Int_Int_goMux1_select_d );
  logic [1:0] \call_f''''''''_f''''''''_Int_Int_goMux1_emit_q ;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \call_f''''''''_f''''''''_Int_Int_goMux1_emit_q  <= 2'd0;
    else
      \call_f''''''''_f''''''''_Int_Int_goMux1_emit_q  <= (\call_f''''''''_f''''''''_Int_Int_goMux1_done  ? 2'd0 :
                                                           \call_f''''''''_f''''''''_Int_Int_goMux1_emit_d );
  logic [1:0] \call_f''''''''_f''''''''_Int_Int_goMux1_emit_d ;
  assign \call_f''''''''_f''''''''_Int_Int_goMux1_emit_d  = (\call_f''''''''_f''''''''_Int_Int_goMux1_emit_q  | ({go_11_goMux_choice_d[0],
                                                                                                                  go_11_goMux_data_d[0]} & {go_11_goMux_choice_r,
                                                                                                                                            go_11_goMux_data_r}));
  logic \call_f''''''''_f''''''''_Int_Int_goMux1_done ;
  assign \call_f''''''''_f''''''''_Int_Int_goMux1_done  = (& \call_f''''''''_f''''''''_Int_Int_goMux1_emit_d );
  assign {lizzieLet6_3QNode_Int_1_argbuf_r,
          \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int1_1_argbuf_r ,
          \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int2_1_argbuf_r ,
          \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int3_1_argbuf_r ,
          \call_f''''''''_f''''''''_Int_Int_goMux1_r } = (\call_f''''''''_f''''''''_Int_Int_goMux1_done  ? \call_f''''''''_f''''''''_Int_Int_goMux1_select_d  :
                                                          5'd0);
  assign go_11_goMux_data_d = ((\call_f''''''''_f''''''''_Int_Int_goMux1_select_d [0] && (! \call_f''''''''_f''''''''_Int_Int_goMux1_emit_q [0])) ? \call_f''''''''_f''''''''_Int_Int_goMux1_d  :
                               ((\call_f''''''''_f''''''''_Int_Int_goMux1_select_d [1] && (! \call_f''''''''_f''''''''_Int_Int_goMux1_emit_q [0])) ? \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int3_1_argbuf_d  :
                                ((\call_f''''''''_f''''''''_Int_Int_goMux1_select_d [2] && (! \call_f''''''''_f''''''''_Int_Int_goMux1_emit_q [0])) ? \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int2_1_argbuf_d  :
                                 ((\call_f''''''''_f''''''''_Int_Int_goMux1_select_d [3] && (! \call_f''''''''_f''''''''_Int_Int_goMux1_emit_q [0])) ? \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int1_1_argbuf_d  :
                                  ((\call_f''''''''_f''''''''_Int_Int_goMux1_select_d [4] && (! \call_f''''''''_f''''''''_Int_Int_goMux1_emit_q [0])) ? lizzieLet6_3QNode_Int_1_argbuf_d :
                                   1'd0)))));
  assign go_11_goMux_choice_d = ((\call_f''''''''_f''''''''_Int_Int_goMux1_select_d [0] && (! \call_f''''''''_f''''''''_Int_Int_goMux1_emit_q [1])) ? C1_5_dc(1'd1) :
                                 ((\call_f''''''''_f''''''''_Int_Int_goMux1_select_d [1] && (! \call_f''''''''_f''''''''_Int_Int_goMux1_emit_q [1])) ? C2_5_dc(1'd1) :
                                  ((\call_f''''''''_f''''''''_Int_Int_goMux1_select_d [2] && (! \call_f''''''''_f''''''''_Int_Int_goMux1_emit_q [1])) ? C3_5_dc(1'd1) :
                                   ((\call_f''''''''_f''''''''_Int_Int_goMux1_select_d [3] && (! \call_f''''''''_f''''''''_Int_Int_goMux1_emit_q [1])) ? C4_5_dc(1'd1) :
                                    ((\call_f''''''''_f''''''''_Int_Int_goMux1_select_d [4] && (! \call_f''''''''_f''''''''_Int_Int_goMux1_emit_q [1])) ? C5_5_dc(1'd1) :
                                     {3'd0, 1'd0})))));
  
  /* fork (Ty Go) : (call_f''''''''_f''''''''_Int_Int_initBuf,Go) > [(call_f''''''''_f''''''''_Int_Int_unlockFork1,Go),
                                                                (call_f''''''''_f''''''''_Int_Int_unlockFork2,Go),
                                                                (call_f''''''''_f''''''''_Int_Int_unlockFork3,Go),
                                                                (call_f''''''''_f''''''''_Int_Int_unlockFork4,Go),
                                                                (call_f''''''''_f''''''''_Int_Int_unlockFork5,Go)] */
  logic [4:0] \call_f''''''''_f''''''''_Int_Int_initBuf_emitted ;
  logic [4:0] \call_f''''''''_f''''''''_Int_Int_initBuf_done ;
  assign \call_f''''''''_f''''''''_Int_Int_unlockFork1_d  = (\call_f''''''''_f''''''''_Int_Int_initBuf_d [0] && (! \call_f''''''''_f''''''''_Int_Int_initBuf_emitted [0]));
  assign \call_f''''''''_f''''''''_Int_Int_unlockFork2_d  = (\call_f''''''''_f''''''''_Int_Int_initBuf_d [0] && (! \call_f''''''''_f''''''''_Int_Int_initBuf_emitted [1]));
  assign \call_f''''''''_f''''''''_Int_Int_unlockFork3_d  = (\call_f''''''''_f''''''''_Int_Int_initBuf_d [0] && (! \call_f''''''''_f''''''''_Int_Int_initBuf_emitted [2]));
  assign \call_f''''''''_f''''''''_Int_Int_unlockFork4_d  = (\call_f''''''''_f''''''''_Int_Int_initBuf_d [0] && (! \call_f''''''''_f''''''''_Int_Int_initBuf_emitted [3]));
  assign \call_f''''''''_f''''''''_Int_Int_unlockFork5_d  = (\call_f''''''''_f''''''''_Int_Int_initBuf_d [0] && (! \call_f''''''''_f''''''''_Int_Int_initBuf_emitted [4]));
  assign \call_f''''''''_f''''''''_Int_Int_initBuf_done  = (\call_f''''''''_f''''''''_Int_Int_initBuf_emitted  | ({\call_f''''''''_f''''''''_Int_Int_unlockFork5_d [0],
                                                                                                                   \call_f''''''''_f''''''''_Int_Int_unlockFork4_d [0],
                                                                                                                   \call_f''''''''_f''''''''_Int_Int_unlockFork3_d [0],
                                                                                                                   \call_f''''''''_f''''''''_Int_Int_unlockFork2_d [0],
                                                                                                                   \call_f''''''''_f''''''''_Int_Int_unlockFork1_d [0]} & {\call_f''''''''_f''''''''_Int_Int_unlockFork5_r ,
                                                                                                                                                                           \call_f''''''''_f''''''''_Int_Int_unlockFork4_r ,
                                                                                                                                                                           \call_f''''''''_f''''''''_Int_Int_unlockFork3_r ,
                                                                                                                                                                           \call_f''''''''_f''''''''_Int_Int_unlockFork2_r ,
                                                                                                                                                                           \call_f''''''''_f''''''''_Int_Int_unlockFork1_r }));
  assign \call_f''''''''_f''''''''_Int_Int_initBuf_r  = (& \call_f''''''''_f''''''''_Int_Int_initBuf_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \call_f''''''''_f''''''''_Int_Int_initBuf_emitted  <= 5'd0;
    else
      \call_f''''''''_f''''''''_Int_Int_initBuf_emitted  <= (\call_f''''''''_f''''''''_Int_Int_initBuf_r  ? 5'd0 :
                                                             \call_f''''''''_f''''''''_Int_Int_initBuf_done );
  
  /* initbuf (Ty Go,
         Dcon Go) : (call_f''''''''_f''''''''_Int_Int_initBufi,Go) > (call_f''''''''_f''''''''_Int_Int_initBuf,Go) */
  assign \call_f''''''''_f''''''''_Int_Int_initBufi_r  = ((! \call_f''''''''_f''''''''_Int_Int_initBuf_d [0]) || \call_f''''''''_f''''''''_Int_Int_initBuf_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \call_f''''''''_f''''''''_Int_Int_initBuf_d  <= Go_dc(1'd1);
    else
      if (\call_f''''''''_f''''''''_Int_Int_initBufi_r )
        \call_f''''''''_f''''''''_Int_Int_initBuf_d  <= \call_f''''''''_f''''''''_Int_Int_initBufi_d ;
  
  /* mux (Ty Go,
     Ty Go) : (call_f''''''''_f''''''''_Int_Int_unlockFork1,Go) [(call_f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf''''''''_f''''''''_Int_Intgo_11,Go)] > (call_f''''''''_f''''''''_Int_Int_goMux1,Go) */
  assign \call_f''''''''_f''''''''_Int_Int_goMux1_d  = (\call_f''''''''_f''''''''_Int_Int_unlockFork1_d [0] && \call_f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf''''''''_f''''''''_Int_Intgo_11_d [0]);
  assign \call_f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf''''''''_f''''''''_Int_Intgo_11_r  = (\call_f''''''''_f''''''''_Int_Int_goMux1_r  && (\call_f''''''''_f''''''''_Int_Int_unlockFork1_d [0] && \call_f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf''''''''_f''''''''_Int_Intgo_11_d [0]));
  assign \call_f''''''''_f''''''''_Int_Int_unlockFork1_r  = (\call_f''''''''_f''''''''_Int_Int_goMux1_r  && (\call_f''''''''_f''''''''_Int_Int_unlockFork1_d [0] && \call_f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf''''''''_f''''''''_Int_Intgo_11_d [0]));
  
  /* mux (Ty Go,
     Ty Pointer_QTree_Int) : (call_f''''''''_f''''''''_Int_Int_unlockFork2,Go) [(call_f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf''''''''_f''''''''_Int_Intq4a8u,Pointer_QTree_Int)] > (call_f''''''''_f''''''''_Int_Int_goMux2,Pointer_QTree_Int) */
  assign \call_f''''''''_f''''''''_Int_Int_goMux2_d  = {\call_f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf''''''''_f''''''''_Int_Intq4a8u_d [16:1],
                                                        (\call_f''''''''_f''''''''_Int_Int_unlockFork2_d [0] && \call_f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf''''''''_f''''''''_Int_Intq4a8u_d [0])};
  assign \call_f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf''''''''_f''''''''_Int_Intq4a8u_r  = (\call_f''''''''_f''''''''_Int_Int_goMux2_r  && (\call_f''''''''_f''''''''_Int_Int_unlockFork2_d [0] && \call_f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf''''''''_f''''''''_Int_Intq4a8u_d [0]));
  assign \call_f''''''''_f''''''''_Int_Int_unlockFork2_r  = (\call_f''''''''_f''''''''_Int_Int_goMux2_r  && (\call_f''''''''_f''''''''_Int_Int_unlockFork2_d [0] && \call_f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf''''''''_f''''''''_Int_Intq4a8u_d [0]));
  
  /* mux (Ty Go,
     Ty MyDTInt_Bool) : (call_f''''''''_f''''''''_Int_Int_unlockFork3,Go) [(call_f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf''''''''_f''''''''_Int_Intis_z_mapa8v,MyDTInt_Bool)] > (call_f''''''''_f''''''''_Int_Int_goMux3,MyDTInt_Bool) */
  assign \call_f''''''''_f''''''''_Int_Int_goMux3_d  = (\call_f''''''''_f''''''''_Int_Int_unlockFork3_d [0] && \call_f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf''''''''_f''''''''_Int_Intis_z_mapa8v_d [0]);
  assign \call_f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf''''''''_f''''''''_Int_Intis_z_mapa8v_r  = (\call_f''''''''_f''''''''_Int_Int_goMux3_r  && (\call_f''''''''_f''''''''_Int_Int_unlockFork3_d [0] && \call_f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf''''''''_f''''''''_Int_Intis_z_mapa8v_d [0]));
  assign \call_f''''''''_f''''''''_Int_Int_unlockFork3_r  = (\call_f''''''''_f''''''''_Int_Int_goMux3_r  && (\call_f''''''''_f''''''''_Int_Int_unlockFork3_d [0] && \call_f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf''''''''_f''''''''_Int_Intis_z_mapa8v_d [0]));
  
  /* mux (Ty Go,
     Ty MyDTInt_Int) : (call_f''''''''_f''''''''_Int_Int_unlockFork4,Go) [(call_f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf''''''''_f''''''''_Int_Intop_mapa8w,MyDTInt_Int)] > (call_f''''''''_f''''''''_Int_Int_goMux4,MyDTInt_Int) */
  assign \call_f''''''''_f''''''''_Int_Int_goMux4_d  = (\call_f''''''''_f''''''''_Int_Int_unlockFork4_d [0] && \call_f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf''''''''_f''''''''_Int_Intop_mapa8w_d [0]);
  assign \call_f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf''''''''_f''''''''_Int_Intop_mapa8w_r  = (\call_f''''''''_f''''''''_Int_Int_goMux4_r  && (\call_f''''''''_f''''''''_Int_Int_unlockFork4_d [0] && \call_f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf''''''''_f''''''''_Int_Intop_mapa8w_d [0]));
  assign \call_f''''''''_f''''''''_Int_Int_unlockFork4_r  = (\call_f''''''''_f''''''''_Int_Int_goMux4_r  && (\call_f''''''''_f''''''''_Int_Int_unlockFork4_d [0] && \call_f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf''''''''_f''''''''_Int_Intop_mapa8w_d [0]));
  
  /* mux (Ty Go,
     Ty Pointer_CTf''''''''_f''''''''_Int_Int) : (call_f''''''''_f''''''''_Int_Int_unlockFork5,Go) [(call_f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf''''''''_f''''''''_Int_Intsc_0_1,Pointer_CTf''''''''_f''''''''_Int_Int)] > (call_f''''''''_f''''''''_Int_Int_goMux5,Pointer_CTf''''''''_f''''''''_Int_Int) */
  assign \call_f''''''''_f''''''''_Int_Int_goMux5_d  = {\call_f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf''''''''_f''''''''_Int_Intsc_0_1_d [16:1],
                                                        (\call_f''''''''_f''''''''_Int_Int_unlockFork5_d [0] && \call_f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf''''''''_f''''''''_Int_Intsc_0_1_d [0])};
  assign \call_f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf''''''''_f''''''''_Int_Intsc_0_1_r  = (\call_f''''''''_f''''''''_Int_Int_goMux5_r  && (\call_f''''''''_f''''''''_Int_Int_unlockFork5_d [0] && \call_f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf''''''''_f''''''''_Int_Intsc_0_1_d [0]));
  assign \call_f''''''''_f''''''''_Int_Int_unlockFork5_r  = (\call_f''''''''_f''''''''_Int_Int_goMux5_r  && (\call_f''''''''_f''''''''_Int_Int_unlockFork5_d [0] && \call_f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf''''''''_f''''''''_Int_Intsc_0_1_d [0]));
  
  /* destruct (Ty TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Int,
          Dcon TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Int) : (call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Int_1,TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Int) > [(call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Intgo_12,Go),
                                                                                                                                                                                                                                                                                                                                                                                                                                                     (call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Intm1a8C,Pointer_QTree_Int),
                                                                                                                                                                                                                                                                                                                                                                                                                                                     (call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Intm2a8D,Pointer_QTree_Int),
                                                                                                                                                                                                                                                                                                                                                                                                                                                     (call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Intis_z_mapa8E,MyDTInt_Bool),
                                                                                                                                                                                                                                                                                                                                                                                                                                                     (call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Intop_mapa8F,MyDTInt_Int),
                                                                                                                                                                                                                                                                                                                                                                                                                                                     (call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Intis_z_adda8G,MyDTInt_Bool),
                                                                                                                                                                                                                                                                                                                                                                                                                                                     (call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Intop_adda8H,MyDTInt_Int_Int),
                                                                                                                                                                                                                                                                                                                                                                                                                                                     (call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Intsc_0_2,Pointer_CTf_f_Int_Int)] */
  logic [7:0] call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Int_1_emitted;
  logic [7:0] call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Int_1_done;
  assign call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Intgo_12_d = (call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Int_1_d[0] && (! call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Int_1_emitted[0]));
  assign call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Intm1a8C_d = {call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Int_1_d[16:1],
                                                                                                                                                                       (call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Int_1_d[0] && (! call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Int_1_emitted[1]))};
  assign call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Intm2a8D_d = {call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Int_1_d[32:17],
                                                                                                                                                                       (call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Int_1_d[0] && (! call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Int_1_emitted[2]))};
  assign call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Intis_z_mapa8E_d = (call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Int_1_d[0] && (! call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Int_1_emitted[3]));
  assign call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Intop_mapa8F_d = (call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Int_1_d[0] && (! call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Int_1_emitted[4]));
  assign call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Intis_z_adda8G_d = (call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Int_1_d[0] && (! call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Int_1_emitted[5]));
  assign call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Intop_adda8H_d = (call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Int_1_d[0] && (! call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Int_1_emitted[6]));
  assign call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Intsc_0_2_d = {call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Int_1_d[48:33],
                                                                                                                                                                        (call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Int_1_d[0] && (! call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Int_1_emitted[7]))};
  assign call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Int_1_done = (call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Int_1_emitted | ({call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Intsc_0_2_d[0],
                                                                                                                                                                                                                                                                                                                                         call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Intop_adda8H_d[0],
                                                                                                                                                                                                                                                                                                                                         call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Intis_z_adda8G_d[0],
                                                                                                                                                                                                                                                                                                                                         call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Intop_mapa8F_d[0],
                                                                                                                                                                                                                                                                                                                                         call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Intis_z_mapa8E_d[0],
                                                                                                                                                                                                                                                                                                                                         call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Intm2a8D_d[0],
                                                                                                                                                                                                                                                                                                                                         call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Intm1a8C_d[0],
                                                                                                                                                                                                                                                                                                                                         call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Intgo_12_d[0]} & {call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Intsc_0_2_r,
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Intop_adda8H_r,
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Intis_z_adda8G_r,
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Intop_mapa8F_r,
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Intis_z_mapa8E_r,
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Intm2a8D_r,
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Intm1a8C_r,
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Intgo_12_r}));
  assign call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Int_1_r = (& call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Int_1_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Int_1_emitted <= 8'd0;
    else
      call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Int_1_emitted <= (call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Int_1_r ? 8'd0 :
                                                                                                                                                                        call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Int_1_done);
  
  /* rbuf (Ty Go) : (call_f_f_Int_Int_goConst,Go) > (call_f_f_Int_Int_initBufi,Go) */
  Go_t call_f_f_Int_Int_goConst_buf;
  assign call_f_f_Int_Int_goConst_r = (! call_f_f_Int_Int_goConst_buf[0]);
  assign call_f_f_Int_Int_initBufi_d = (call_f_f_Int_Int_goConst_buf[0] ? call_f_f_Int_Int_goConst_buf :
                                        call_f_f_Int_Int_goConst_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_f_f_Int_Int_goConst_buf <= 1'd0;
    else
      if ((call_f_f_Int_Int_initBufi_r && call_f_f_Int_Int_goConst_buf[0]))
        call_f_f_Int_Int_goConst_buf <= 1'd0;
      else if (((! call_f_f_Int_Int_initBufi_r) && (! call_f_f_Int_Int_goConst_buf[0])))
        call_f_f_Int_Int_goConst_buf <= call_f_f_Int_Int_goConst_d;
  
  /* mergectrl (Ty C5,Ty Go) : [(call_f_f_Int_Int_goMux1,Go),
                           (lizzieLet44_3Lcall_f_f_Int_Int3_1_argbuf,Go),
                           (lizzieLet44_3Lcall_f_f_Int_Int2_1_argbuf,Go),
                           (lizzieLet44_3Lcall_f_f_Int_Int1_1_argbuf,Go),
                           (lizzieLet12_6QNode_Int_3QNode_Int_1_argbuf,Go)] > (go_12_goMux_choice,C5) (go_12_goMux_data,Go) */
  logic [4:0] call_f_f_Int_Int_goMux1_select_d;
  assign call_f_f_Int_Int_goMux1_select_d = ((| call_f_f_Int_Int_goMux1_select_q) ? call_f_f_Int_Int_goMux1_select_q :
                                             (call_f_f_Int_Int_goMux1_d[0] ? 5'd1 :
                                              (lizzieLet44_3Lcall_f_f_Int_Int3_1_argbuf_d[0] ? 5'd2 :
                                               (lizzieLet44_3Lcall_f_f_Int_Int2_1_argbuf_d[0] ? 5'd4 :
                                                (lizzieLet44_3Lcall_f_f_Int_Int1_1_argbuf_d[0] ? 5'd8 :
                                                 (lizzieLet12_6QNode_Int_3QNode_Int_1_argbuf_d[0] ? 5'd16 :
                                                  5'd0))))));
  logic [4:0] call_f_f_Int_Int_goMux1_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_f_f_Int_Int_goMux1_select_q <= 5'd0;
    else
      call_f_f_Int_Int_goMux1_select_q <= (call_f_f_Int_Int_goMux1_done ? 5'd0 :
                                           call_f_f_Int_Int_goMux1_select_d);
  logic [1:0] call_f_f_Int_Int_goMux1_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_f_f_Int_Int_goMux1_emit_q <= 2'd0;
    else
      call_f_f_Int_Int_goMux1_emit_q <= (call_f_f_Int_Int_goMux1_done ? 2'd0 :
                                         call_f_f_Int_Int_goMux1_emit_d);
  logic [1:0] call_f_f_Int_Int_goMux1_emit_d;
  assign call_f_f_Int_Int_goMux1_emit_d = (call_f_f_Int_Int_goMux1_emit_q | ({go_12_goMux_choice_d[0],
                                                                              go_12_goMux_data_d[0]} & {go_12_goMux_choice_r,
                                                                                                        go_12_goMux_data_r}));
  logic call_f_f_Int_Int_goMux1_done;
  assign call_f_f_Int_Int_goMux1_done = (& call_f_f_Int_Int_goMux1_emit_d);
  assign {lizzieLet12_6QNode_Int_3QNode_Int_1_argbuf_r,
          lizzieLet44_3Lcall_f_f_Int_Int1_1_argbuf_r,
          lizzieLet44_3Lcall_f_f_Int_Int2_1_argbuf_r,
          lizzieLet44_3Lcall_f_f_Int_Int3_1_argbuf_r,
          call_f_f_Int_Int_goMux1_r} = (call_f_f_Int_Int_goMux1_done ? call_f_f_Int_Int_goMux1_select_d :
                                        5'd0);
  assign go_12_goMux_data_d = ((call_f_f_Int_Int_goMux1_select_d[0] && (! call_f_f_Int_Int_goMux1_emit_q[0])) ? call_f_f_Int_Int_goMux1_d :
                               ((call_f_f_Int_Int_goMux1_select_d[1] && (! call_f_f_Int_Int_goMux1_emit_q[0])) ? lizzieLet44_3Lcall_f_f_Int_Int3_1_argbuf_d :
                                ((call_f_f_Int_Int_goMux1_select_d[2] && (! call_f_f_Int_Int_goMux1_emit_q[0])) ? lizzieLet44_3Lcall_f_f_Int_Int2_1_argbuf_d :
                                 ((call_f_f_Int_Int_goMux1_select_d[3] && (! call_f_f_Int_Int_goMux1_emit_q[0])) ? lizzieLet44_3Lcall_f_f_Int_Int1_1_argbuf_d :
                                  ((call_f_f_Int_Int_goMux1_select_d[4] && (! call_f_f_Int_Int_goMux1_emit_q[0])) ? lizzieLet12_6QNode_Int_3QNode_Int_1_argbuf_d :
                                   1'd0)))));
  assign go_12_goMux_choice_d = ((call_f_f_Int_Int_goMux1_select_d[0] && (! call_f_f_Int_Int_goMux1_emit_q[1])) ? C1_5_dc(1'd1) :
                                 ((call_f_f_Int_Int_goMux1_select_d[1] && (! call_f_f_Int_Int_goMux1_emit_q[1])) ? C2_5_dc(1'd1) :
                                  ((call_f_f_Int_Int_goMux1_select_d[2] && (! call_f_f_Int_Int_goMux1_emit_q[1])) ? C3_5_dc(1'd1) :
                                   ((call_f_f_Int_Int_goMux1_select_d[3] && (! call_f_f_Int_Int_goMux1_emit_q[1])) ? C4_5_dc(1'd1) :
                                    ((call_f_f_Int_Int_goMux1_select_d[4] && (! call_f_f_Int_Int_goMux1_emit_q[1])) ? C5_5_dc(1'd1) :
                                     {3'd0, 1'd0})))));
  
  /* fork (Ty Go) : (call_f_f_Int_Int_initBuf,Go) > [(call_f_f_Int_Int_unlockFork1,Go),
                                                (call_f_f_Int_Int_unlockFork2,Go),
                                                (call_f_f_Int_Int_unlockFork3,Go),
                                                (call_f_f_Int_Int_unlockFork4,Go),
                                                (call_f_f_Int_Int_unlockFork5,Go),
                                                (call_f_f_Int_Int_unlockFork6,Go),
                                                (call_f_f_Int_Int_unlockFork7,Go),
                                                (call_f_f_Int_Int_unlockFork8,Go)] */
  logic [7:0] call_f_f_Int_Int_initBuf_emitted;
  logic [7:0] call_f_f_Int_Int_initBuf_done;
  assign call_f_f_Int_Int_unlockFork1_d = (call_f_f_Int_Int_initBuf_d[0] && (! call_f_f_Int_Int_initBuf_emitted[0]));
  assign call_f_f_Int_Int_unlockFork2_d = (call_f_f_Int_Int_initBuf_d[0] && (! call_f_f_Int_Int_initBuf_emitted[1]));
  assign call_f_f_Int_Int_unlockFork3_d = (call_f_f_Int_Int_initBuf_d[0] && (! call_f_f_Int_Int_initBuf_emitted[2]));
  assign call_f_f_Int_Int_unlockFork4_d = (call_f_f_Int_Int_initBuf_d[0] && (! call_f_f_Int_Int_initBuf_emitted[3]));
  assign call_f_f_Int_Int_unlockFork5_d = (call_f_f_Int_Int_initBuf_d[0] && (! call_f_f_Int_Int_initBuf_emitted[4]));
  assign call_f_f_Int_Int_unlockFork6_d = (call_f_f_Int_Int_initBuf_d[0] && (! call_f_f_Int_Int_initBuf_emitted[5]));
  assign call_f_f_Int_Int_unlockFork7_d = (call_f_f_Int_Int_initBuf_d[0] && (! call_f_f_Int_Int_initBuf_emitted[6]));
  assign call_f_f_Int_Int_unlockFork8_d = (call_f_f_Int_Int_initBuf_d[0] && (! call_f_f_Int_Int_initBuf_emitted[7]));
  assign call_f_f_Int_Int_initBuf_done = (call_f_f_Int_Int_initBuf_emitted | ({call_f_f_Int_Int_unlockFork8_d[0],
                                                                               call_f_f_Int_Int_unlockFork7_d[0],
                                                                               call_f_f_Int_Int_unlockFork6_d[0],
                                                                               call_f_f_Int_Int_unlockFork5_d[0],
                                                                               call_f_f_Int_Int_unlockFork4_d[0],
                                                                               call_f_f_Int_Int_unlockFork3_d[0],
                                                                               call_f_f_Int_Int_unlockFork2_d[0],
                                                                               call_f_f_Int_Int_unlockFork1_d[0]} & {call_f_f_Int_Int_unlockFork8_r,
                                                                                                                     call_f_f_Int_Int_unlockFork7_r,
                                                                                                                     call_f_f_Int_Int_unlockFork6_r,
                                                                                                                     call_f_f_Int_Int_unlockFork5_r,
                                                                                                                     call_f_f_Int_Int_unlockFork4_r,
                                                                                                                     call_f_f_Int_Int_unlockFork3_r,
                                                                                                                     call_f_f_Int_Int_unlockFork2_r,
                                                                                                                     call_f_f_Int_Int_unlockFork1_r}));
  assign call_f_f_Int_Int_initBuf_r = (& call_f_f_Int_Int_initBuf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_f_f_Int_Int_initBuf_emitted <= 8'd0;
    else
      call_f_f_Int_Int_initBuf_emitted <= (call_f_f_Int_Int_initBuf_r ? 8'd0 :
                                           call_f_f_Int_Int_initBuf_done);
  
  /* initbuf (Ty Go,
         Dcon Go) : (call_f_f_Int_Int_initBufi,Go) > (call_f_f_Int_Int_initBuf,Go) */
  assign call_f_f_Int_Int_initBufi_r = ((! call_f_f_Int_Int_initBuf_d[0]) || call_f_f_Int_Int_initBuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_f_f_Int_Int_initBuf_d <= Go_dc(1'd1);
    else
      if (call_f_f_Int_Int_initBufi_r)
        call_f_f_Int_Int_initBuf_d <= call_f_f_Int_Int_initBufi_d;
  
  /* mux (Ty Go,
     Ty Go) : (call_f_f_Int_Int_unlockFork1,Go) [(call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Intgo_12,Go)] > (call_f_f_Int_Int_goMux1,Go) */
  assign call_f_f_Int_Int_goMux1_d = (call_f_f_Int_Int_unlockFork1_d[0] && call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Intgo_12_d[0]);
  assign call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Intgo_12_r = (call_f_f_Int_Int_goMux1_r && (call_f_f_Int_Int_unlockFork1_d[0] && call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Intgo_12_d[0]));
  assign call_f_f_Int_Int_unlockFork1_r = (call_f_f_Int_Int_goMux1_r && (call_f_f_Int_Int_unlockFork1_d[0] && call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Intgo_12_d[0]));
  
  /* mux (Ty Go,
     Ty Pointer_QTree_Int) : (call_f_f_Int_Int_unlockFork2,Go) [(call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Intm1a8C,Pointer_QTree_Int)] > (call_f_f_Int_Int_goMux2,Pointer_QTree_Int) */
  assign call_f_f_Int_Int_goMux2_d = {call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Intm1a8C_d[16:1],
                                      (call_f_f_Int_Int_unlockFork2_d[0] && call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Intm1a8C_d[0])};
  assign call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Intm1a8C_r = (call_f_f_Int_Int_goMux2_r && (call_f_f_Int_Int_unlockFork2_d[0] && call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Intm1a8C_d[0]));
  assign call_f_f_Int_Int_unlockFork2_r = (call_f_f_Int_Int_goMux2_r && (call_f_f_Int_Int_unlockFork2_d[0] && call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Intm1a8C_d[0]));
  
  /* mux (Ty Go,
     Ty Pointer_QTree_Int) : (call_f_f_Int_Int_unlockFork3,Go) [(call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Intm2a8D,Pointer_QTree_Int)] > (call_f_f_Int_Int_goMux3,Pointer_QTree_Int) */
  assign call_f_f_Int_Int_goMux3_d = {call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Intm2a8D_d[16:1],
                                      (call_f_f_Int_Int_unlockFork3_d[0] && call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Intm2a8D_d[0])};
  assign call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Intm2a8D_r = (call_f_f_Int_Int_goMux3_r && (call_f_f_Int_Int_unlockFork3_d[0] && call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Intm2a8D_d[0]));
  assign call_f_f_Int_Int_unlockFork3_r = (call_f_f_Int_Int_goMux3_r && (call_f_f_Int_Int_unlockFork3_d[0] && call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Intm2a8D_d[0]));
  
  /* mux (Ty Go,
     Ty MyDTInt_Bool) : (call_f_f_Int_Int_unlockFork4,Go) [(call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Intis_z_mapa8E,MyDTInt_Bool)] > (call_f_f_Int_Int_goMux4,MyDTInt_Bool) */
  assign call_f_f_Int_Int_goMux4_d = (call_f_f_Int_Int_unlockFork4_d[0] && call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Intis_z_mapa8E_d[0]);
  assign call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Intis_z_mapa8E_r = (call_f_f_Int_Int_goMux4_r && (call_f_f_Int_Int_unlockFork4_d[0] && call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Intis_z_mapa8E_d[0]));
  assign call_f_f_Int_Int_unlockFork4_r = (call_f_f_Int_Int_goMux4_r && (call_f_f_Int_Int_unlockFork4_d[0] && call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Intis_z_mapa8E_d[0]));
  
  /* mux (Ty Go,
     Ty MyDTInt_Int) : (call_f_f_Int_Int_unlockFork5,Go) [(call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Intop_mapa8F,MyDTInt_Int)] > (call_f_f_Int_Int_goMux5,MyDTInt_Int) */
  assign call_f_f_Int_Int_goMux5_d = (call_f_f_Int_Int_unlockFork5_d[0] && call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Intop_mapa8F_d[0]);
  assign call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Intop_mapa8F_r = (call_f_f_Int_Int_goMux5_r && (call_f_f_Int_Int_unlockFork5_d[0] && call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Intop_mapa8F_d[0]));
  assign call_f_f_Int_Int_unlockFork5_r = (call_f_f_Int_Int_goMux5_r && (call_f_f_Int_Int_unlockFork5_d[0] && call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Intop_mapa8F_d[0]));
  
  /* mux (Ty Go,
     Ty MyDTInt_Bool) : (call_f_f_Int_Int_unlockFork6,Go) [(call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Intis_z_adda8G,MyDTInt_Bool)] > (call_f_f_Int_Int_goMux6,MyDTInt_Bool) */
  assign call_f_f_Int_Int_goMux6_d = (call_f_f_Int_Int_unlockFork6_d[0] && call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Intis_z_adda8G_d[0]);
  assign call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Intis_z_adda8G_r = (call_f_f_Int_Int_goMux6_r && (call_f_f_Int_Int_unlockFork6_d[0] && call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Intis_z_adda8G_d[0]));
  assign call_f_f_Int_Int_unlockFork6_r = (call_f_f_Int_Int_goMux6_r && (call_f_f_Int_Int_unlockFork6_d[0] && call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Intis_z_adda8G_d[0]));
  
  /* mux (Ty Go,
     Ty MyDTInt_Int_Int) : (call_f_f_Int_Int_unlockFork7,Go) [(call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Intop_adda8H,MyDTInt_Int_Int)] > (call_f_f_Int_Int_goMux7,MyDTInt_Int_Int) */
  assign call_f_f_Int_Int_goMux7_d = (call_f_f_Int_Int_unlockFork7_d[0] && call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Intop_adda8H_d[0]);
  assign call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Intop_adda8H_r = (call_f_f_Int_Int_goMux7_r && (call_f_f_Int_Int_unlockFork7_d[0] && call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Intop_adda8H_d[0]));
  assign call_f_f_Int_Int_unlockFork7_r = (call_f_f_Int_Int_goMux7_r && (call_f_f_Int_Int_unlockFork7_d[0] && call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Intop_adda8H_d[0]));
  
  /* mux (Ty Go,
     Ty Pointer_CTf_f_Int_Int) : (call_f_f_Int_Int_unlockFork8,Go) [(call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Intsc_0_2,Pointer_CTf_f_Int_Int)] > (call_f_f_Int_Int_goMux8,Pointer_CTf_f_Int_Int) */
  assign call_f_f_Int_Int_goMux8_d = {call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Intsc_0_2_d[16:1],
                                      (call_f_f_Int_Int_unlockFork8_d[0] && call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Intsc_0_2_d[0])};
  assign call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Intsc_0_2_r = (call_f_f_Int_Int_goMux8_r && (call_f_f_Int_Int_unlockFork8_d[0] && call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Intsc_0_2_d[0]));
  assign call_f_f_Int_Int_unlockFork8_r = (call_f_f_Int_Int_goMux8_r && (call_f_f_Int_Int_unlockFork8_d[0] && call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Intsc_0_2_d[0]));
  
  /* demux (Ty MyBool,
       Ty Go) : (es_10_1,MyBool) (lizzieLet12_6QVal_Int_3QNone_Int_3,Go) > [(es_10_1MyFalse,Go),
                                                                            (es_10_1MyTrue,Go)] */
  logic [1:0] lizzieLet12_6QVal_Int_3QNone_Int_3_onehotd;
  always_comb
    if ((es_10_1_d[0] && lizzieLet12_6QVal_Int_3QNone_Int_3_d[0]))
      unique case (es_10_1_d[1:1])
        1'd0: lizzieLet12_6QVal_Int_3QNone_Int_3_onehotd = 2'd1;
        1'd1: lizzieLet12_6QVal_Int_3QNone_Int_3_onehotd = 2'd2;
        default: lizzieLet12_6QVal_Int_3QNone_Int_3_onehotd = 2'd0;
      endcase
    else lizzieLet12_6QVal_Int_3QNone_Int_3_onehotd = 2'd0;
  assign es_10_1MyFalse_d = lizzieLet12_6QVal_Int_3QNone_Int_3_onehotd[0];
  assign es_10_1MyTrue_d = lizzieLet12_6QVal_Int_3QNone_Int_3_onehotd[1];
  assign lizzieLet12_6QVal_Int_3QNone_Int_3_r = (| (lizzieLet12_6QVal_Int_3QNone_Int_3_onehotd & {es_10_1MyTrue_r,
                                                                                                  es_10_1MyFalse_r}));
  assign es_10_1_r = lizzieLet12_6QVal_Int_3QNone_Int_3_r;
  
  /* fork (Ty Go) : (es_10_1MyFalse,Go) > [(es_10_1MyFalse_1,Go),
                                      (es_10_1MyFalse_2,Go)] */
  logic [1:0] es_10_1MyFalse_emitted;
  logic [1:0] es_10_1MyFalse_done;
  assign es_10_1MyFalse_1_d = (es_10_1MyFalse_d[0] && (! es_10_1MyFalse_emitted[0]));
  assign es_10_1MyFalse_2_d = (es_10_1MyFalse_d[0] && (! es_10_1MyFalse_emitted[1]));
  assign es_10_1MyFalse_done = (es_10_1MyFalse_emitted | ({es_10_1MyFalse_2_d[0],
                                                           es_10_1MyFalse_1_d[0]} & {es_10_1MyFalse_2_r,
                                                                                     es_10_1MyFalse_1_r}));
  assign es_10_1MyFalse_r = (& es_10_1MyFalse_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_10_1MyFalse_emitted <= 2'd0;
    else
      es_10_1MyFalse_emitted <= (es_10_1MyFalse_r ? 2'd0 :
                                 es_10_1MyFalse_done);
  
  /* buf (Ty Go) : (es_10_1MyFalse_1,Go) > (es_10_1MyFalse_1_argbuf,Go) */
  Go_t es_10_1MyFalse_1_bufchan_d;
  logic es_10_1MyFalse_1_bufchan_r;
  assign es_10_1MyFalse_1_r = ((! es_10_1MyFalse_1_bufchan_d[0]) || es_10_1MyFalse_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_10_1MyFalse_1_bufchan_d <= 1'd0;
    else
      if (es_10_1MyFalse_1_r)
        es_10_1MyFalse_1_bufchan_d <= es_10_1MyFalse_1_d;
  Go_t es_10_1MyFalse_1_bufchan_buf;
  assign es_10_1MyFalse_1_bufchan_r = (! es_10_1MyFalse_1_bufchan_buf[0]);
  assign es_10_1MyFalse_1_argbuf_d = (es_10_1MyFalse_1_bufchan_buf[0] ? es_10_1MyFalse_1_bufchan_buf :
                                      es_10_1MyFalse_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_10_1MyFalse_1_bufchan_buf <= 1'd0;
    else
      if ((es_10_1MyFalse_1_argbuf_r && es_10_1MyFalse_1_bufchan_buf[0]))
        es_10_1MyFalse_1_bufchan_buf <= 1'd0;
      else if (((! es_10_1MyFalse_1_argbuf_r) && (! es_10_1MyFalse_1_bufchan_buf[0])))
        es_10_1MyFalse_1_bufchan_buf <= es_10_1MyFalse_1_bufchan_d;
  
  /* dcon (Ty TupGo___MyDTInt_Int___Int,
      Dcon TupGo___MyDTInt_Int___Int) : [(es_10_1MyFalse_1_argbuf,Go),
                                         (es_10_2MyFalse_1_argbuf,MyDTInt_Int),
                                         (es_10_4MyFalse_1_argbuf,Int)] > (applyfnInt_Int_5TupGo___MyDTInt_Int___Int6,TupGo___MyDTInt_Int___Int) */
  assign applyfnInt_Int_5TupGo___MyDTInt_Int___Int6_d = TupGo___MyDTInt_Int___Int_dc((& {es_10_1MyFalse_1_argbuf_d[0],
                                                                                         es_10_2MyFalse_1_argbuf_d[0],
                                                                                         es_10_4MyFalse_1_argbuf_d[0]}), es_10_1MyFalse_1_argbuf_d, es_10_2MyFalse_1_argbuf_d, es_10_4MyFalse_1_argbuf_d);
  assign {es_10_1MyFalse_1_argbuf_r,
          es_10_2MyFalse_1_argbuf_r,
          es_10_4MyFalse_1_argbuf_r} = {3 {(applyfnInt_Int_5TupGo___MyDTInt_Int___Int6_r && applyfnInt_Int_5TupGo___MyDTInt_Int___Int6_d[0])}};
  
  /* buf (Ty Go) : (es_10_1MyFalse_2,Go) > (es_10_1MyFalse_2_argbuf,Go) */
  Go_t es_10_1MyFalse_2_bufchan_d;
  logic es_10_1MyFalse_2_bufchan_r;
  assign es_10_1MyFalse_2_r = ((! es_10_1MyFalse_2_bufchan_d[0]) || es_10_1MyFalse_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_10_1MyFalse_2_bufchan_d <= 1'd0;
    else
      if (es_10_1MyFalse_2_r)
        es_10_1MyFalse_2_bufchan_d <= es_10_1MyFalse_2_d;
  Go_t es_10_1MyFalse_2_bufchan_buf;
  assign es_10_1MyFalse_2_bufchan_r = (! es_10_1MyFalse_2_bufchan_buf[0]);
  assign es_10_1MyFalse_2_argbuf_d = (es_10_1MyFalse_2_bufchan_buf[0] ? es_10_1MyFalse_2_bufchan_buf :
                                      es_10_1MyFalse_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_10_1MyFalse_2_bufchan_buf <= 1'd0;
    else
      if ((es_10_1MyFalse_2_argbuf_r && es_10_1MyFalse_2_bufchan_buf[0]))
        es_10_1MyFalse_2_bufchan_buf <= 1'd0;
      else if (((! es_10_1MyFalse_2_argbuf_r) && (! es_10_1MyFalse_2_bufchan_buf[0])))
        es_10_1MyFalse_2_bufchan_buf <= es_10_1MyFalse_2_bufchan_d;
  
  /* fork (Ty Go) : (es_10_1MyTrue,Go) > [(es_10_1MyTrue_1,Go),
                                     (es_10_1MyTrue_2,Go)] */
  logic [1:0] es_10_1MyTrue_emitted;
  logic [1:0] es_10_1MyTrue_done;
  assign es_10_1MyTrue_1_d = (es_10_1MyTrue_d[0] && (! es_10_1MyTrue_emitted[0]));
  assign es_10_1MyTrue_2_d = (es_10_1MyTrue_d[0] && (! es_10_1MyTrue_emitted[1]));
  assign es_10_1MyTrue_done = (es_10_1MyTrue_emitted | ({es_10_1MyTrue_2_d[0],
                                                         es_10_1MyTrue_1_d[0]} & {es_10_1MyTrue_2_r,
                                                                                  es_10_1MyTrue_1_r}));
  assign es_10_1MyTrue_r = (& es_10_1MyTrue_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_10_1MyTrue_emitted <= 2'd0;
    else
      es_10_1MyTrue_emitted <= (es_10_1MyTrue_r ? 2'd0 :
                                es_10_1MyTrue_done);
  
  /* dcon (Ty QTree_Int,
      Dcon QNone_Int) : [(es_10_1MyTrue_1,Go)] > (es_10_1MyTrue_1QNone_Int,QTree_Int) */
  assign es_10_1MyTrue_1QNone_Int_d = QNone_Int_dc((& {es_10_1MyTrue_1_d[0]}), es_10_1MyTrue_1_d);
  assign {es_10_1MyTrue_1_r} = {1 {(es_10_1MyTrue_1QNone_Int_r && es_10_1MyTrue_1QNone_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (es_10_1MyTrue_1QNone_Int,QTree_Int) > (lizzieLet21_1_argbuf,QTree_Int) */
  QTree_Int_t es_10_1MyTrue_1QNone_Int_bufchan_d;
  logic es_10_1MyTrue_1QNone_Int_bufchan_r;
  assign es_10_1MyTrue_1QNone_Int_r = ((! es_10_1MyTrue_1QNone_Int_bufchan_d[0]) || es_10_1MyTrue_1QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_10_1MyTrue_1QNone_Int_bufchan_d <= {66'd0, 1'd0};
    else
      if (es_10_1MyTrue_1QNone_Int_r)
        es_10_1MyTrue_1QNone_Int_bufchan_d <= es_10_1MyTrue_1QNone_Int_d;
  QTree_Int_t es_10_1MyTrue_1QNone_Int_bufchan_buf;
  assign es_10_1MyTrue_1QNone_Int_bufchan_r = (! es_10_1MyTrue_1QNone_Int_bufchan_buf[0]);
  assign lizzieLet21_1_argbuf_d = (es_10_1MyTrue_1QNone_Int_bufchan_buf[0] ? es_10_1MyTrue_1QNone_Int_bufchan_buf :
                                   es_10_1MyTrue_1QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_10_1MyTrue_1QNone_Int_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((lizzieLet21_1_argbuf_r && es_10_1MyTrue_1QNone_Int_bufchan_buf[0]))
        es_10_1MyTrue_1QNone_Int_bufchan_buf <= {66'd0, 1'd0};
      else if (((! lizzieLet21_1_argbuf_r) && (! es_10_1MyTrue_1QNone_Int_bufchan_buf[0])))
        es_10_1MyTrue_1QNone_Int_bufchan_buf <= es_10_1MyTrue_1QNone_Int_bufchan_d;
  
  /* buf (Ty Go) : (es_10_1MyTrue_2,Go) > (es_10_1MyTrue_2_argbuf,Go) */
  Go_t es_10_1MyTrue_2_bufchan_d;
  logic es_10_1MyTrue_2_bufchan_r;
  assign es_10_1MyTrue_2_r = ((! es_10_1MyTrue_2_bufchan_d[0]) || es_10_1MyTrue_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_10_1MyTrue_2_bufchan_d <= 1'd0;
    else
      if (es_10_1MyTrue_2_r)
        es_10_1MyTrue_2_bufchan_d <= es_10_1MyTrue_2_d;
  Go_t es_10_1MyTrue_2_bufchan_buf;
  assign es_10_1MyTrue_2_bufchan_r = (! es_10_1MyTrue_2_bufchan_buf[0]);
  assign es_10_1MyTrue_2_argbuf_d = (es_10_1MyTrue_2_bufchan_buf[0] ? es_10_1MyTrue_2_bufchan_buf :
                                     es_10_1MyTrue_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_10_1MyTrue_2_bufchan_buf <= 1'd0;
    else
      if ((es_10_1MyTrue_2_argbuf_r && es_10_1MyTrue_2_bufchan_buf[0]))
        es_10_1MyTrue_2_bufchan_buf <= 1'd0;
      else if (((! es_10_1MyTrue_2_argbuf_r) && (! es_10_1MyTrue_2_bufchan_buf[0])))
        es_10_1MyTrue_2_bufchan_buf <= es_10_1MyTrue_2_bufchan_d;
  
  /* demux (Ty MyBool,
       Ty MyDTInt_Int) : (es_10_2,MyBool) (lizzieLet12_6QVal_Int_7QNone_Int_2,MyDTInt_Int) > [(es_10_2MyFalse,MyDTInt_Int),
                                                                                              (_80,MyDTInt_Int)] */
  logic [1:0] lizzieLet12_6QVal_Int_7QNone_Int_2_onehotd;
  always_comb
    if ((es_10_2_d[0] && lizzieLet12_6QVal_Int_7QNone_Int_2_d[0]))
      unique case (es_10_2_d[1:1])
        1'd0: lizzieLet12_6QVal_Int_7QNone_Int_2_onehotd = 2'd1;
        1'd1: lizzieLet12_6QVal_Int_7QNone_Int_2_onehotd = 2'd2;
        default: lizzieLet12_6QVal_Int_7QNone_Int_2_onehotd = 2'd0;
      endcase
    else lizzieLet12_6QVal_Int_7QNone_Int_2_onehotd = 2'd0;
  assign es_10_2MyFalse_d = lizzieLet12_6QVal_Int_7QNone_Int_2_onehotd[0];
  assign _80_d = lizzieLet12_6QVal_Int_7QNone_Int_2_onehotd[1];
  assign lizzieLet12_6QVal_Int_7QNone_Int_2_r = (| (lizzieLet12_6QVal_Int_7QNone_Int_2_onehotd & {_80_r,
                                                                                                  es_10_2MyFalse_r}));
  assign es_10_2_r = lizzieLet12_6QVal_Int_7QNone_Int_2_r;
  
  /* buf (Ty MyDTInt_Int) : (es_10_2MyFalse,MyDTInt_Int) > (es_10_2MyFalse_1_argbuf,MyDTInt_Int) */
  MyDTInt_Int_t es_10_2MyFalse_bufchan_d;
  logic es_10_2MyFalse_bufchan_r;
  assign es_10_2MyFalse_r = ((! es_10_2MyFalse_bufchan_d[0]) || es_10_2MyFalse_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_10_2MyFalse_bufchan_d <= 1'd0;
    else
      if (es_10_2MyFalse_r) es_10_2MyFalse_bufchan_d <= es_10_2MyFalse_d;
  MyDTInt_Int_t es_10_2MyFalse_bufchan_buf;
  assign es_10_2MyFalse_bufchan_r = (! es_10_2MyFalse_bufchan_buf[0]);
  assign es_10_2MyFalse_1_argbuf_d = (es_10_2MyFalse_bufchan_buf[0] ? es_10_2MyFalse_bufchan_buf :
                                      es_10_2MyFalse_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_10_2MyFalse_bufchan_buf <= 1'd0;
    else
      if ((es_10_2MyFalse_1_argbuf_r && es_10_2MyFalse_bufchan_buf[0]))
        es_10_2MyFalse_bufchan_buf <= 1'd0;
      else if (((! es_10_2MyFalse_1_argbuf_r) && (! es_10_2MyFalse_bufchan_buf[0])))
        es_10_2MyFalse_bufchan_buf <= es_10_2MyFalse_bufchan_d;
  
  /* demux (Ty MyBool,
       Ty Pointer_CTf_f_Int_Int) : (es_10_3,MyBool) (lizzieLet12_6QVal_Int_8QNone_Int,Pointer_CTf_f_Int_Int) > [(es_10_3MyFalse,Pointer_CTf_f_Int_Int),
                                                                                                                (es_10_3MyTrue,Pointer_CTf_f_Int_Int)] */
  logic [1:0] lizzieLet12_6QVal_Int_8QNone_Int_onehotd;
  always_comb
    if ((es_10_3_d[0] && lizzieLet12_6QVal_Int_8QNone_Int_d[0]))
      unique case (es_10_3_d[1:1])
        1'd0: lizzieLet12_6QVal_Int_8QNone_Int_onehotd = 2'd1;
        1'd1: lizzieLet12_6QVal_Int_8QNone_Int_onehotd = 2'd2;
        default: lizzieLet12_6QVal_Int_8QNone_Int_onehotd = 2'd0;
      endcase
    else lizzieLet12_6QVal_Int_8QNone_Int_onehotd = 2'd0;
  assign es_10_3MyFalse_d = {lizzieLet12_6QVal_Int_8QNone_Int_d[16:1],
                             lizzieLet12_6QVal_Int_8QNone_Int_onehotd[0]};
  assign es_10_3MyTrue_d = {lizzieLet12_6QVal_Int_8QNone_Int_d[16:1],
                            lizzieLet12_6QVal_Int_8QNone_Int_onehotd[1]};
  assign lizzieLet12_6QVal_Int_8QNone_Int_r = (| (lizzieLet12_6QVal_Int_8QNone_Int_onehotd & {es_10_3MyTrue_r,
                                                                                              es_10_3MyFalse_r}));
  assign es_10_3_r = lizzieLet12_6QVal_Int_8QNone_Int_r;
  
  /* buf (Ty Pointer_CTf_f_Int_Int) : (es_10_3MyFalse,Pointer_CTf_f_Int_Int) > (es_10_3MyFalse_1_argbuf,Pointer_CTf_f_Int_Int) */
  Pointer_CTf_f_Int_Int_t es_10_3MyFalse_bufchan_d;
  logic es_10_3MyFalse_bufchan_r;
  assign es_10_3MyFalse_r = ((! es_10_3MyFalse_bufchan_d[0]) || es_10_3MyFalse_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_10_3MyFalse_bufchan_d <= {16'd0, 1'd0};
    else
      if (es_10_3MyFalse_r) es_10_3MyFalse_bufchan_d <= es_10_3MyFalse_d;
  Pointer_CTf_f_Int_Int_t es_10_3MyFalse_bufchan_buf;
  assign es_10_3MyFalse_bufchan_r = (! es_10_3MyFalse_bufchan_buf[0]);
  assign es_10_3MyFalse_1_argbuf_d = (es_10_3MyFalse_bufchan_buf[0] ? es_10_3MyFalse_bufchan_buf :
                                      es_10_3MyFalse_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_10_3MyFalse_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((es_10_3MyFalse_1_argbuf_r && es_10_3MyFalse_bufchan_buf[0]))
        es_10_3MyFalse_bufchan_buf <= {16'd0, 1'd0};
      else if (((! es_10_3MyFalse_1_argbuf_r) && (! es_10_3MyFalse_bufchan_buf[0])))
        es_10_3MyFalse_bufchan_buf <= es_10_3MyFalse_bufchan_d;
  
  /* buf (Ty Pointer_CTf_f_Int_Int) : (es_10_3MyTrue,Pointer_CTf_f_Int_Int) > (es_10_3MyTrue_1_argbuf,Pointer_CTf_f_Int_Int) */
  Pointer_CTf_f_Int_Int_t es_10_3MyTrue_bufchan_d;
  logic es_10_3MyTrue_bufchan_r;
  assign es_10_3MyTrue_r = ((! es_10_3MyTrue_bufchan_d[0]) || es_10_3MyTrue_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_10_3MyTrue_bufchan_d <= {16'd0, 1'd0};
    else
      if (es_10_3MyTrue_r) es_10_3MyTrue_bufchan_d <= es_10_3MyTrue_d;
  Pointer_CTf_f_Int_Int_t es_10_3MyTrue_bufchan_buf;
  assign es_10_3MyTrue_bufchan_r = (! es_10_3MyTrue_bufchan_buf[0]);
  assign es_10_3MyTrue_1_argbuf_d = (es_10_3MyTrue_bufchan_buf[0] ? es_10_3MyTrue_bufchan_buf :
                                     es_10_3MyTrue_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_10_3MyTrue_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((es_10_3MyTrue_1_argbuf_r && es_10_3MyTrue_bufchan_buf[0]))
        es_10_3MyTrue_bufchan_buf <= {16'd0, 1'd0};
      else if (((! es_10_3MyTrue_1_argbuf_r) && (! es_10_3MyTrue_bufchan_buf[0])))
        es_10_3MyTrue_bufchan_buf <= es_10_3MyTrue_bufchan_d;
  
  /* demux (Ty MyBool,
       Ty Int) : (es_10_4,MyBool) (lizzieLet12_6QVal_Int_9QNone_Int_2,Int) > [(es_10_4MyFalse,Int),
                                                                              (_79,Int)] */
  logic [1:0] lizzieLet12_6QVal_Int_9QNone_Int_2_onehotd;
  always_comb
    if ((es_10_4_d[0] && lizzieLet12_6QVal_Int_9QNone_Int_2_d[0]))
      unique case (es_10_4_d[1:1])
        1'd0: lizzieLet12_6QVal_Int_9QNone_Int_2_onehotd = 2'd1;
        1'd1: lizzieLet12_6QVal_Int_9QNone_Int_2_onehotd = 2'd2;
        default: lizzieLet12_6QVal_Int_9QNone_Int_2_onehotd = 2'd0;
      endcase
    else lizzieLet12_6QVal_Int_9QNone_Int_2_onehotd = 2'd0;
  assign es_10_4MyFalse_d = {lizzieLet12_6QVal_Int_9QNone_Int_2_d[32:1],
                             lizzieLet12_6QVal_Int_9QNone_Int_2_onehotd[0]};
  assign _79_d = {lizzieLet12_6QVal_Int_9QNone_Int_2_d[32:1],
                  lizzieLet12_6QVal_Int_9QNone_Int_2_onehotd[1]};
  assign lizzieLet12_6QVal_Int_9QNone_Int_2_r = (| (lizzieLet12_6QVal_Int_9QNone_Int_2_onehotd & {_79_r,
                                                                                                  es_10_4MyFalse_r}));
  assign es_10_4_r = lizzieLet12_6QVal_Int_9QNone_Int_2_r;
  
  /* buf (Ty Int) : (es_10_4MyFalse,Int) > (es_10_4MyFalse_1_argbuf,Int) */
  Int_t es_10_4MyFalse_bufchan_d;
  logic es_10_4MyFalse_bufchan_r;
  assign es_10_4MyFalse_r = ((! es_10_4MyFalse_bufchan_d[0]) || es_10_4MyFalse_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_10_4MyFalse_bufchan_d <= {32'd0, 1'd0};
    else
      if (es_10_4MyFalse_r) es_10_4MyFalse_bufchan_d <= es_10_4MyFalse_d;
  Int_t es_10_4MyFalse_bufchan_buf;
  assign es_10_4MyFalse_bufchan_r = (! es_10_4MyFalse_bufchan_buf[0]);
  assign es_10_4MyFalse_1_argbuf_d = (es_10_4MyFalse_bufchan_buf[0] ? es_10_4MyFalse_bufchan_buf :
                                      es_10_4MyFalse_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_10_4MyFalse_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((es_10_4MyFalse_1_argbuf_r && es_10_4MyFalse_bufchan_buf[0]))
        es_10_4MyFalse_bufchan_buf <= {32'd0, 1'd0};
      else if (((! es_10_4MyFalse_1_argbuf_r) && (! es_10_4MyFalse_bufchan_buf[0])))
        es_10_4MyFalse_bufchan_buf <= es_10_4MyFalse_bufchan_d;
  
  /* buf (Ty QTree_Int) : (es_11_1QVal_Int,QTree_Int) > (lizzieLet20_1_argbuf,QTree_Int) */
  QTree_Int_t es_11_1QVal_Int_bufchan_d;
  logic es_11_1QVal_Int_bufchan_r;
  assign es_11_1QVal_Int_r = ((! es_11_1QVal_Int_bufchan_d[0]) || es_11_1QVal_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_11_1QVal_Int_bufchan_d <= {66'd0, 1'd0};
    else
      if (es_11_1QVal_Int_r)
        es_11_1QVal_Int_bufchan_d <= es_11_1QVal_Int_d;
  QTree_Int_t es_11_1QVal_Int_bufchan_buf;
  assign es_11_1QVal_Int_bufchan_r = (! es_11_1QVal_Int_bufchan_buf[0]);
  assign lizzieLet20_1_argbuf_d = (es_11_1QVal_Int_bufchan_buf[0] ? es_11_1QVal_Int_bufchan_buf :
                                   es_11_1QVal_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_11_1QVal_Int_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((lizzieLet20_1_argbuf_r && es_11_1QVal_Int_bufchan_buf[0]))
        es_11_1QVal_Int_bufchan_buf <= {66'd0, 1'd0};
      else if (((! lizzieLet20_1_argbuf_r) && (! es_11_1QVal_Int_bufchan_buf[0])))
        es_11_1QVal_Int_bufchan_buf <= es_11_1QVal_Int_bufchan_d;
  
  /* demux (Ty MyBool,
       Ty Go) : (es_14_1,MyBool) (lizzieLet12_6QVal_Int_3QVal_Int_2,Go) > [(es_14_1MyFalse,Go),
                                                                           (es_14_1MyTrue,Go)] */
  logic [1:0] lizzieLet12_6QVal_Int_3QVal_Int_2_onehotd;
  always_comb
    if ((es_14_1_d[0] && lizzieLet12_6QVal_Int_3QVal_Int_2_d[0]))
      unique case (es_14_1_d[1:1])
        1'd0: lizzieLet12_6QVal_Int_3QVal_Int_2_onehotd = 2'd1;
        1'd1: lizzieLet12_6QVal_Int_3QVal_Int_2_onehotd = 2'd2;
        default: lizzieLet12_6QVal_Int_3QVal_Int_2_onehotd = 2'd0;
      endcase
    else lizzieLet12_6QVal_Int_3QVal_Int_2_onehotd = 2'd0;
  assign es_14_1MyFalse_d = lizzieLet12_6QVal_Int_3QVal_Int_2_onehotd[0];
  assign es_14_1MyTrue_d = lizzieLet12_6QVal_Int_3QVal_Int_2_onehotd[1];
  assign lizzieLet12_6QVal_Int_3QVal_Int_2_r = (| (lizzieLet12_6QVal_Int_3QVal_Int_2_onehotd & {es_14_1MyTrue_r,
                                                                                                es_14_1MyFalse_r}));
  assign es_14_1_r = lizzieLet12_6QVal_Int_3QVal_Int_2_r;
  
  /* fork (Ty Go) : (es_14_1MyFalse,Go) > [(es_14_1MyFalse_1,Go),
                                      (es_14_1MyFalse_2,Go),
                                      (es_14_1MyFalse_3,Go)] */
  logic [2:0] es_14_1MyFalse_emitted;
  logic [2:0] es_14_1MyFalse_done;
  assign es_14_1MyFalse_1_d = (es_14_1MyFalse_d[0] && (! es_14_1MyFalse_emitted[0]));
  assign es_14_1MyFalse_2_d = (es_14_1MyFalse_d[0] && (! es_14_1MyFalse_emitted[1]));
  assign es_14_1MyFalse_3_d = (es_14_1MyFalse_d[0] && (! es_14_1MyFalse_emitted[2]));
  assign es_14_1MyFalse_done = (es_14_1MyFalse_emitted | ({es_14_1MyFalse_3_d[0],
                                                           es_14_1MyFalse_2_d[0],
                                                           es_14_1MyFalse_1_d[0]} & {es_14_1MyFalse_3_r,
                                                                                     es_14_1MyFalse_2_r,
                                                                                     es_14_1MyFalse_1_r}));
  assign es_14_1MyFalse_r = (& es_14_1MyFalse_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_14_1MyFalse_emitted <= 3'd0;
    else
      es_14_1MyFalse_emitted <= (es_14_1MyFalse_r ? 3'd0 :
                                 es_14_1MyFalse_done);
  
  /* buf (Ty Go) : (es_14_1MyFalse_1,Go) > (es_14_1MyFalse_1_argbuf,Go) */
  Go_t es_14_1MyFalse_1_bufchan_d;
  logic es_14_1MyFalse_1_bufchan_r;
  assign es_14_1MyFalse_1_r = ((! es_14_1MyFalse_1_bufchan_d[0]) || es_14_1MyFalse_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_14_1MyFalse_1_bufchan_d <= 1'd0;
    else
      if (es_14_1MyFalse_1_r)
        es_14_1MyFalse_1_bufchan_d <= es_14_1MyFalse_1_d;
  Go_t es_14_1MyFalse_1_bufchan_buf;
  assign es_14_1MyFalse_1_bufchan_r = (! es_14_1MyFalse_1_bufchan_buf[0]);
  assign es_14_1MyFalse_1_argbuf_d = (es_14_1MyFalse_1_bufchan_buf[0] ? es_14_1MyFalse_1_bufchan_buf :
                                      es_14_1MyFalse_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_14_1MyFalse_1_bufchan_buf <= 1'd0;
    else
      if ((es_14_1MyFalse_1_argbuf_r && es_14_1MyFalse_1_bufchan_buf[0]))
        es_14_1MyFalse_1_bufchan_buf <= 1'd0;
      else if (((! es_14_1MyFalse_1_argbuf_r) && (! es_14_1MyFalse_1_bufchan_buf[0])))
        es_14_1MyFalse_1_bufchan_buf <= es_14_1MyFalse_1_bufchan_d;
  
  /* dcon (Ty TupGo___MyDTInt_Int___Int,
      Dcon TupGo___MyDTInt_Int___Int) : [(es_14_1MyFalse_1_argbuf,Go),
                                         (es_14_4MyFalse_1_argbuf,MyDTInt_Int),
                                         (es_18_1_argbuf,Int)] > (applyfnInt_Int_5TupGo___MyDTInt_Int___Int7,TupGo___MyDTInt_Int___Int) */
  assign applyfnInt_Int_5TupGo___MyDTInt_Int___Int7_d = TupGo___MyDTInt_Int___Int_dc((& {es_14_1MyFalse_1_argbuf_d[0],
                                                                                         es_14_4MyFalse_1_argbuf_d[0],
                                                                                         es_18_1_argbuf_d[0]}), es_14_1MyFalse_1_argbuf_d, es_14_4MyFalse_1_argbuf_d, es_18_1_argbuf_d);
  assign {es_14_1MyFalse_1_argbuf_r,
          es_14_4MyFalse_1_argbuf_r,
          es_18_1_argbuf_r} = {3 {(applyfnInt_Int_5TupGo___MyDTInt_Int___Int7_r && applyfnInt_Int_5TupGo___MyDTInt_Int___Int7_d[0])}};
  
  /* buf (Ty Go) : (es_14_1MyFalse_2,Go) > (es_14_1MyFalse_2_argbuf,Go) */
  Go_t es_14_1MyFalse_2_bufchan_d;
  logic es_14_1MyFalse_2_bufchan_r;
  assign es_14_1MyFalse_2_r = ((! es_14_1MyFalse_2_bufchan_d[0]) || es_14_1MyFalse_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_14_1MyFalse_2_bufchan_d <= 1'd0;
    else
      if (es_14_1MyFalse_2_r)
        es_14_1MyFalse_2_bufchan_d <= es_14_1MyFalse_2_d;
  Go_t es_14_1MyFalse_2_bufchan_buf;
  assign es_14_1MyFalse_2_bufchan_r = (! es_14_1MyFalse_2_bufchan_buf[0]);
  assign es_14_1MyFalse_2_argbuf_d = (es_14_1MyFalse_2_bufchan_buf[0] ? es_14_1MyFalse_2_bufchan_buf :
                                      es_14_1MyFalse_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_14_1MyFalse_2_bufchan_buf <= 1'd0;
    else
      if ((es_14_1MyFalse_2_argbuf_r && es_14_1MyFalse_2_bufchan_buf[0]))
        es_14_1MyFalse_2_bufchan_buf <= 1'd0;
      else if (((! es_14_1MyFalse_2_argbuf_r) && (! es_14_1MyFalse_2_bufchan_buf[0])))
        es_14_1MyFalse_2_bufchan_buf <= es_14_1MyFalse_2_bufchan_d;
  
  /* dcon (Ty TupGo___MyDTInt_Bool___Int,
      Dcon TupGo___MyDTInt_Bool___Int) : [(es_14_1MyFalse_2_argbuf,Go),
                                          (es_14_2MyFalse_1_argbuf,MyDTInt_Bool),
                                          (es_16_1_argbuf,Int)] > (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int5,TupGo___MyDTInt_Bool___Int) */
  assign applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int5_d = TupGo___MyDTInt_Bool___Int_dc((& {es_14_1MyFalse_2_argbuf_d[0],
                                                                                            es_14_2MyFalse_1_argbuf_d[0],
                                                                                            es_16_1_argbuf_d[0]}), es_14_1MyFalse_2_argbuf_d, es_14_2MyFalse_1_argbuf_d, es_16_1_argbuf_d);
  assign {es_14_1MyFalse_2_argbuf_r,
          es_14_2MyFalse_1_argbuf_r,
          es_16_1_argbuf_r} = {3 {(applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int5_r && applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int5_d[0])}};
  
  /* fork (Ty Go) : (es_14_1MyTrue,Go) > [(es_14_1MyTrue_1,Go),
                                     (es_14_1MyTrue_2,Go)] */
  logic [1:0] es_14_1MyTrue_emitted;
  logic [1:0] es_14_1MyTrue_done;
  assign es_14_1MyTrue_1_d = (es_14_1MyTrue_d[0] && (! es_14_1MyTrue_emitted[0]));
  assign es_14_1MyTrue_2_d = (es_14_1MyTrue_d[0] && (! es_14_1MyTrue_emitted[1]));
  assign es_14_1MyTrue_done = (es_14_1MyTrue_emitted | ({es_14_1MyTrue_2_d[0],
                                                         es_14_1MyTrue_1_d[0]} & {es_14_1MyTrue_2_r,
                                                                                  es_14_1MyTrue_1_r}));
  assign es_14_1MyTrue_r = (& es_14_1MyTrue_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_14_1MyTrue_emitted <= 2'd0;
    else
      es_14_1MyTrue_emitted <= (es_14_1MyTrue_r ? 2'd0 :
                                es_14_1MyTrue_done);
  
  /* dcon (Ty QTree_Int,
      Dcon QNone_Int) : [(es_14_1MyTrue_1,Go)] > (es_14_1MyTrue_1QNone_Int,QTree_Int) */
  assign es_14_1MyTrue_1QNone_Int_d = QNone_Int_dc((& {es_14_1MyTrue_1_d[0]}), es_14_1MyTrue_1_d);
  assign {es_14_1MyTrue_1_r} = {1 {(es_14_1MyTrue_1QNone_Int_r && es_14_1MyTrue_1QNone_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (es_14_1MyTrue_1QNone_Int,QTree_Int) > (lizzieLet24_1_1_argbuf,QTree_Int) */
  QTree_Int_t es_14_1MyTrue_1QNone_Int_bufchan_d;
  logic es_14_1MyTrue_1QNone_Int_bufchan_r;
  assign es_14_1MyTrue_1QNone_Int_r = ((! es_14_1MyTrue_1QNone_Int_bufchan_d[0]) || es_14_1MyTrue_1QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_14_1MyTrue_1QNone_Int_bufchan_d <= {66'd0, 1'd0};
    else
      if (es_14_1MyTrue_1QNone_Int_r)
        es_14_1MyTrue_1QNone_Int_bufchan_d <= es_14_1MyTrue_1QNone_Int_d;
  QTree_Int_t es_14_1MyTrue_1QNone_Int_bufchan_buf;
  assign es_14_1MyTrue_1QNone_Int_bufchan_r = (! es_14_1MyTrue_1QNone_Int_bufchan_buf[0]);
  assign lizzieLet24_1_1_argbuf_d = (es_14_1MyTrue_1QNone_Int_bufchan_buf[0] ? es_14_1MyTrue_1QNone_Int_bufchan_buf :
                                     es_14_1MyTrue_1QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_14_1MyTrue_1QNone_Int_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((lizzieLet24_1_1_argbuf_r && es_14_1MyTrue_1QNone_Int_bufchan_buf[0]))
        es_14_1MyTrue_1QNone_Int_bufchan_buf <= {66'd0, 1'd0};
      else if (((! lizzieLet24_1_1_argbuf_r) && (! es_14_1MyTrue_1QNone_Int_bufchan_buf[0])))
        es_14_1MyTrue_1QNone_Int_bufchan_buf <= es_14_1MyTrue_1QNone_Int_bufchan_d;
  
  /* buf (Ty Go) : (es_14_1MyTrue_2,Go) > (es_14_1MyTrue_2_argbuf,Go) */
  Go_t es_14_1MyTrue_2_bufchan_d;
  logic es_14_1MyTrue_2_bufchan_r;
  assign es_14_1MyTrue_2_r = ((! es_14_1MyTrue_2_bufchan_d[0]) || es_14_1MyTrue_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_14_1MyTrue_2_bufchan_d <= 1'd0;
    else
      if (es_14_1MyTrue_2_r)
        es_14_1MyTrue_2_bufchan_d <= es_14_1MyTrue_2_d;
  Go_t es_14_1MyTrue_2_bufchan_buf;
  assign es_14_1MyTrue_2_bufchan_r = (! es_14_1MyTrue_2_bufchan_buf[0]);
  assign es_14_1MyTrue_2_argbuf_d = (es_14_1MyTrue_2_bufchan_buf[0] ? es_14_1MyTrue_2_bufchan_buf :
                                     es_14_1MyTrue_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_14_1MyTrue_2_bufchan_buf <= 1'd0;
    else
      if ((es_14_1MyTrue_2_argbuf_r && es_14_1MyTrue_2_bufchan_buf[0]))
        es_14_1MyTrue_2_bufchan_buf <= 1'd0;
      else if (((! es_14_1MyTrue_2_argbuf_r) && (! es_14_1MyTrue_2_bufchan_buf[0])))
        es_14_1MyTrue_2_bufchan_buf <= es_14_1MyTrue_2_bufchan_d;
  
  /* demux (Ty MyBool,
       Ty MyDTInt_Bool) : (es_14_2,MyBool) (lizzieLet12_6QVal_Int_5QVal_Int,MyDTInt_Bool) > [(es_14_2MyFalse,MyDTInt_Bool),
                                                                                             (_78,MyDTInt_Bool)] */
  logic [1:0] lizzieLet12_6QVal_Int_5QVal_Int_onehotd;
  always_comb
    if ((es_14_2_d[0] && lizzieLet12_6QVal_Int_5QVal_Int_d[0]))
      unique case (es_14_2_d[1:1])
        1'd0: lizzieLet12_6QVal_Int_5QVal_Int_onehotd = 2'd1;
        1'd1: lizzieLet12_6QVal_Int_5QVal_Int_onehotd = 2'd2;
        default: lizzieLet12_6QVal_Int_5QVal_Int_onehotd = 2'd0;
      endcase
    else lizzieLet12_6QVal_Int_5QVal_Int_onehotd = 2'd0;
  assign es_14_2MyFalse_d = lizzieLet12_6QVal_Int_5QVal_Int_onehotd[0];
  assign _78_d = lizzieLet12_6QVal_Int_5QVal_Int_onehotd[1];
  assign lizzieLet12_6QVal_Int_5QVal_Int_r = (| (lizzieLet12_6QVal_Int_5QVal_Int_onehotd & {_78_r,
                                                                                            es_14_2MyFalse_r}));
  assign es_14_2_r = lizzieLet12_6QVal_Int_5QVal_Int_r;
  
  /* buf (Ty MyDTInt_Bool) : (es_14_2MyFalse,MyDTInt_Bool) > (es_14_2MyFalse_1_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t es_14_2MyFalse_bufchan_d;
  logic es_14_2MyFalse_bufchan_r;
  assign es_14_2MyFalse_r = ((! es_14_2MyFalse_bufchan_d[0]) || es_14_2MyFalse_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_14_2MyFalse_bufchan_d <= 1'd0;
    else
      if (es_14_2MyFalse_r) es_14_2MyFalse_bufchan_d <= es_14_2MyFalse_d;
  MyDTInt_Bool_t es_14_2MyFalse_bufchan_buf;
  assign es_14_2MyFalse_bufchan_r = (! es_14_2MyFalse_bufchan_buf[0]);
  assign es_14_2MyFalse_1_argbuf_d = (es_14_2MyFalse_bufchan_buf[0] ? es_14_2MyFalse_bufchan_buf :
                                      es_14_2MyFalse_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_14_2MyFalse_bufchan_buf <= 1'd0;
    else
      if ((es_14_2MyFalse_1_argbuf_r && es_14_2MyFalse_bufchan_buf[0]))
        es_14_2MyFalse_bufchan_buf <= 1'd0;
      else if (((! es_14_2MyFalse_1_argbuf_r) && (! es_14_2MyFalse_bufchan_buf[0])))
        es_14_2MyFalse_bufchan_buf <= es_14_2MyFalse_bufchan_d;
  
  /* demux (Ty MyBool,
       Ty MyDTInt_Int_Int) : (es_14_3,MyBool) (lizzieLet12_6QVal_Int_6QVal_Int_2,MyDTInt_Int_Int) > [(es_14_3MyFalse,MyDTInt_Int_Int),
                                                                                                     (_77,MyDTInt_Int_Int)] */
  logic [1:0] lizzieLet12_6QVal_Int_6QVal_Int_2_onehotd;
  always_comb
    if ((es_14_3_d[0] && lizzieLet12_6QVal_Int_6QVal_Int_2_d[0]))
      unique case (es_14_3_d[1:1])
        1'd0: lizzieLet12_6QVal_Int_6QVal_Int_2_onehotd = 2'd1;
        1'd1: lizzieLet12_6QVal_Int_6QVal_Int_2_onehotd = 2'd2;
        default: lizzieLet12_6QVal_Int_6QVal_Int_2_onehotd = 2'd0;
      endcase
    else lizzieLet12_6QVal_Int_6QVal_Int_2_onehotd = 2'd0;
  assign es_14_3MyFalse_d = lizzieLet12_6QVal_Int_6QVal_Int_2_onehotd[0];
  assign _77_d = lizzieLet12_6QVal_Int_6QVal_Int_2_onehotd[1];
  assign lizzieLet12_6QVal_Int_6QVal_Int_2_r = (| (lizzieLet12_6QVal_Int_6QVal_Int_2_onehotd & {_77_r,
                                                                                                es_14_3MyFalse_r}));
  assign es_14_3_r = lizzieLet12_6QVal_Int_6QVal_Int_2_r;
  
  /* fork (Ty MyDTInt_Int_Int) : (es_14_3MyFalse,MyDTInt_Int_Int) > [(es_14_3MyFalse_1,MyDTInt_Int_Int),
                                                                (es_14_3MyFalse_2,MyDTInt_Int_Int)] */
  logic [1:0] es_14_3MyFalse_emitted;
  logic [1:0] es_14_3MyFalse_done;
  assign es_14_3MyFalse_1_d = (es_14_3MyFalse_d[0] && (! es_14_3MyFalse_emitted[0]));
  assign es_14_3MyFalse_2_d = (es_14_3MyFalse_d[0] && (! es_14_3MyFalse_emitted[1]));
  assign es_14_3MyFalse_done = (es_14_3MyFalse_emitted | ({es_14_3MyFalse_2_d[0],
                                                           es_14_3MyFalse_1_d[0]} & {es_14_3MyFalse_2_r,
                                                                                     es_14_3MyFalse_1_r}));
  assign es_14_3MyFalse_r = (& es_14_3MyFalse_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_14_3MyFalse_emitted <= 2'd0;
    else
      es_14_3MyFalse_emitted <= (es_14_3MyFalse_r ? 2'd0 :
                                 es_14_3MyFalse_done);
  
  /* buf (Ty MyDTInt_Int_Int) : (es_14_3MyFalse_1,MyDTInt_Int_Int) > (es_14_3MyFalse_1_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t es_14_3MyFalse_1_bufchan_d;
  logic es_14_3MyFalse_1_bufchan_r;
  assign es_14_3MyFalse_1_r = ((! es_14_3MyFalse_1_bufchan_d[0]) || es_14_3MyFalse_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_14_3MyFalse_1_bufchan_d <= 1'd0;
    else
      if (es_14_3MyFalse_1_r)
        es_14_3MyFalse_1_bufchan_d <= es_14_3MyFalse_1_d;
  MyDTInt_Int_Int_t es_14_3MyFalse_1_bufchan_buf;
  assign es_14_3MyFalse_1_bufchan_r = (! es_14_3MyFalse_1_bufchan_buf[0]);
  assign es_14_3MyFalse_1_argbuf_d = (es_14_3MyFalse_1_bufchan_buf[0] ? es_14_3MyFalse_1_bufchan_buf :
                                      es_14_3MyFalse_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_14_3MyFalse_1_bufchan_buf <= 1'd0;
    else
      if ((es_14_3MyFalse_1_argbuf_r && es_14_3MyFalse_1_bufchan_buf[0]))
        es_14_3MyFalse_1_bufchan_buf <= 1'd0;
      else if (((! es_14_3MyFalse_1_argbuf_r) && (! es_14_3MyFalse_1_bufchan_buf[0])))
        es_14_3MyFalse_1_bufchan_buf <= es_14_3MyFalse_1_bufchan_d;
  
  /* dcon (Ty TupMyDTInt_Int_Int___Int___Int,
      Dcon TupMyDTInt_Int_Int___Int___Int) : [(es_14_3MyFalse_1_argbuf,MyDTInt_Int_Int),
                                              (es_14_6MyFalse_1_argbuf,Int),
                                              (es_14_7MyFalse_1_argbuf,Int)] > (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int2,TupMyDTInt_Int_Int___Int___Int) */
  assign applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int2_d = TupMyDTInt_Int_Int___Int___Int_dc((& {es_14_3MyFalse_1_argbuf_d[0],
                                                                                                       es_14_6MyFalse_1_argbuf_d[0],
                                                                                                       es_14_7MyFalse_1_argbuf_d[0]}), es_14_3MyFalse_1_argbuf_d, es_14_6MyFalse_1_argbuf_d, es_14_7MyFalse_1_argbuf_d);
  assign {es_14_3MyFalse_1_argbuf_r,
          es_14_6MyFalse_1_argbuf_r,
          es_14_7MyFalse_1_argbuf_r} = {3 {(applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int2_r && applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int2_d[0])}};
  
  /* demux (Ty MyBool,
       Ty MyDTInt_Int) : (es_14_4,MyBool) (lizzieLet12_6QVal_Int_7QVal_Int,MyDTInt_Int) > [(es_14_4MyFalse,MyDTInt_Int),
                                                                                           (_76,MyDTInt_Int)] */
  logic [1:0] lizzieLet12_6QVal_Int_7QVal_Int_onehotd;
  always_comb
    if ((es_14_4_d[0] && lizzieLet12_6QVal_Int_7QVal_Int_d[0]))
      unique case (es_14_4_d[1:1])
        1'd0: lizzieLet12_6QVal_Int_7QVal_Int_onehotd = 2'd1;
        1'd1: lizzieLet12_6QVal_Int_7QVal_Int_onehotd = 2'd2;
        default: lizzieLet12_6QVal_Int_7QVal_Int_onehotd = 2'd0;
      endcase
    else lizzieLet12_6QVal_Int_7QVal_Int_onehotd = 2'd0;
  assign es_14_4MyFalse_d = lizzieLet12_6QVal_Int_7QVal_Int_onehotd[0];
  assign _76_d = lizzieLet12_6QVal_Int_7QVal_Int_onehotd[1];
  assign lizzieLet12_6QVal_Int_7QVal_Int_r = (| (lizzieLet12_6QVal_Int_7QVal_Int_onehotd & {_76_r,
                                                                                            es_14_4MyFalse_r}));
  assign es_14_4_r = lizzieLet12_6QVal_Int_7QVal_Int_r;
  
  /* fork (Ty MyDTInt_Int) : (es_14_4MyFalse,MyDTInt_Int) > [(es_14_4MyFalse_1,MyDTInt_Int),
                                                        (es_14_4MyFalse_2,MyDTInt_Int)] */
  logic [1:0] es_14_4MyFalse_emitted;
  logic [1:0] es_14_4MyFalse_done;
  assign es_14_4MyFalse_1_d = (es_14_4MyFalse_d[0] && (! es_14_4MyFalse_emitted[0]));
  assign es_14_4MyFalse_2_d = (es_14_4MyFalse_d[0] && (! es_14_4MyFalse_emitted[1]));
  assign es_14_4MyFalse_done = (es_14_4MyFalse_emitted | ({es_14_4MyFalse_2_d[0],
                                                           es_14_4MyFalse_1_d[0]} & {es_14_4MyFalse_2_r,
                                                                                     es_14_4MyFalse_1_r}));
  assign es_14_4MyFalse_r = (& es_14_4MyFalse_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_14_4MyFalse_emitted <= 2'd0;
    else
      es_14_4MyFalse_emitted <= (es_14_4MyFalse_r ? 2'd0 :
                                 es_14_4MyFalse_done);
  
  /* buf (Ty MyDTInt_Int) : (es_14_4MyFalse_1,MyDTInt_Int) > (es_14_4MyFalse_1_argbuf,MyDTInt_Int) */
  MyDTInt_Int_t es_14_4MyFalse_1_bufchan_d;
  logic es_14_4MyFalse_1_bufchan_r;
  assign es_14_4MyFalse_1_r = ((! es_14_4MyFalse_1_bufchan_d[0]) || es_14_4MyFalse_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_14_4MyFalse_1_bufchan_d <= 1'd0;
    else
      if (es_14_4MyFalse_1_r)
        es_14_4MyFalse_1_bufchan_d <= es_14_4MyFalse_1_d;
  MyDTInt_Int_t es_14_4MyFalse_1_bufchan_buf;
  assign es_14_4MyFalse_1_bufchan_r = (! es_14_4MyFalse_1_bufchan_buf[0]);
  assign es_14_4MyFalse_1_argbuf_d = (es_14_4MyFalse_1_bufchan_buf[0] ? es_14_4MyFalse_1_bufchan_buf :
                                      es_14_4MyFalse_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_14_4MyFalse_1_bufchan_buf <= 1'd0;
    else
      if ((es_14_4MyFalse_1_argbuf_r && es_14_4MyFalse_1_bufchan_buf[0]))
        es_14_4MyFalse_1_bufchan_buf <= 1'd0;
      else if (((! es_14_4MyFalse_1_argbuf_r) && (! es_14_4MyFalse_1_bufchan_buf[0])))
        es_14_4MyFalse_1_bufchan_buf <= es_14_4MyFalse_1_bufchan_d;
  
  /* demux (Ty MyBool,
       Ty Pointer_CTf_f_Int_Int) : (es_14_5,MyBool) (lizzieLet12_6QVal_Int_8QVal_Int,Pointer_CTf_f_Int_Int) > [(es_14_5MyFalse,Pointer_CTf_f_Int_Int),
                                                                                                               (es_14_5MyTrue,Pointer_CTf_f_Int_Int)] */
  logic [1:0] lizzieLet12_6QVal_Int_8QVal_Int_onehotd;
  always_comb
    if ((es_14_5_d[0] && lizzieLet12_6QVal_Int_8QVal_Int_d[0]))
      unique case (es_14_5_d[1:1])
        1'd0: lizzieLet12_6QVal_Int_8QVal_Int_onehotd = 2'd1;
        1'd1: lizzieLet12_6QVal_Int_8QVal_Int_onehotd = 2'd2;
        default: lizzieLet12_6QVal_Int_8QVal_Int_onehotd = 2'd0;
      endcase
    else lizzieLet12_6QVal_Int_8QVal_Int_onehotd = 2'd0;
  assign es_14_5MyFalse_d = {lizzieLet12_6QVal_Int_8QVal_Int_d[16:1],
                             lizzieLet12_6QVal_Int_8QVal_Int_onehotd[0]};
  assign es_14_5MyTrue_d = {lizzieLet12_6QVal_Int_8QVal_Int_d[16:1],
                            lizzieLet12_6QVal_Int_8QVal_Int_onehotd[1]};
  assign lizzieLet12_6QVal_Int_8QVal_Int_r = (| (lizzieLet12_6QVal_Int_8QVal_Int_onehotd & {es_14_5MyTrue_r,
                                                                                            es_14_5MyFalse_r}));
  assign es_14_5_r = lizzieLet12_6QVal_Int_8QVal_Int_r;
  
  /* buf (Ty Pointer_CTf_f_Int_Int) : (es_14_5MyTrue,Pointer_CTf_f_Int_Int) > (es_14_5MyTrue_1_argbuf,Pointer_CTf_f_Int_Int) */
  Pointer_CTf_f_Int_Int_t es_14_5MyTrue_bufchan_d;
  logic es_14_5MyTrue_bufchan_r;
  assign es_14_5MyTrue_r = ((! es_14_5MyTrue_bufchan_d[0]) || es_14_5MyTrue_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_14_5MyTrue_bufchan_d <= {16'd0, 1'd0};
    else
      if (es_14_5MyTrue_r) es_14_5MyTrue_bufchan_d <= es_14_5MyTrue_d;
  Pointer_CTf_f_Int_Int_t es_14_5MyTrue_bufchan_buf;
  assign es_14_5MyTrue_bufchan_r = (! es_14_5MyTrue_bufchan_buf[0]);
  assign es_14_5MyTrue_1_argbuf_d = (es_14_5MyTrue_bufchan_buf[0] ? es_14_5MyTrue_bufchan_buf :
                                     es_14_5MyTrue_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_14_5MyTrue_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((es_14_5MyTrue_1_argbuf_r && es_14_5MyTrue_bufchan_buf[0]))
        es_14_5MyTrue_bufchan_buf <= {16'd0, 1'd0};
      else if (((! es_14_5MyTrue_1_argbuf_r) && (! es_14_5MyTrue_bufchan_buf[0])))
        es_14_5MyTrue_bufchan_buf <= es_14_5MyTrue_bufchan_d;
  
  /* demux (Ty MyBool,
       Ty Int) : (es_14_6,MyBool) (lizzieLet12_6QVal_Int_9QVal_Int_2,Int) > [(es_14_6MyFalse,Int),
                                                                             (_75,Int)] */
  logic [1:0] lizzieLet12_6QVal_Int_9QVal_Int_2_onehotd;
  always_comb
    if ((es_14_6_d[0] && lizzieLet12_6QVal_Int_9QVal_Int_2_d[0]))
      unique case (es_14_6_d[1:1])
        1'd0: lizzieLet12_6QVal_Int_9QVal_Int_2_onehotd = 2'd1;
        1'd1: lizzieLet12_6QVal_Int_9QVal_Int_2_onehotd = 2'd2;
        default: lizzieLet12_6QVal_Int_9QVal_Int_2_onehotd = 2'd0;
      endcase
    else lizzieLet12_6QVal_Int_9QVal_Int_2_onehotd = 2'd0;
  assign es_14_6MyFalse_d = {lizzieLet12_6QVal_Int_9QVal_Int_2_d[32:1],
                             lizzieLet12_6QVal_Int_9QVal_Int_2_onehotd[0]};
  assign _75_d = {lizzieLet12_6QVal_Int_9QVal_Int_2_d[32:1],
                  lizzieLet12_6QVal_Int_9QVal_Int_2_onehotd[1]};
  assign lizzieLet12_6QVal_Int_9QVal_Int_2_r = (| (lizzieLet12_6QVal_Int_9QVal_Int_2_onehotd & {_75_r,
                                                                                                es_14_6MyFalse_r}));
  assign es_14_6_r = lizzieLet12_6QVal_Int_9QVal_Int_2_r;
  
  /* fork (Ty Int) : (es_14_6MyFalse,Int) > [(es_14_6MyFalse_1,Int),
                                        (es_14_6MyFalse_2,Int)] */
  logic [1:0] es_14_6MyFalse_emitted;
  logic [1:0] es_14_6MyFalse_done;
  assign es_14_6MyFalse_1_d = {es_14_6MyFalse_d[32:1],
                               (es_14_6MyFalse_d[0] && (! es_14_6MyFalse_emitted[0]))};
  assign es_14_6MyFalse_2_d = {es_14_6MyFalse_d[32:1],
                               (es_14_6MyFalse_d[0] && (! es_14_6MyFalse_emitted[1]))};
  assign es_14_6MyFalse_done = (es_14_6MyFalse_emitted | ({es_14_6MyFalse_2_d[0],
                                                           es_14_6MyFalse_1_d[0]} & {es_14_6MyFalse_2_r,
                                                                                     es_14_6MyFalse_1_r}));
  assign es_14_6MyFalse_r = (& es_14_6MyFalse_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_14_6MyFalse_emitted <= 2'd0;
    else
      es_14_6MyFalse_emitted <= (es_14_6MyFalse_r ? 2'd0 :
                                 es_14_6MyFalse_done);
  
  /* buf (Ty Int) : (es_14_6MyFalse_1,Int) > (es_14_6MyFalse_1_argbuf,Int) */
  Int_t es_14_6MyFalse_1_bufchan_d;
  logic es_14_6MyFalse_1_bufchan_r;
  assign es_14_6MyFalse_1_r = ((! es_14_6MyFalse_1_bufchan_d[0]) || es_14_6MyFalse_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_14_6MyFalse_1_bufchan_d <= {32'd0, 1'd0};
    else
      if (es_14_6MyFalse_1_r)
        es_14_6MyFalse_1_bufchan_d <= es_14_6MyFalse_1_d;
  Int_t es_14_6MyFalse_1_bufchan_buf;
  assign es_14_6MyFalse_1_bufchan_r = (! es_14_6MyFalse_1_bufchan_buf[0]);
  assign es_14_6MyFalse_1_argbuf_d = (es_14_6MyFalse_1_bufchan_buf[0] ? es_14_6MyFalse_1_bufchan_buf :
                                      es_14_6MyFalse_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_14_6MyFalse_1_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((es_14_6MyFalse_1_argbuf_r && es_14_6MyFalse_1_bufchan_buf[0]))
        es_14_6MyFalse_1_bufchan_buf <= {32'd0, 1'd0};
      else if (((! es_14_6MyFalse_1_argbuf_r) && (! es_14_6MyFalse_1_bufchan_buf[0])))
        es_14_6MyFalse_1_bufchan_buf <= es_14_6MyFalse_1_bufchan_d;
  
  /* demux (Ty MyBool,
       Ty Int) : (es_14_7,MyBool) (va8O_2,Int) > [(es_14_7MyFalse,Int),
                                                  (_74,Int)] */
  logic [1:0] va8O_2_onehotd;
  always_comb
    if ((es_14_7_d[0] && va8O_2_d[0]))
      unique case (es_14_7_d[1:1])
        1'd0: va8O_2_onehotd = 2'd1;
        1'd1: va8O_2_onehotd = 2'd2;
        default: va8O_2_onehotd = 2'd0;
      endcase
    else va8O_2_onehotd = 2'd0;
  assign es_14_7MyFalse_d = {va8O_2_d[32:1], va8O_2_onehotd[0]};
  assign _74_d = {va8O_2_d[32:1], va8O_2_onehotd[1]};
  assign va8O_2_r = (| (va8O_2_onehotd & {_74_r, es_14_7MyFalse_r}));
  assign es_14_7_r = va8O_2_r;
  
  /* fork (Ty Int) : (es_14_7MyFalse,Int) > [(es_14_7MyFalse_1,Int),
                                        (es_14_7MyFalse_2,Int)] */
  logic [1:0] es_14_7MyFalse_emitted;
  logic [1:0] es_14_7MyFalse_done;
  assign es_14_7MyFalse_1_d = {es_14_7MyFalse_d[32:1],
                               (es_14_7MyFalse_d[0] && (! es_14_7MyFalse_emitted[0]))};
  assign es_14_7MyFalse_2_d = {es_14_7MyFalse_d[32:1],
                               (es_14_7MyFalse_d[0] && (! es_14_7MyFalse_emitted[1]))};
  assign es_14_7MyFalse_done = (es_14_7MyFalse_emitted | ({es_14_7MyFalse_2_d[0],
                                                           es_14_7MyFalse_1_d[0]} & {es_14_7MyFalse_2_r,
                                                                                     es_14_7MyFalse_1_r}));
  assign es_14_7MyFalse_r = (& es_14_7MyFalse_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_14_7MyFalse_emitted <= 2'd0;
    else
      es_14_7MyFalse_emitted <= (es_14_7MyFalse_r ? 2'd0 :
                                 es_14_7MyFalse_done);
  
  /* buf (Ty Int) : (es_14_7MyFalse_1,Int) > (es_14_7MyFalse_1_argbuf,Int) */
  Int_t es_14_7MyFalse_1_bufchan_d;
  logic es_14_7MyFalse_1_bufchan_r;
  assign es_14_7MyFalse_1_r = ((! es_14_7MyFalse_1_bufchan_d[0]) || es_14_7MyFalse_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_14_7MyFalse_1_bufchan_d <= {32'd0, 1'd0};
    else
      if (es_14_7MyFalse_1_r)
        es_14_7MyFalse_1_bufchan_d <= es_14_7MyFalse_1_d;
  Int_t es_14_7MyFalse_1_bufchan_buf;
  assign es_14_7MyFalse_1_bufchan_r = (! es_14_7MyFalse_1_bufchan_buf[0]);
  assign es_14_7MyFalse_1_argbuf_d = (es_14_7MyFalse_1_bufchan_buf[0] ? es_14_7MyFalse_1_bufchan_buf :
                                      es_14_7MyFalse_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_14_7MyFalse_1_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((es_14_7MyFalse_1_argbuf_r && es_14_7MyFalse_1_bufchan_buf[0]))
        es_14_7MyFalse_1_bufchan_buf <= {32'd0, 1'd0};
      else if (((! es_14_7MyFalse_1_argbuf_r) && (! es_14_7MyFalse_1_bufchan_buf[0])))
        es_14_7MyFalse_1_bufchan_buf <= es_14_7MyFalse_1_bufchan_d;
  
  /* demux (Ty MyBool,
       Ty Go) : (es_19_1,MyBool) (es_14_1MyFalse_3,Go) > [(es_19_1MyFalse,Go),
                                                          (es_19_1MyTrue,Go)] */
  logic [1:0] es_14_1MyFalse_3_onehotd;
  always_comb
    if ((es_19_1_d[0] && es_14_1MyFalse_3_d[0]))
      unique case (es_19_1_d[1:1])
        1'd0: es_14_1MyFalse_3_onehotd = 2'd1;
        1'd1: es_14_1MyFalse_3_onehotd = 2'd2;
        default: es_14_1MyFalse_3_onehotd = 2'd0;
      endcase
    else es_14_1MyFalse_3_onehotd = 2'd0;
  assign es_19_1MyFalse_d = es_14_1MyFalse_3_onehotd[0];
  assign es_19_1MyTrue_d = es_14_1MyFalse_3_onehotd[1];
  assign es_14_1MyFalse_3_r = (| (es_14_1MyFalse_3_onehotd & {es_19_1MyTrue_r,
                                                              es_19_1MyFalse_r}));
  assign es_19_1_r = es_14_1MyFalse_3_r;
  
  /* fork (Ty Go) : (es_19_1MyFalse,Go) > [(es_19_1MyFalse_1,Go),
                                      (es_19_1MyFalse_2,Go)] */
  logic [1:0] es_19_1MyFalse_emitted;
  logic [1:0] es_19_1MyFalse_done;
  assign es_19_1MyFalse_1_d = (es_19_1MyFalse_d[0] && (! es_19_1MyFalse_emitted[0]));
  assign es_19_1MyFalse_2_d = (es_19_1MyFalse_d[0] && (! es_19_1MyFalse_emitted[1]));
  assign es_19_1MyFalse_done = (es_19_1MyFalse_emitted | ({es_19_1MyFalse_2_d[0],
                                                           es_19_1MyFalse_1_d[0]} & {es_19_1MyFalse_2_r,
                                                                                     es_19_1MyFalse_1_r}));
  assign es_19_1MyFalse_r = (& es_19_1MyFalse_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_19_1MyFalse_emitted <= 2'd0;
    else
      es_19_1MyFalse_emitted <= (es_19_1MyFalse_r ? 2'd0 :
                                 es_19_1MyFalse_done);
  
  /* buf (Ty Go) : (es_19_1MyFalse_1,Go) > (es_19_1MyFalse_1_argbuf,Go) */
  Go_t es_19_1MyFalse_1_bufchan_d;
  logic es_19_1MyFalse_1_bufchan_r;
  assign es_19_1MyFalse_1_r = ((! es_19_1MyFalse_1_bufchan_d[0]) || es_19_1MyFalse_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_19_1MyFalse_1_bufchan_d <= 1'd0;
    else
      if (es_19_1MyFalse_1_r)
        es_19_1MyFalse_1_bufchan_d <= es_19_1MyFalse_1_d;
  Go_t es_19_1MyFalse_1_bufchan_buf;
  assign es_19_1MyFalse_1_bufchan_r = (! es_19_1MyFalse_1_bufchan_buf[0]);
  assign es_19_1MyFalse_1_argbuf_d = (es_19_1MyFalse_1_bufchan_buf[0] ? es_19_1MyFalse_1_bufchan_buf :
                                      es_19_1MyFalse_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_19_1MyFalse_1_bufchan_buf <= 1'd0;
    else
      if ((es_19_1MyFalse_1_argbuf_r && es_19_1MyFalse_1_bufchan_buf[0]))
        es_19_1MyFalse_1_bufchan_buf <= 1'd0;
      else if (((! es_19_1MyFalse_1_argbuf_r) && (! es_19_1MyFalse_1_bufchan_buf[0])))
        es_19_1MyFalse_1_bufchan_buf <= es_19_1MyFalse_1_bufchan_d;
  
  /* dcon (Ty TupGo___MyDTInt_Int___Int,
      Dcon TupGo___MyDTInt_Int___Int) : [(es_19_1MyFalse_1_argbuf,Go),
                                         (es_19_3MyFalse_1_argbuf,MyDTInt_Int),
                                         (es_22_1_argbuf,Int)] > (applyfnInt_Int_5TupGo___MyDTInt_Int___Int8,TupGo___MyDTInt_Int___Int) */
  assign applyfnInt_Int_5TupGo___MyDTInt_Int___Int8_d = TupGo___MyDTInt_Int___Int_dc((& {es_19_1MyFalse_1_argbuf_d[0],
                                                                                         es_19_3MyFalse_1_argbuf_d[0],
                                                                                         es_22_1_argbuf_d[0]}), es_19_1MyFalse_1_argbuf_d, es_19_3MyFalse_1_argbuf_d, es_22_1_argbuf_d);
  assign {es_19_1MyFalse_1_argbuf_r,
          es_19_3MyFalse_1_argbuf_r,
          es_22_1_argbuf_r} = {3 {(applyfnInt_Int_5TupGo___MyDTInt_Int___Int8_r && applyfnInt_Int_5TupGo___MyDTInt_Int___Int8_d[0])}};
  
  /* buf (Ty Go) : (es_19_1MyFalse_2,Go) > (es_19_1MyFalse_2_argbuf,Go) */
  Go_t es_19_1MyFalse_2_bufchan_d;
  logic es_19_1MyFalse_2_bufchan_r;
  assign es_19_1MyFalse_2_r = ((! es_19_1MyFalse_2_bufchan_d[0]) || es_19_1MyFalse_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_19_1MyFalse_2_bufchan_d <= 1'd0;
    else
      if (es_19_1MyFalse_2_r)
        es_19_1MyFalse_2_bufchan_d <= es_19_1MyFalse_2_d;
  Go_t es_19_1MyFalse_2_bufchan_buf;
  assign es_19_1MyFalse_2_bufchan_r = (! es_19_1MyFalse_2_bufchan_buf[0]);
  assign es_19_1MyFalse_2_argbuf_d = (es_19_1MyFalse_2_bufchan_buf[0] ? es_19_1MyFalse_2_bufchan_buf :
                                      es_19_1MyFalse_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_19_1MyFalse_2_bufchan_buf <= 1'd0;
    else
      if ((es_19_1MyFalse_2_argbuf_r && es_19_1MyFalse_2_bufchan_buf[0]))
        es_19_1MyFalse_2_bufchan_buf <= 1'd0;
      else if (((! es_19_1MyFalse_2_argbuf_r) && (! es_19_1MyFalse_2_bufchan_buf[0])))
        es_19_1MyFalse_2_bufchan_buf <= es_19_1MyFalse_2_bufchan_d;
  
  /* fork (Ty Go) : (es_19_1MyTrue,Go) > [(es_19_1MyTrue_1,Go),
                                     (es_19_1MyTrue_2,Go)] */
  logic [1:0] es_19_1MyTrue_emitted;
  logic [1:0] es_19_1MyTrue_done;
  assign es_19_1MyTrue_1_d = (es_19_1MyTrue_d[0] && (! es_19_1MyTrue_emitted[0]));
  assign es_19_1MyTrue_2_d = (es_19_1MyTrue_d[0] && (! es_19_1MyTrue_emitted[1]));
  assign es_19_1MyTrue_done = (es_19_1MyTrue_emitted | ({es_19_1MyTrue_2_d[0],
                                                         es_19_1MyTrue_1_d[0]} & {es_19_1MyTrue_2_r,
                                                                                  es_19_1MyTrue_1_r}));
  assign es_19_1MyTrue_r = (& es_19_1MyTrue_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_19_1MyTrue_emitted <= 2'd0;
    else
      es_19_1MyTrue_emitted <= (es_19_1MyTrue_r ? 2'd0 :
                                es_19_1MyTrue_done);
  
  /* dcon (Ty QTree_Int,
      Dcon QNone_Int) : [(es_19_1MyTrue_1,Go)] > (es_19_1MyTrue_1QNone_Int,QTree_Int) */
  assign es_19_1MyTrue_1QNone_Int_d = QNone_Int_dc((& {es_19_1MyTrue_1_d[0]}), es_19_1MyTrue_1_d);
  assign {es_19_1MyTrue_1_r} = {1 {(es_19_1MyTrue_1QNone_Int_r && es_19_1MyTrue_1QNone_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (es_19_1MyTrue_1QNone_Int,QTree_Int) > (lizzieLet23_2_1_argbuf,QTree_Int) */
  QTree_Int_t es_19_1MyTrue_1QNone_Int_bufchan_d;
  logic es_19_1MyTrue_1QNone_Int_bufchan_r;
  assign es_19_1MyTrue_1QNone_Int_r = ((! es_19_1MyTrue_1QNone_Int_bufchan_d[0]) || es_19_1MyTrue_1QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_19_1MyTrue_1QNone_Int_bufchan_d <= {66'd0, 1'd0};
    else
      if (es_19_1MyTrue_1QNone_Int_r)
        es_19_1MyTrue_1QNone_Int_bufchan_d <= es_19_1MyTrue_1QNone_Int_d;
  QTree_Int_t es_19_1MyTrue_1QNone_Int_bufchan_buf;
  assign es_19_1MyTrue_1QNone_Int_bufchan_r = (! es_19_1MyTrue_1QNone_Int_bufchan_buf[0]);
  assign lizzieLet23_2_1_argbuf_d = (es_19_1MyTrue_1QNone_Int_bufchan_buf[0] ? es_19_1MyTrue_1QNone_Int_bufchan_buf :
                                     es_19_1MyTrue_1QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_19_1MyTrue_1QNone_Int_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((lizzieLet23_2_1_argbuf_r && es_19_1MyTrue_1QNone_Int_bufchan_buf[0]))
        es_19_1MyTrue_1QNone_Int_bufchan_buf <= {66'd0, 1'd0};
      else if (((! lizzieLet23_2_1_argbuf_r) && (! es_19_1MyTrue_1QNone_Int_bufchan_buf[0])))
        es_19_1MyTrue_1QNone_Int_bufchan_buf <= es_19_1MyTrue_1QNone_Int_bufchan_d;
  
  /* buf (Ty Go) : (es_19_1MyTrue_2,Go) > (es_19_1MyTrue_2_argbuf,Go) */
  Go_t es_19_1MyTrue_2_bufchan_d;
  logic es_19_1MyTrue_2_bufchan_r;
  assign es_19_1MyTrue_2_r = ((! es_19_1MyTrue_2_bufchan_d[0]) || es_19_1MyTrue_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_19_1MyTrue_2_bufchan_d <= 1'd0;
    else
      if (es_19_1MyTrue_2_r)
        es_19_1MyTrue_2_bufchan_d <= es_19_1MyTrue_2_d;
  Go_t es_19_1MyTrue_2_bufchan_buf;
  assign es_19_1MyTrue_2_bufchan_r = (! es_19_1MyTrue_2_bufchan_buf[0]);
  assign es_19_1MyTrue_2_argbuf_d = (es_19_1MyTrue_2_bufchan_buf[0] ? es_19_1MyTrue_2_bufchan_buf :
                                     es_19_1MyTrue_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_19_1MyTrue_2_bufchan_buf <= 1'd0;
    else
      if ((es_19_1MyTrue_2_argbuf_r && es_19_1MyTrue_2_bufchan_buf[0]))
        es_19_1MyTrue_2_bufchan_buf <= 1'd0;
      else if (((! es_19_1MyTrue_2_argbuf_r) && (! es_19_1MyTrue_2_bufchan_buf[0])))
        es_19_1MyTrue_2_bufchan_buf <= es_19_1MyTrue_2_bufchan_d;
  
  /* demux (Ty MyBool,
       Ty MyDTInt_Int_Int) : (es_19_2,MyBool) (es_14_3MyFalse_2,MyDTInt_Int_Int) > [(es_19_2MyFalse,MyDTInt_Int_Int),
                                                                                    (_73,MyDTInt_Int_Int)] */
  logic [1:0] es_14_3MyFalse_2_onehotd;
  always_comb
    if ((es_19_2_d[0] && es_14_3MyFalse_2_d[0]))
      unique case (es_19_2_d[1:1])
        1'd0: es_14_3MyFalse_2_onehotd = 2'd1;
        1'd1: es_14_3MyFalse_2_onehotd = 2'd2;
        default: es_14_3MyFalse_2_onehotd = 2'd0;
      endcase
    else es_14_3MyFalse_2_onehotd = 2'd0;
  assign es_19_2MyFalse_d = es_14_3MyFalse_2_onehotd[0];
  assign _73_d = es_14_3MyFalse_2_onehotd[1];
  assign es_14_3MyFalse_2_r = (| (es_14_3MyFalse_2_onehotd & {_73_r,
                                                              es_19_2MyFalse_r}));
  assign es_19_2_r = es_14_3MyFalse_2_r;
  
  /* buf (Ty MyDTInt_Int_Int) : (es_19_2MyFalse,MyDTInt_Int_Int) > (es_19_2MyFalse_1_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t es_19_2MyFalse_bufchan_d;
  logic es_19_2MyFalse_bufchan_r;
  assign es_19_2MyFalse_r = ((! es_19_2MyFalse_bufchan_d[0]) || es_19_2MyFalse_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_19_2MyFalse_bufchan_d <= 1'd0;
    else
      if (es_19_2MyFalse_r) es_19_2MyFalse_bufchan_d <= es_19_2MyFalse_d;
  MyDTInt_Int_Int_t es_19_2MyFalse_bufchan_buf;
  assign es_19_2MyFalse_bufchan_r = (! es_19_2MyFalse_bufchan_buf[0]);
  assign es_19_2MyFalse_1_argbuf_d = (es_19_2MyFalse_bufchan_buf[0] ? es_19_2MyFalse_bufchan_buf :
                                      es_19_2MyFalse_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_19_2MyFalse_bufchan_buf <= 1'd0;
    else
      if ((es_19_2MyFalse_1_argbuf_r && es_19_2MyFalse_bufchan_buf[0]))
        es_19_2MyFalse_bufchan_buf <= 1'd0;
      else if (((! es_19_2MyFalse_1_argbuf_r) && (! es_19_2MyFalse_bufchan_buf[0])))
        es_19_2MyFalse_bufchan_buf <= es_19_2MyFalse_bufchan_d;
  
  /* dcon (Ty TupMyDTInt_Int_Int___Int___Int,
      Dcon TupMyDTInt_Int_Int___Int___Int) : [(es_19_2MyFalse_1_argbuf,MyDTInt_Int_Int),
                                              (es_19_5MyFalse_1_argbuf,Int),
                                              (es_19_6MyFalse_1_argbuf,Int)] > (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int3,TupMyDTInt_Int_Int___Int___Int) */
  assign applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int3_d = TupMyDTInt_Int_Int___Int___Int_dc((& {es_19_2MyFalse_1_argbuf_d[0],
                                                                                                       es_19_5MyFalse_1_argbuf_d[0],
                                                                                                       es_19_6MyFalse_1_argbuf_d[0]}), es_19_2MyFalse_1_argbuf_d, es_19_5MyFalse_1_argbuf_d, es_19_6MyFalse_1_argbuf_d);
  assign {es_19_2MyFalse_1_argbuf_r,
          es_19_5MyFalse_1_argbuf_r,
          es_19_6MyFalse_1_argbuf_r} = {3 {(applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int3_r && applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int3_d[0])}};
  
  /* demux (Ty MyBool,
       Ty MyDTInt_Int) : (es_19_3,MyBool) (es_14_4MyFalse_2,MyDTInt_Int) > [(es_19_3MyFalse,MyDTInt_Int),
                                                                            (_72,MyDTInt_Int)] */
  logic [1:0] es_14_4MyFalse_2_onehotd;
  always_comb
    if ((es_19_3_d[0] && es_14_4MyFalse_2_d[0]))
      unique case (es_19_3_d[1:1])
        1'd0: es_14_4MyFalse_2_onehotd = 2'd1;
        1'd1: es_14_4MyFalse_2_onehotd = 2'd2;
        default: es_14_4MyFalse_2_onehotd = 2'd0;
      endcase
    else es_14_4MyFalse_2_onehotd = 2'd0;
  assign es_19_3MyFalse_d = es_14_4MyFalse_2_onehotd[0];
  assign _72_d = es_14_4MyFalse_2_onehotd[1];
  assign es_14_4MyFalse_2_r = (| (es_14_4MyFalse_2_onehotd & {_72_r,
                                                              es_19_3MyFalse_r}));
  assign es_19_3_r = es_14_4MyFalse_2_r;
  
  /* buf (Ty MyDTInt_Int) : (es_19_3MyFalse,MyDTInt_Int) > (es_19_3MyFalse_1_argbuf,MyDTInt_Int) */
  MyDTInt_Int_t es_19_3MyFalse_bufchan_d;
  logic es_19_3MyFalse_bufchan_r;
  assign es_19_3MyFalse_r = ((! es_19_3MyFalse_bufchan_d[0]) || es_19_3MyFalse_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_19_3MyFalse_bufchan_d <= 1'd0;
    else
      if (es_19_3MyFalse_r) es_19_3MyFalse_bufchan_d <= es_19_3MyFalse_d;
  MyDTInt_Int_t es_19_3MyFalse_bufchan_buf;
  assign es_19_3MyFalse_bufchan_r = (! es_19_3MyFalse_bufchan_buf[0]);
  assign es_19_3MyFalse_1_argbuf_d = (es_19_3MyFalse_bufchan_buf[0] ? es_19_3MyFalse_bufchan_buf :
                                      es_19_3MyFalse_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_19_3MyFalse_bufchan_buf <= 1'd0;
    else
      if ((es_19_3MyFalse_1_argbuf_r && es_19_3MyFalse_bufchan_buf[0]))
        es_19_3MyFalse_bufchan_buf <= 1'd0;
      else if (((! es_19_3MyFalse_1_argbuf_r) && (! es_19_3MyFalse_bufchan_buf[0])))
        es_19_3MyFalse_bufchan_buf <= es_19_3MyFalse_bufchan_d;
  
  /* demux (Ty MyBool,
       Ty Pointer_CTf_f_Int_Int) : (es_19_4,MyBool) (es_14_5MyFalse,Pointer_CTf_f_Int_Int) > [(es_19_4MyFalse,Pointer_CTf_f_Int_Int),
                                                                                              (es_19_4MyTrue,Pointer_CTf_f_Int_Int)] */
  logic [1:0] es_14_5MyFalse_onehotd;
  always_comb
    if ((es_19_4_d[0] && es_14_5MyFalse_d[0]))
      unique case (es_19_4_d[1:1])
        1'd0: es_14_5MyFalse_onehotd = 2'd1;
        1'd1: es_14_5MyFalse_onehotd = 2'd2;
        default: es_14_5MyFalse_onehotd = 2'd0;
      endcase
    else es_14_5MyFalse_onehotd = 2'd0;
  assign es_19_4MyFalse_d = {es_14_5MyFalse_d[16:1],
                             es_14_5MyFalse_onehotd[0]};
  assign es_19_4MyTrue_d = {es_14_5MyFalse_d[16:1],
                            es_14_5MyFalse_onehotd[1]};
  assign es_14_5MyFalse_r = (| (es_14_5MyFalse_onehotd & {es_19_4MyTrue_r,
                                                          es_19_4MyFalse_r}));
  assign es_19_4_r = es_14_5MyFalse_r;
  
  /* buf (Ty Pointer_CTf_f_Int_Int) : (es_19_4MyFalse,Pointer_CTf_f_Int_Int) > (es_19_4MyFalse_1_argbuf,Pointer_CTf_f_Int_Int) */
  Pointer_CTf_f_Int_Int_t es_19_4MyFalse_bufchan_d;
  logic es_19_4MyFalse_bufchan_r;
  assign es_19_4MyFalse_r = ((! es_19_4MyFalse_bufchan_d[0]) || es_19_4MyFalse_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_19_4MyFalse_bufchan_d <= {16'd0, 1'd0};
    else
      if (es_19_4MyFalse_r) es_19_4MyFalse_bufchan_d <= es_19_4MyFalse_d;
  Pointer_CTf_f_Int_Int_t es_19_4MyFalse_bufchan_buf;
  assign es_19_4MyFalse_bufchan_r = (! es_19_4MyFalse_bufchan_buf[0]);
  assign es_19_4MyFalse_1_argbuf_d = (es_19_4MyFalse_bufchan_buf[0] ? es_19_4MyFalse_bufchan_buf :
                                      es_19_4MyFalse_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_19_4MyFalse_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((es_19_4MyFalse_1_argbuf_r && es_19_4MyFalse_bufchan_buf[0]))
        es_19_4MyFalse_bufchan_buf <= {16'd0, 1'd0};
      else if (((! es_19_4MyFalse_1_argbuf_r) && (! es_19_4MyFalse_bufchan_buf[0])))
        es_19_4MyFalse_bufchan_buf <= es_19_4MyFalse_bufchan_d;
  
  /* buf (Ty Pointer_CTf_f_Int_Int) : (es_19_4MyTrue,Pointer_CTf_f_Int_Int) > (es_19_4MyTrue_1_argbuf,Pointer_CTf_f_Int_Int) */
  Pointer_CTf_f_Int_Int_t es_19_4MyTrue_bufchan_d;
  logic es_19_4MyTrue_bufchan_r;
  assign es_19_4MyTrue_r = ((! es_19_4MyTrue_bufchan_d[0]) || es_19_4MyTrue_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_19_4MyTrue_bufchan_d <= {16'd0, 1'd0};
    else
      if (es_19_4MyTrue_r) es_19_4MyTrue_bufchan_d <= es_19_4MyTrue_d;
  Pointer_CTf_f_Int_Int_t es_19_4MyTrue_bufchan_buf;
  assign es_19_4MyTrue_bufchan_r = (! es_19_4MyTrue_bufchan_buf[0]);
  assign es_19_4MyTrue_1_argbuf_d = (es_19_4MyTrue_bufchan_buf[0] ? es_19_4MyTrue_bufchan_buf :
                                     es_19_4MyTrue_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_19_4MyTrue_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((es_19_4MyTrue_1_argbuf_r && es_19_4MyTrue_bufchan_buf[0]))
        es_19_4MyTrue_bufchan_buf <= {16'd0, 1'd0};
      else if (((! es_19_4MyTrue_1_argbuf_r) && (! es_19_4MyTrue_bufchan_buf[0])))
        es_19_4MyTrue_bufchan_buf <= es_19_4MyTrue_bufchan_d;
  
  /* demux (Ty MyBool,
       Ty Int) : (es_19_5,MyBool) (es_14_6MyFalse_2,Int) > [(es_19_5MyFalse,Int),
                                                            (_71,Int)] */
  logic [1:0] es_14_6MyFalse_2_onehotd;
  always_comb
    if ((es_19_5_d[0] && es_14_6MyFalse_2_d[0]))
      unique case (es_19_5_d[1:1])
        1'd0: es_14_6MyFalse_2_onehotd = 2'd1;
        1'd1: es_14_6MyFalse_2_onehotd = 2'd2;
        default: es_14_6MyFalse_2_onehotd = 2'd0;
      endcase
    else es_14_6MyFalse_2_onehotd = 2'd0;
  assign es_19_5MyFalse_d = {es_14_6MyFalse_2_d[32:1],
                             es_14_6MyFalse_2_onehotd[0]};
  assign _71_d = {es_14_6MyFalse_2_d[32:1],
                  es_14_6MyFalse_2_onehotd[1]};
  assign es_14_6MyFalse_2_r = (| (es_14_6MyFalse_2_onehotd & {_71_r,
                                                              es_19_5MyFalse_r}));
  assign es_19_5_r = es_14_6MyFalse_2_r;
  
  /* buf (Ty Int) : (es_19_5MyFalse,Int) > (es_19_5MyFalse_1_argbuf,Int) */
  Int_t es_19_5MyFalse_bufchan_d;
  logic es_19_5MyFalse_bufchan_r;
  assign es_19_5MyFalse_r = ((! es_19_5MyFalse_bufchan_d[0]) || es_19_5MyFalse_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_19_5MyFalse_bufchan_d <= {32'd0, 1'd0};
    else
      if (es_19_5MyFalse_r) es_19_5MyFalse_bufchan_d <= es_19_5MyFalse_d;
  Int_t es_19_5MyFalse_bufchan_buf;
  assign es_19_5MyFalse_bufchan_r = (! es_19_5MyFalse_bufchan_buf[0]);
  assign es_19_5MyFalse_1_argbuf_d = (es_19_5MyFalse_bufchan_buf[0] ? es_19_5MyFalse_bufchan_buf :
                                      es_19_5MyFalse_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_19_5MyFalse_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((es_19_5MyFalse_1_argbuf_r && es_19_5MyFalse_bufchan_buf[0]))
        es_19_5MyFalse_bufchan_buf <= {32'd0, 1'd0};
      else if (((! es_19_5MyFalse_1_argbuf_r) && (! es_19_5MyFalse_bufchan_buf[0])))
        es_19_5MyFalse_bufchan_buf <= es_19_5MyFalse_bufchan_d;
  
  /* demux (Ty MyBool,
       Ty Int) : (es_19_6,MyBool) (es_14_7MyFalse_2,Int) > [(es_19_6MyFalse,Int),
                                                            (_70,Int)] */
  logic [1:0] es_14_7MyFalse_2_onehotd;
  always_comb
    if ((es_19_6_d[0] && es_14_7MyFalse_2_d[0]))
      unique case (es_19_6_d[1:1])
        1'd0: es_14_7MyFalse_2_onehotd = 2'd1;
        1'd1: es_14_7MyFalse_2_onehotd = 2'd2;
        default: es_14_7MyFalse_2_onehotd = 2'd0;
      endcase
    else es_14_7MyFalse_2_onehotd = 2'd0;
  assign es_19_6MyFalse_d = {es_14_7MyFalse_2_d[32:1],
                             es_14_7MyFalse_2_onehotd[0]};
  assign _70_d = {es_14_7MyFalse_2_d[32:1],
                  es_14_7MyFalse_2_onehotd[1]};
  assign es_14_7MyFalse_2_r = (| (es_14_7MyFalse_2_onehotd & {_70_r,
                                                              es_19_6MyFalse_r}));
  assign es_19_6_r = es_14_7MyFalse_2_r;
  
  /* buf (Ty Int) : (es_19_6MyFalse,Int) > (es_19_6MyFalse_1_argbuf,Int) */
  Int_t es_19_6MyFalse_bufchan_d;
  logic es_19_6MyFalse_bufchan_r;
  assign es_19_6MyFalse_r = ((! es_19_6MyFalse_bufchan_d[0]) || es_19_6MyFalse_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_19_6MyFalse_bufchan_d <= {32'd0, 1'd0};
    else
      if (es_19_6MyFalse_r) es_19_6MyFalse_bufchan_d <= es_19_6MyFalse_d;
  Int_t es_19_6MyFalse_bufchan_buf;
  assign es_19_6MyFalse_bufchan_r = (! es_19_6MyFalse_bufchan_buf[0]);
  assign es_19_6MyFalse_1_argbuf_d = (es_19_6MyFalse_bufchan_buf[0] ? es_19_6MyFalse_bufchan_buf :
                                      es_19_6MyFalse_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_19_6MyFalse_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((es_19_6MyFalse_1_argbuf_r && es_19_6MyFalse_bufchan_buf[0]))
        es_19_6MyFalse_bufchan_buf <= {32'd0, 1'd0};
      else if (((! es_19_6MyFalse_1_argbuf_r) && (! es_19_6MyFalse_bufchan_buf[0])))
        es_19_6MyFalse_bufchan_buf <= es_19_6MyFalse_bufchan_d;
  
  /* buf (Ty QTree_Int) : (es_20_1QVal_Int,QTree_Int) > (lizzieLet22_1_argbuf,QTree_Int) */
  QTree_Int_t es_20_1QVal_Int_bufchan_d;
  logic es_20_1QVal_Int_bufchan_r;
  assign es_20_1QVal_Int_r = ((! es_20_1QVal_Int_bufchan_d[0]) || es_20_1QVal_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_20_1QVal_Int_bufchan_d <= {66'd0, 1'd0};
    else
      if (es_20_1QVal_Int_r)
        es_20_1QVal_Int_bufchan_d <= es_20_1QVal_Int_d;
  QTree_Int_t es_20_1QVal_Int_bufchan_buf;
  assign es_20_1QVal_Int_bufchan_r = (! es_20_1QVal_Int_bufchan_buf[0]);
  assign lizzieLet22_1_argbuf_d = (es_20_1QVal_Int_bufchan_buf[0] ? es_20_1QVal_Int_bufchan_buf :
                                   es_20_1QVal_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_20_1QVal_Int_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((lizzieLet22_1_argbuf_r && es_20_1QVal_Int_bufchan_buf[0]))
        es_20_1QVal_Int_bufchan_buf <= {66'd0, 1'd0};
      else if (((! lizzieLet22_1_argbuf_r) && (! es_20_1QVal_Int_bufchan_buf[0])))
        es_20_1QVal_Int_bufchan_buf <= es_20_1QVal_Int_bufchan_d;
  
  /* buf (Ty QTree_Int) : (es_23_1es_24_1es_25_1es_26_1QNode_Int,QTree_Int) > (lizzieLet28_1_argbuf,QTree_Int) */
  QTree_Int_t es_23_1es_24_1es_25_1es_26_1QNode_Int_bufchan_d;
  logic es_23_1es_24_1es_25_1es_26_1QNode_Int_bufchan_r;
  assign es_23_1es_24_1es_25_1es_26_1QNode_Int_r = ((! es_23_1es_24_1es_25_1es_26_1QNode_Int_bufchan_d[0]) || es_23_1es_24_1es_25_1es_26_1QNode_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_23_1es_24_1es_25_1es_26_1QNode_Int_bufchan_d <= {66'd0, 1'd0};
    else
      if (es_23_1es_24_1es_25_1es_26_1QNode_Int_r)
        es_23_1es_24_1es_25_1es_26_1QNode_Int_bufchan_d <= es_23_1es_24_1es_25_1es_26_1QNode_Int_d;
  QTree_Int_t es_23_1es_24_1es_25_1es_26_1QNode_Int_bufchan_buf;
  assign es_23_1es_24_1es_25_1es_26_1QNode_Int_bufchan_r = (! es_23_1es_24_1es_25_1es_26_1QNode_Int_bufchan_buf[0]);
  assign lizzieLet28_1_argbuf_d = (es_23_1es_24_1es_25_1es_26_1QNode_Int_bufchan_buf[0] ? es_23_1es_24_1es_25_1es_26_1QNode_Int_bufchan_buf :
                                   es_23_1es_24_1es_25_1es_26_1QNode_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_23_1es_24_1es_25_1es_26_1QNode_Int_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((lizzieLet28_1_argbuf_r && es_23_1es_24_1es_25_1es_26_1QNode_Int_bufchan_buf[0]))
        es_23_1es_24_1es_25_1es_26_1QNode_Int_bufchan_buf <= {66'd0, 1'd0};
      else if (((! lizzieLet28_1_argbuf_r) && (! es_23_1es_24_1es_25_1es_26_1QNode_Int_bufchan_buf[0])))
        es_23_1es_24_1es_25_1es_26_1QNode_Int_bufchan_buf <= es_23_1es_24_1es_25_1es_26_1QNode_Int_bufchan_d;
  
  /* demux (Ty MyBool,
       Ty Go) : (es_2_1,MyBool) (lizzieLet6_3QVal_Int_3,Go) > [(es_2_1MyFalse,Go),
                                                               (es_2_1MyTrue,Go)] */
  logic [1:0] lizzieLet6_3QVal_Int_3_onehotd;
  always_comb
    if ((es_2_1_d[0] && lizzieLet6_3QVal_Int_3_d[0]))
      unique case (es_2_1_d[1:1])
        1'd0: lizzieLet6_3QVal_Int_3_onehotd = 2'd1;
        1'd1: lizzieLet6_3QVal_Int_3_onehotd = 2'd2;
        default: lizzieLet6_3QVal_Int_3_onehotd = 2'd0;
      endcase
    else lizzieLet6_3QVal_Int_3_onehotd = 2'd0;
  assign es_2_1MyFalse_d = lizzieLet6_3QVal_Int_3_onehotd[0];
  assign es_2_1MyTrue_d = lizzieLet6_3QVal_Int_3_onehotd[1];
  assign lizzieLet6_3QVal_Int_3_r = (| (lizzieLet6_3QVal_Int_3_onehotd & {es_2_1MyTrue_r,
                                                                          es_2_1MyFalse_r}));
  assign es_2_1_r = lizzieLet6_3QVal_Int_3_r;
  
  /* fork (Ty Go) : (es_2_1MyFalse,Go) > [(es_2_1MyFalse_1,Go),
                                     (es_2_1MyFalse_2,Go)] */
  logic [1:0] es_2_1MyFalse_emitted;
  logic [1:0] es_2_1MyFalse_done;
  assign es_2_1MyFalse_1_d = (es_2_1MyFalse_d[0] && (! es_2_1MyFalse_emitted[0]));
  assign es_2_1MyFalse_2_d = (es_2_1MyFalse_d[0] && (! es_2_1MyFalse_emitted[1]));
  assign es_2_1MyFalse_done = (es_2_1MyFalse_emitted | ({es_2_1MyFalse_2_d[0],
                                                         es_2_1MyFalse_1_d[0]} & {es_2_1MyFalse_2_r,
                                                                                  es_2_1MyFalse_1_r}));
  assign es_2_1MyFalse_r = (& es_2_1MyFalse_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_2_1MyFalse_emitted <= 2'd0;
    else
      es_2_1MyFalse_emitted <= (es_2_1MyFalse_r ? 2'd0 :
                                es_2_1MyFalse_done);
  
  /* buf (Ty Go) : (es_2_1MyFalse_1,Go) > (es_2_1MyFalse_1_argbuf,Go) */
  Go_t es_2_1MyFalse_1_bufchan_d;
  logic es_2_1MyFalse_1_bufchan_r;
  assign es_2_1MyFalse_1_r = ((! es_2_1MyFalse_1_bufchan_d[0]) || es_2_1MyFalse_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_2_1MyFalse_1_bufchan_d <= 1'd0;
    else
      if (es_2_1MyFalse_1_r)
        es_2_1MyFalse_1_bufchan_d <= es_2_1MyFalse_1_d;
  Go_t es_2_1MyFalse_1_bufchan_buf;
  assign es_2_1MyFalse_1_bufchan_r = (! es_2_1MyFalse_1_bufchan_buf[0]);
  assign es_2_1MyFalse_1_argbuf_d = (es_2_1MyFalse_1_bufchan_buf[0] ? es_2_1MyFalse_1_bufchan_buf :
                                     es_2_1MyFalse_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_2_1MyFalse_1_bufchan_buf <= 1'd0;
    else
      if ((es_2_1MyFalse_1_argbuf_r && es_2_1MyFalse_1_bufchan_buf[0]))
        es_2_1MyFalse_1_bufchan_buf <= 1'd0;
      else if (((! es_2_1MyFalse_1_argbuf_r) && (! es_2_1MyFalse_1_bufchan_buf[0])))
        es_2_1MyFalse_1_bufchan_buf <= es_2_1MyFalse_1_bufchan_d;
  
  /* dcon (Ty TupGo___MyDTInt_Int___Int,
      Dcon TupGo___MyDTInt_Int___Int) : [(es_2_1MyFalse_1_argbuf,Go),
                                         (es_2_2MyFalse_1_argbuf,MyDTInt_Int),
                                         (es_2_4MyFalse_1_argbuf,Int)] > (applyfnInt_Int_5TupGo___MyDTInt_Int___Int4,TupGo___MyDTInt_Int___Int) */
  assign applyfnInt_Int_5TupGo___MyDTInt_Int___Int4_d = TupGo___MyDTInt_Int___Int_dc((& {es_2_1MyFalse_1_argbuf_d[0],
                                                                                         es_2_2MyFalse_1_argbuf_d[0],
                                                                                         es_2_4MyFalse_1_argbuf_d[0]}), es_2_1MyFalse_1_argbuf_d, es_2_2MyFalse_1_argbuf_d, es_2_4MyFalse_1_argbuf_d);
  assign {es_2_1MyFalse_1_argbuf_r,
          es_2_2MyFalse_1_argbuf_r,
          es_2_4MyFalse_1_argbuf_r} = {3 {(applyfnInt_Int_5TupGo___MyDTInt_Int___Int4_r && applyfnInt_Int_5TupGo___MyDTInt_Int___Int4_d[0])}};
  
  /* buf (Ty Go) : (es_2_1MyFalse_2,Go) > (es_2_1MyFalse_2_argbuf,Go) */
  Go_t es_2_1MyFalse_2_bufchan_d;
  logic es_2_1MyFalse_2_bufchan_r;
  assign es_2_1MyFalse_2_r = ((! es_2_1MyFalse_2_bufchan_d[0]) || es_2_1MyFalse_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_2_1MyFalse_2_bufchan_d <= 1'd0;
    else
      if (es_2_1MyFalse_2_r)
        es_2_1MyFalse_2_bufchan_d <= es_2_1MyFalse_2_d;
  Go_t es_2_1MyFalse_2_bufchan_buf;
  assign es_2_1MyFalse_2_bufchan_r = (! es_2_1MyFalse_2_bufchan_buf[0]);
  assign es_2_1MyFalse_2_argbuf_d = (es_2_1MyFalse_2_bufchan_buf[0] ? es_2_1MyFalse_2_bufchan_buf :
                                     es_2_1MyFalse_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_2_1MyFalse_2_bufchan_buf <= 1'd0;
    else
      if ((es_2_1MyFalse_2_argbuf_r && es_2_1MyFalse_2_bufchan_buf[0]))
        es_2_1MyFalse_2_bufchan_buf <= 1'd0;
      else if (((! es_2_1MyFalse_2_argbuf_r) && (! es_2_1MyFalse_2_bufchan_buf[0])))
        es_2_1MyFalse_2_bufchan_buf <= es_2_1MyFalse_2_bufchan_d;
  
  /* fork (Ty Go) : (es_2_1MyTrue,Go) > [(es_2_1MyTrue_1,Go),
                                    (es_2_1MyTrue_2,Go)] */
  logic [1:0] es_2_1MyTrue_emitted;
  logic [1:0] es_2_1MyTrue_done;
  assign es_2_1MyTrue_1_d = (es_2_1MyTrue_d[0] && (! es_2_1MyTrue_emitted[0]));
  assign es_2_1MyTrue_2_d = (es_2_1MyTrue_d[0] && (! es_2_1MyTrue_emitted[1]));
  assign es_2_1MyTrue_done = (es_2_1MyTrue_emitted | ({es_2_1MyTrue_2_d[0],
                                                       es_2_1MyTrue_1_d[0]} & {es_2_1MyTrue_2_r,
                                                                               es_2_1MyTrue_1_r}));
  assign es_2_1MyTrue_r = (& es_2_1MyTrue_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_2_1MyTrue_emitted <= 2'd0;
    else
      es_2_1MyTrue_emitted <= (es_2_1MyTrue_r ? 2'd0 :
                               es_2_1MyTrue_done);
  
  /* dcon (Ty QTree_Int,
      Dcon QNone_Int) : [(es_2_1MyTrue_1,Go)] > (es_2_1MyTrue_1QNone_Int,QTree_Int) */
  assign es_2_1MyTrue_1QNone_Int_d = QNone_Int_dc((& {es_2_1MyTrue_1_d[0]}), es_2_1MyTrue_1_d);
  assign {es_2_1MyTrue_1_r} = {1 {(es_2_1MyTrue_1QNone_Int_r && es_2_1MyTrue_1QNone_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (es_2_1MyTrue_1QNone_Int,QTree_Int) > (lizzieLet9_1_argbuf,QTree_Int) */
  QTree_Int_t es_2_1MyTrue_1QNone_Int_bufchan_d;
  logic es_2_1MyTrue_1QNone_Int_bufchan_r;
  assign es_2_1MyTrue_1QNone_Int_r = ((! es_2_1MyTrue_1QNone_Int_bufchan_d[0]) || es_2_1MyTrue_1QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_2_1MyTrue_1QNone_Int_bufchan_d <= {66'd0, 1'd0};
    else
      if (es_2_1MyTrue_1QNone_Int_r)
        es_2_1MyTrue_1QNone_Int_bufchan_d <= es_2_1MyTrue_1QNone_Int_d;
  QTree_Int_t es_2_1MyTrue_1QNone_Int_bufchan_buf;
  assign es_2_1MyTrue_1QNone_Int_bufchan_r = (! es_2_1MyTrue_1QNone_Int_bufchan_buf[0]);
  assign lizzieLet9_1_argbuf_d = (es_2_1MyTrue_1QNone_Int_bufchan_buf[0] ? es_2_1MyTrue_1QNone_Int_bufchan_buf :
                                  es_2_1MyTrue_1QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_2_1MyTrue_1QNone_Int_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((lizzieLet9_1_argbuf_r && es_2_1MyTrue_1QNone_Int_bufchan_buf[0]))
        es_2_1MyTrue_1QNone_Int_bufchan_buf <= {66'd0, 1'd0};
      else if (((! lizzieLet9_1_argbuf_r) && (! es_2_1MyTrue_1QNone_Int_bufchan_buf[0])))
        es_2_1MyTrue_1QNone_Int_bufchan_buf <= es_2_1MyTrue_1QNone_Int_bufchan_d;
  
  /* buf (Ty Go) : (es_2_1MyTrue_2,Go) > (es_2_1MyTrue_2_argbuf,Go) */
  Go_t es_2_1MyTrue_2_bufchan_d;
  logic es_2_1MyTrue_2_bufchan_r;
  assign es_2_1MyTrue_2_r = ((! es_2_1MyTrue_2_bufchan_d[0]) || es_2_1MyTrue_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_2_1MyTrue_2_bufchan_d <= 1'd0;
    else
      if (es_2_1MyTrue_2_r) es_2_1MyTrue_2_bufchan_d <= es_2_1MyTrue_2_d;
  Go_t es_2_1MyTrue_2_bufchan_buf;
  assign es_2_1MyTrue_2_bufchan_r = (! es_2_1MyTrue_2_bufchan_buf[0]);
  assign es_2_1MyTrue_2_argbuf_d = (es_2_1MyTrue_2_bufchan_buf[0] ? es_2_1MyTrue_2_bufchan_buf :
                                    es_2_1MyTrue_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_2_1MyTrue_2_bufchan_buf <= 1'd0;
    else
      if ((es_2_1MyTrue_2_argbuf_r && es_2_1MyTrue_2_bufchan_buf[0]))
        es_2_1MyTrue_2_bufchan_buf <= 1'd0;
      else if (((! es_2_1MyTrue_2_argbuf_r) && (! es_2_1MyTrue_2_bufchan_buf[0])))
        es_2_1MyTrue_2_bufchan_buf <= es_2_1MyTrue_2_bufchan_d;
  
  /* demux (Ty MyBool,
       Ty Go) : (es_2_1_1,MyBool) (lizzieLet12_6QNone_Int_3QVal_Int_3,Go) > [(es_2_1_1MyFalse,Go),
                                                                             (es_2_1_1MyTrue,Go)] */
  logic [1:0] lizzieLet12_6QNone_Int_3QVal_Int_3_onehotd;
  always_comb
    if ((es_2_1_1_d[0] && lizzieLet12_6QNone_Int_3QVal_Int_3_d[0]))
      unique case (es_2_1_1_d[1:1])
        1'd0: lizzieLet12_6QNone_Int_3QVal_Int_3_onehotd = 2'd1;
        1'd1: lizzieLet12_6QNone_Int_3QVal_Int_3_onehotd = 2'd2;
        default: lizzieLet12_6QNone_Int_3QVal_Int_3_onehotd = 2'd0;
      endcase
    else lizzieLet12_6QNone_Int_3QVal_Int_3_onehotd = 2'd0;
  assign es_2_1_1MyFalse_d = lizzieLet12_6QNone_Int_3QVal_Int_3_onehotd[0];
  assign es_2_1_1MyTrue_d = lizzieLet12_6QNone_Int_3QVal_Int_3_onehotd[1];
  assign lizzieLet12_6QNone_Int_3QVal_Int_3_r = (| (lizzieLet12_6QNone_Int_3QVal_Int_3_onehotd & {es_2_1_1MyTrue_r,
                                                                                                  es_2_1_1MyFalse_r}));
  assign es_2_1_1_r = lizzieLet12_6QNone_Int_3QVal_Int_3_r;
  
  /* fork (Ty Go) : (es_2_1_1MyFalse,Go) > [(es_2_1_1MyFalse_1,Go),
                                       (es_2_1_1MyFalse_2,Go)] */
  logic [1:0] es_2_1_1MyFalse_emitted;
  logic [1:0] es_2_1_1MyFalse_done;
  assign es_2_1_1MyFalse_1_d = (es_2_1_1MyFalse_d[0] && (! es_2_1_1MyFalse_emitted[0]));
  assign es_2_1_1MyFalse_2_d = (es_2_1_1MyFalse_d[0] && (! es_2_1_1MyFalse_emitted[1]));
  assign es_2_1_1MyFalse_done = (es_2_1_1MyFalse_emitted | ({es_2_1_1MyFalse_2_d[0],
                                                             es_2_1_1MyFalse_1_d[0]} & {es_2_1_1MyFalse_2_r,
                                                                                        es_2_1_1MyFalse_1_r}));
  assign es_2_1_1MyFalse_r = (& es_2_1_1MyFalse_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_2_1_1MyFalse_emitted <= 2'd0;
    else
      es_2_1_1MyFalse_emitted <= (es_2_1_1MyFalse_r ? 2'd0 :
                                  es_2_1_1MyFalse_done);
  
  /* buf (Ty Go) : (es_2_1_1MyFalse_1,Go) > (es_2_1_1MyFalse_1_argbuf,Go) */
  Go_t es_2_1_1MyFalse_1_bufchan_d;
  logic es_2_1_1MyFalse_1_bufchan_r;
  assign es_2_1_1MyFalse_1_r = ((! es_2_1_1MyFalse_1_bufchan_d[0]) || es_2_1_1MyFalse_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_2_1_1MyFalse_1_bufchan_d <= 1'd0;
    else
      if (es_2_1_1MyFalse_1_r)
        es_2_1_1MyFalse_1_bufchan_d <= es_2_1_1MyFalse_1_d;
  Go_t es_2_1_1MyFalse_1_bufchan_buf;
  assign es_2_1_1MyFalse_1_bufchan_r = (! es_2_1_1MyFalse_1_bufchan_buf[0]);
  assign es_2_1_1MyFalse_1_argbuf_d = (es_2_1_1MyFalse_1_bufchan_buf[0] ? es_2_1_1MyFalse_1_bufchan_buf :
                                       es_2_1_1MyFalse_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_2_1_1MyFalse_1_bufchan_buf <= 1'd0;
    else
      if ((es_2_1_1MyFalse_1_argbuf_r && es_2_1_1MyFalse_1_bufchan_buf[0]))
        es_2_1_1MyFalse_1_bufchan_buf <= 1'd0;
      else if (((! es_2_1_1MyFalse_1_argbuf_r) && (! es_2_1_1MyFalse_1_bufchan_buf[0])))
        es_2_1_1MyFalse_1_bufchan_buf <= es_2_1_1MyFalse_1_bufchan_d;
  
  /* dcon (Ty TupGo___MyDTInt_Int___Int,
      Dcon TupGo___MyDTInt_Int___Int) : [(es_2_1_1MyFalse_1_argbuf,Go),
                                         (es_2_1_2MyFalse_1_argbuf,MyDTInt_Int),
                                         (es_2_1_4MyFalse_1_argbuf,Int)] > (applyfnInt_Int_5TupGo___MyDTInt_Int___Int2,TupGo___MyDTInt_Int___Int) */
  assign applyfnInt_Int_5TupGo___MyDTInt_Int___Int2_d = TupGo___MyDTInt_Int___Int_dc((& {es_2_1_1MyFalse_1_argbuf_d[0],
                                                                                         es_2_1_2MyFalse_1_argbuf_d[0],
                                                                                         es_2_1_4MyFalse_1_argbuf_d[0]}), es_2_1_1MyFalse_1_argbuf_d, es_2_1_2MyFalse_1_argbuf_d, es_2_1_4MyFalse_1_argbuf_d);
  assign {es_2_1_1MyFalse_1_argbuf_r,
          es_2_1_2MyFalse_1_argbuf_r,
          es_2_1_4MyFalse_1_argbuf_r} = {3 {(applyfnInt_Int_5TupGo___MyDTInt_Int___Int2_r && applyfnInt_Int_5TupGo___MyDTInt_Int___Int2_d[0])}};
  
  /* buf (Ty Go) : (es_2_1_1MyFalse_2,Go) > (es_2_1_1MyFalse_2_argbuf,Go) */
  Go_t es_2_1_1MyFalse_2_bufchan_d;
  logic es_2_1_1MyFalse_2_bufchan_r;
  assign es_2_1_1MyFalse_2_r = ((! es_2_1_1MyFalse_2_bufchan_d[0]) || es_2_1_1MyFalse_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_2_1_1MyFalse_2_bufchan_d <= 1'd0;
    else
      if (es_2_1_1MyFalse_2_r)
        es_2_1_1MyFalse_2_bufchan_d <= es_2_1_1MyFalse_2_d;
  Go_t es_2_1_1MyFalse_2_bufchan_buf;
  assign es_2_1_1MyFalse_2_bufchan_r = (! es_2_1_1MyFalse_2_bufchan_buf[0]);
  assign es_2_1_1MyFalse_2_argbuf_d = (es_2_1_1MyFalse_2_bufchan_buf[0] ? es_2_1_1MyFalse_2_bufchan_buf :
                                       es_2_1_1MyFalse_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_2_1_1MyFalse_2_bufchan_buf <= 1'd0;
    else
      if ((es_2_1_1MyFalse_2_argbuf_r && es_2_1_1MyFalse_2_bufchan_buf[0]))
        es_2_1_1MyFalse_2_bufchan_buf <= 1'd0;
      else if (((! es_2_1_1MyFalse_2_argbuf_r) && (! es_2_1_1MyFalse_2_bufchan_buf[0])))
        es_2_1_1MyFalse_2_bufchan_buf <= es_2_1_1MyFalse_2_bufchan_d;
  
  /* fork (Ty Go) : (es_2_1_1MyTrue,Go) > [(es_2_1_1MyTrue_1,Go),
                                      (es_2_1_1MyTrue_2,Go)] */
  logic [1:0] es_2_1_1MyTrue_emitted;
  logic [1:0] es_2_1_1MyTrue_done;
  assign es_2_1_1MyTrue_1_d = (es_2_1_1MyTrue_d[0] && (! es_2_1_1MyTrue_emitted[0]));
  assign es_2_1_1MyTrue_2_d = (es_2_1_1MyTrue_d[0] && (! es_2_1_1MyTrue_emitted[1]));
  assign es_2_1_1MyTrue_done = (es_2_1_1MyTrue_emitted | ({es_2_1_1MyTrue_2_d[0],
                                                           es_2_1_1MyTrue_1_d[0]} & {es_2_1_1MyTrue_2_r,
                                                                                     es_2_1_1MyTrue_1_r}));
  assign es_2_1_1MyTrue_r = (& es_2_1_1MyTrue_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_2_1_1MyTrue_emitted <= 2'd0;
    else
      es_2_1_1MyTrue_emitted <= (es_2_1_1MyTrue_r ? 2'd0 :
                                 es_2_1_1MyTrue_done);
  
  /* dcon (Ty QTree_Int,
      Dcon QNone_Int) : [(es_2_1_1MyTrue_1,Go)] > (es_2_1_1MyTrue_1QNone_Int,QTree_Int) */
  assign es_2_1_1MyTrue_1QNone_Int_d = QNone_Int_dc((& {es_2_1_1MyTrue_1_d[0]}), es_2_1_1MyTrue_1_d);
  assign {es_2_1_1MyTrue_1_r} = {1 {(es_2_1_1MyTrue_1QNone_Int_r && es_2_1_1MyTrue_1QNone_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (es_2_1_1MyTrue_1QNone_Int,QTree_Int) > (lizzieLet16_1_argbuf,QTree_Int) */
  QTree_Int_t es_2_1_1MyTrue_1QNone_Int_bufchan_d;
  logic es_2_1_1MyTrue_1QNone_Int_bufchan_r;
  assign es_2_1_1MyTrue_1QNone_Int_r = ((! es_2_1_1MyTrue_1QNone_Int_bufchan_d[0]) || es_2_1_1MyTrue_1QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_2_1_1MyTrue_1QNone_Int_bufchan_d <= {66'd0, 1'd0};
    else
      if (es_2_1_1MyTrue_1QNone_Int_r)
        es_2_1_1MyTrue_1QNone_Int_bufchan_d <= es_2_1_1MyTrue_1QNone_Int_d;
  QTree_Int_t es_2_1_1MyTrue_1QNone_Int_bufchan_buf;
  assign es_2_1_1MyTrue_1QNone_Int_bufchan_r = (! es_2_1_1MyTrue_1QNone_Int_bufchan_buf[0]);
  assign lizzieLet16_1_argbuf_d = (es_2_1_1MyTrue_1QNone_Int_bufchan_buf[0] ? es_2_1_1MyTrue_1QNone_Int_bufchan_buf :
                                   es_2_1_1MyTrue_1QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_2_1_1MyTrue_1QNone_Int_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((lizzieLet16_1_argbuf_r && es_2_1_1MyTrue_1QNone_Int_bufchan_buf[0]))
        es_2_1_1MyTrue_1QNone_Int_bufchan_buf <= {66'd0, 1'd0};
      else if (((! lizzieLet16_1_argbuf_r) && (! es_2_1_1MyTrue_1QNone_Int_bufchan_buf[0])))
        es_2_1_1MyTrue_1QNone_Int_bufchan_buf <= es_2_1_1MyTrue_1QNone_Int_bufchan_d;
  
  /* buf (Ty Go) : (es_2_1_1MyTrue_2,Go) > (es_2_1_1MyTrue_2_argbuf,Go) */
  Go_t es_2_1_1MyTrue_2_bufchan_d;
  logic es_2_1_1MyTrue_2_bufchan_r;
  assign es_2_1_1MyTrue_2_r = ((! es_2_1_1MyTrue_2_bufchan_d[0]) || es_2_1_1MyTrue_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_2_1_1MyTrue_2_bufchan_d <= 1'd0;
    else
      if (es_2_1_1MyTrue_2_r)
        es_2_1_1MyTrue_2_bufchan_d <= es_2_1_1MyTrue_2_d;
  Go_t es_2_1_1MyTrue_2_bufchan_buf;
  assign es_2_1_1MyTrue_2_bufchan_r = (! es_2_1_1MyTrue_2_bufchan_buf[0]);
  assign es_2_1_1MyTrue_2_argbuf_d = (es_2_1_1MyTrue_2_bufchan_buf[0] ? es_2_1_1MyTrue_2_bufchan_buf :
                                      es_2_1_1MyTrue_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_2_1_1MyTrue_2_bufchan_buf <= 1'd0;
    else
      if ((es_2_1_1MyTrue_2_argbuf_r && es_2_1_1MyTrue_2_bufchan_buf[0]))
        es_2_1_1MyTrue_2_bufchan_buf <= 1'd0;
      else if (((! es_2_1_1MyTrue_2_argbuf_r) && (! es_2_1_1MyTrue_2_bufchan_buf[0])))
        es_2_1_1MyTrue_2_bufchan_buf <= es_2_1_1MyTrue_2_bufchan_d;
  
  /* demux (Ty MyBool,
       Ty MyDTInt_Int) : (es_2_1_2,MyBool) (lizzieLet12_6QNone_Int_5QVal_Int_2,MyDTInt_Int) > [(es_2_1_2MyFalse,MyDTInt_Int),
                                                                                               (_69,MyDTInt_Int)] */
  logic [1:0] lizzieLet12_6QNone_Int_5QVal_Int_2_onehotd;
  always_comb
    if ((es_2_1_2_d[0] && lizzieLet12_6QNone_Int_5QVal_Int_2_d[0]))
      unique case (es_2_1_2_d[1:1])
        1'd0: lizzieLet12_6QNone_Int_5QVal_Int_2_onehotd = 2'd1;
        1'd1: lizzieLet12_6QNone_Int_5QVal_Int_2_onehotd = 2'd2;
        default: lizzieLet12_6QNone_Int_5QVal_Int_2_onehotd = 2'd0;
      endcase
    else lizzieLet12_6QNone_Int_5QVal_Int_2_onehotd = 2'd0;
  assign es_2_1_2MyFalse_d = lizzieLet12_6QNone_Int_5QVal_Int_2_onehotd[0];
  assign _69_d = lizzieLet12_6QNone_Int_5QVal_Int_2_onehotd[1];
  assign lizzieLet12_6QNone_Int_5QVal_Int_2_r = (| (lizzieLet12_6QNone_Int_5QVal_Int_2_onehotd & {_69_r,
                                                                                                  es_2_1_2MyFalse_r}));
  assign es_2_1_2_r = lizzieLet12_6QNone_Int_5QVal_Int_2_r;
  
  /* buf (Ty MyDTInt_Int) : (es_2_1_2MyFalse,MyDTInt_Int) > (es_2_1_2MyFalse_1_argbuf,MyDTInt_Int) */
  MyDTInt_Int_t es_2_1_2MyFalse_bufchan_d;
  logic es_2_1_2MyFalse_bufchan_r;
  assign es_2_1_2MyFalse_r = ((! es_2_1_2MyFalse_bufchan_d[0]) || es_2_1_2MyFalse_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_2_1_2MyFalse_bufchan_d <= 1'd0;
    else
      if (es_2_1_2MyFalse_r)
        es_2_1_2MyFalse_bufchan_d <= es_2_1_2MyFalse_d;
  MyDTInt_Int_t es_2_1_2MyFalse_bufchan_buf;
  assign es_2_1_2MyFalse_bufchan_r = (! es_2_1_2MyFalse_bufchan_buf[0]);
  assign es_2_1_2MyFalse_1_argbuf_d = (es_2_1_2MyFalse_bufchan_buf[0] ? es_2_1_2MyFalse_bufchan_buf :
                                       es_2_1_2MyFalse_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_2_1_2MyFalse_bufchan_buf <= 1'd0;
    else
      if ((es_2_1_2MyFalse_1_argbuf_r && es_2_1_2MyFalse_bufchan_buf[0]))
        es_2_1_2MyFalse_bufchan_buf <= 1'd0;
      else if (((! es_2_1_2MyFalse_1_argbuf_r) && (! es_2_1_2MyFalse_bufchan_buf[0])))
        es_2_1_2MyFalse_bufchan_buf <= es_2_1_2MyFalse_bufchan_d;
  
  /* demux (Ty MyBool,
       Ty Pointer_CTf_f_Int_Int) : (es_2_1_3,MyBool) (lizzieLet12_6QNone_Int_6QVal_Int,Pointer_CTf_f_Int_Int) > [(es_2_1_3MyFalse,Pointer_CTf_f_Int_Int),
                                                                                                                 (es_2_1_3MyTrue,Pointer_CTf_f_Int_Int)] */
  logic [1:0] lizzieLet12_6QNone_Int_6QVal_Int_onehotd;
  always_comb
    if ((es_2_1_3_d[0] && lizzieLet12_6QNone_Int_6QVal_Int_d[0]))
      unique case (es_2_1_3_d[1:1])
        1'd0: lizzieLet12_6QNone_Int_6QVal_Int_onehotd = 2'd1;
        1'd1: lizzieLet12_6QNone_Int_6QVal_Int_onehotd = 2'd2;
        default: lizzieLet12_6QNone_Int_6QVal_Int_onehotd = 2'd0;
      endcase
    else lizzieLet12_6QNone_Int_6QVal_Int_onehotd = 2'd0;
  assign es_2_1_3MyFalse_d = {lizzieLet12_6QNone_Int_6QVal_Int_d[16:1],
                              lizzieLet12_6QNone_Int_6QVal_Int_onehotd[0]};
  assign es_2_1_3MyTrue_d = {lizzieLet12_6QNone_Int_6QVal_Int_d[16:1],
                             lizzieLet12_6QNone_Int_6QVal_Int_onehotd[1]};
  assign lizzieLet12_6QNone_Int_6QVal_Int_r = (| (lizzieLet12_6QNone_Int_6QVal_Int_onehotd & {es_2_1_3MyTrue_r,
                                                                                              es_2_1_3MyFalse_r}));
  assign es_2_1_3_r = lizzieLet12_6QNone_Int_6QVal_Int_r;
  
  /* buf (Ty Pointer_CTf_f_Int_Int) : (es_2_1_3MyFalse,Pointer_CTf_f_Int_Int) > (es_2_1_3MyFalse_1_argbuf,Pointer_CTf_f_Int_Int) */
  Pointer_CTf_f_Int_Int_t es_2_1_3MyFalse_bufchan_d;
  logic es_2_1_3MyFalse_bufchan_r;
  assign es_2_1_3MyFalse_r = ((! es_2_1_3MyFalse_bufchan_d[0]) || es_2_1_3MyFalse_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_2_1_3MyFalse_bufchan_d <= {16'd0, 1'd0};
    else
      if (es_2_1_3MyFalse_r)
        es_2_1_3MyFalse_bufchan_d <= es_2_1_3MyFalse_d;
  Pointer_CTf_f_Int_Int_t es_2_1_3MyFalse_bufchan_buf;
  assign es_2_1_3MyFalse_bufchan_r = (! es_2_1_3MyFalse_bufchan_buf[0]);
  assign es_2_1_3MyFalse_1_argbuf_d = (es_2_1_3MyFalse_bufchan_buf[0] ? es_2_1_3MyFalse_bufchan_buf :
                                       es_2_1_3MyFalse_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_2_1_3MyFalse_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((es_2_1_3MyFalse_1_argbuf_r && es_2_1_3MyFalse_bufchan_buf[0]))
        es_2_1_3MyFalse_bufchan_buf <= {16'd0, 1'd0};
      else if (((! es_2_1_3MyFalse_1_argbuf_r) && (! es_2_1_3MyFalse_bufchan_buf[0])))
        es_2_1_3MyFalse_bufchan_buf <= es_2_1_3MyFalse_bufchan_d;
  
  /* buf (Ty Pointer_CTf_f_Int_Int) : (es_2_1_3MyTrue,Pointer_CTf_f_Int_Int) > (es_2_1_3MyTrue_1_argbuf,Pointer_CTf_f_Int_Int) */
  Pointer_CTf_f_Int_Int_t es_2_1_3MyTrue_bufchan_d;
  logic es_2_1_3MyTrue_bufchan_r;
  assign es_2_1_3MyTrue_r = ((! es_2_1_3MyTrue_bufchan_d[0]) || es_2_1_3MyTrue_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_2_1_3MyTrue_bufchan_d <= {16'd0, 1'd0};
    else
      if (es_2_1_3MyTrue_r) es_2_1_3MyTrue_bufchan_d <= es_2_1_3MyTrue_d;
  Pointer_CTf_f_Int_Int_t es_2_1_3MyTrue_bufchan_buf;
  assign es_2_1_3MyTrue_bufchan_r = (! es_2_1_3MyTrue_bufchan_buf[0]);
  assign es_2_1_3MyTrue_1_argbuf_d = (es_2_1_3MyTrue_bufchan_buf[0] ? es_2_1_3MyTrue_bufchan_buf :
                                      es_2_1_3MyTrue_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_2_1_3MyTrue_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((es_2_1_3MyTrue_1_argbuf_r && es_2_1_3MyTrue_bufchan_buf[0]))
        es_2_1_3MyTrue_bufchan_buf <= {16'd0, 1'd0};
      else if (((! es_2_1_3MyTrue_1_argbuf_r) && (! es_2_1_3MyTrue_bufchan_buf[0])))
        es_2_1_3MyTrue_bufchan_buf <= es_2_1_3MyTrue_bufchan_d;
  
  /* demux (Ty MyBool,
       Ty Int) : (es_2_1_4,MyBool) (va8I_2,Int) > [(es_2_1_4MyFalse,Int),
                                                   (_68,Int)] */
  logic [1:0] va8I_2_onehotd;
  always_comb
    if ((es_2_1_4_d[0] && va8I_2_d[0]))
      unique case (es_2_1_4_d[1:1])
        1'd0: va8I_2_onehotd = 2'd1;
        1'd1: va8I_2_onehotd = 2'd2;
        default: va8I_2_onehotd = 2'd0;
      endcase
    else va8I_2_onehotd = 2'd0;
  assign es_2_1_4MyFalse_d = {va8I_2_d[32:1], va8I_2_onehotd[0]};
  assign _68_d = {va8I_2_d[32:1], va8I_2_onehotd[1]};
  assign va8I_2_r = (| (va8I_2_onehotd & {_68_r,
                                          es_2_1_4MyFalse_r}));
  assign es_2_1_4_r = va8I_2_r;
  
  /* buf (Ty Int) : (es_2_1_4MyFalse,Int) > (es_2_1_4MyFalse_1_argbuf,Int) */
  Int_t es_2_1_4MyFalse_bufchan_d;
  logic es_2_1_4MyFalse_bufchan_r;
  assign es_2_1_4MyFalse_r = ((! es_2_1_4MyFalse_bufchan_d[0]) || es_2_1_4MyFalse_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_2_1_4MyFalse_bufchan_d <= {32'd0, 1'd0};
    else
      if (es_2_1_4MyFalse_r)
        es_2_1_4MyFalse_bufchan_d <= es_2_1_4MyFalse_d;
  Int_t es_2_1_4MyFalse_bufchan_buf;
  assign es_2_1_4MyFalse_bufchan_r = (! es_2_1_4MyFalse_bufchan_buf[0]);
  assign es_2_1_4MyFalse_1_argbuf_d = (es_2_1_4MyFalse_bufchan_buf[0] ? es_2_1_4MyFalse_bufchan_buf :
                                       es_2_1_4MyFalse_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_2_1_4MyFalse_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((es_2_1_4MyFalse_1_argbuf_r && es_2_1_4MyFalse_bufchan_buf[0]))
        es_2_1_4MyFalse_bufchan_buf <= {32'd0, 1'd0};
      else if (((! es_2_1_4MyFalse_1_argbuf_r) && (! es_2_1_4MyFalse_bufchan_buf[0])))
        es_2_1_4MyFalse_bufchan_buf <= es_2_1_4MyFalse_bufchan_d;
  
  /* demux (Ty MyBool,
       Ty MyDTInt_Int) : (es_2_2,MyBool) (lizzieLet6_5QVal_Int_2,MyDTInt_Int) > [(es_2_2MyFalse,MyDTInt_Int),
                                                                                 (_67,MyDTInt_Int)] */
  logic [1:0] lizzieLet6_5QVal_Int_2_onehotd;
  always_comb
    if ((es_2_2_d[0] && lizzieLet6_5QVal_Int_2_d[0]))
      unique case (es_2_2_d[1:1])
        1'd0: lizzieLet6_5QVal_Int_2_onehotd = 2'd1;
        1'd1: lizzieLet6_5QVal_Int_2_onehotd = 2'd2;
        default: lizzieLet6_5QVal_Int_2_onehotd = 2'd0;
      endcase
    else lizzieLet6_5QVal_Int_2_onehotd = 2'd0;
  assign es_2_2MyFalse_d = lizzieLet6_5QVal_Int_2_onehotd[0];
  assign _67_d = lizzieLet6_5QVal_Int_2_onehotd[1];
  assign lizzieLet6_5QVal_Int_2_r = (| (lizzieLet6_5QVal_Int_2_onehotd & {_67_r,
                                                                          es_2_2MyFalse_r}));
  assign es_2_2_r = lizzieLet6_5QVal_Int_2_r;
  
  /* buf (Ty MyDTInt_Int) : (es_2_2MyFalse,MyDTInt_Int) > (es_2_2MyFalse_1_argbuf,MyDTInt_Int) */
  MyDTInt_Int_t es_2_2MyFalse_bufchan_d;
  logic es_2_2MyFalse_bufchan_r;
  assign es_2_2MyFalse_r = ((! es_2_2MyFalse_bufchan_d[0]) || es_2_2MyFalse_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_2_2MyFalse_bufchan_d <= 1'd0;
    else
      if (es_2_2MyFalse_r) es_2_2MyFalse_bufchan_d <= es_2_2MyFalse_d;
  MyDTInt_Int_t es_2_2MyFalse_bufchan_buf;
  assign es_2_2MyFalse_bufchan_r = (! es_2_2MyFalse_bufchan_buf[0]);
  assign es_2_2MyFalse_1_argbuf_d = (es_2_2MyFalse_bufchan_buf[0] ? es_2_2MyFalse_bufchan_buf :
                                     es_2_2MyFalse_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_2_2MyFalse_bufchan_buf <= 1'd0;
    else
      if ((es_2_2MyFalse_1_argbuf_r && es_2_2MyFalse_bufchan_buf[0]))
        es_2_2MyFalse_bufchan_buf <= 1'd0;
      else if (((! es_2_2MyFalse_1_argbuf_r) && (! es_2_2MyFalse_bufchan_buf[0])))
        es_2_2MyFalse_bufchan_buf <= es_2_2MyFalse_bufchan_d;
  
  /* demux (Ty MyBool,
       Ty Pointer_CTf''''''''_f''''''''_Int_Int) : (es_2_3,MyBool) (lizzieLet6_6QVal_Int,Pointer_CTf''''''''_f''''''''_Int_Int) > [(es_2_3MyFalse,Pointer_CTf''''''''_f''''''''_Int_Int),
                                                                                                                                   (es_2_3MyTrue,Pointer_CTf''''''''_f''''''''_Int_Int)] */
  logic [1:0] lizzieLet6_6QVal_Int_onehotd;
  always_comb
    if ((es_2_3_d[0] && lizzieLet6_6QVal_Int_d[0]))
      unique case (es_2_3_d[1:1])
        1'd0: lizzieLet6_6QVal_Int_onehotd = 2'd1;
        1'd1: lizzieLet6_6QVal_Int_onehotd = 2'd2;
        default: lizzieLet6_6QVal_Int_onehotd = 2'd0;
      endcase
    else lizzieLet6_6QVal_Int_onehotd = 2'd0;
  assign es_2_3MyFalse_d = {lizzieLet6_6QVal_Int_d[16:1],
                            lizzieLet6_6QVal_Int_onehotd[0]};
  assign es_2_3MyTrue_d = {lizzieLet6_6QVal_Int_d[16:1],
                           lizzieLet6_6QVal_Int_onehotd[1]};
  assign lizzieLet6_6QVal_Int_r = (| (lizzieLet6_6QVal_Int_onehotd & {es_2_3MyTrue_r,
                                                                      es_2_3MyFalse_r}));
  assign es_2_3_r = lizzieLet6_6QVal_Int_r;
  
  /* buf (Ty Pointer_CTf''''''''_f''''''''_Int_Int) : (es_2_3MyFalse,Pointer_CTf''''''''_f''''''''_Int_Int) > (es_2_3MyFalse_1_argbuf,Pointer_CTf''''''''_f''''''''_Int_Int) */
  \Pointer_CTf''''''''_f''''''''_Int_Int_t  es_2_3MyFalse_bufchan_d;
  logic es_2_3MyFalse_bufchan_r;
  assign es_2_3MyFalse_r = ((! es_2_3MyFalse_bufchan_d[0]) || es_2_3MyFalse_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_2_3MyFalse_bufchan_d <= {16'd0, 1'd0};
    else
      if (es_2_3MyFalse_r) es_2_3MyFalse_bufchan_d <= es_2_3MyFalse_d;
  \Pointer_CTf''''''''_f''''''''_Int_Int_t  es_2_3MyFalse_bufchan_buf;
  assign es_2_3MyFalse_bufchan_r = (! es_2_3MyFalse_bufchan_buf[0]);
  assign es_2_3MyFalse_1_argbuf_d = (es_2_3MyFalse_bufchan_buf[0] ? es_2_3MyFalse_bufchan_buf :
                                     es_2_3MyFalse_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_2_3MyFalse_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((es_2_3MyFalse_1_argbuf_r && es_2_3MyFalse_bufchan_buf[0]))
        es_2_3MyFalse_bufchan_buf <= {16'd0, 1'd0};
      else if (((! es_2_3MyFalse_1_argbuf_r) && (! es_2_3MyFalse_bufchan_buf[0])))
        es_2_3MyFalse_bufchan_buf <= es_2_3MyFalse_bufchan_d;
  
  /* buf (Ty Pointer_CTf''''''''_f''''''''_Int_Int) : (es_2_3MyTrue,Pointer_CTf''''''''_f''''''''_Int_Int) > (es_2_3MyTrue_1_argbuf,Pointer_CTf''''''''_f''''''''_Int_Int) */
  \Pointer_CTf''''''''_f''''''''_Int_Int_t  es_2_3MyTrue_bufchan_d;
  logic es_2_3MyTrue_bufchan_r;
  assign es_2_3MyTrue_r = ((! es_2_3MyTrue_bufchan_d[0]) || es_2_3MyTrue_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_2_3MyTrue_bufchan_d <= {16'd0, 1'd0};
    else if (es_2_3MyTrue_r) es_2_3MyTrue_bufchan_d <= es_2_3MyTrue_d;
  \Pointer_CTf''''''''_f''''''''_Int_Int_t  es_2_3MyTrue_bufchan_buf;
  assign es_2_3MyTrue_bufchan_r = (! es_2_3MyTrue_bufchan_buf[0]);
  assign es_2_3MyTrue_1_argbuf_d = (es_2_3MyTrue_bufchan_buf[0] ? es_2_3MyTrue_bufchan_buf :
                                    es_2_3MyTrue_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_2_3MyTrue_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((es_2_3MyTrue_1_argbuf_r && es_2_3MyTrue_bufchan_buf[0]))
        es_2_3MyTrue_bufchan_buf <= {16'd0, 1'd0};
      else if (((! es_2_3MyTrue_1_argbuf_r) && (! es_2_3MyTrue_bufchan_buf[0])))
        es_2_3MyTrue_bufchan_buf <= es_2_3MyTrue_bufchan_d;
  
  /* demux (Ty MyBool,
       Ty Int) : (es_2_4,MyBool) (va8x_2,Int) > [(es_2_4MyFalse,Int),
                                                 (_66,Int)] */
  logic [1:0] va8x_2_onehotd;
  always_comb
    if ((es_2_4_d[0] && va8x_2_d[0]))
      unique case (es_2_4_d[1:1])
        1'd0: va8x_2_onehotd = 2'd1;
        1'd1: va8x_2_onehotd = 2'd2;
        default: va8x_2_onehotd = 2'd0;
      endcase
    else va8x_2_onehotd = 2'd0;
  assign es_2_4MyFalse_d = {va8x_2_d[32:1], va8x_2_onehotd[0]};
  assign _66_d = {va8x_2_d[32:1], va8x_2_onehotd[1]};
  assign va8x_2_r = (| (va8x_2_onehotd & {_66_r, es_2_4MyFalse_r}));
  assign es_2_4_r = va8x_2_r;
  
  /* buf (Ty Int) : (es_2_4MyFalse,Int) > (es_2_4MyFalse_1_argbuf,Int) */
  Int_t es_2_4MyFalse_bufchan_d;
  logic es_2_4MyFalse_bufchan_r;
  assign es_2_4MyFalse_r = ((! es_2_4MyFalse_bufchan_d[0]) || es_2_4MyFalse_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_2_4MyFalse_bufchan_d <= {32'd0, 1'd0};
    else
      if (es_2_4MyFalse_r) es_2_4MyFalse_bufchan_d <= es_2_4MyFalse_d;
  Int_t es_2_4MyFalse_bufchan_buf;
  assign es_2_4MyFalse_bufchan_r = (! es_2_4MyFalse_bufchan_buf[0]);
  assign es_2_4MyFalse_1_argbuf_d = (es_2_4MyFalse_bufchan_buf[0] ? es_2_4MyFalse_bufchan_buf :
                                     es_2_4MyFalse_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_2_4MyFalse_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((es_2_4MyFalse_1_argbuf_r && es_2_4MyFalse_bufchan_buf[0]))
        es_2_4MyFalse_bufchan_buf <= {32'd0, 1'd0};
      else if (((! es_2_4MyFalse_1_argbuf_r) && (! es_2_4MyFalse_bufchan_buf[0])))
        es_2_4MyFalse_bufchan_buf <= es_2_4MyFalse_bufchan_d;
  
  /* buf (Ty QTree_Int) : (es_3_1_1QVal_Int,QTree_Int) > (lizzieLet8_1_argbuf,QTree_Int) */
  QTree_Int_t es_3_1_1QVal_Int_bufchan_d;
  logic es_3_1_1QVal_Int_bufchan_r;
  assign es_3_1_1QVal_Int_r = ((! es_3_1_1QVal_Int_bufchan_d[0]) || es_3_1_1QVal_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_3_1_1QVal_Int_bufchan_d <= {66'd0, 1'd0};
    else
      if (es_3_1_1QVal_Int_r)
        es_3_1_1QVal_Int_bufchan_d <= es_3_1_1QVal_Int_d;
  QTree_Int_t es_3_1_1QVal_Int_bufchan_buf;
  assign es_3_1_1QVal_Int_bufchan_r = (! es_3_1_1QVal_Int_bufchan_buf[0]);
  assign lizzieLet8_1_argbuf_d = (es_3_1_1QVal_Int_bufchan_buf[0] ? es_3_1_1QVal_Int_bufchan_buf :
                                  es_3_1_1QVal_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_3_1_1QVal_Int_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((lizzieLet8_1_argbuf_r && es_3_1_1QVal_Int_bufchan_buf[0]))
        es_3_1_1QVal_Int_bufchan_buf <= {66'd0, 1'd0};
      else if (((! lizzieLet8_1_argbuf_r) && (! es_3_1_1QVal_Int_bufchan_buf[0])))
        es_3_1_1QVal_Int_bufchan_buf <= es_3_1_1QVal_Int_bufchan_d;
  
  /* buf (Ty QTree_Int) : (es_3_2_1QVal_Int,QTree_Int) > (lizzieLet15_1_argbuf,QTree_Int) */
  QTree_Int_t es_3_2_1QVal_Int_bufchan_d;
  logic es_3_2_1QVal_Int_bufchan_r;
  assign es_3_2_1QVal_Int_r = ((! es_3_2_1QVal_Int_bufchan_d[0]) || es_3_2_1QVal_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_3_2_1QVal_Int_bufchan_d <= {66'd0, 1'd0};
    else
      if (es_3_2_1QVal_Int_r)
        es_3_2_1QVal_Int_bufchan_d <= es_3_2_1QVal_Int_d;
  QTree_Int_t es_3_2_1QVal_Int_bufchan_buf;
  assign es_3_2_1QVal_Int_bufchan_r = (! es_3_2_1QVal_Int_bufchan_buf[0]);
  assign lizzieLet15_1_argbuf_d = (es_3_2_1QVal_Int_bufchan_buf[0] ? es_3_2_1QVal_Int_bufchan_buf :
                                   es_3_2_1QVal_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_3_2_1QVal_Int_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((lizzieLet15_1_argbuf_r && es_3_2_1QVal_Int_bufchan_buf[0]))
        es_3_2_1QVal_Int_bufchan_buf <= {66'd0, 1'd0};
      else if (((! lizzieLet15_1_argbuf_r) && (! es_3_2_1QVal_Int_bufchan_buf[0])))
        es_3_2_1QVal_Int_bufchan_buf <= es_3_2_1QVal_Int_bufchan_d;
  
  /* buf (Ty QTree_Int) : (es_4_1_1es_5_1_1es_6_1_1es_7_1_1QNode_Int,QTree_Int) > (lizzieLet17_1_argbuf,QTree_Int) */
  QTree_Int_t es_4_1_1es_5_1_1es_6_1_1es_7_1_1QNode_Int_bufchan_d;
  logic es_4_1_1es_5_1_1es_6_1_1es_7_1_1QNode_Int_bufchan_r;
  assign es_4_1_1es_5_1_1es_6_1_1es_7_1_1QNode_Int_r = ((! es_4_1_1es_5_1_1es_6_1_1es_7_1_1QNode_Int_bufchan_d[0]) || es_4_1_1es_5_1_1es_6_1_1es_7_1_1QNode_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_4_1_1es_5_1_1es_6_1_1es_7_1_1QNode_Int_bufchan_d <= {66'd0,
                                                              1'd0};
    else
      if (es_4_1_1es_5_1_1es_6_1_1es_7_1_1QNode_Int_r)
        es_4_1_1es_5_1_1es_6_1_1es_7_1_1QNode_Int_bufchan_d <= es_4_1_1es_5_1_1es_6_1_1es_7_1_1QNode_Int_d;
  QTree_Int_t es_4_1_1es_5_1_1es_6_1_1es_7_1_1QNode_Int_bufchan_buf;
  assign es_4_1_1es_5_1_1es_6_1_1es_7_1_1QNode_Int_bufchan_r = (! es_4_1_1es_5_1_1es_6_1_1es_7_1_1QNode_Int_bufchan_buf[0]);
  assign lizzieLet17_1_argbuf_d = (es_4_1_1es_5_1_1es_6_1_1es_7_1_1QNode_Int_bufchan_buf[0] ? es_4_1_1es_5_1_1es_6_1_1es_7_1_1QNode_Int_bufchan_buf :
                                   es_4_1_1es_5_1_1es_6_1_1es_7_1_1QNode_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_4_1_1es_5_1_1es_6_1_1es_7_1_1QNode_Int_bufchan_buf <= {66'd0,
                                                                1'd0};
    else
      if ((lizzieLet17_1_argbuf_r && es_4_1_1es_5_1_1es_6_1_1es_7_1_1QNode_Int_bufchan_buf[0]))
        es_4_1_1es_5_1_1es_6_1_1es_7_1_1QNode_Int_bufchan_buf <= {66'd0,
                                                                  1'd0};
      else if (((! lizzieLet17_1_argbuf_r) && (! es_4_1_1es_5_1_1es_6_1_1es_7_1_1QNode_Int_bufchan_buf[0])))
        es_4_1_1es_5_1_1es_6_1_1es_7_1_1QNode_Int_bufchan_buf <= es_4_1_1es_5_1_1es_6_1_1es_7_1_1QNode_Int_bufchan_d;
  
  /* buf (Ty Int#) : (es_4_2_1lizzieLet35_4Lcall_$wnnz0_1_Add32,Int#) > (contRet_0_1_argbuf,Int#) */
  \Int#_t  es_4_2_1lizzieLet35_4Lcall_$wnnz0_1_Add32_bufchan_d;
  logic es_4_2_1lizzieLet35_4Lcall_$wnnz0_1_Add32_bufchan_r;
  assign es_4_2_1lizzieLet35_4Lcall_$wnnz0_1_Add32_r = ((! es_4_2_1lizzieLet35_4Lcall_$wnnz0_1_Add32_bufchan_d[0]) || es_4_2_1lizzieLet35_4Lcall_$wnnz0_1_Add32_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_4_2_1lizzieLet35_4Lcall_$wnnz0_1_Add32_bufchan_d <= {32'd0,
                                                              1'd0};
    else
      if (es_4_2_1lizzieLet35_4Lcall_$wnnz0_1_Add32_r)
        es_4_2_1lizzieLet35_4Lcall_$wnnz0_1_Add32_bufchan_d <= es_4_2_1lizzieLet35_4Lcall_$wnnz0_1_Add32_d;
  \Int#_t  es_4_2_1lizzieLet35_4Lcall_$wnnz0_1_Add32_bufchan_buf;
  assign es_4_2_1lizzieLet35_4Lcall_$wnnz0_1_Add32_bufchan_r = (! es_4_2_1lizzieLet35_4Lcall_$wnnz0_1_Add32_bufchan_buf[0]);
  assign contRet_0_1_argbuf_d = (es_4_2_1lizzieLet35_4Lcall_$wnnz0_1_Add32_bufchan_buf[0] ? es_4_2_1lizzieLet35_4Lcall_$wnnz0_1_Add32_bufchan_buf :
                                 es_4_2_1lizzieLet35_4Lcall_$wnnz0_1_Add32_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_4_2_1lizzieLet35_4Lcall_$wnnz0_1_Add32_bufchan_buf <= {32'd0,
                                                                1'd0};
    else
      if ((contRet_0_1_argbuf_r && es_4_2_1lizzieLet35_4Lcall_$wnnz0_1_Add32_bufchan_buf[0]))
        es_4_2_1lizzieLet35_4Lcall_$wnnz0_1_Add32_bufchan_buf <= {32'd0,
                                                                  1'd0};
      else if (((! contRet_0_1_argbuf_r) && (! es_4_2_1lizzieLet35_4Lcall_$wnnz0_1_Add32_bufchan_buf[0])))
        es_4_2_1lizzieLet35_4Lcall_$wnnz0_1_Add32_bufchan_buf <= es_4_2_1lizzieLet35_4Lcall_$wnnz0_1_Add32_bufchan_d;
  
  /* op_add (Ty Int#) : (es_6_2_1ww2Xjx_1_1_Add32,Int#) (lizzieLet35_4Lcall_$wnnz0,Int#) > (es_4_2_1lizzieLet35_4Lcall_$wnnz0_1_Add32,Int#) */
  assign es_4_2_1lizzieLet35_4Lcall_$wnnz0_1_Add32_d = {(es_6_2_1ww2Xjx_1_1_Add32_d[32:1] + lizzieLet35_4Lcall_$wnnz0_d[32:1]),
                                                        (es_6_2_1ww2Xjx_1_1_Add32_d[0] && lizzieLet35_4Lcall_$wnnz0_d[0])};
  assign {es_6_2_1ww2Xjx_1_1_Add32_r,
          lizzieLet35_4Lcall_$wnnz0_r} = {2 {(es_4_2_1lizzieLet35_4Lcall_$wnnz0_1_Add32_r && es_4_2_1lizzieLet35_4Lcall_$wnnz0_1_Add32_d[0])}};
  
  /* sink (Ty Int) : (es_7_1I#,Int) > */
  assign {\es_7_1I#_r , \es_7_1I#_dout } = {\es_7_1I#_rout ,
                                            \es_7_1I#_d };
  
  /* mergectrl (Ty C8,
           Ty TupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int) : [(f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_1,TupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int),
                                                                         (f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int2,TupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int),
                                                                         (f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int3,TupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int),
                                                                         (f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int4,TupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int),
                                                                         (f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int5,TupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int),
                                                                         (f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int6,TupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int),
                                                                         (f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int7,TupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int),
                                                                         (f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int8,TupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int)] > (f''''''''_f''''''''_Int_Int_choice,C8) (f''''''''_f''''''''_Int_Int_data,TupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int) */
  logic [7:0] \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_1_select_d ;
  assign \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_1_select_d  = ((| \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_1_select_q ) ? \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_1_select_q  :
                                                                                                           (\f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_1_d [0] ? 8'd1 :
                                                                                                            (\f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int2_d [0] ? 8'd2 :
                                                                                                             (\f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int3_d [0] ? 8'd4 :
                                                                                                              (\f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int4_d [0] ? 8'd8 :
                                                                                                               (\f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int5_d [0] ? 8'd16 :
                                                                                                                (\f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int6_d [0] ? 8'd32 :
                                                                                                                 (\f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int7_d [0] ? 8'd64 :
                                                                                                                  (\f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int8_d [0] ? 8'd128 :
                                                                                                                   8'd0)))))))));
  logic [7:0] \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_1_select_q ;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_1_select_q  <= 8'd0;
    else
      \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_1_select_q  <= (\f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_1_done  ? 8'd0 :
                                                                                                         \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_1_select_d );
  logic [1:0] \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_1_emit_q ;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_1_emit_q  <= 2'd0;
    else
      \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_1_emit_q  <= (\f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_1_done  ? 2'd0 :
                                                                                                       \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_1_emit_d );
  logic [1:0] \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_1_emit_d ;
  assign \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_1_emit_d  = (\f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_1_emit_q  | ({\f''''''''_f''''''''_Int_Int_choice_d [0],
                                                                                                                                                                                                          \f''''''''_f''''''''_Int_Int_data_d [0]} & {\f''''''''_f''''''''_Int_Int_choice_r ,
                                                                                                                                                                                                                                                      \f''''''''_f''''''''_Int_Int_data_r }));
  logic \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_1_done ;
  assign \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_1_done  = (& \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_1_emit_d );
  assign {\f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int8_r ,
          \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int7_r ,
          \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int6_r ,
          \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int5_r ,
          \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int4_r ,
          \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int3_r ,
          \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int2_r ,
          \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_1_r } = (\f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_1_done  ? \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_1_select_d  :
                                                                                                      8'd0);
  assign \f''''''''_f''''''''_Int_Int_data_d  = ((\f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_1_select_d [0] && (! \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_1_emit_q [0])) ? \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_1_d  :
                                                 ((\f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_1_select_d [1] && (! \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_1_emit_q [0])) ? \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int2_d  :
                                                  ((\f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_1_select_d [2] && (! \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_1_emit_q [0])) ? \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int3_d  :
                                                   ((\f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_1_select_d [3] && (! \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_1_emit_q [0])) ? \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int4_d  :
                                                    ((\f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_1_select_d [4] && (! \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_1_emit_q [0])) ? \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int5_d  :
                                                     ((\f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_1_select_d [5] && (! \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_1_emit_q [0])) ? \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int6_d  :
                                                      ((\f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_1_select_d [6] && (! \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_1_emit_q [0])) ? \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int7_d  :
                                                       ((\f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_1_select_d [7] && (! \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_1_emit_q [0])) ? \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int8_d  :
                                                        {16'd0, 1'd0}))))))));
  assign \f''''''''_f''''''''_Int_Int_choice_d  = ((\f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_1_select_d [0] && (! \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_1_emit_q [1])) ? C1_8_dc(1'd1) :
                                                   ((\f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_1_select_d [1] && (! \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_1_emit_q [1])) ? C2_8_dc(1'd1) :
                                                    ((\f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_1_select_d [2] && (! \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_1_emit_q [1])) ? C3_8_dc(1'd1) :
                                                     ((\f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_1_select_d [3] && (! \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_1_emit_q [1])) ? C4_8_dc(1'd1) :
                                                      ((\f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_1_select_d [4] && (! \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_1_emit_q [1])) ? C5_8_dc(1'd1) :
                                                       ((\f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_1_select_d [5] && (! \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_1_emit_q [1])) ? C6_8_dc(1'd1) :
                                                        ((\f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_1_select_d [6] && (! \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_1_emit_q [1])) ? C7_8_dc(1'd1) :
                                                         ((\f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_1_select_d [7] && (! \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_1_emit_q [1])) ? C8_8_dc(1'd1) :
                                                          {3'd0, 1'd0}))))))));
  
  /* fork (Ty Go) : (f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Intgo_13,Go) > [(go_13_1,Go),
                                                                                                              (go_13_2,Go)] */
  logic [1:0] \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Intgo_13_emitted ;
  logic [1:0] \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Intgo_13_done ;
  assign go_13_1_d = (\f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Intgo_13_d [0] && (! \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Intgo_13_emitted [0]));
  assign go_13_2_d = (\f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Intgo_13_d [0] && (! \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Intgo_13_emitted [1]));
  assign \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Intgo_13_done  = (\f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Intgo_13_emitted  | ({go_13_2_d[0],
                                                                                                                                                                                                               go_13_1_d[0]} & {go_13_2_r,
                                                                                                                                                                                                                                go_13_1_r}));
  assign \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Intgo_13_r  = (& \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Intgo_13_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Intgo_13_emitted  <= 2'd0;
    else
      \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Intgo_13_emitted  <= (\f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Intgo_13_r  ? 2'd0 :
                                                                                                           \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Intgo_13_done );
  
  /* buf (Ty MyDTInt_Bool) : (f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Intis_z_mapa8v_1,MyDTInt_Bool) > (is_z_mapa8v_1_1_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Intis_z_mapa8v_1_bufchan_d ;
  logic \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Intis_z_mapa8v_1_bufchan_r ;
  assign \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Intis_z_mapa8v_1_r  = ((! \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Intis_z_mapa8v_1_bufchan_d [0]) || \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Intis_z_mapa8v_1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Intis_z_mapa8v_1_bufchan_d  <= 1'd0;
    else
      if (\f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Intis_z_mapa8v_1_r )
        \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Intis_z_mapa8v_1_bufchan_d  <= \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Intis_z_mapa8v_1_d ;
  MyDTInt_Bool_t \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Intis_z_mapa8v_1_bufchan_buf ;
  assign \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Intis_z_mapa8v_1_bufchan_r  = (! \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Intis_z_mapa8v_1_bufchan_buf [0]);
  assign is_z_mapa8v_1_1_argbuf_d = (\f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Intis_z_mapa8v_1_bufchan_buf [0] ? \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Intis_z_mapa8v_1_bufchan_buf  :
                                     \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Intis_z_mapa8v_1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Intis_z_mapa8v_1_bufchan_buf  <= 1'd0;
    else
      if ((is_z_mapa8v_1_1_argbuf_r && \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Intis_z_mapa8v_1_bufchan_buf [0]))
        \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Intis_z_mapa8v_1_bufchan_buf  <= 1'd0;
      else if (((! is_z_mapa8v_1_1_argbuf_r) && (! \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Intis_z_mapa8v_1_bufchan_buf [0])))
        \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Intis_z_mapa8v_1_bufchan_buf  <= \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Intis_z_mapa8v_1_bufchan_d ;
  
  /* buf (Ty MyDTInt_Int) : (f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Intop_mapa8w_1,MyDTInt_Int) > (op_mapa8w_1_1_argbuf,MyDTInt_Int) */
  MyDTInt_Int_t \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Intop_mapa8w_1_bufchan_d ;
  logic \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Intop_mapa8w_1_bufchan_r ;
  assign \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Intop_mapa8w_1_r  = ((! \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Intop_mapa8w_1_bufchan_d [0]) || \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Intop_mapa8w_1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Intop_mapa8w_1_bufchan_d  <= 1'd0;
    else
      if (\f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Intop_mapa8w_1_r )
        \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Intop_mapa8w_1_bufchan_d  <= \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Intop_mapa8w_1_d ;
  MyDTInt_Int_t \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Intop_mapa8w_1_bufchan_buf ;
  assign \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Intop_mapa8w_1_bufchan_r  = (! \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Intop_mapa8w_1_bufchan_buf [0]);
  assign op_mapa8w_1_1_argbuf_d = (\f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Intop_mapa8w_1_bufchan_buf [0] ? \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Intop_mapa8w_1_bufchan_buf  :
                                   \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Intop_mapa8w_1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Intop_mapa8w_1_bufchan_buf  <= 1'd0;
    else
      if ((op_mapa8w_1_1_argbuf_r && \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Intop_mapa8w_1_bufchan_buf [0]))
        \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Intop_mapa8w_1_bufchan_buf  <= 1'd0;
      else if (((! op_mapa8w_1_1_argbuf_r) && (! \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Intop_mapa8w_1_bufchan_buf [0])))
        \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Intop_mapa8w_1_bufchan_buf  <= \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Intop_mapa8w_1_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Int) : (f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Intq4a8u_1,Pointer_QTree_Int) > (q4a8u_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Intq4a8u_1_bufchan_d ;
  logic \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Intq4a8u_1_bufchan_r ;
  assign \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Intq4a8u_1_r  = ((! \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Intq4a8u_1_bufchan_d [0]) || \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Intq4a8u_1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Intq4a8u_1_bufchan_d  <= {16'd0,
                                                                                                               1'd0};
    else
      if (\f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Intq4a8u_1_r )
        \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Intq4a8u_1_bufchan_d  <= \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Intq4a8u_1_d ;
  Pointer_QTree_Int_t \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Intq4a8u_1_bufchan_buf ;
  assign \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Intq4a8u_1_bufchan_r  = (! \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Intq4a8u_1_bufchan_buf [0]);
  assign q4a8u_1_1_argbuf_d = (\f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Intq4a8u_1_bufchan_buf [0] ? \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Intq4a8u_1_bufchan_buf  :
                               \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Intq4a8u_1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Intq4a8u_1_bufchan_buf  <= {16'd0,
                                                                                                                 1'd0};
    else
      if ((q4a8u_1_1_argbuf_r && \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Intq4a8u_1_bufchan_buf [0]))
        \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Intq4a8u_1_bufchan_buf  <= {16'd0,
                                                                                                                   1'd0};
      else if (((! q4a8u_1_1_argbuf_r) && (! \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Intq4a8u_1_bufchan_buf [0])))
        \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Intq4a8u_1_bufchan_buf  <= \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Intq4a8u_1_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Int) : (f''''''''_f''''''''_Int_Int_1,Pointer_QTree_Int) > (f''''''''_f''''''''_Int_Int_resbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t \f''''''''_f''''''''_Int_Int_1_bufchan_d ;
  logic \f''''''''_f''''''''_Int_Int_1_bufchan_r ;
  assign \f''''''''_f''''''''_Int_Int_1_r  = ((! \f''''''''_f''''''''_Int_Int_1_bufchan_d [0]) || \f''''''''_f''''''''_Int_Int_1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''_f''''''''_Int_Int_1_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\f''''''''_f''''''''_Int_Int_1_r )
        \f''''''''_f''''''''_Int_Int_1_bufchan_d  <= \f''''''''_f''''''''_Int_Int_1_d ;
  Pointer_QTree_Int_t \f''''''''_f''''''''_Int_Int_1_bufchan_buf ;
  assign \f''''''''_f''''''''_Int_Int_1_bufchan_r  = (! \f''''''''_f''''''''_Int_Int_1_bufchan_buf [0]);
  assign \f''''''''_f''''''''_Int_Int_resbuf_d  = (\f''''''''_f''''''''_Int_Int_1_bufchan_buf [0] ? \f''''''''_f''''''''_Int_Int_1_bufchan_buf  :
                                                   \f''''''''_f''''''''_Int_Int_1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''_f''''''''_Int_Int_1_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((\f''''''''_f''''''''_Int_Int_resbuf_r  && \f''''''''_f''''''''_Int_Int_1_bufchan_buf [0]))
        \f''''''''_f''''''''_Int_Int_1_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! \f''''''''_f''''''''_Int_Int_resbuf_r ) && (! \f''''''''_f''''''''_Int_Int_1_bufchan_buf [0])))
        \f''''''''_f''''''''_Int_Int_1_bufchan_buf  <= \f''''''''_f''''''''_Int_Int_1_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Int) : (f''''''''_f''''''''_Int_Int_2,Pointer_QTree_Int) > (f''''''''_f''''''''_Int_Int_2_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t \f''''''''_f''''''''_Int_Int_2_bufchan_d ;
  logic \f''''''''_f''''''''_Int_Int_2_bufchan_r ;
  assign \f''''''''_f''''''''_Int_Int_2_r  = ((! \f''''''''_f''''''''_Int_Int_2_bufchan_d [0]) || \f''''''''_f''''''''_Int_Int_2_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''_f''''''''_Int_Int_2_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\f''''''''_f''''''''_Int_Int_2_r )
        \f''''''''_f''''''''_Int_Int_2_bufchan_d  <= \f''''''''_f''''''''_Int_Int_2_d ;
  Pointer_QTree_Int_t \f''''''''_f''''''''_Int_Int_2_bufchan_buf ;
  assign \f''''''''_f''''''''_Int_Int_2_bufchan_r  = (! \f''''''''_f''''''''_Int_Int_2_bufchan_buf [0]);
  assign \f''''''''_f''''''''_Int_Int_2_argbuf_d  = (\f''''''''_f''''''''_Int_Int_2_bufchan_buf [0] ? \f''''''''_f''''''''_Int_Int_2_bufchan_buf  :
                                                     \f''''''''_f''''''''_Int_Int_2_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''_f''''''''_Int_Int_2_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((\f''''''''_f''''''''_Int_Int_2_argbuf_r  && \f''''''''_f''''''''_Int_Int_2_bufchan_buf [0]))
        \f''''''''_f''''''''_Int_Int_2_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! \f''''''''_f''''''''_Int_Int_2_argbuf_r ) && (! \f''''''''_f''''''''_Int_Int_2_bufchan_buf [0])))
        \f''''''''_f''''''''_Int_Int_2_bufchan_buf  <= \f''''''''_f''''''''_Int_Int_2_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Int) : (f''''''''_f''''''''_Int_Int_3,Pointer_QTree_Int) > (f''''''''_f''''''''_Int_Int_3_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t \f''''''''_f''''''''_Int_Int_3_bufchan_d ;
  logic \f''''''''_f''''''''_Int_Int_3_bufchan_r ;
  assign \f''''''''_f''''''''_Int_Int_3_r  = ((! \f''''''''_f''''''''_Int_Int_3_bufchan_d [0]) || \f''''''''_f''''''''_Int_Int_3_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''_f''''''''_Int_Int_3_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\f''''''''_f''''''''_Int_Int_3_r )
        \f''''''''_f''''''''_Int_Int_3_bufchan_d  <= \f''''''''_f''''''''_Int_Int_3_d ;
  Pointer_QTree_Int_t \f''''''''_f''''''''_Int_Int_3_bufchan_buf ;
  assign \f''''''''_f''''''''_Int_Int_3_bufchan_r  = (! \f''''''''_f''''''''_Int_Int_3_bufchan_buf [0]);
  assign \f''''''''_f''''''''_Int_Int_3_argbuf_d  = (\f''''''''_f''''''''_Int_Int_3_bufchan_buf [0] ? \f''''''''_f''''''''_Int_Int_3_bufchan_buf  :
                                                     \f''''''''_f''''''''_Int_Int_3_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''_f''''''''_Int_Int_3_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((\f''''''''_f''''''''_Int_Int_3_argbuf_r  && \f''''''''_f''''''''_Int_Int_3_bufchan_buf [0]))
        \f''''''''_f''''''''_Int_Int_3_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! \f''''''''_f''''''''_Int_Int_3_argbuf_r ) && (! \f''''''''_f''''''''_Int_Int_3_bufchan_buf [0])))
        \f''''''''_f''''''''_Int_Int_3_bufchan_buf  <= \f''''''''_f''''''''_Int_Int_3_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Int) : (f''''''''_f''''''''_Int_Int_4,Pointer_QTree_Int) > (f''''''''_f''''''''_Int_Int_4_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t \f''''''''_f''''''''_Int_Int_4_bufchan_d ;
  logic \f''''''''_f''''''''_Int_Int_4_bufchan_r ;
  assign \f''''''''_f''''''''_Int_Int_4_r  = ((! \f''''''''_f''''''''_Int_Int_4_bufchan_d [0]) || \f''''''''_f''''''''_Int_Int_4_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''_f''''''''_Int_Int_4_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\f''''''''_f''''''''_Int_Int_4_r )
        \f''''''''_f''''''''_Int_Int_4_bufchan_d  <= \f''''''''_f''''''''_Int_Int_4_d ;
  Pointer_QTree_Int_t \f''''''''_f''''''''_Int_Int_4_bufchan_buf ;
  assign \f''''''''_f''''''''_Int_Int_4_bufchan_r  = (! \f''''''''_f''''''''_Int_Int_4_bufchan_buf [0]);
  assign \f''''''''_f''''''''_Int_Int_4_argbuf_d  = (\f''''''''_f''''''''_Int_Int_4_bufchan_buf [0] ? \f''''''''_f''''''''_Int_Int_4_bufchan_buf  :
                                                     \f''''''''_f''''''''_Int_Int_4_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''_f''''''''_Int_Int_4_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((\f''''''''_f''''''''_Int_Int_4_argbuf_r  && \f''''''''_f''''''''_Int_Int_4_bufchan_buf [0]))
        \f''''''''_f''''''''_Int_Int_4_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! \f''''''''_f''''''''_Int_Int_4_argbuf_r ) && (! \f''''''''_f''''''''_Int_Int_4_bufchan_buf [0])))
        \f''''''''_f''''''''_Int_Int_4_bufchan_buf  <= \f''''''''_f''''''''_Int_Int_4_bufchan_d ;
  
  /* dcon (Ty QTree_Int,
      Dcon QNode_Int) : [(f''''''''_f''''''''_Int_Int_4_argbuf,Pointer_QTree_Int),
                         (f''''''''_f''''''''_Int_Int_3_argbuf,Pointer_QTree_Int),
                         (f''''''''_f''''''''_Int_Int_2_argbuf,Pointer_QTree_Int),
                         (f''''''''_f''''''''_Int_Int_resbuf,Pointer_QTree_Int)] > (es_4_1_1es_5_1_1es_6_1_1es_7_1_1QNode_Int,QTree_Int) */
  assign es_4_1_1es_5_1_1es_6_1_1es_7_1_1QNode_Int_d = QNode_Int_dc((& {\f''''''''_f''''''''_Int_Int_4_argbuf_d [0],
                                                                        \f''''''''_f''''''''_Int_Int_3_argbuf_d [0],
                                                                        \f''''''''_f''''''''_Int_Int_2_argbuf_d [0],
                                                                        \f''''''''_f''''''''_Int_Int_resbuf_d [0]}), \f''''''''_f''''''''_Int_Int_4_argbuf_d , \f''''''''_f''''''''_Int_Int_3_argbuf_d , \f''''''''_f''''''''_Int_Int_2_argbuf_d , \f''''''''_f''''''''_Int_Int_resbuf_d );
  assign {\f''''''''_f''''''''_Int_Int_4_argbuf_r ,
          \f''''''''_f''''''''_Int_Int_3_argbuf_r ,
          \f''''''''_f''''''''_Int_Int_2_argbuf_r ,
          \f''''''''_f''''''''_Int_Int_resbuf_r } = {4 {(es_4_1_1es_5_1_1es_6_1_1es_7_1_1QNode_Int_r && es_4_1_1es_5_1_1es_6_1_1es_7_1_1QNode_Int_d[0])}};
  
  /* buf (Ty Pointer_QTree_Int) : (f''''''''_f''''''''_Int_Int_5,Pointer_QTree_Int) > (f''''''''_f''''''''_Int_Int_5_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t \f''''''''_f''''''''_Int_Int_5_bufchan_d ;
  logic \f''''''''_f''''''''_Int_Int_5_bufchan_r ;
  assign \f''''''''_f''''''''_Int_Int_5_r  = ((! \f''''''''_f''''''''_Int_Int_5_bufchan_d [0]) || \f''''''''_f''''''''_Int_Int_5_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''_f''''''''_Int_Int_5_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\f''''''''_f''''''''_Int_Int_5_r )
        \f''''''''_f''''''''_Int_Int_5_bufchan_d  <= \f''''''''_f''''''''_Int_Int_5_d ;
  Pointer_QTree_Int_t \f''''''''_f''''''''_Int_Int_5_bufchan_buf ;
  assign \f''''''''_f''''''''_Int_Int_5_bufchan_r  = (! \f''''''''_f''''''''_Int_Int_5_bufchan_buf [0]);
  assign \f''''''''_f''''''''_Int_Int_5_argbuf_d  = (\f''''''''_f''''''''_Int_Int_5_bufchan_buf [0] ? \f''''''''_f''''''''_Int_Int_5_bufchan_buf  :
                                                     \f''''''''_f''''''''_Int_Int_5_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''_f''''''''_Int_Int_5_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((\f''''''''_f''''''''_Int_Int_5_argbuf_r  && \f''''''''_f''''''''_Int_Int_5_bufchan_buf [0]))
        \f''''''''_f''''''''_Int_Int_5_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! \f''''''''_f''''''''_Int_Int_5_argbuf_r ) && (! \f''''''''_f''''''''_Int_Int_5_bufchan_buf [0])))
        \f''''''''_f''''''''_Int_Int_5_bufchan_buf  <= \f''''''''_f''''''''_Int_Int_5_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Int) : (f''''''''_f''''''''_Int_Int_6,Pointer_QTree_Int) > (f''''''''_f''''''''_Int_Int_6_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t \f''''''''_f''''''''_Int_Int_6_bufchan_d ;
  logic \f''''''''_f''''''''_Int_Int_6_bufchan_r ;
  assign \f''''''''_f''''''''_Int_Int_6_r  = ((! \f''''''''_f''''''''_Int_Int_6_bufchan_d [0]) || \f''''''''_f''''''''_Int_Int_6_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''_f''''''''_Int_Int_6_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\f''''''''_f''''''''_Int_Int_6_r )
        \f''''''''_f''''''''_Int_Int_6_bufchan_d  <= \f''''''''_f''''''''_Int_Int_6_d ;
  Pointer_QTree_Int_t \f''''''''_f''''''''_Int_Int_6_bufchan_buf ;
  assign \f''''''''_f''''''''_Int_Int_6_bufchan_r  = (! \f''''''''_f''''''''_Int_Int_6_bufchan_buf [0]);
  assign \f''''''''_f''''''''_Int_Int_6_argbuf_d  = (\f''''''''_f''''''''_Int_Int_6_bufchan_buf [0] ? \f''''''''_f''''''''_Int_Int_6_bufchan_buf  :
                                                     \f''''''''_f''''''''_Int_Int_6_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''_f''''''''_Int_Int_6_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((\f''''''''_f''''''''_Int_Int_6_argbuf_r  && \f''''''''_f''''''''_Int_Int_6_bufchan_buf [0]))
        \f''''''''_f''''''''_Int_Int_6_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! \f''''''''_f''''''''_Int_Int_6_argbuf_r ) && (! \f''''''''_f''''''''_Int_Int_6_bufchan_buf [0])))
        \f''''''''_f''''''''_Int_Int_6_bufchan_buf  <= \f''''''''_f''''''''_Int_Int_6_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Int) : (f''''''''_f''''''''_Int_Int_7,Pointer_QTree_Int) > (f''''''''_f''''''''_Int_Int_7_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t \f''''''''_f''''''''_Int_Int_7_bufchan_d ;
  logic \f''''''''_f''''''''_Int_Int_7_bufchan_r ;
  assign \f''''''''_f''''''''_Int_Int_7_r  = ((! \f''''''''_f''''''''_Int_Int_7_bufchan_d [0]) || \f''''''''_f''''''''_Int_Int_7_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''_f''''''''_Int_Int_7_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\f''''''''_f''''''''_Int_Int_7_r )
        \f''''''''_f''''''''_Int_Int_7_bufchan_d  <= \f''''''''_f''''''''_Int_Int_7_d ;
  Pointer_QTree_Int_t \f''''''''_f''''''''_Int_Int_7_bufchan_buf ;
  assign \f''''''''_f''''''''_Int_Int_7_bufchan_r  = (! \f''''''''_f''''''''_Int_Int_7_bufchan_buf [0]);
  assign \f''''''''_f''''''''_Int_Int_7_argbuf_d  = (\f''''''''_f''''''''_Int_Int_7_bufchan_buf [0] ? \f''''''''_f''''''''_Int_Int_7_bufchan_buf  :
                                                     \f''''''''_f''''''''_Int_Int_7_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''_f''''''''_Int_Int_7_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((\f''''''''_f''''''''_Int_Int_7_argbuf_r  && \f''''''''_f''''''''_Int_Int_7_bufchan_buf [0]))
        \f''''''''_f''''''''_Int_Int_7_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! \f''''''''_f''''''''_Int_Int_7_argbuf_r ) && (! \f''''''''_f''''''''_Int_Int_7_bufchan_buf [0])))
        \f''''''''_f''''''''_Int_Int_7_bufchan_buf  <= \f''''''''_f''''''''_Int_Int_7_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Int) : (f''''''''_f''''''''_Int_Int_8,Pointer_QTree_Int) > (f''''''''_f''''''''_Int_Int_8_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t \f''''''''_f''''''''_Int_Int_8_bufchan_d ;
  logic \f''''''''_f''''''''_Int_Int_8_bufchan_r ;
  assign \f''''''''_f''''''''_Int_Int_8_r  = ((! \f''''''''_f''''''''_Int_Int_8_bufchan_d [0]) || \f''''''''_f''''''''_Int_Int_8_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''_f''''''''_Int_Int_8_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\f''''''''_f''''''''_Int_Int_8_r )
        \f''''''''_f''''''''_Int_Int_8_bufchan_d  <= \f''''''''_f''''''''_Int_Int_8_d ;
  Pointer_QTree_Int_t \f''''''''_f''''''''_Int_Int_8_bufchan_buf ;
  assign \f''''''''_f''''''''_Int_Int_8_bufchan_r  = (! \f''''''''_f''''''''_Int_Int_8_bufchan_buf [0]);
  assign \f''''''''_f''''''''_Int_Int_8_argbuf_d  = (\f''''''''_f''''''''_Int_Int_8_bufchan_buf [0] ? \f''''''''_f''''''''_Int_Int_8_bufchan_buf  :
                                                     \f''''''''_f''''''''_Int_Int_8_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''_f''''''''_Int_Int_8_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((\f''''''''_f''''''''_Int_Int_8_argbuf_r  && \f''''''''_f''''''''_Int_Int_8_bufchan_buf [0]))
        \f''''''''_f''''''''_Int_Int_8_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! \f''''''''_f''''''''_Int_Int_8_argbuf_r ) && (! \f''''''''_f''''''''_Int_Int_8_bufchan_buf [0])))
        \f''''''''_f''''''''_Int_Int_8_bufchan_buf  <= \f''''''''_f''''''''_Int_Int_8_bufchan_d ;
  
  /* dcon (Ty QTree_Int,
      Dcon QNode_Int) : [(f''''''''_f''''''''_Int_Int_8_argbuf,Pointer_QTree_Int),
                         (f''''''''_f''''''''_Int_Int_7_argbuf,Pointer_QTree_Int),
                         (f''''''''_f''''''''_Int_Int_6_argbuf,Pointer_QTree_Int),
                         (f''''''''_f''''''''_Int_Int_5_argbuf,Pointer_QTree_Int)] > (es_23_1es_24_1es_25_1es_26_1QNode_Int,QTree_Int) */
  assign es_23_1es_24_1es_25_1es_26_1QNode_Int_d = QNode_Int_dc((& {\f''''''''_f''''''''_Int_Int_8_argbuf_d [0],
                                                                    \f''''''''_f''''''''_Int_Int_7_argbuf_d [0],
                                                                    \f''''''''_f''''''''_Int_Int_6_argbuf_d [0],
                                                                    \f''''''''_f''''''''_Int_Int_5_argbuf_d [0]}), \f''''''''_f''''''''_Int_Int_8_argbuf_d , \f''''''''_f''''''''_Int_Int_7_argbuf_d , \f''''''''_f''''''''_Int_Int_6_argbuf_d , \f''''''''_f''''''''_Int_Int_5_argbuf_d );
  assign {\f''''''''_f''''''''_Int_Int_8_argbuf_r ,
          \f''''''''_f''''''''_Int_Int_7_argbuf_r ,
          \f''''''''_f''''''''_Int_Int_6_argbuf_r ,
          \f''''''''_f''''''''_Int_Int_5_argbuf_r } = {4 {(es_23_1es_24_1es_25_1es_26_1QNode_Int_r && es_23_1es_24_1es_25_1es_26_1QNode_Int_d[0])}};
  
  /* demux (Ty C8,
       Ty Pointer_QTree_Int) : (f''''''''_f''''''''_Int_Int_choice,C8) (lizzieLet39_4Lf''''''''_f''''''''_Int_Intsbos_1_merge_merge_fork_2,Pointer_QTree_Int) > [(f''''''''_f''''''''_Int_Int_1,Pointer_QTree_Int),
                                                                                                                                                                 (f''''''''_f''''''''_Int_Int_2,Pointer_QTree_Int),
                                                                                                                                                                 (f''''''''_f''''''''_Int_Int_3,Pointer_QTree_Int),
                                                                                                                                                                 (f''''''''_f''''''''_Int_Int_4,Pointer_QTree_Int),
                                                                                                                                                                 (f''''''''_f''''''''_Int_Int_5,Pointer_QTree_Int),
                                                                                                                                                                 (f''''''''_f''''''''_Int_Int_6,Pointer_QTree_Int),
                                                                                                                                                                 (f''''''''_f''''''''_Int_Int_7,Pointer_QTree_Int),
                                                                                                                                                                 (f''''''''_f''''''''_Int_Int_8,Pointer_QTree_Int)] */
  logic [7:0] \lizzieLet39_4Lf''''''''_f''''''''_Int_Intsbos_1_merge_merge_fork_2_onehotd ;
  always_comb
    if ((\f''''''''_f''''''''_Int_Int_choice_d [0] && \lizzieLet39_4Lf''''''''_f''''''''_Int_Intsbos_1_merge_merge_fork_2_d [0]))
      unique case (\f''''''''_f''''''''_Int_Int_choice_d [3:1])
        3'd0:
          \lizzieLet39_4Lf''''''''_f''''''''_Int_Intsbos_1_merge_merge_fork_2_onehotd  = 8'd1;
        3'd1:
          \lizzieLet39_4Lf''''''''_f''''''''_Int_Intsbos_1_merge_merge_fork_2_onehotd  = 8'd2;
        3'd2:
          \lizzieLet39_4Lf''''''''_f''''''''_Int_Intsbos_1_merge_merge_fork_2_onehotd  = 8'd4;
        3'd3:
          \lizzieLet39_4Lf''''''''_f''''''''_Int_Intsbos_1_merge_merge_fork_2_onehotd  = 8'd8;
        3'd4:
          \lizzieLet39_4Lf''''''''_f''''''''_Int_Intsbos_1_merge_merge_fork_2_onehotd  = 8'd16;
        3'd5:
          \lizzieLet39_4Lf''''''''_f''''''''_Int_Intsbos_1_merge_merge_fork_2_onehotd  = 8'd32;
        3'd6:
          \lizzieLet39_4Lf''''''''_f''''''''_Int_Intsbos_1_merge_merge_fork_2_onehotd  = 8'd64;
        3'd7:
          \lizzieLet39_4Lf''''''''_f''''''''_Int_Intsbos_1_merge_merge_fork_2_onehotd  = 8'd128;
        default:
          \lizzieLet39_4Lf''''''''_f''''''''_Int_Intsbos_1_merge_merge_fork_2_onehotd  = 8'd0;
      endcase
    else
      \lizzieLet39_4Lf''''''''_f''''''''_Int_Intsbos_1_merge_merge_fork_2_onehotd  = 8'd0;
  assign \f''''''''_f''''''''_Int_Int_1_d  = {\lizzieLet39_4Lf''''''''_f''''''''_Int_Intsbos_1_merge_merge_fork_2_d [16:1],
                                              \lizzieLet39_4Lf''''''''_f''''''''_Int_Intsbos_1_merge_merge_fork_2_onehotd [0]};
  assign \f''''''''_f''''''''_Int_Int_2_d  = {\lizzieLet39_4Lf''''''''_f''''''''_Int_Intsbos_1_merge_merge_fork_2_d [16:1],
                                              \lizzieLet39_4Lf''''''''_f''''''''_Int_Intsbos_1_merge_merge_fork_2_onehotd [1]};
  assign \f''''''''_f''''''''_Int_Int_3_d  = {\lizzieLet39_4Lf''''''''_f''''''''_Int_Intsbos_1_merge_merge_fork_2_d [16:1],
                                              \lizzieLet39_4Lf''''''''_f''''''''_Int_Intsbos_1_merge_merge_fork_2_onehotd [2]};
  assign \f''''''''_f''''''''_Int_Int_4_d  = {\lizzieLet39_4Lf''''''''_f''''''''_Int_Intsbos_1_merge_merge_fork_2_d [16:1],
                                              \lizzieLet39_4Lf''''''''_f''''''''_Int_Intsbos_1_merge_merge_fork_2_onehotd [3]};
  assign \f''''''''_f''''''''_Int_Int_5_d  = {\lizzieLet39_4Lf''''''''_f''''''''_Int_Intsbos_1_merge_merge_fork_2_d [16:1],
                                              \lizzieLet39_4Lf''''''''_f''''''''_Int_Intsbos_1_merge_merge_fork_2_onehotd [4]};
  assign \f''''''''_f''''''''_Int_Int_6_d  = {\lizzieLet39_4Lf''''''''_f''''''''_Int_Intsbos_1_merge_merge_fork_2_d [16:1],
                                              \lizzieLet39_4Lf''''''''_f''''''''_Int_Intsbos_1_merge_merge_fork_2_onehotd [5]};
  assign \f''''''''_f''''''''_Int_Int_7_d  = {\lizzieLet39_4Lf''''''''_f''''''''_Int_Intsbos_1_merge_merge_fork_2_d [16:1],
                                              \lizzieLet39_4Lf''''''''_f''''''''_Int_Intsbos_1_merge_merge_fork_2_onehotd [6]};
  assign \f''''''''_f''''''''_Int_Int_8_d  = {\lizzieLet39_4Lf''''''''_f''''''''_Int_Intsbos_1_merge_merge_fork_2_d [16:1],
                                              \lizzieLet39_4Lf''''''''_f''''''''_Int_Intsbos_1_merge_merge_fork_2_onehotd [7]};
  assign \lizzieLet39_4Lf''''''''_f''''''''_Int_Intsbos_1_merge_merge_fork_2_r  = (| (\lizzieLet39_4Lf''''''''_f''''''''_Int_Intsbos_1_merge_merge_fork_2_onehotd  & {\f''''''''_f''''''''_Int_Int_8_r ,
                                                                                                                                                                      \f''''''''_f''''''''_Int_Int_7_r ,
                                                                                                                                                                      \f''''''''_f''''''''_Int_Int_6_r ,
                                                                                                                                                                      \f''''''''_f''''''''_Int_Int_5_r ,
                                                                                                                                                                      \f''''''''_f''''''''_Int_Int_4_r ,
                                                                                                                                                                      \f''''''''_f''''''''_Int_Int_3_r ,
                                                                                                                                                                      \f''''''''_f''''''''_Int_Int_2_r ,
                                                                                                                                                                      \f''''''''_f''''''''_Int_Int_1_r }));
  assign \f''''''''_f''''''''_Int_Int_choice_r  = \lizzieLet39_4Lf''''''''_f''''''''_Int_Intsbos_1_merge_merge_fork_2_r ;
  
  /* destruct (Ty TupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int,
          Dcon TupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int) : (f''''''''_f''''''''_Int_Int_data,TupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int) > [(f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Intgo_13,Go),
                                                                                                                                                                      (f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Intq4a8u_1,Pointer_QTree_Int),
                                                                                                                                                                      (f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Intis_z_mapa8v_1,MyDTInt_Bool),
                                                                                                                                                                      (f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Intop_mapa8w_1,MyDTInt_Int)] */
  logic [3:0] \f''''''''_f''''''''_Int_Int_data_emitted ;
  logic [3:0] \f''''''''_f''''''''_Int_Int_data_done ;
  assign \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Intgo_13_d  = (\f''''''''_f''''''''_Int_Int_data_d [0] && (! \f''''''''_f''''''''_Int_Int_data_emitted [0]));
  assign \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Intq4a8u_1_d  = {\f''''''''_f''''''''_Int_Int_data_d [16:1],
                                                                                                         (\f''''''''_f''''''''_Int_Int_data_d [0] && (! \f''''''''_f''''''''_Int_Int_data_emitted [1]))};
  assign \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Intis_z_mapa8v_1_d  = (\f''''''''_f''''''''_Int_Int_data_d [0] && (! \f''''''''_f''''''''_Int_Int_data_emitted [2]));
  assign \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Intop_mapa8w_1_d  = (\f''''''''_f''''''''_Int_Int_data_d [0] && (! \f''''''''_f''''''''_Int_Int_data_emitted [3]));
  assign \f''''''''_f''''''''_Int_Int_data_done  = (\f''''''''_f''''''''_Int_Int_data_emitted  | ({\f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Intop_mapa8w_1_d [0],
                                                                                                   \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Intis_z_mapa8v_1_d [0],
                                                                                                   \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Intq4a8u_1_d [0],
                                                                                                   \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Intgo_13_d [0]} & {\f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Intop_mapa8w_1_r ,
                                                                                                                                                                                                     \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Intis_z_mapa8v_1_r ,
                                                                                                                                                                                                     \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Intq4a8u_1_r ,
                                                                                                                                                                                                     \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Intgo_13_r }));
  assign \f''''''''_f''''''''_Int_Int_data_r  = (& \f''''''''_f''''''''_Int_Int_data_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''_f''''''''_Int_Int_data_emitted  <= 4'd0;
    else
      \f''''''''_f''''''''_Int_Int_data_emitted  <= (\f''''''''_f''''''''_Int_Int_data_r  ? 4'd0 :
                                                     \f''''''''_f''''''''_Int_Int_data_done );
  
  /* destruct (Ty TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int,
          Dcon TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int) : (f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int_1,TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int) > [(f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intgo_14,Go),
                                                                                                                                                                                                                                                                                                                                                                        (f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intm1a8C_1,Pointer_QTree_Int),
                                                                                                                                                                                                                                                                                                                                                                        (f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intm2a8D_1,Pointer_QTree_Int),
                                                                                                                                                                                                                                                                                                                                                                        (f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intis_z_mapa8E_1,MyDTInt_Bool),
                                                                                                                                                                                                                                                                                                                                                                        (f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intop_mapa8F_1,MyDTInt_Int),
                                                                                                                                                                                                                                                                                                                                                                        (f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intis_z_adda8G_1,MyDTInt_Bool),
                                                                                                                                                                                                                                                                                                                                                                        (f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intop_adda8H_1,MyDTInt_Int_Int)] */
  logic [6:0] f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_emitted;
  logic [6:0] f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_done;
  assign f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intgo_14_d = (f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_d[0] && (! f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_emitted[0]));
  assign f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intm1a8C_1_d = {f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_d[16:1],
                                                                                                                                            (f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_d[0] && (! f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_emitted[1]))};
  assign f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intm2a8D_1_d = {f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_d[32:17],
                                                                                                                                            (f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_d[0] && (! f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_emitted[2]))};
  assign f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intis_z_mapa8E_1_d = (f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_d[0] && (! f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_emitted[3]));
  assign f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intop_mapa8F_1_d = (f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_d[0] && (! f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_emitted[4]));
  assign f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intis_z_adda8G_1_d = (f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_d[0] && (! f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_emitted[5]));
  assign f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intop_adda8H_1_d = (f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_d[0] && (! f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_emitted[6]));
  assign f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_done = (f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_emitted | ({f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intop_adda8H_1_d[0],
                                                                                                                                                                                                                                                                               f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intis_z_adda8G_1_d[0],
                                                                                                                                                                                                                                                                               f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intop_mapa8F_1_d[0],
                                                                                                                                                                                                                                                                               f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intis_z_mapa8E_1_d[0],
                                                                                                                                                                                                                                                                               f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intm2a8D_1_d[0],
                                                                                                                                                                                                                                                                               f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intm1a8C_1_d[0],
                                                                                                                                                                                                                                                                               f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intgo_14_d[0]} & {f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intop_adda8H_1_r,
                                                                                                                                                                                                                                                                                                                                                                                                                    f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intis_z_adda8G_1_r,
                                                                                                                                                                                                                                                                                                                                                                                                                    f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intop_mapa8F_1_r,
                                                                                                                                                                                                                                                                                                                                                                                                                    f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intis_z_mapa8E_1_r,
                                                                                                                                                                                                                                                                                                                                                                                                                    f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intm2a8D_1_r,
                                                                                                                                                                                                                                                                                                                                                                                                                    f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intm1a8C_1_r,
                                                                                                                                                                                                                                                                                                                                                                                                                    f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intgo_14_r}));
  assign f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_r = (& f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_emitted <= 7'd0;
    else
      f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_emitted <= (f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_r ? 7'd0 :
                                                                                                                                           f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_done);
  
  /* fork (Ty Go) : (f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intgo_14,Go) > [(go_14_1,Go),
                                                                                                                                                   (go_14_2,Go)] */
  logic [1:0] f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intgo_14_emitted;
  logic [1:0] f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intgo_14_done;
  assign go_14_1_d = (f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intgo_14_d[0] && (! f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intgo_14_emitted[0]));
  assign go_14_2_d = (f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intgo_14_d[0] && (! f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intgo_14_emitted[1]));
  assign f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intgo_14_done = (f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intgo_14_emitted | ({go_14_2_d[0],
                                                                                                                                                                                                                                                                                     go_14_1_d[0]} & {go_14_2_r,
                                                                                                                                                                                                                                                                                                      go_14_1_r}));
  assign f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intgo_14_r = (& f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intgo_14_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intgo_14_emitted <= 2'd0;
    else
      f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intgo_14_emitted <= (f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intgo_14_r ? 2'd0 :
                                                                                                                                              f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intgo_14_done);
  
  /* buf (Ty MyDTInt_Bool) : (f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intis_z_adda8G_1,MyDTInt_Bool) > (is_z_adda8G_1_1_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intis_z_adda8G_1_bufchan_d;
  logic f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intis_z_adda8G_1_bufchan_r;
  assign f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intis_z_adda8G_1_r = ((! f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intis_z_adda8G_1_bufchan_d[0]) || f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intis_z_adda8G_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intis_z_adda8G_1_bufchan_d <= 1'd0;
    else
      if (f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intis_z_adda8G_1_r)
        f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intis_z_adda8G_1_bufchan_d <= f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intis_z_adda8G_1_d;
  MyDTInt_Bool_t f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intis_z_adda8G_1_bufchan_buf;
  assign f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intis_z_adda8G_1_bufchan_r = (! f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intis_z_adda8G_1_bufchan_buf[0]);
  assign is_z_adda8G_1_1_argbuf_d = (f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intis_z_adda8G_1_bufchan_buf[0] ? f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intis_z_adda8G_1_bufchan_buf :
                                     f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intis_z_adda8G_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intis_z_adda8G_1_bufchan_buf <= 1'd0;
    else
      if ((is_z_adda8G_1_1_argbuf_r && f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intis_z_adda8G_1_bufchan_buf[0]))
        f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intis_z_adda8G_1_bufchan_buf <= 1'd0;
      else if (((! is_z_adda8G_1_1_argbuf_r) && (! f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intis_z_adda8G_1_bufchan_buf[0])))
        f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intis_z_adda8G_1_bufchan_buf <= f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intis_z_adda8G_1_bufchan_d;
  
  /* buf (Ty MyDTInt_Bool) : (f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intis_z_mapa8E_1,MyDTInt_Bool) > (is_z_mapa8E_1_1_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intis_z_mapa8E_1_bufchan_d;
  logic f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intis_z_mapa8E_1_bufchan_r;
  assign f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intis_z_mapa8E_1_r = ((! f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intis_z_mapa8E_1_bufchan_d[0]) || f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intis_z_mapa8E_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intis_z_mapa8E_1_bufchan_d <= 1'd0;
    else
      if (f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intis_z_mapa8E_1_r)
        f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intis_z_mapa8E_1_bufchan_d <= f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intis_z_mapa8E_1_d;
  MyDTInt_Bool_t f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intis_z_mapa8E_1_bufchan_buf;
  assign f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intis_z_mapa8E_1_bufchan_r = (! f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intis_z_mapa8E_1_bufchan_buf[0]);
  assign is_z_mapa8E_1_1_argbuf_d = (f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intis_z_mapa8E_1_bufchan_buf[0] ? f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intis_z_mapa8E_1_bufchan_buf :
                                     f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intis_z_mapa8E_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intis_z_mapa8E_1_bufchan_buf <= 1'd0;
    else
      if ((is_z_mapa8E_1_1_argbuf_r && f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intis_z_mapa8E_1_bufchan_buf[0]))
        f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intis_z_mapa8E_1_bufchan_buf <= 1'd0;
      else if (((! is_z_mapa8E_1_1_argbuf_r) && (! f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intis_z_mapa8E_1_bufchan_buf[0])))
        f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intis_z_mapa8E_1_bufchan_buf <= f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intis_z_mapa8E_1_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intm1a8C_1,Pointer_QTree_Int) > (m1a8C_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intm1a8C_1_bufchan_d;
  logic f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intm1a8C_1_bufchan_r;
  assign f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intm1a8C_1_r = ((! f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intm1a8C_1_bufchan_d[0]) || f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intm1a8C_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intm1a8C_1_bufchan_d <= {16'd0,
                                                                                                                                                  1'd0};
    else
      if (f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intm1a8C_1_r)
        f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intm1a8C_1_bufchan_d <= f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intm1a8C_1_d;
  Pointer_QTree_Int_t f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intm1a8C_1_bufchan_buf;
  assign f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intm1a8C_1_bufchan_r = (! f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intm1a8C_1_bufchan_buf[0]);
  assign m1a8C_1_1_argbuf_d = (f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intm1a8C_1_bufchan_buf[0] ? f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intm1a8C_1_bufchan_buf :
                               f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intm1a8C_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intm1a8C_1_bufchan_buf <= {16'd0,
                                                                                                                                                    1'd0};
    else
      if ((m1a8C_1_1_argbuf_r && f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intm1a8C_1_bufchan_buf[0]))
        f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intm1a8C_1_bufchan_buf <= {16'd0,
                                                                                                                                                      1'd0};
      else if (((! m1a8C_1_1_argbuf_r) && (! f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intm1a8C_1_bufchan_buf[0])))
        f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intm1a8C_1_bufchan_buf <= f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intm1a8C_1_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intm2a8D_1,Pointer_QTree_Int) > (m2a8D_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intm2a8D_1_bufchan_d;
  logic f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intm2a8D_1_bufchan_r;
  assign f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intm2a8D_1_r = ((! f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intm2a8D_1_bufchan_d[0]) || f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intm2a8D_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intm2a8D_1_bufchan_d <= {16'd0,
                                                                                                                                                  1'd0};
    else
      if (f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intm2a8D_1_r)
        f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intm2a8D_1_bufchan_d <= f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intm2a8D_1_d;
  Pointer_QTree_Int_t f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intm2a8D_1_bufchan_buf;
  assign f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intm2a8D_1_bufchan_r = (! f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intm2a8D_1_bufchan_buf[0]);
  assign m2a8D_1_1_argbuf_d = (f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intm2a8D_1_bufchan_buf[0] ? f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intm2a8D_1_bufchan_buf :
                               f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intm2a8D_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intm2a8D_1_bufchan_buf <= {16'd0,
                                                                                                                                                    1'd0};
    else
      if ((m2a8D_1_1_argbuf_r && f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intm2a8D_1_bufchan_buf[0]))
        f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intm2a8D_1_bufchan_buf <= {16'd0,
                                                                                                                                                      1'd0};
      else if (((! m2a8D_1_1_argbuf_r) && (! f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intm2a8D_1_bufchan_buf[0])))
        f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intm2a8D_1_bufchan_buf <= f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intm2a8D_1_bufchan_d;
  
  /* buf (Ty MyDTInt_Int_Int) : (f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intop_adda8H_1,MyDTInt_Int_Int) > (op_adda8H_1_1_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intop_adda8H_1_bufchan_d;
  logic f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intop_adda8H_1_bufchan_r;
  assign f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intop_adda8H_1_r = ((! f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intop_adda8H_1_bufchan_d[0]) || f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intop_adda8H_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intop_adda8H_1_bufchan_d <= 1'd0;
    else
      if (f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intop_adda8H_1_r)
        f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intop_adda8H_1_bufchan_d <= f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intop_adda8H_1_d;
  MyDTInt_Int_Int_t f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intop_adda8H_1_bufchan_buf;
  assign f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intop_adda8H_1_bufchan_r = (! f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intop_adda8H_1_bufchan_buf[0]);
  assign op_adda8H_1_1_argbuf_d = (f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intop_adda8H_1_bufchan_buf[0] ? f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intop_adda8H_1_bufchan_buf :
                                   f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intop_adda8H_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intop_adda8H_1_bufchan_buf <= 1'd0;
    else
      if ((op_adda8H_1_1_argbuf_r && f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intop_adda8H_1_bufchan_buf[0]))
        f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intop_adda8H_1_bufchan_buf <= 1'd0;
      else if (((! op_adda8H_1_1_argbuf_r) && (! f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intop_adda8H_1_bufchan_buf[0])))
        f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intop_adda8H_1_bufchan_buf <= f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intop_adda8H_1_bufchan_d;
  
  /* buf (Ty MyDTInt_Int) : (f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intop_mapa8F_1,MyDTInt_Int) > (op_mapa8F_1_1_argbuf,MyDTInt_Int) */
  MyDTInt_Int_t f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intop_mapa8F_1_bufchan_d;
  logic f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intop_mapa8F_1_bufchan_r;
  assign f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intop_mapa8F_1_r = ((! f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intop_mapa8F_1_bufchan_d[0]) || f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intop_mapa8F_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intop_mapa8F_1_bufchan_d <= 1'd0;
    else
      if (f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intop_mapa8F_1_r)
        f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intop_mapa8F_1_bufchan_d <= f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intop_mapa8F_1_d;
  MyDTInt_Int_t f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intop_mapa8F_1_bufchan_buf;
  assign f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intop_mapa8F_1_bufchan_r = (! f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intop_mapa8F_1_bufchan_buf[0]);
  assign op_mapa8F_1_1_argbuf_d = (f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intop_mapa8F_1_bufchan_buf[0] ? f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intop_mapa8F_1_bufchan_buf :
                                   f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intop_mapa8F_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intop_mapa8F_1_bufchan_buf <= 1'd0;
    else
      if ((op_mapa8F_1_1_argbuf_r && f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intop_mapa8F_1_bufchan_buf[0]))
        f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intop_mapa8F_1_bufchan_buf <= 1'd0;
      else if (((! op_mapa8F_1_1_argbuf_r) && (! f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intop_mapa8F_1_bufchan_buf[0])))
        f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intop_mapa8F_1_bufchan_buf <= f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Intop_mapa8F_1_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (f_f_Int_Int_resbuf,Pointer_QTree_Int) > (es_0_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t f_f_Int_Int_resbuf_bufchan_d;
  logic f_f_Int_Int_resbuf_bufchan_r;
  assign f_f_Int_Int_resbuf_r = ((! f_f_Int_Int_resbuf_bufchan_d[0]) || f_f_Int_Int_resbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) f_f_Int_Int_resbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (f_f_Int_Int_resbuf_r)
        f_f_Int_Int_resbuf_bufchan_d <= f_f_Int_Int_resbuf_d;
  Pointer_QTree_Int_t f_f_Int_Int_resbuf_bufchan_buf;
  assign f_f_Int_Int_resbuf_bufchan_r = (! f_f_Int_Int_resbuf_bufchan_buf[0]);
  assign es_0_1_argbuf_d = (f_f_Int_Int_resbuf_bufchan_buf[0] ? f_f_Int_Int_resbuf_bufchan_buf :
                            f_f_Int_Int_resbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      f_f_Int_Int_resbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((es_0_1_argbuf_r && f_f_Int_Int_resbuf_bufchan_buf[0]))
        f_f_Int_Int_resbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! es_0_1_argbuf_r) && (! f_f_Int_Int_resbuf_bufchan_buf[0])))
        f_f_Int_Int_resbuf_bufchan_buf <= f_f_Int_Int_resbuf_bufchan_d;
  
  /* dcon (Ty MyDTInt_Int_Int,
      Dcon Dcon_$fNumInt_$c+) : [(go_1,Go)] > (go_1Dcon_$fNumInt_$c+,MyDTInt_Int_Int) */
  assign \go_1Dcon_$fNumInt_$c+_d  = \Dcon_$fNumInt_$c+_dc ((& {go_1_d[0]}), go_1_d);
  assign {go_1_r} = {1 {(\go_1Dcon_$fNumInt_$c+_r  && \go_1Dcon_$fNumInt_$c+_d [0])}};
  
  /* fork (Ty C5) : (go_10_goMux_choice,C5) > [(go_10_goMux_choice_1,C5),
                                          (go_10_goMux_choice_2,C5)] */
  logic [1:0] go_10_goMux_choice_emitted;
  logic [1:0] go_10_goMux_choice_done;
  assign go_10_goMux_choice_1_d = {go_10_goMux_choice_d[3:1],
                                   (go_10_goMux_choice_d[0] && (! go_10_goMux_choice_emitted[0]))};
  assign go_10_goMux_choice_2_d = {go_10_goMux_choice_d[3:1],
                                   (go_10_goMux_choice_d[0] && (! go_10_goMux_choice_emitted[1]))};
  assign go_10_goMux_choice_done = (go_10_goMux_choice_emitted | ({go_10_goMux_choice_2_d[0],
                                                                   go_10_goMux_choice_1_d[0]} & {go_10_goMux_choice_2_r,
                                                                                                 go_10_goMux_choice_1_r}));
  assign go_10_goMux_choice_r = (& go_10_goMux_choice_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_10_goMux_choice_emitted <= 2'd0;
    else
      go_10_goMux_choice_emitted <= (go_10_goMux_choice_r ? 2'd0 :
                                     go_10_goMux_choice_done);
  
  /* mux (Ty C5,
     Ty Pointer_QTree_Int) : (go_10_goMux_choice_1,C5) [(call_$wnnz_goMux2,Pointer_QTree_Int),
                                                        (q2a85_1_1_argbuf,Pointer_QTree_Int),
                                                        (q3a86_2_1_argbuf,Pointer_QTree_Int),
                                                        (q4a87_3_1_argbuf,Pointer_QTree_Int),
                                                        (q1a84_1_argbuf,Pointer_QTree_Int)] > (wsiX_1_goMux_mux,Pointer_QTree_Int) */
  logic [16:0] wsiX_1_goMux_mux_mux;
  logic [4:0] wsiX_1_goMux_mux_onehot;
  always_comb
    unique case (go_10_goMux_choice_1_d[3:1])
      3'd0:
        {wsiX_1_goMux_mux_onehot, wsiX_1_goMux_mux_mux} = {5'd1,
                                                           call_$wnnz_goMux2_d};
      3'd1:
        {wsiX_1_goMux_mux_onehot, wsiX_1_goMux_mux_mux} = {5'd2,
                                                           q2a85_1_1_argbuf_d};
      3'd2:
        {wsiX_1_goMux_mux_onehot, wsiX_1_goMux_mux_mux} = {5'd4,
                                                           q3a86_2_1_argbuf_d};
      3'd3:
        {wsiX_1_goMux_mux_onehot, wsiX_1_goMux_mux_mux} = {5'd8,
                                                           q4a87_3_1_argbuf_d};
      3'd4:
        {wsiX_1_goMux_mux_onehot, wsiX_1_goMux_mux_mux} = {5'd16,
                                                           q1a84_1_argbuf_d};
      default:
        {wsiX_1_goMux_mux_onehot, wsiX_1_goMux_mux_mux} = {5'd0,
                                                           {16'd0, 1'd0}};
    endcase
  assign wsiX_1_goMux_mux_d = {wsiX_1_goMux_mux_mux[16:1],
                               (wsiX_1_goMux_mux_mux[0] && go_10_goMux_choice_1_d[0])};
  assign go_10_goMux_choice_1_r = (wsiX_1_goMux_mux_d[0] && wsiX_1_goMux_mux_r);
  assign {q1a84_1_argbuf_r,
          q4a87_3_1_argbuf_r,
          q3a86_2_1_argbuf_r,
          q2a85_1_1_argbuf_r,
          call_$wnnz_goMux2_r} = (go_10_goMux_choice_1_r ? wsiX_1_goMux_mux_onehot :
                                  5'd0);
  
  /* mux (Ty C5,
     Ty Pointer_CT$wnnz) : (go_10_goMux_choice_2,C5) [(call_$wnnz_goMux3,Pointer_CT$wnnz),
                                                      (sca2_1_argbuf,Pointer_CT$wnnz),
                                                      (sca1_1_argbuf,Pointer_CT$wnnz),
                                                      (sca0_1_argbuf,Pointer_CT$wnnz),
                                                      (sca3_1_argbuf,Pointer_CT$wnnz)] > (sc_0_goMux_mux,Pointer_CT$wnnz) */
  logic [16:0] sc_0_goMux_mux_mux;
  logic [4:0] sc_0_goMux_mux_onehot;
  always_comb
    unique case (go_10_goMux_choice_2_d[3:1])
      3'd0:
        {sc_0_goMux_mux_onehot, sc_0_goMux_mux_mux} = {5'd1,
                                                       call_$wnnz_goMux3_d};
      3'd1:
        {sc_0_goMux_mux_onehot, sc_0_goMux_mux_mux} = {5'd2,
                                                       sca2_1_argbuf_d};
      3'd2:
        {sc_0_goMux_mux_onehot, sc_0_goMux_mux_mux} = {5'd4,
                                                       sca1_1_argbuf_d};
      3'd3:
        {sc_0_goMux_mux_onehot, sc_0_goMux_mux_mux} = {5'd8,
                                                       sca0_1_argbuf_d};
      3'd4:
        {sc_0_goMux_mux_onehot, sc_0_goMux_mux_mux} = {5'd16,
                                                       sca3_1_argbuf_d};
      default:
        {sc_0_goMux_mux_onehot, sc_0_goMux_mux_mux} = {5'd0,
                                                       {16'd0, 1'd0}};
    endcase
  assign sc_0_goMux_mux_d = {sc_0_goMux_mux_mux[16:1],
                             (sc_0_goMux_mux_mux[0] && go_10_goMux_choice_2_d[0])};
  assign go_10_goMux_choice_2_r = (sc_0_goMux_mux_d[0] && sc_0_goMux_mux_r);
  assign {sca3_1_argbuf_r,
          sca0_1_argbuf_r,
          sca1_1_argbuf_r,
          sca2_1_argbuf_r,
          call_$wnnz_goMux3_r} = (go_10_goMux_choice_2_r ? sc_0_goMux_mux_onehot :
                                  5'd0);
  
  /* fork (Ty C5) : (go_11_goMux_choice,C5) > [(go_11_goMux_choice_1,C5),
                                          (go_11_goMux_choice_2,C5),
                                          (go_11_goMux_choice_3,C5),
                                          (go_11_goMux_choice_4,C5)] */
  logic [3:0] go_11_goMux_choice_emitted;
  logic [3:0] go_11_goMux_choice_done;
  assign go_11_goMux_choice_1_d = {go_11_goMux_choice_d[3:1],
                                   (go_11_goMux_choice_d[0] && (! go_11_goMux_choice_emitted[0]))};
  assign go_11_goMux_choice_2_d = {go_11_goMux_choice_d[3:1],
                                   (go_11_goMux_choice_d[0] && (! go_11_goMux_choice_emitted[1]))};
  assign go_11_goMux_choice_3_d = {go_11_goMux_choice_d[3:1],
                                   (go_11_goMux_choice_d[0] && (! go_11_goMux_choice_emitted[2]))};
  assign go_11_goMux_choice_4_d = {go_11_goMux_choice_d[3:1],
                                   (go_11_goMux_choice_d[0] && (! go_11_goMux_choice_emitted[3]))};
  assign go_11_goMux_choice_done = (go_11_goMux_choice_emitted | ({go_11_goMux_choice_4_d[0],
                                                                   go_11_goMux_choice_3_d[0],
                                                                   go_11_goMux_choice_2_d[0],
                                                                   go_11_goMux_choice_1_d[0]} & {go_11_goMux_choice_4_r,
                                                                                                 go_11_goMux_choice_3_r,
                                                                                                 go_11_goMux_choice_2_r,
                                                                                                 go_11_goMux_choice_1_r}));
  assign go_11_goMux_choice_r = (& go_11_goMux_choice_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_11_goMux_choice_emitted <= 4'd0;
    else
      go_11_goMux_choice_emitted <= (go_11_goMux_choice_r ? 4'd0 :
                                     go_11_goMux_choice_done);
  
  /* mux (Ty C5,
     Ty Pointer_QTree_Int) : (go_11_goMux_choice_1,C5) [(call_f''''''''_f''''''''_Int_Int_goMux2,Pointer_QTree_Int),
                                                        (bla8A_1_1_argbuf,Pointer_QTree_Int),
                                                        (tra8z_2_1_argbuf,Pointer_QTree_Int),
                                                        (tla8y_3_1_argbuf,Pointer_QTree_Int),
                                                        (bra8B_1_argbuf,Pointer_QTree_Int)] > (q4a8u_goMux_mux,Pointer_QTree_Int) */
  logic [16:0] q4a8u_goMux_mux_mux;
  logic [4:0] q4a8u_goMux_mux_onehot;
  always_comb
    unique case (go_11_goMux_choice_1_d[3:1])
      3'd0:
        {q4a8u_goMux_mux_onehot, q4a8u_goMux_mux_mux} = {5'd1,
                                                         \call_f''''''''_f''''''''_Int_Int_goMux2_d };
      3'd1:
        {q4a8u_goMux_mux_onehot, q4a8u_goMux_mux_mux} = {5'd2,
                                                         bla8A_1_1_argbuf_d};
      3'd2:
        {q4a8u_goMux_mux_onehot, q4a8u_goMux_mux_mux} = {5'd4,
                                                         tra8z_2_1_argbuf_d};
      3'd3:
        {q4a8u_goMux_mux_onehot, q4a8u_goMux_mux_mux} = {5'd8,
                                                         tla8y_3_1_argbuf_d};
      3'd4:
        {q4a8u_goMux_mux_onehot, q4a8u_goMux_mux_mux} = {5'd16,
                                                         bra8B_1_argbuf_d};
      default:
        {q4a8u_goMux_mux_onehot, q4a8u_goMux_mux_mux} = {5'd0,
                                                         {16'd0, 1'd0}};
    endcase
  assign q4a8u_goMux_mux_d = {q4a8u_goMux_mux_mux[16:1],
                              (q4a8u_goMux_mux_mux[0] && go_11_goMux_choice_1_d[0])};
  assign go_11_goMux_choice_1_r = (q4a8u_goMux_mux_d[0] && q4a8u_goMux_mux_r);
  assign {bra8B_1_argbuf_r,
          tla8y_3_1_argbuf_r,
          tra8z_2_1_argbuf_r,
          bla8A_1_1_argbuf_r,
          \call_f''''''''_f''''''''_Int_Int_goMux2_r } = (go_11_goMux_choice_1_r ? q4a8u_goMux_mux_onehot :
                                                          5'd0);
  
  /* mux (Ty C5,
     Ty MyDTInt_Bool) : (go_11_goMux_choice_2,C5) [(call_f''''''''_f''''''''_Int_Int_goMux3,MyDTInt_Bool),
                                                   (is_z_mapa8v_2_2_argbuf,MyDTInt_Bool),
                                                   (is_z_mapa8v_3_2_argbuf,MyDTInt_Bool),
                                                   (is_z_mapa8v_4_1_argbuf,MyDTInt_Bool),
                                                   (lizzieLet6_4QNode_Int_2_argbuf,MyDTInt_Bool)] > (is_z_mapa8v_goMux_mux,MyDTInt_Bool) */
  logic [0:0] is_z_mapa8v_goMux_mux_mux;
  logic [4:0] is_z_mapa8v_goMux_mux_onehot;
  always_comb
    unique case (go_11_goMux_choice_2_d[3:1])
      3'd0:
        {is_z_mapa8v_goMux_mux_onehot, is_z_mapa8v_goMux_mux_mux} = {5'd1,
                                                                     \call_f''''''''_f''''''''_Int_Int_goMux3_d };
      3'd1:
        {is_z_mapa8v_goMux_mux_onehot, is_z_mapa8v_goMux_mux_mux} = {5'd2,
                                                                     is_z_mapa8v_2_2_argbuf_d};
      3'd2:
        {is_z_mapa8v_goMux_mux_onehot, is_z_mapa8v_goMux_mux_mux} = {5'd4,
                                                                     is_z_mapa8v_3_2_argbuf_d};
      3'd3:
        {is_z_mapa8v_goMux_mux_onehot, is_z_mapa8v_goMux_mux_mux} = {5'd8,
                                                                     is_z_mapa8v_4_1_argbuf_d};
      3'd4:
        {is_z_mapa8v_goMux_mux_onehot, is_z_mapa8v_goMux_mux_mux} = {5'd16,
                                                                     lizzieLet6_4QNode_Int_2_argbuf_d};
      default:
        {is_z_mapa8v_goMux_mux_onehot, is_z_mapa8v_goMux_mux_mux} = {5'd0,
                                                                     1'd0};
    endcase
  assign is_z_mapa8v_goMux_mux_d = (is_z_mapa8v_goMux_mux_mux[0] && go_11_goMux_choice_2_d[0]);
  assign go_11_goMux_choice_2_r = (is_z_mapa8v_goMux_mux_d[0] && is_z_mapa8v_goMux_mux_r);
  assign {lizzieLet6_4QNode_Int_2_argbuf_r,
          is_z_mapa8v_4_1_argbuf_r,
          is_z_mapa8v_3_2_argbuf_r,
          is_z_mapa8v_2_2_argbuf_r,
          \call_f''''''''_f''''''''_Int_Int_goMux3_r } = (go_11_goMux_choice_2_r ? is_z_mapa8v_goMux_mux_onehot :
                                                          5'd0);
  
  /* mux (Ty C5,
     Ty MyDTInt_Int) : (go_11_goMux_choice_3,C5) [(call_f''''''''_f''''''''_Int_Int_goMux4,MyDTInt_Int),
                                                  (op_mapa8w_2_2_argbuf,MyDTInt_Int),
                                                  (op_mapa8w_3_2_argbuf,MyDTInt_Int),
                                                  (op_mapa8w_4_1_argbuf,MyDTInt_Int),
                                                  (lizzieLet6_5QNode_Int_2_argbuf,MyDTInt_Int)] > (op_mapa8w_goMux_mux,MyDTInt_Int) */
  logic [0:0] op_mapa8w_goMux_mux_mux;
  logic [4:0] op_mapa8w_goMux_mux_onehot;
  always_comb
    unique case (go_11_goMux_choice_3_d[3:1])
      3'd0:
        {op_mapa8w_goMux_mux_onehot, op_mapa8w_goMux_mux_mux} = {5'd1,
                                                                 \call_f''''''''_f''''''''_Int_Int_goMux4_d };
      3'd1:
        {op_mapa8w_goMux_mux_onehot, op_mapa8w_goMux_mux_mux} = {5'd2,
                                                                 op_mapa8w_2_2_argbuf_d};
      3'd2:
        {op_mapa8w_goMux_mux_onehot, op_mapa8w_goMux_mux_mux} = {5'd4,
                                                                 op_mapa8w_3_2_argbuf_d};
      3'd3:
        {op_mapa8w_goMux_mux_onehot, op_mapa8w_goMux_mux_mux} = {5'd8,
                                                                 op_mapa8w_4_1_argbuf_d};
      3'd4:
        {op_mapa8w_goMux_mux_onehot, op_mapa8w_goMux_mux_mux} = {5'd16,
                                                                 lizzieLet6_5QNode_Int_2_argbuf_d};
      default:
        {op_mapa8w_goMux_mux_onehot, op_mapa8w_goMux_mux_mux} = {5'd0,
                                                                 1'd0};
    endcase
  assign op_mapa8w_goMux_mux_d = (op_mapa8w_goMux_mux_mux[0] && go_11_goMux_choice_3_d[0]);
  assign go_11_goMux_choice_3_r = (op_mapa8w_goMux_mux_d[0] && op_mapa8w_goMux_mux_r);
  assign {lizzieLet6_5QNode_Int_2_argbuf_r,
          op_mapa8w_4_1_argbuf_r,
          op_mapa8w_3_2_argbuf_r,
          op_mapa8w_2_2_argbuf_r,
          \call_f''''''''_f''''''''_Int_Int_goMux4_r } = (go_11_goMux_choice_3_r ? op_mapa8w_goMux_mux_onehot :
                                                          5'd0);
  
  /* mux (Ty C5,
     Ty Pointer_CTf''''''''_f''''''''_Int_Int) : (go_11_goMux_choice_4,C5) [(call_f''''''''_f''''''''_Int_Int_goMux5,Pointer_CTf''''''''_f''''''''_Int_Int),
                                                                            (sca2_1_1_argbuf,Pointer_CTf''''''''_f''''''''_Int_Int),
                                                                            (sca1_1_1_argbuf,Pointer_CTf''''''''_f''''''''_Int_Int),
                                                                            (sca0_1_1_argbuf,Pointer_CTf''''''''_f''''''''_Int_Int),
                                                                            (sca3_1_1_argbuf,Pointer_CTf''''''''_f''''''''_Int_Int)] > (sc_0_1_goMux_mux,Pointer_CTf''''''''_f''''''''_Int_Int) */
  logic [16:0] sc_0_1_goMux_mux_mux;
  logic [4:0] sc_0_1_goMux_mux_onehot;
  always_comb
    unique case (go_11_goMux_choice_4_d[3:1])
      3'd0:
        {sc_0_1_goMux_mux_onehot, sc_0_1_goMux_mux_mux} = {5'd1,
                                                           \call_f''''''''_f''''''''_Int_Int_goMux5_d };
      3'd1:
        {sc_0_1_goMux_mux_onehot, sc_0_1_goMux_mux_mux} = {5'd2,
                                                           sca2_1_1_argbuf_d};
      3'd2:
        {sc_0_1_goMux_mux_onehot, sc_0_1_goMux_mux_mux} = {5'd4,
                                                           sca1_1_1_argbuf_d};
      3'd3:
        {sc_0_1_goMux_mux_onehot, sc_0_1_goMux_mux_mux} = {5'd8,
                                                           sca0_1_1_argbuf_d};
      3'd4:
        {sc_0_1_goMux_mux_onehot, sc_0_1_goMux_mux_mux} = {5'd16,
                                                           sca3_1_1_argbuf_d};
      default:
        {sc_0_1_goMux_mux_onehot, sc_0_1_goMux_mux_mux} = {5'd0,
                                                           {16'd0, 1'd0}};
    endcase
  assign sc_0_1_goMux_mux_d = {sc_0_1_goMux_mux_mux[16:1],
                               (sc_0_1_goMux_mux_mux[0] && go_11_goMux_choice_4_d[0])};
  assign go_11_goMux_choice_4_r = (sc_0_1_goMux_mux_d[0] && sc_0_1_goMux_mux_r);
  assign {sca3_1_1_argbuf_r,
          sca0_1_1_argbuf_r,
          sca1_1_1_argbuf_r,
          sca2_1_1_argbuf_r,
          \call_f''''''''_f''''''''_Int_Int_goMux5_r } = (go_11_goMux_choice_4_r ? sc_0_1_goMux_mux_onehot :
                                                          5'd0);
  
  /* fork (Ty C5) : (go_12_goMux_choice,C5) > [(go_12_goMux_choice_1,C5),
                                          (go_12_goMux_choice_2,C5),
                                          (go_12_goMux_choice_3,C5),
                                          (go_12_goMux_choice_4,C5),
                                          (go_12_goMux_choice_5,C5),
                                          (go_12_goMux_choice_6,C5),
                                          (go_12_goMux_choice_7,C5)] */
  logic [6:0] go_12_goMux_choice_emitted;
  logic [6:0] go_12_goMux_choice_done;
  assign go_12_goMux_choice_1_d = {go_12_goMux_choice_d[3:1],
                                   (go_12_goMux_choice_d[0] && (! go_12_goMux_choice_emitted[0]))};
  assign go_12_goMux_choice_2_d = {go_12_goMux_choice_d[3:1],
                                   (go_12_goMux_choice_d[0] && (! go_12_goMux_choice_emitted[1]))};
  assign go_12_goMux_choice_3_d = {go_12_goMux_choice_d[3:1],
                                   (go_12_goMux_choice_d[0] && (! go_12_goMux_choice_emitted[2]))};
  assign go_12_goMux_choice_4_d = {go_12_goMux_choice_d[3:1],
                                   (go_12_goMux_choice_d[0] && (! go_12_goMux_choice_emitted[3]))};
  assign go_12_goMux_choice_5_d = {go_12_goMux_choice_d[3:1],
                                   (go_12_goMux_choice_d[0] && (! go_12_goMux_choice_emitted[4]))};
  assign go_12_goMux_choice_6_d = {go_12_goMux_choice_d[3:1],
                                   (go_12_goMux_choice_d[0] && (! go_12_goMux_choice_emitted[5]))};
  assign go_12_goMux_choice_7_d = {go_12_goMux_choice_d[3:1],
                                   (go_12_goMux_choice_d[0] && (! go_12_goMux_choice_emitted[6]))};
  assign go_12_goMux_choice_done = (go_12_goMux_choice_emitted | ({go_12_goMux_choice_7_d[0],
                                                                   go_12_goMux_choice_6_d[0],
                                                                   go_12_goMux_choice_5_d[0],
                                                                   go_12_goMux_choice_4_d[0],
                                                                   go_12_goMux_choice_3_d[0],
                                                                   go_12_goMux_choice_2_d[0],
                                                                   go_12_goMux_choice_1_d[0]} & {go_12_goMux_choice_7_r,
                                                                                                 go_12_goMux_choice_6_r,
                                                                                                 go_12_goMux_choice_5_r,
                                                                                                 go_12_goMux_choice_4_r,
                                                                                                 go_12_goMux_choice_3_r,
                                                                                                 go_12_goMux_choice_2_r,
                                                                                                 go_12_goMux_choice_1_r}));
  assign go_12_goMux_choice_r = (& go_12_goMux_choice_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_12_goMux_choice_emitted <= 7'd0;
    else
      go_12_goMux_choice_emitted <= (go_12_goMux_choice_r ? 7'd0 :
                                     go_12_goMux_choice_done);
  
  /* mux (Ty C5,
     Ty Pointer_QTree_Int) : (go_12_goMux_choice_1,C5) [(call_f_f_Int_Int_goMux2,Pointer_QTree_Int),
                                                        (q3a8V_1_1_argbuf,Pointer_QTree_Int),
                                                        (q2a8U_2_1_argbuf,Pointer_QTree_Int),
                                                        (q1a8T_3_1_argbuf,Pointer_QTree_Int),
                                                        (lizzieLet12_6QNode_Int_12QNode_Int_1_argbuf,Pointer_QTree_Int)] > (m1a8C_goMux_mux,Pointer_QTree_Int) */
  logic [16:0] m1a8C_goMux_mux_mux;
  logic [4:0] m1a8C_goMux_mux_onehot;
  always_comb
    unique case (go_12_goMux_choice_1_d[3:1])
      3'd0:
        {m1a8C_goMux_mux_onehot, m1a8C_goMux_mux_mux} = {5'd1,
                                                         call_f_f_Int_Int_goMux2_d};
      3'd1:
        {m1a8C_goMux_mux_onehot, m1a8C_goMux_mux_mux} = {5'd2,
                                                         q3a8V_1_1_argbuf_d};
      3'd2:
        {m1a8C_goMux_mux_onehot, m1a8C_goMux_mux_mux} = {5'd4,
                                                         q2a8U_2_1_argbuf_d};
      3'd3:
        {m1a8C_goMux_mux_onehot, m1a8C_goMux_mux_mux} = {5'd8,
                                                         q1a8T_3_1_argbuf_d};
      3'd4:
        {m1a8C_goMux_mux_onehot, m1a8C_goMux_mux_mux} = {5'd16,
                                                         lizzieLet12_6QNode_Int_12QNode_Int_1_argbuf_d};
      default:
        {m1a8C_goMux_mux_onehot, m1a8C_goMux_mux_mux} = {5'd0,
                                                         {16'd0, 1'd0}};
    endcase
  assign m1a8C_goMux_mux_d = {m1a8C_goMux_mux_mux[16:1],
                              (m1a8C_goMux_mux_mux[0] && go_12_goMux_choice_1_d[0])};
  assign go_12_goMux_choice_1_r = (m1a8C_goMux_mux_d[0] && m1a8C_goMux_mux_r);
  assign {lizzieLet12_6QNode_Int_12QNode_Int_1_argbuf_r,
          q1a8T_3_1_argbuf_r,
          q2a8U_2_1_argbuf_r,
          q3a8V_1_1_argbuf_r,
          call_f_f_Int_Int_goMux2_r} = (go_12_goMux_choice_1_r ? m1a8C_goMux_mux_onehot :
                                        5'd0);
  
  /* mux (Ty C5,
     Ty Pointer_QTree_Int) : (go_12_goMux_choice_2,C5) [(call_f_f_Int_Int_goMux3,Pointer_QTree_Int),
                                                        (t3a90_1_1_argbuf,Pointer_QTree_Int),
                                                        (t2a8Z_2_1_argbuf,Pointer_QTree_Int),
                                                        (t1a8Y_3_1_argbuf,Pointer_QTree_Int),
                                                        (t4a91_1_argbuf,Pointer_QTree_Int)] > (m2a8D_goMux_mux,Pointer_QTree_Int) */
  logic [16:0] m2a8D_goMux_mux_mux;
  logic [4:0] m2a8D_goMux_mux_onehot;
  always_comb
    unique case (go_12_goMux_choice_2_d[3:1])
      3'd0:
        {m2a8D_goMux_mux_onehot, m2a8D_goMux_mux_mux} = {5'd1,
                                                         call_f_f_Int_Int_goMux3_d};
      3'd1:
        {m2a8D_goMux_mux_onehot, m2a8D_goMux_mux_mux} = {5'd2,
                                                         t3a90_1_1_argbuf_d};
      3'd2:
        {m2a8D_goMux_mux_onehot, m2a8D_goMux_mux_mux} = {5'd4,
                                                         t2a8Z_2_1_argbuf_d};
      3'd3:
        {m2a8D_goMux_mux_onehot, m2a8D_goMux_mux_mux} = {5'd8,
                                                         t1a8Y_3_1_argbuf_d};
      3'd4:
        {m2a8D_goMux_mux_onehot, m2a8D_goMux_mux_mux} = {5'd16,
                                                         t4a91_1_argbuf_d};
      default:
        {m2a8D_goMux_mux_onehot, m2a8D_goMux_mux_mux} = {5'd0,
                                                         {16'd0, 1'd0}};
    endcase
  assign m2a8D_goMux_mux_d = {m2a8D_goMux_mux_mux[16:1],
                              (m2a8D_goMux_mux_mux[0] && go_12_goMux_choice_2_d[0])};
  assign go_12_goMux_choice_2_r = (m2a8D_goMux_mux_d[0] && m2a8D_goMux_mux_r);
  assign {t4a91_1_argbuf_r,
          t1a8Y_3_1_argbuf_r,
          t2a8Z_2_1_argbuf_r,
          t3a90_1_1_argbuf_r,
          call_f_f_Int_Int_goMux3_r} = (go_12_goMux_choice_2_r ? m2a8D_goMux_mux_onehot :
                                        5'd0);
  
  /* mux (Ty C5,
     Ty MyDTInt_Bool) : (go_12_goMux_choice_3,C5) [(call_f_f_Int_Int_goMux4,MyDTInt_Bool),
                                                   (is_z_mapa8E_2_2_argbuf,MyDTInt_Bool),
                                                   (is_z_mapa8E_3_2_argbuf,MyDTInt_Bool),
                                                   (is_z_mapa8E_4_1_argbuf,MyDTInt_Bool),
                                                   (lizzieLet12_6QNode_Int_5QNode_Int_2_argbuf,MyDTInt_Bool)] > (is_z_mapa8E_goMux_mux,MyDTInt_Bool) */
  logic [0:0] is_z_mapa8E_goMux_mux_mux;
  logic [4:0] is_z_mapa8E_goMux_mux_onehot;
  always_comb
    unique case (go_12_goMux_choice_3_d[3:1])
      3'd0:
        {is_z_mapa8E_goMux_mux_onehot, is_z_mapa8E_goMux_mux_mux} = {5'd1,
                                                                     call_f_f_Int_Int_goMux4_d};
      3'd1:
        {is_z_mapa8E_goMux_mux_onehot, is_z_mapa8E_goMux_mux_mux} = {5'd2,
                                                                     is_z_mapa8E_2_2_argbuf_d};
      3'd2:
        {is_z_mapa8E_goMux_mux_onehot, is_z_mapa8E_goMux_mux_mux} = {5'd4,
                                                                     is_z_mapa8E_3_2_argbuf_d};
      3'd3:
        {is_z_mapa8E_goMux_mux_onehot, is_z_mapa8E_goMux_mux_mux} = {5'd8,
                                                                     is_z_mapa8E_4_1_argbuf_d};
      3'd4:
        {is_z_mapa8E_goMux_mux_onehot, is_z_mapa8E_goMux_mux_mux} = {5'd16,
                                                                     lizzieLet12_6QNode_Int_5QNode_Int_2_argbuf_d};
      default:
        {is_z_mapa8E_goMux_mux_onehot, is_z_mapa8E_goMux_mux_mux} = {5'd0,
                                                                     1'd0};
    endcase
  assign is_z_mapa8E_goMux_mux_d = (is_z_mapa8E_goMux_mux_mux[0] && go_12_goMux_choice_3_d[0]);
  assign go_12_goMux_choice_3_r = (is_z_mapa8E_goMux_mux_d[0] && is_z_mapa8E_goMux_mux_r);
  assign {lizzieLet12_6QNode_Int_5QNode_Int_2_argbuf_r,
          is_z_mapa8E_4_1_argbuf_r,
          is_z_mapa8E_3_2_argbuf_r,
          is_z_mapa8E_2_2_argbuf_r,
          call_f_f_Int_Int_goMux4_r} = (go_12_goMux_choice_3_r ? is_z_mapa8E_goMux_mux_onehot :
                                        5'd0);
  
  /* mux (Ty C5,
     Ty MyDTInt_Int) : (go_12_goMux_choice_4,C5) [(call_f_f_Int_Int_goMux5,MyDTInt_Int),
                                                  (op_mapa8F_2_2_argbuf,MyDTInt_Int),
                                                  (op_mapa8F_3_2_argbuf,MyDTInt_Int),
                                                  (op_mapa8F_4_1_argbuf,MyDTInt_Int),
                                                  (lizzieLet12_6QNode_Int_7QNode_Int_2_argbuf,MyDTInt_Int)] > (op_mapa8F_goMux_mux,MyDTInt_Int) */
  logic [0:0] op_mapa8F_goMux_mux_mux;
  logic [4:0] op_mapa8F_goMux_mux_onehot;
  always_comb
    unique case (go_12_goMux_choice_4_d[3:1])
      3'd0:
        {op_mapa8F_goMux_mux_onehot, op_mapa8F_goMux_mux_mux} = {5'd1,
                                                                 call_f_f_Int_Int_goMux5_d};
      3'd1:
        {op_mapa8F_goMux_mux_onehot, op_mapa8F_goMux_mux_mux} = {5'd2,
                                                                 op_mapa8F_2_2_argbuf_d};
      3'd2:
        {op_mapa8F_goMux_mux_onehot, op_mapa8F_goMux_mux_mux} = {5'd4,
                                                                 op_mapa8F_3_2_argbuf_d};
      3'd3:
        {op_mapa8F_goMux_mux_onehot, op_mapa8F_goMux_mux_mux} = {5'd8,
                                                                 op_mapa8F_4_1_argbuf_d};
      3'd4:
        {op_mapa8F_goMux_mux_onehot, op_mapa8F_goMux_mux_mux} = {5'd16,
                                                                 lizzieLet12_6QNode_Int_7QNode_Int_2_argbuf_d};
      default:
        {op_mapa8F_goMux_mux_onehot, op_mapa8F_goMux_mux_mux} = {5'd0,
                                                                 1'd0};
    endcase
  assign op_mapa8F_goMux_mux_d = (op_mapa8F_goMux_mux_mux[0] && go_12_goMux_choice_4_d[0]);
  assign go_12_goMux_choice_4_r = (op_mapa8F_goMux_mux_d[0] && op_mapa8F_goMux_mux_r);
  assign {lizzieLet12_6QNode_Int_7QNode_Int_2_argbuf_r,
          op_mapa8F_4_1_argbuf_r,
          op_mapa8F_3_2_argbuf_r,
          op_mapa8F_2_2_argbuf_r,
          call_f_f_Int_Int_goMux5_r} = (go_12_goMux_choice_4_r ? op_mapa8F_goMux_mux_onehot :
                                        5'd0);
  
  /* mux (Ty C5,
     Ty MyDTInt_Bool) : (go_12_goMux_choice_5,C5) [(call_f_f_Int_Int_goMux6,MyDTInt_Bool),
                                                   (is_z_adda8G_2_2_argbuf,MyDTInt_Bool),
                                                   (is_z_adda8G_3_2_argbuf,MyDTInt_Bool),
                                                   (is_z_adda8G_4_1_argbuf,MyDTInt_Bool),
                                                   (lizzieLet12_6QNode_Int_4QNode_Int_2_argbuf,MyDTInt_Bool)] > (is_z_adda8G_goMux_mux,MyDTInt_Bool) */
  logic [0:0] is_z_adda8G_goMux_mux_mux;
  logic [4:0] is_z_adda8G_goMux_mux_onehot;
  always_comb
    unique case (go_12_goMux_choice_5_d[3:1])
      3'd0:
        {is_z_adda8G_goMux_mux_onehot, is_z_adda8G_goMux_mux_mux} = {5'd1,
                                                                     call_f_f_Int_Int_goMux6_d};
      3'd1:
        {is_z_adda8G_goMux_mux_onehot, is_z_adda8G_goMux_mux_mux} = {5'd2,
                                                                     is_z_adda8G_2_2_argbuf_d};
      3'd2:
        {is_z_adda8G_goMux_mux_onehot, is_z_adda8G_goMux_mux_mux} = {5'd4,
                                                                     is_z_adda8G_3_2_argbuf_d};
      3'd3:
        {is_z_adda8G_goMux_mux_onehot, is_z_adda8G_goMux_mux_mux} = {5'd8,
                                                                     is_z_adda8G_4_1_argbuf_d};
      3'd4:
        {is_z_adda8G_goMux_mux_onehot, is_z_adda8G_goMux_mux_mux} = {5'd16,
                                                                     lizzieLet12_6QNode_Int_4QNode_Int_2_argbuf_d};
      default:
        {is_z_adda8G_goMux_mux_onehot, is_z_adda8G_goMux_mux_mux} = {5'd0,
                                                                     1'd0};
    endcase
  assign is_z_adda8G_goMux_mux_d = (is_z_adda8G_goMux_mux_mux[0] && go_12_goMux_choice_5_d[0]);
  assign go_12_goMux_choice_5_r = (is_z_adda8G_goMux_mux_d[0] && is_z_adda8G_goMux_mux_r);
  assign {lizzieLet12_6QNode_Int_4QNode_Int_2_argbuf_r,
          is_z_adda8G_4_1_argbuf_r,
          is_z_adda8G_3_2_argbuf_r,
          is_z_adda8G_2_2_argbuf_r,
          call_f_f_Int_Int_goMux6_r} = (go_12_goMux_choice_5_r ? is_z_adda8G_goMux_mux_onehot :
                                        5'd0);
  
  /* mux (Ty C5,
     Ty MyDTInt_Int_Int) : (go_12_goMux_choice_6,C5) [(call_f_f_Int_Int_goMux7,MyDTInt_Int_Int),
                                                      (op_adda8H_2_2_argbuf,MyDTInt_Int_Int),
                                                      (op_adda8H_3_2_argbuf,MyDTInt_Int_Int),
                                                      (op_adda8H_4_1_argbuf,MyDTInt_Int_Int),
                                                      (lizzieLet12_6QNode_Int_6QNode_Int_2_argbuf,MyDTInt_Int_Int)] > (op_adda8H_goMux_mux,MyDTInt_Int_Int) */
  logic [0:0] op_adda8H_goMux_mux_mux;
  logic [4:0] op_adda8H_goMux_mux_onehot;
  always_comb
    unique case (go_12_goMux_choice_6_d[3:1])
      3'd0:
        {op_adda8H_goMux_mux_onehot, op_adda8H_goMux_mux_mux} = {5'd1,
                                                                 call_f_f_Int_Int_goMux7_d};
      3'd1:
        {op_adda8H_goMux_mux_onehot, op_adda8H_goMux_mux_mux} = {5'd2,
                                                                 op_adda8H_2_2_argbuf_d};
      3'd2:
        {op_adda8H_goMux_mux_onehot, op_adda8H_goMux_mux_mux} = {5'd4,
                                                                 op_adda8H_3_2_argbuf_d};
      3'd3:
        {op_adda8H_goMux_mux_onehot, op_adda8H_goMux_mux_mux} = {5'd8,
                                                                 op_adda8H_4_1_argbuf_d};
      3'd4:
        {op_adda8H_goMux_mux_onehot, op_adda8H_goMux_mux_mux} = {5'd16,
                                                                 lizzieLet12_6QNode_Int_6QNode_Int_2_argbuf_d};
      default:
        {op_adda8H_goMux_mux_onehot, op_adda8H_goMux_mux_mux} = {5'd0,
                                                                 1'd0};
    endcase
  assign op_adda8H_goMux_mux_d = (op_adda8H_goMux_mux_mux[0] && go_12_goMux_choice_6_d[0]);
  assign go_12_goMux_choice_6_r = (op_adda8H_goMux_mux_d[0] && op_adda8H_goMux_mux_r);
  assign {lizzieLet12_6QNode_Int_6QNode_Int_2_argbuf_r,
          op_adda8H_4_1_argbuf_r,
          op_adda8H_3_2_argbuf_r,
          op_adda8H_2_2_argbuf_r,
          call_f_f_Int_Int_goMux7_r} = (go_12_goMux_choice_6_r ? op_adda8H_goMux_mux_onehot :
                                        5'd0);
  
  /* mux (Ty C5,
     Ty Pointer_CTf_f_Int_Int) : (go_12_goMux_choice_7,C5) [(call_f_f_Int_Int_goMux8,Pointer_CTf_f_Int_Int),
                                                            (sca2_2_1_argbuf,Pointer_CTf_f_Int_Int),
                                                            (sca1_2_1_argbuf,Pointer_CTf_f_Int_Int),
                                                            (sca0_2_1_argbuf,Pointer_CTf_f_Int_Int),
                                                            (sca3_2_1_argbuf,Pointer_CTf_f_Int_Int)] > (sc_0_2_goMux_mux,Pointer_CTf_f_Int_Int) */
  logic [16:0] sc_0_2_goMux_mux_mux;
  logic [4:0] sc_0_2_goMux_mux_onehot;
  always_comb
    unique case (go_12_goMux_choice_7_d[3:1])
      3'd0:
        {sc_0_2_goMux_mux_onehot, sc_0_2_goMux_mux_mux} = {5'd1,
                                                           call_f_f_Int_Int_goMux8_d};
      3'd1:
        {sc_0_2_goMux_mux_onehot, sc_0_2_goMux_mux_mux} = {5'd2,
                                                           sca2_2_1_argbuf_d};
      3'd2:
        {sc_0_2_goMux_mux_onehot, sc_0_2_goMux_mux_mux} = {5'd4,
                                                           sca1_2_1_argbuf_d};
      3'd3:
        {sc_0_2_goMux_mux_onehot, sc_0_2_goMux_mux_mux} = {5'd8,
                                                           sca0_2_1_argbuf_d};
      3'd4:
        {sc_0_2_goMux_mux_onehot, sc_0_2_goMux_mux_mux} = {5'd16,
                                                           sca3_2_1_argbuf_d};
      default:
        {sc_0_2_goMux_mux_onehot, sc_0_2_goMux_mux_mux} = {5'd0,
                                                           {16'd0, 1'd0}};
    endcase
  assign sc_0_2_goMux_mux_d = {sc_0_2_goMux_mux_mux[16:1],
                               (sc_0_2_goMux_mux_mux[0] && go_12_goMux_choice_7_d[0])};
  assign go_12_goMux_choice_7_r = (sc_0_2_goMux_mux_d[0] && sc_0_2_goMux_mux_r);
  assign {sca3_2_1_argbuf_r,
          sca0_2_1_argbuf_r,
          sca1_2_1_argbuf_r,
          sca2_2_1_argbuf_r,
          call_f_f_Int_Int_goMux8_r} = (go_12_goMux_choice_7_r ? sc_0_2_goMux_mux_onehot :
                                        5'd0);
  
  /* dcon (Ty CTf''''''''_f''''''''_Int_Int,
      Dcon Lf''''''''_f''''''''_Int_Intsbos) : [(go_13_1,Go)] > (go_13_1Lf''''''''_f''''''''_Int_Intsbos,CTf''''''''_f''''''''_Int_Int) */
  assign \go_13_1Lf''''''''_f''''''''_Int_Intsbos_d  = \Lf''''''''_f''''''''_Int_Intsbos_dc ((& {go_13_1_d[0]}), go_13_1_d);
  assign {go_13_1_r} = {1 {(\go_13_1Lf''''''''_f''''''''_Int_Intsbos_r  && \go_13_1Lf''''''''_f''''''''_Int_Intsbos_d [0])}};
  
  /* buf (Ty CTf''''''''_f''''''''_Int_Int) : (go_13_1Lf''''''''_f''''''''_Int_Intsbos,CTf''''''''_f''''''''_Int_Int) > (lizzieLet33_1_argbuf,CTf''''''''_f''''''''_Int_Int) */
  \CTf''''''''_f''''''''_Int_Int_t  \go_13_1Lf''''''''_f''''''''_Int_Intsbos_bufchan_d ;
  logic \go_13_1Lf''''''''_f''''''''_Int_Intsbos_bufchan_r ;
  assign \go_13_1Lf''''''''_f''''''''_Int_Intsbos_r  = ((! \go_13_1Lf''''''''_f''''''''_Int_Intsbos_bufchan_d [0]) || \go_13_1Lf''''''''_f''''''''_Int_Intsbos_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \go_13_1Lf''''''''_f''''''''_Int_Intsbos_bufchan_d  <= {67'd0,
                                                              1'd0};
    else
      if (\go_13_1Lf''''''''_f''''''''_Int_Intsbos_r )
        \go_13_1Lf''''''''_f''''''''_Int_Intsbos_bufchan_d  <= \go_13_1Lf''''''''_f''''''''_Int_Intsbos_d ;
  \CTf''''''''_f''''''''_Int_Int_t  \go_13_1Lf''''''''_f''''''''_Int_Intsbos_bufchan_buf ;
  assign \go_13_1Lf''''''''_f''''''''_Int_Intsbos_bufchan_r  = (! \go_13_1Lf''''''''_f''''''''_Int_Intsbos_bufchan_buf [0]);
  assign lizzieLet33_1_argbuf_d = (\go_13_1Lf''''''''_f''''''''_Int_Intsbos_bufchan_buf [0] ? \go_13_1Lf''''''''_f''''''''_Int_Intsbos_bufchan_buf  :
                                   \go_13_1Lf''''''''_f''''''''_Int_Intsbos_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \go_13_1Lf''''''''_f''''''''_Int_Intsbos_bufchan_buf  <= {67'd0,
                                                                1'd0};
    else
      if ((lizzieLet33_1_argbuf_r && \go_13_1Lf''''''''_f''''''''_Int_Intsbos_bufchan_buf [0]))
        \go_13_1Lf''''''''_f''''''''_Int_Intsbos_bufchan_buf  <= {67'd0,
                                                                  1'd0};
      else if (((! lizzieLet33_1_argbuf_r) && (! \go_13_1Lf''''''''_f''''''''_Int_Intsbos_bufchan_buf [0])))
        \go_13_1Lf''''''''_f''''''''_Int_Intsbos_bufchan_buf  <= \go_13_1Lf''''''''_f''''''''_Int_Intsbos_bufchan_d ;
  
  /* buf (Ty Go) : (go_13_2,Go) > (go_13_2_argbuf,Go) */
  Go_t go_13_2_bufchan_d;
  logic go_13_2_bufchan_r;
  assign go_13_2_r = ((! go_13_2_bufchan_d[0]) || go_13_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_13_2_bufchan_d <= 1'd0;
    else if (go_13_2_r) go_13_2_bufchan_d <= go_13_2_d;
  Go_t go_13_2_bufchan_buf;
  assign go_13_2_bufchan_r = (! go_13_2_bufchan_buf[0]);
  assign go_13_2_argbuf_d = (go_13_2_bufchan_buf[0] ? go_13_2_bufchan_buf :
                             go_13_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_13_2_bufchan_buf <= 1'd0;
    else
      if ((go_13_2_argbuf_r && go_13_2_bufchan_buf[0]))
        go_13_2_bufchan_buf <= 1'd0;
      else if (((! go_13_2_argbuf_r) && (! go_13_2_bufchan_buf[0])))
        go_13_2_bufchan_buf <= go_13_2_bufchan_d;
  
  /* dcon (Ty TupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf''''''''_f''''''''_Int_Int,
      Dcon TupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf''''''''_f''''''''_Int_Int) : [(go_13_2_argbuf,Go),
                                                                                                              (q4a8u_1_1_argbuf,Pointer_QTree_Int),
                                                                                                              (is_z_mapa8v_1_1_argbuf,MyDTInt_Bool),
                                                                                                              (op_mapa8w_1_1_argbuf,MyDTInt_Int),
                                                                                                              (lizzieLet5_1_1_argbuf,Pointer_CTf''''''''_f''''''''_Int_Int)] > (call_f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf''''''''_f''''''''_Int_Int_1,TupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf''''''''_f''''''''_Int_Int) */
  assign \call_f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf''''''''_f''''''''_Int_Int_1_d  = \TupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf''''''''_f''''''''_Int_Int_dc ((& {go_13_2_argbuf_d[0],
                                                                                                                                                                                                                                                        q4a8u_1_1_argbuf_d[0],
                                                                                                                                                                                                                                                        is_z_mapa8v_1_1_argbuf_d[0],
                                                                                                                                                                                                                                                        op_mapa8w_1_1_argbuf_d[0],
                                                                                                                                                                                                                                                        lizzieLet5_1_1_argbuf_d[0]}), go_13_2_argbuf_d, q4a8u_1_1_argbuf_d, is_z_mapa8v_1_1_argbuf_d, op_mapa8w_1_1_argbuf_d, lizzieLet5_1_1_argbuf_d);
  assign {go_13_2_argbuf_r,
          q4a8u_1_1_argbuf_r,
          is_z_mapa8v_1_1_argbuf_r,
          op_mapa8w_1_1_argbuf_r,
          lizzieLet5_1_1_argbuf_r} = {5 {(\call_f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf''''''''_f''''''''_Int_Int_1_r  && \call_f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf''''''''_f''''''''_Int_Int_1_d [0])}};
  
  /* dcon (Ty CTf_f_Int_Int,
      Dcon Lf_f_Int_Intsbos) : [(go_14_1,Go)] > (go_14_1Lf_f_Int_Intsbos,CTf_f_Int_Int) */
  assign go_14_1Lf_f_Int_Intsbos_d = Lf_f_Int_Intsbos_dc((& {go_14_1_d[0]}), go_14_1_d);
  assign {go_14_1_r} = {1 {(go_14_1Lf_f_Int_Intsbos_r && go_14_1Lf_f_Int_Intsbos_d[0])}};
  
  /* buf (Ty CTf_f_Int_Int) : (go_14_1Lf_f_Int_Intsbos,CTf_f_Int_Int) > (lizzieLet34_1_argbuf,CTf_f_Int_Int) */
  CTf_f_Int_Int_t go_14_1Lf_f_Int_Intsbos_bufchan_d;
  logic go_14_1Lf_f_Int_Intsbos_bufchan_r;
  assign go_14_1Lf_f_Int_Intsbos_r = ((! go_14_1Lf_f_Int_Intsbos_bufchan_d[0]) || go_14_1Lf_f_Int_Intsbos_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      go_14_1Lf_f_Int_Intsbos_bufchan_d <= {115'd0, 1'd0};
    else
      if (go_14_1Lf_f_Int_Intsbos_r)
        go_14_1Lf_f_Int_Intsbos_bufchan_d <= go_14_1Lf_f_Int_Intsbos_d;
  CTf_f_Int_Int_t go_14_1Lf_f_Int_Intsbos_bufchan_buf;
  assign go_14_1Lf_f_Int_Intsbos_bufchan_r = (! go_14_1Lf_f_Int_Intsbos_bufchan_buf[0]);
  assign lizzieLet34_1_argbuf_d = (go_14_1Lf_f_Int_Intsbos_bufchan_buf[0] ? go_14_1Lf_f_Int_Intsbos_bufchan_buf :
                                   go_14_1Lf_f_Int_Intsbos_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      go_14_1Lf_f_Int_Intsbos_bufchan_buf <= {115'd0, 1'd0};
    else
      if ((lizzieLet34_1_argbuf_r && go_14_1Lf_f_Int_Intsbos_bufchan_buf[0]))
        go_14_1Lf_f_Int_Intsbos_bufchan_buf <= {115'd0, 1'd0};
      else if (((! lizzieLet34_1_argbuf_r) && (! go_14_1Lf_f_Int_Intsbos_bufchan_buf[0])))
        go_14_1Lf_f_Int_Intsbos_bufchan_buf <= go_14_1Lf_f_Int_Intsbos_bufchan_d;
  
  /* buf (Ty Go) : (go_14_2,Go) > (go_14_2_argbuf,Go) */
  Go_t go_14_2_bufchan_d;
  logic go_14_2_bufchan_r;
  assign go_14_2_r = ((! go_14_2_bufchan_d[0]) || go_14_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_14_2_bufchan_d <= 1'd0;
    else if (go_14_2_r) go_14_2_bufchan_d <= go_14_2_d;
  Go_t go_14_2_bufchan_buf;
  assign go_14_2_bufchan_r = (! go_14_2_bufchan_buf[0]);
  assign go_14_2_argbuf_d = (go_14_2_bufchan_buf[0] ? go_14_2_bufchan_buf :
                             go_14_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_14_2_bufchan_buf <= 1'd0;
    else
      if ((go_14_2_argbuf_r && go_14_2_bufchan_buf[0]))
        go_14_2_bufchan_buf <= 1'd0;
      else if (((! go_14_2_argbuf_r) && (! go_14_2_bufchan_buf[0])))
        go_14_2_bufchan_buf <= go_14_2_bufchan_d;
  
  /* dcon (Ty TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Int,
      Dcon TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Int) : [(go_14_2_argbuf,Go),
                                                                                                                                                   (m1a8C_1_1_argbuf,Pointer_QTree_Int),
                                                                                                                                                   (m2a8D_1_1_argbuf,Pointer_QTree_Int),
                                                                                                                                                   (is_z_mapa8E_1_1_argbuf,MyDTInt_Bool),
                                                                                                                                                   (op_mapa8F_1_1_argbuf,MyDTInt_Int),
                                                                                                                                                   (is_z_adda8G_1_1_argbuf,MyDTInt_Bool),
                                                                                                                                                   (op_adda8H_1_1_argbuf,MyDTInt_Int_Int),
                                                                                                                                                   (lizzieLet22_1_1_argbuf,Pointer_CTf_f_Int_Int)] > (call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Int_1,TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Int) */
  assign call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Int_1_d = TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Int_dc((& {go_14_2_argbuf_d[0],
                                                                                                                                                                                                                                                                                                              m1a8C_1_1_argbuf_d[0],
                                                                                                                                                                                                                                                                                                              m2a8D_1_1_argbuf_d[0],
                                                                                                                                                                                                                                                                                                              is_z_mapa8E_1_1_argbuf_d[0],
                                                                                                                                                                                                                                                                                                              op_mapa8F_1_1_argbuf_d[0],
                                                                                                                                                                                                                                                                                                              is_z_adda8G_1_1_argbuf_d[0],
                                                                                                                                                                                                                                                                                                              op_adda8H_1_1_argbuf_d[0],
                                                                                                                                                                                                                                                                                                              lizzieLet22_1_1_argbuf_d[0]}), go_14_2_argbuf_d, m1a8C_1_1_argbuf_d, m2a8D_1_1_argbuf_d, is_z_mapa8E_1_1_argbuf_d, op_mapa8F_1_1_argbuf_d, is_z_adda8G_1_1_argbuf_d, op_adda8H_1_1_argbuf_d, lizzieLet22_1_1_argbuf_d);
  assign {go_14_2_argbuf_r,
          m1a8C_1_1_argbuf_r,
          m2a8D_1_1_argbuf_r,
          is_z_mapa8E_1_1_argbuf_r,
          op_mapa8F_1_1_argbuf_r,
          is_z_adda8G_1_1_argbuf_r,
          op_adda8H_1_1_argbuf_r,
          lizzieLet22_1_1_argbuf_r} = {8 {(call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Int_1_r && call_f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_Int_1_d[0])}};
  
  /* fork (Ty C4) : (go_15_goMux_choice,C4) > [(go_15_goMux_choice_1,C4),
                                          (go_15_goMux_choice_2,C4)] */
  logic [1:0] go_15_goMux_choice_emitted;
  logic [1:0] go_15_goMux_choice_done;
  assign go_15_goMux_choice_1_d = {go_15_goMux_choice_d[2:1],
                                   (go_15_goMux_choice_d[0] && (! go_15_goMux_choice_emitted[0]))};
  assign go_15_goMux_choice_2_d = {go_15_goMux_choice_d[2:1],
                                   (go_15_goMux_choice_d[0] && (! go_15_goMux_choice_emitted[1]))};
  assign go_15_goMux_choice_done = (go_15_goMux_choice_emitted | ({go_15_goMux_choice_2_d[0],
                                                                   go_15_goMux_choice_1_d[0]} & {go_15_goMux_choice_2_r,
                                                                                                 go_15_goMux_choice_1_r}));
  assign go_15_goMux_choice_r = (& go_15_goMux_choice_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_15_goMux_choice_emitted <= 2'd0;
    else
      go_15_goMux_choice_emitted <= (go_15_goMux_choice_r ? 2'd0 :
                                     go_15_goMux_choice_done);
  
  /* mux (Ty C4,
     Ty Int#) : (go_15_goMux_choice_1,C4) [(lizzieLet23_1_argbuf,Int#),
                                           (contRet_0_1_argbuf,Int#),
                                           (lizzieLet24_1_argbuf,Int#),
                                           (lizzieLet23_1_1_argbuf,Int#)] > (srtarg_0_goMux_mux,Int#) */
  logic [32:0] srtarg_0_goMux_mux_mux;
  logic [3:0] srtarg_0_goMux_mux_onehot;
  always_comb
    unique case (go_15_goMux_choice_1_d[2:1])
      2'd0:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {4'd1,
                                                               lizzieLet23_1_argbuf_d};
      2'd1:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {4'd2,
                                                               contRet_0_1_argbuf_d};
      2'd2:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {4'd4,
                                                               lizzieLet24_1_argbuf_d};
      2'd3:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {4'd8,
                                                               lizzieLet23_1_1_argbuf_d};
      default:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {4'd0,
                                                               {32'd0, 1'd0}};
    endcase
  assign srtarg_0_goMux_mux_d = {srtarg_0_goMux_mux_mux[32:1],
                                 (srtarg_0_goMux_mux_mux[0] && go_15_goMux_choice_1_d[0])};
  assign go_15_goMux_choice_1_r = (srtarg_0_goMux_mux_d[0] && srtarg_0_goMux_mux_r);
  assign {lizzieLet23_1_1_argbuf_r,
          lizzieLet24_1_argbuf_r,
          contRet_0_1_argbuf_r,
          lizzieLet23_1_argbuf_r} = (go_15_goMux_choice_1_r ? srtarg_0_goMux_mux_onehot :
                                     4'd0);
  
  /* mux (Ty C4,
     Ty Pointer_CT$wnnz) : (go_15_goMux_choice_2,C4) [(lizzieLet4_4QNone_Int_1_argbuf,Pointer_CT$wnnz),
                                                      (sc_0_6_1_argbuf,Pointer_CT$wnnz),
                                                      (lizzieLet4_4QVal_Int_1_argbuf,Pointer_CT$wnnz),
                                                      (lizzieLet4_4QError_Int_1_argbuf,Pointer_CT$wnnz)] > (scfarg_0_goMux_mux,Pointer_CT$wnnz) */
  logic [16:0] scfarg_0_goMux_mux_mux;
  logic [3:0] scfarg_0_goMux_mux_onehot;
  always_comb
    unique case (go_15_goMux_choice_2_d[2:1])
      2'd0:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {4'd1,
                                                               lizzieLet4_4QNone_Int_1_argbuf_d};
      2'd1:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {4'd2,
                                                               sc_0_6_1_argbuf_d};
      2'd2:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {4'd4,
                                                               lizzieLet4_4QVal_Int_1_argbuf_d};
      2'd3:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {4'd8,
                                                               lizzieLet4_4QError_Int_1_argbuf_d};
      default:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {4'd0,
                                                               {16'd0, 1'd0}};
    endcase
  assign scfarg_0_goMux_mux_d = {scfarg_0_goMux_mux_mux[16:1],
                                 (scfarg_0_goMux_mux_mux[0] && go_15_goMux_choice_2_d[0])};
  assign go_15_goMux_choice_2_r = (scfarg_0_goMux_mux_d[0] && scfarg_0_goMux_mux_r);
  assign {lizzieLet4_4QError_Int_1_argbuf_r,
          lizzieLet4_4QVal_Int_1_argbuf_r,
          sc_0_6_1_argbuf_r,
          lizzieLet4_4QNone_Int_1_argbuf_r} = (go_15_goMux_choice_2_r ? scfarg_0_goMux_mux_onehot :
                                               4'd0);
  
  /* fork (Ty C5) : (go_16_goMux_choice,C5) > [(go_16_goMux_choice_1,C5),
                                          (go_16_goMux_choice_2,C5)] */
  logic [1:0] go_16_goMux_choice_emitted;
  logic [1:0] go_16_goMux_choice_done;
  assign go_16_goMux_choice_1_d = {go_16_goMux_choice_d[3:1],
                                   (go_16_goMux_choice_d[0] && (! go_16_goMux_choice_emitted[0]))};
  assign go_16_goMux_choice_2_d = {go_16_goMux_choice_d[3:1],
                                   (go_16_goMux_choice_d[0] && (! go_16_goMux_choice_emitted[1]))};
  assign go_16_goMux_choice_done = (go_16_goMux_choice_emitted | ({go_16_goMux_choice_2_d[0],
                                                                   go_16_goMux_choice_1_d[0]} & {go_16_goMux_choice_2_r,
                                                                                                 go_16_goMux_choice_1_r}));
  assign go_16_goMux_choice_r = (& go_16_goMux_choice_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_16_goMux_choice_emitted <= 2'd0;
    else
      go_16_goMux_choice_emitted <= (go_16_goMux_choice_r ? 2'd0 :
                                     go_16_goMux_choice_done);
  
  /* mux (Ty C5,
     Ty Pointer_QTree_Int) : (go_16_goMux_choice_1,C5) [(lizzieLet1_1_1_argbuf,Pointer_QTree_Int),
                                                        (contRet_0_1_1_argbuf,Pointer_QTree_Int),
                                                        (lizzieLet2_1_1_argbuf,Pointer_QTree_Int),
                                                        (lizzieLet3_1_1_argbuf,Pointer_QTree_Int),
                                                        (lizzieLet4_1_1_argbuf,Pointer_QTree_Int)] > (srtarg_0_1_goMux_mux,Pointer_QTree_Int) */
  logic [16:0] srtarg_0_1_goMux_mux_mux;
  logic [4:0] srtarg_0_1_goMux_mux_onehot;
  always_comb
    unique case (go_16_goMux_choice_1_d[3:1])
      3'd0:
        {srtarg_0_1_goMux_mux_onehot, srtarg_0_1_goMux_mux_mux} = {5'd1,
                                                                   lizzieLet1_1_1_argbuf_d};
      3'd1:
        {srtarg_0_1_goMux_mux_onehot, srtarg_0_1_goMux_mux_mux} = {5'd2,
                                                                   contRet_0_1_1_argbuf_d};
      3'd2:
        {srtarg_0_1_goMux_mux_onehot, srtarg_0_1_goMux_mux_mux} = {5'd4,
                                                                   lizzieLet2_1_1_argbuf_d};
      3'd3:
        {srtarg_0_1_goMux_mux_onehot, srtarg_0_1_goMux_mux_mux} = {5'd8,
                                                                   lizzieLet3_1_1_argbuf_d};
      3'd4:
        {srtarg_0_1_goMux_mux_onehot, srtarg_0_1_goMux_mux_mux} = {5'd16,
                                                                   lizzieLet4_1_1_argbuf_d};
      default:
        {srtarg_0_1_goMux_mux_onehot, srtarg_0_1_goMux_mux_mux} = {5'd0,
                                                                   {16'd0, 1'd0}};
    endcase
  assign srtarg_0_1_goMux_mux_d = {srtarg_0_1_goMux_mux_mux[16:1],
                                   (srtarg_0_1_goMux_mux_mux[0] && go_16_goMux_choice_1_d[0])};
  assign go_16_goMux_choice_1_r = (srtarg_0_1_goMux_mux_d[0] && srtarg_0_1_goMux_mux_r);
  assign {lizzieLet4_1_1_argbuf_r,
          lizzieLet3_1_1_argbuf_r,
          lizzieLet2_1_1_argbuf_r,
          contRet_0_1_1_argbuf_r,
          lizzieLet1_1_1_argbuf_r} = (go_16_goMux_choice_1_r ? srtarg_0_1_goMux_mux_onehot :
                                      5'd0);
  
  /* mux (Ty C5,
     Ty Pointer_CTf''''''''_f''''''''_Int_Int) : (go_16_goMux_choice_2,C5) [(lizzieLet6_6QNone_Int_1_argbuf,Pointer_CTf''''''''_f''''''''_Int_Int),
                                                                            (sc_0_10_1_argbuf,Pointer_CTf''''''''_f''''''''_Int_Int),
                                                                            (es_2_3MyFalse_1_argbuf,Pointer_CTf''''''''_f''''''''_Int_Int),
                                                                            (es_2_3MyTrue_1_argbuf,Pointer_CTf''''''''_f''''''''_Int_Int),
                                                                            (lizzieLet6_6QError_Int_1_argbuf,Pointer_CTf''''''''_f''''''''_Int_Int)] > (scfarg_0_1_goMux_mux,Pointer_CTf''''''''_f''''''''_Int_Int) */
  logic [16:0] scfarg_0_1_goMux_mux_mux;
  logic [4:0] scfarg_0_1_goMux_mux_onehot;
  always_comb
    unique case (go_16_goMux_choice_2_d[3:1])
      3'd0:
        {scfarg_0_1_goMux_mux_onehot, scfarg_0_1_goMux_mux_mux} = {5'd1,
                                                                   lizzieLet6_6QNone_Int_1_argbuf_d};
      3'd1:
        {scfarg_0_1_goMux_mux_onehot, scfarg_0_1_goMux_mux_mux} = {5'd2,
                                                                   sc_0_10_1_argbuf_d};
      3'd2:
        {scfarg_0_1_goMux_mux_onehot, scfarg_0_1_goMux_mux_mux} = {5'd4,
                                                                   es_2_3MyFalse_1_argbuf_d};
      3'd3:
        {scfarg_0_1_goMux_mux_onehot, scfarg_0_1_goMux_mux_mux} = {5'd8,
                                                                   es_2_3MyTrue_1_argbuf_d};
      3'd4:
        {scfarg_0_1_goMux_mux_onehot, scfarg_0_1_goMux_mux_mux} = {5'd16,
                                                                   lizzieLet6_6QError_Int_1_argbuf_d};
      default:
        {scfarg_0_1_goMux_mux_onehot, scfarg_0_1_goMux_mux_mux} = {5'd0,
                                                                   {16'd0, 1'd0}};
    endcase
  assign scfarg_0_1_goMux_mux_d = {scfarg_0_1_goMux_mux_mux[16:1],
                                   (scfarg_0_1_goMux_mux_mux[0] && go_16_goMux_choice_2_d[0])};
  assign go_16_goMux_choice_2_r = (scfarg_0_1_goMux_mux_d[0] && scfarg_0_1_goMux_mux_r);
  assign {lizzieLet6_6QError_Int_1_argbuf_r,
          es_2_3MyTrue_1_argbuf_r,
          es_2_3MyFalse_1_argbuf_r,
          sc_0_10_1_argbuf_r,
          lizzieLet6_6QNone_Int_1_argbuf_r} = (go_16_goMux_choice_2_r ? scfarg_0_1_goMux_mux_onehot :
                                               5'd0);
  
  /* fork (Ty C17) : (go_17_goMux_choice,C17) > [(go_17_goMux_choice_1,C17),
                                            (go_17_goMux_choice_2,C17)] */
  logic [1:0] go_17_goMux_choice_emitted;
  logic [1:0] go_17_goMux_choice_done;
  assign go_17_goMux_choice_1_d = {go_17_goMux_choice_d[5:1],
                                   (go_17_goMux_choice_d[0] && (! go_17_goMux_choice_emitted[0]))};
  assign go_17_goMux_choice_2_d = {go_17_goMux_choice_d[5:1],
                                   (go_17_goMux_choice_d[0] && (! go_17_goMux_choice_emitted[1]))};
  assign go_17_goMux_choice_done = (go_17_goMux_choice_emitted | ({go_17_goMux_choice_2_d[0],
                                                                   go_17_goMux_choice_1_d[0]} & {go_17_goMux_choice_2_r,
                                                                                                 go_17_goMux_choice_1_r}));
  assign go_17_goMux_choice_r = (& go_17_goMux_choice_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_17_goMux_choice_emitted <= 2'd0;
    else
      go_17_goMux_choice_emitted <= (go_17_goMux_choice_r ? 2'd0 :
                                     go_17_goMux_choice_done);
  
  /* mux (Ty C17,
     Ty Pointer_QTree_Int) : (go_17_goMux_choice_1,C17) [(lizzieLet6_1_1_argbuf,Pointer_QTree_Int),
                                                         (contRet_0_2_1_argbuf,Pointer_QTree_Int),
                                                         (lizzieLet7_1_1_argbuf,Pointer_QTree_Int),
                                                         (lizzieLet8_1_1_argbuf,Pointer_QTree_Int),
                                                         (lizzieLet9_1_1_argbuf,Pointer_QTree_Int),
                                                         (lizzieLet10_1_1_argbuf,Pointer_QTree_Int),
                                                         (lizzieLet11_1_1_argbuf,Pointer_QTree_Int),
                                                         (lizzieLet12_1_1_argbuf,Pointer_QTree_Int),
                                                         (lizzieLet13_1_1_argbuf,Pointer_QTree_Int),
                                                         (lizzieLet14_1_1_argbuf,Pointer_QTree_Int),
                                                         (lizzieLet15_1_1_argbuf,Pointer_QTree_Int),
                                                         (lizzieLet16_1_1_argbuf,Pointer_QTree_Int),
                                                         (lizzieLet17_1_1_argbuf,Pointer_QTree_Int),
                                                         (lizzieLet18_1_1_argbuf,Pointer_QTree_Int),
                                                         (lizzieLet19_1_argbuf,Pointer_QTree_Int),
                                                         (lizzieLet20_1_1_argbuf,Pointer_QTree_Int),
                                                         (lizzieLet21_1_1_argbuf,Pointer_QTree_Int)] > (srtarg_0_2_goMux_mux,Pointer_QTree_Int) */
  logic [16:0] srtarg_0_2_goMux_mux_mux;
  logic [16:0] srtarg_0_2_goMux_mux_onehot;
  always_comb
    unique case (go_17_goMux_choice_1_d[5:1])
      5'd0:
        {srtarg_0_2_goMux_mux_onehot, srtarg_0_2_goMux_mux_mux} = {17'd1,
                                                                   lizzieLet6_1_1_argbuf_d};
      5'd1:
        {srtarg_0_2_goMux_mux_onehot, srtarg_0_2_goMux_mux_mux} = {17'd2,
                                                                   contRet_0_2_1_argbuf_d};
      5'd2:
        {srtarg_0_2_goMux_mux_onehot, srtarg_0_2_goMux_mux_mux} = {17'd4,
                                                                   lizzieLet7_1_1_argbuf_d};
      5'd3:
        {srtarg_0_2_goMux_mux_onehot, srtarg_0_2_goMux_mux_mux} = {17'd8,
                                                                   lizzieLet8_1_1_argbuf_d};
      5'd4:
        {srtarg_0_2_goMux_mux_onehot, srtarg_0_2_goMux_mux_mux} = {17'd16,
                                                                   lizzieLet9_1_1_argbuf_d};
      5'd5:
        {srtarg_0_2_goMux_mux_onehot, srtarg_0_2_goMux_mux_mux} = {17'd32,
                                                                   lizzieLet10_1_1_argbuf_d};
      5'd6:
        {srtarg_0_2_goMux_mux_onehot, srtarg_0_2_goMux_mux_mux} = {17'd64,
                                                                   lizzieLet11_1_1_argbuf_d};
      5'd7:
        {srtarg_0_2_goMux_mux_onehot, srtarg_0_2_goMux_mux_mux} = {17'd128,
                                                                   lizzieLet12_1_1_argbuf_d};
      5'd8:
        {srtarg_0_2_goMux_mux_onehot, srtarg_0_2_goMux_mux_mux} = {17'd256,
                                                                   lizzieLet13_1_1_argbuf_d};
      5'd9:
        {srtarg_0_2_goMux_mux_onehot, srtarg_0_2_goMux_mux_mux} = {17'd512,
                                                                   lizzieLet14_1_1_argbuf_d};
      5'd10:
        {srtarg_0_2_goMux_mux_onehot,
         srtarg_0_2_goMux_mux_mux} = {17'd1024, lizzieLet15_1_1_argbuf_d};
      5'd11:
        {srtarg_0_2_goMux_mux_onehot,
         srtarg_0_2_goMux_mux_mux} = {17'd2048, lizzieLet16_1_1_argbuf_d};
      5'd12:
        {srtarg_0_2_goMux_mux_onehot,
         srtarg_0_2_goMux_mux_mux} = {17'd4096, lizzieLet17_1_1_argbuf_d};
      5'd13:
        {srtarg_0_2_goMux_mux_onehot,
         srtarg_0_2_goMux_mux_mux} = {17'd8192, lizzieLet18_1_1_argbuf_d};
      5'd14:
        {srtarg_0_2_goMux_mux_onehot,
         srtarg_0_2_goMux_mux_mux} = {17'd16384, lizzieLet19_1_argbuf_d};
      5'd15:
        {srtarg_0_2_goMux_mux_onehot,
         srtarg_0_2_goMux_mux_mux} = {17'd32768, lizzieLet20_1_1_argbuf_d};
      5'd16:
        {srtarg_0_2_goMux_mux_onehot,
         srtarg_0_2_goMux_mux_mux} = {17'd65536, lizzieLet21_1_1_argbuf_d};
      default:
        {srtarg_0_2_goMux_mux_onehot, srtarg_0_2_goMux_mux_mux} = {17'd0,
                                                                   {16'd0, 1'd0}};
    endcase
  assign srtarg_0_2_goMux_mux_d = {srtarg_0_2_goMux_mux_mux[16:1],
                                   (srtarg_0_2_goMux_mux_mux[0] && go_17_goMux_choice_1_d[0])};
  assign go_17_goMux_choice_1_r = (srtarg_0_2_goMux_mux_d[0] && srtarg_0_2_goMux_mux_r);
  assign {lizzieLet21_1_1_argbuf_r,
          lizzieLet20_1_1_argbuf_r,
          lizzieLet19_1_argbuf_r,
          lizzieLet18_1_1_argbuf_r,
          lizzieLet17_1_1_argbuf_r,
          lizzieLet16_1_1_argbuf_r,
          lizzieLet15_1_1_argbuf_r,
          lizzieLet14_1_1_argbuf_r,
          lizzieLet13_1_1_argbuf_r,
          lizzieLet12_1_1_argbuf_r,
          lizzieLet11_1_1_argbuf_r,
          lizzieLet10_1_1_argbuf_r,
          lizzieLet9_1_1_argbuf_r,
          lizzieLet8_1_1_argbuf_r,
          lizzieLet7_1_1_argbuf_r,
          contRet_0_2_1_argbuf_r,
          lizzieLet6_1_1_argbuf_r} = (go_17_goMux_choice_1_r ? srtarg_0_2_goMux_mux_onehot :
                                      17'd0);
  
  /* mux (Ty C17,
     Ty Pointer_CTf_f_Int_Int) : (go_17_goMux_choice_2,C17) [(lizzieLet12_6QNone_Int_6QNone_Int_1_argbuf,Pointer_CTf_f_Int_Int),
                                                             (sc_0_14_1_argbuf,Pointer_CTf_f_Int_Int),
                                                             (es_2_1_3MyFalse_1_argbuf,Pointer_CTf_f_Int_Int),
                                                             (es_2_1_3MyTrue_1_argbuf,Pointer_CTf_f_Int_Int),
                                                             (lizzieLet12_6QNone_Int_6QNode_Int_1_argbuf,Pointer_CTf_f_Int_Int),
                                                             (lizzieLet12_6QNone_Int_6QError_Int_1_argbuf,Pointer_CTf_f_Int_Int),
                                                             (es_10_3MyFalse_1_argbuf,Pointer_CTf_f_Int_Int),
                                                             (es_10_3MyTrue_1_argbuf,Pointer_CTf_f_Int_Int),
                                                             (es_19_4MyFalse_1_argbuf,Pointer_CTf_f_Int_Int),
                                                             (es_19_4MyTrue_1_argbuf,Pointer_CTf_f_Int_Int),
                                                             (es_14_5MyTrue_1_argbuf,Pointer_CTf_f_Int_Int),
                                                             (lizzieLet12_6QVal_Int_8QNode_Int_1_argbuf,Pointer_CTf_f_Int_Int),
                                                             (lizzieLet12_6QVal_Int_8QError_Int_1_argbuf,Pointer_CTf_f_Int_Int),
                                                             (lizzieLet12_6QNode_Int_8QNone_Int_1_argbuf,Pointer_CTf_f_Int_Int),
                                                             (lizzieLet12_6QNode_Int_8QVal_Int_1_argbuf,Pointer_CTf_f_Int_Int),
                                                             (lizzieLet12_6QNode_Int_8QError_Int_1_argbuf,Pointer_CTf_f_Int_Int),
                                                             (lizzieLet12_9QError_Int_1_argbuf,Pointer_CTf_f_Int_Int)] > (scfarg_0_2_goMux_mux,Pointer_CTf_f_Int_Int) */
  logic [16:0] scfarg_0_2_goMux_mux_mux;
  logic [16:0] scfarg_0_2_goMux_mux_onehot;
  always_comb
    unique case (go_17_goMux_choice_2_d[5:1])
      5'd0:
        {scfarg_0_2_goMux_mux_onehot, scfarg_0_2_goMux_mux_mux} = {17'd1,
                                                                   lizzieLet12_6QNone_Int_6QNone_Int_1_argbuf_d};
      5'd1:
        {scfarg_0_2_goMux_mux_onehot, scfarg_0_2_goMux_mux_mux} = {17'd2,
                                                                   sc_0_14_1_argbuf_d};
      5'd2:
        {scfarg_0_2_goMux_mux_onehot, scfarg_0_2_goMux_mux_mux} = {17'd4,
                                                                   es_2_1_3MyFalse_1_argbuf_d};
      5'd3:
        {scfarg_0_2_goMux_mux_onehot, scfarg_0_2_goMux_mux_mux} = {17'd8,
                                                                   es_2_1_3MyTrue_1_argbuf_d};
      5'd4:
        {scfarg_0_2_goMux_mux_onehot, scfarg_0_2_goMux_mux_mux} = {17'd16,
                                                                   lizzieLet12_6QNone_Int_6QNode_Int_1_argbuf_d};
      5'd5:
        {scfarg_0_2_goMux_mux_onehot, scfarg_0_2_goMux_mux_mux} = {17'd32,
                                                                   lizzieLet12_6QNone_Int_6QError_Int_1_argbuf_d};
      5'd6:
        {scfarg_0_2_goMux_mux_onehot, scfarg_0_2_goMux_mux_mux} = {17'd64,
                                                                   es_10_3MyFalse_1_argbuf_d};
      5'd7:
        {scfarg_0_2_goMux_mux_onehot, scfarg_0_2_goMux_mux_mux} = {17'd128,
                                                                   es_10_3MyTrue_1_argbuf_d};
      5'd8:
        {scfarg_0_2_goMux_mux_onehot, scfarg_0_2_goMux_mux_mux} = {17'd256,
                                                                   es_19_4MyFalse_1_argbuf_d};
      5'd9:
        {scfarg_0_2_goMux_mux_onehot, scfarg_0_2_goMux_mux_mux} = {17'd512,
                                                                   es_19_4MyTrue_1_argbuf_d};
      5'd10:
        {scfarg_0_2_goMux_mux_onehot,
         scfarg_0_2_goMux_mux_mux} = {17'd1024, es_14_5MyTrue_1_argbuf_d};
      5'd11:
        {scfarg_0_2_goMux_mux_onehot,
         scfarg_0_2_goMux_mux_mux} = {17'd2048,
                                      lizzieLet12_6QVal_Int_8QNode_Int_1_argbuf_d};
      5'd12:
        {scfarg_0_2_goMux_mux_onehot,
         scfarg_0_2_goMux_mux_mux} = {17'd4096,
                                      lizzieLet12_6QVal_Int_8QError_Int_1_argbuf_d};
      5'd13:
        {scfarg_0_2_goMux_mux_onehot,
         scfarg_0_2_goMux_mux_mux} = {17'd8192,
                                      lizzieLet12_6QNode_Int_8QNone_Int_1_argbuf_d};
      5'd14:
        {scfarg_0_2_goMux_mux_onehot,
         scfarg_0_2_goMux_mux_mux} = {17'd16384,
                                      lizzieLet12_6QNode_Int_8QVal_Int_1_argbuf_d};
      5'd15:
        {scfarg_0_2_goMux_mux_onehot,
         scfarg_0_2_goMux_mux_mux} = {17'd32768,
                                      lizzieLet12_6QNode_Int_8QError_Int_1_argbuf_d};
      5'd16:
        {scfarg_0_2_goMux_mux_onehot,
         scfarg_0_2_goMux_mux_mux} = {17'd65536,
                                      lizzieLet12_9QError_Int_1_argbuf_d};
      default:
        {scfarg_0_2_goMux_mux_onehot, scfarg_0_2_goMux_mux_mux} = {17'd0,
                                                                   {16'd0, 1'd0}};
    endcase
  assign scfarg_0_2_goMux_mux_d = {scfarg_0_2_goMux_mux_mux[16:1],
                                   (scfarg_0_2_goMux_mux_mux[0] && go_17_goMux_choice_2_d[0])};
  assign go_17_goMux_choice_2_r = (scfarg_0_2_goMux_mux_d[0] && scfarg_0_2_goMux_mux_r);
  assign {lizzieLet12_9QError_Int_1_argbuf_r,
          lizzieLet12_6QNode_Int_8QError_Int_1_argbuf_r,
          lizzieLet12_6QNode_Int_8QVal_Int_1_argbuf_r,
          lizzieLet12_6QNode_Int_8QNone_Int_1_argbuf_r,
          lizzieLet12_6QVal_Int_8QError_Int_1_argbuf_r,
          lizzieLet12_6QVal_Int_8QNode_Int_1_argbuf_r,
          es_14_5MyTrue_1_argbuf_r,
          es_19_4MyTrue_1_argbuf_r,
          es_19_4MyFalse_1_argbuf_r,
          es_10_3MyTrue_1_argbuf_r,
          es_10_3MyFalse_1_argbuf_r,
          lizzieLet12_6QNone_Int_6QError_Int_1_argbuf_r,
          lizzieLet12_6QNone_Int_6QNode_Int_1_argbuf_r,
          es_2_1_3MyTrue_1_argbuf_r,
          es_2_1_3MyFalse_1_argbuf_r,
          sc_0_14_1_argbuf_r,
          lizzieLet12_6QNone_Int_6QNone_Int_1_argbuf_r} = (go_17_goMux_choice_2_r ? scfarg_0_2_goMux_mux_onehot :
                                                           17'd0);
  
  /* buf (Ty MyDTInt_Int_Int) : (go_1Dcon_$fNumInt_$c+,MyDTInt_Int_Int) > (es_6_1_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t \go_1Dcon_$fNumInt_$c+_bufchan_d ;
  logic \go_1Dcon_$fNumInt_$c+_bufchan_r ;
  assign \go_1Dcon_$fNumInt_$c+_r  = ((! \go_1Dcon_$fNumInt_$c+_bufchan_d [0]) || \go_1Dcon_$fNumInt_$c+_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \go_1Dcon_$fNumInt_$c+_bufchan_d  <= 1'd0;
    else
      if (\go_1Dcon_$fNumInt_$c+_r )
        \go_1Dcon_$fNumInt_$c+_bufchan_d  <= \go_1Dcon_$fNumInt_$c+_d ;
  MyDTInt_Int_Int_t \go_1Dcon_$fNumInt_$c+_bufchan_buf ;
  assign \go_1Dcon_$fNumInt_$c+_bufchan_r  = (! \go_1Dcon_$fNumInt_$c+_bufchan_buf [0]);
  assign es_6_1_argbuf_d = (\go_1Dcon_$fNumInt_$c+_bufchan_buf [0] ? \go_1Dcon_$fNumInt_$c+_bufchan_buf  :
                            \go_1Dcon_$fNumInt_$c+_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \go_1Dcon_$fNumInt_$c+_bufchan_buf  <= 1'd0;
    else
      if ((es_6_1_argbuf_r && \go_1Dcon_$fNumInt_$c+_bufchan_buf [0]))
        \go_1Dcon_$fNumInt_$c+_bufchan_buf  <= 1'd0;
      else if (((! es_6_1_argbuf_r) && (! \go_1Dcon_$fNumInt_$c+_bufchan_buf [0])))
        \go_1Dcon_$fNumInt_$c+_bufchan_buf  <= \go_1Dcon_$fNumInt_$c+_bufchan_d ;
  
  /* dcon (Ty MyDTInt_Bool,
      Dcon Dcon_is_z_1) : [(go_2,Go)] > (go_2Dcon_is_z_1,MyDTInt_Bool) */
  assign go_2Dcon_is_z_1_d = Dcon_is_z_1_dc((& {go_2_d[0]}), go_2_d);
  assign {go_2_r} = {1 {(go_2Dcon_is_z_1_r && go_2Dcon_is_z_1_d[0])}};
  
  /* buf (Ty MyDTInt_Bool) : (go_2Dcon_is_z_1,MyDTInt_Bool) > (es_5_1_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t go_2Dcon_is_z_1_bufchan_d;
  logic go_2Dcon_is_z_1_bufchan_r;
  assign go_2Dcon_is_z_1_r = ((! go_2Dcon_is_z_1_bufchan_d[0]) || go_2Dcon_is_z_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_2Dcon_is_z_1_bufchan_d <= 1'd0;
    else
      if (go_2Dcon_is_z_1_r)
        go_2Dcon_is_z_1_bufchan_d <= go_2Dcon_is_z_1_d;
  MyDTInt_Bool_t go_2Dcon_is_z_1_bufchan_buf;
  assign go_2Dcon_is_z_1_bufchan_r = (! go_2Dcon_is_z_1_bufchan_buf[0]);
  assign es_5_1_argbuf_d = (go_2Dcon_is_z_1_bufchan_buf[0] ? go_2Dcon_is_z_1_bufchan_buf :
                            go_2Dcon_is_z_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_2Dcon_is_z_1_bufchan_buf <= 1'd0;
    else
      if ((es_5_1_argbuf_r && go_2Dcon_is_z_1_bufchan_buf[0]))
        go_2Dcon_is_z_1_bufchan_buf <= 1'd0;
      else if (((! es_5_1_argbuf_r) && (! go_2Dcon_is_z_1_bufchan_buf[0])))
        go_2Dcon_is_z_1_bufchan_buf <= go_2Dcon_is_z_1_bufchan_d;
  
  /* dcon (Ty MyDTInt_Int,
      Dcon Dcon_main1) : [(go_3,Go)] > (go_3Dcon_main1,MyDTInt_Int) */
  assign go_3Dcon_main1_d = Dcon_main1_dc((& {go_3_d[0]}), go_3_d);
  assign {go_3_r} = {1 {(go_3Dcon_main1_r && go_3Dcon_main1_d[0])}};
  
  /* buf (Ty MyDTInt_Int) : (go_3Dcon_main1,MyDTInt_Int) > (es_4_1_argbuf,MyDTInt_Int) */
  MyDTInt_Int_t go_3Dcon_main1_bufchan_d;
  logic go_3Dcon_main1_bufchan_r;
  assign go_3Dcon_main1_r = ((! go_3Dcon_main1_bufchan_d[0]) || go_3Dcon_main1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_3Dcon_main1_bufchan_d <= 1'd0;
    else
      if (go_3Dcon_main1_r) go_3Dcon_main1_bufchan_d <= go_3Dcon_main1_d;
  MyDTInt_Int_t go_3Dcon_main1_bufchan_buf;
  assign go_3Dcon_main1_bufchan_r = (! go_3Dcon_main1_bufchan_buf[0]);
  assign es_4_1_argbuf_d = (go_3Dcon_main1_bufchan_buf[0] ? go_3Dcon_main1_bufchan_buf :
                            go_3Dcon_main1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_3Dcon_main1_bufchan_buf <= 1'd0;
    else
      if ((es_4_1_argbuf_r && go_3Dcon_main1_bufchan_buf[0]))
        go_3Dcon_main1_bufchan_buf <= 1'd0;
      else if (((! es_4_1_argbuf_r) && (! go_3Dcon_main1_bufchan_buf[0])))
        go_3Dcon_main1_bufchan_buf <= go_3Dcon_main1_bufchan_d;
  
  /* dcon (Ty MyDTInt_Bool,
      Dcon Dcon_is_z_1) : [(go_4,Go)] > (go_4Dcon_is_z_1,MyDTInt_Bool) */
  assign go_4Dcon_is_z_1_d = Dcon_is_z_1_dc((& {go_4_d[0]}), go_4_d);
  assign {go_4_r} = {1 {(go_4Dcon_is_z_1_r && go_4Dcon_is_z_1_d[0])}};
  
  /* buf (Ty MyDTInt_Bool) : (go_4Dcon_is_z_1,MyDTInt_Bool) > (es_3_1_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t go_4Dcon_is_z_1_bufchan_d;
  logic go_4Dcon_is_z_1_bufchan_r;
  assign go_4Dcon_is_z_1_r = ((! go_4Dcon_is_z_1_bufchan_d[0]) || go_4Dcon_is_z_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_4Dcon_is_z_1_bufchan_d <= 1'd0;
    else
      if (go_4Dcon_is_z_1_r)
        go_4Dcon_is_z_1_bufchan_d <= go_4Dcon_is_z_1_d;
  MyDTInt_Bool_t go_4Dcon_is_z_1_bufchan_buf;
  assign go_4Dcon_is_z_1_bufchan_r = (! go_4Dcon_is_z_1_bufchan_buf[0]);
  assign es_3_1_argbuf_d = (go_4Dcon_is_z_1_bufchan_buf[0] ? go_4Dcon_is_z_1_bufchan_buf :
                            go_4Dcon_is_z_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_4Dcon_is_z_1_bufchan_buf <= 1'd0;
    else
      if ((es_3_1_argbuf_r && go_4Dcon_is_z_1_bufchan_buf[0]))
        go_4Dcon_is_z_1_bufchan_buf <= 1'd0;
      else if (((! es_3_1_argbuf_r) && (! go_4Dcon_is_z_1_bufchan_buf[0])))
        go_4Dcon_is_z_1_bufchan_buf <= go_4Dcon_is_z_1_bufchan_d;
  
  /* buf (Ty Go) : (go_5,Go) > (go_5_argbuf,Go) */
  Go_t go_5_bufchan_d;
  logic go_5_bufchan_r;
  assign go_5_r = ((! go_5_bufchan_d[0]) || go_5_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_5_bufchan_d <= 1'd0;
    else if (go_5_r) go_5_bufchan_d <= go_5_d;
  Go_t go_5_bufchan_buf;
  assign go_5_bufchan_r = (! go_5_bufchan_buf[0]);
  assign go_5_argbuf_d = (go_5_bufchan_buf[0] ? go_5_bufchan_buf :
                          go_5_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_5_bufchan_buf <= 1'd0;
    else
      if ((go_5_argbuf_r && go_5_bufchan_buf[0]))
        go_5_bufchan_buf <= 1'd0;
      else if (((! go_5_argbuf_r) && (! go_5_bufchan_buf[0])))
        go_5_bufchan_buf <= go_5_bufchan_d;
  
  /* dcon (Ty TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int,
      Dcon TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int) : [(go_5_argbuf,Go),
                                                                                                                           (m1aey_0,Pointer_QTree_Int),
                                                                                                                           (m2aez_1,Pointer_QTree_Int),
                                                                                                                           (es_3_1_argbuf,MyDTInt_Bool),
                                                                                                                           (es_4_1_argbuf,MyDTInt_Int),
                                                                                                                           (es_5_1_argbuf,MyDTInt_Bool),
                                                                                                                           (es_6_1_argbuf,MyDTInt_Int_Int)] > (f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int_1,TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int) */
  assign f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_d = TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int_dc((& {go_5_argbuf_d[0],
                                                                                                                                                                                                                                                         m1aey_0_d[0],
                                                                                                                                                                                                                                                         m2aez_1_d[0],
                                                                                                                                                                                                                                                         es_3_1_argbuf_d[0],
                                                                                                                                                                                                                                                         es_4_1_argbuf_d[0],
                                                                                                                                                                                                                                                         es_5_1_argbuf_d[0],
                                                                                                                                                                                                                                                         es_6_1_argbuf_d[0]}), go_5_argbuf_d, m1aey_0_d, m2aez_1_d, es_3_1_argbuf_d, es_4_1_argbuf_d, es_5_1_argbuf_d, es_6_1_argbuf_d);
  assign {go_5_argbuf_r,
          m1aey_0_r,
          m2aez_1_r,
          es_3_1_argbuf_r,
          es_4_1_argbuf_r,
          es_5_1_argbuf_r,
          es_6_1_argbuf_r} = {7 {(f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_r && f_f_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_d[0])}};
  
  /* buf (Ty Go) : (go_6,Go) > (go_6_argbuf,Go) */
  Go_t go_6_bufchan_d;
  logic go_6_bufchan_r;
  assign go_6_r = ((! go_6_bufchan_d[0]) || go_6_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_6_bufchan_d <= 1'd0;
    else if (go_6_r) go_6_bufchan_d <= go_6_d;
  Go_t go_6_bufchan_buf;
  assign go_6_bufchan_r = (! go_6_bufchan_buf[0]);
  assign go_6_argbuf_d = (go_6_bufchan_buf[0] ? go_6_bufchan_buf :
                          go_6_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_6_bufchan_buf <= 1'd0;
    else
      if ((go_6_argbuf_r && go_6_bufchan_buf[0]))
        go_6_bufchan_buf <= 1'd0;
      else if (((! go_6_argbuf_r) && (! go_6_bufchan_buf[0])))
        go_6_bufchan_buf <= go_6_bufchan_d;
  
  /* dcon (Ty TupGo___Pointer_QTree_Int,
      Dcon TupGo___Pointer_QTree_Int) : [(go_6_argbuf,Go),
                                         (es_0_1_argbuf,Pointer_QTree_Int)] > ($wnnzTupGo___Pointer_QTree_Int_1,TupGo___Pointer_QTree_Int) */
  assign \$wnnzTupGo___Pointer_QTree_Int_1_d  = TupGo___Pointer_QTree_Int_dc((& {go_6_argbuf_d[0],
                                                                                 es_0_1_argbuf_d[0]}), go_6_argbuf_d, es_0_1_argbuf_d);
  assign {go_6_argbuf_r,
          es_0_1_argbuf_r} = {2 {(\$wnnzTupGo___Pointer_QTree_Int_1_r  && \$wnnzTupGo___Pointer_QTree_Int_1_d [0])}};
  
  /* dcon (Ty CT$wnnz,
      Dcon L$wnnzsbos) : [(go_7_1,Go)] > (go_7_1L$wnnzsbos,CT$wnnz) */
  assign go_7_1L$wnnzsbos_d = L$wnnzsbos_dc((& {go_7_1_d[0]}), go_7_1_d);
  assign {go_7_1_r} = {1 {(go_7_1L$wnnzsbos_r && go_7_1L$wnnzsbos_d[0])}};
  
  /* buf (Ty CT$wnnz) : (go_7_1L$wnnzsbos,CT$wnnz) > (lizzieLet0_1_argbuf,CT$wnnz) */
  CT$wnnz_t go_7_1L$wnnzsbos_bufchan_d;
  logic go_7_1L$wnnzsbos_bufchan_r;
  assign go_7_1L$wnnzsbos_r = ((! go_7_1L$wnnzsbos_bufchan_d[0]) || go_7_1L$wnnzsbos_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_7_1L$wnnzsbos_bufchan_d <= {115'd0, 1'd0};
    else
      if (go_7_1L$wnnzsbos_r)
        go_7_1L$wnnzsbos_bufchan_d <= go_7_1L$wnnzsbos_d;
  CT$wnnz_t go_7_1L$wnnzsbos_bufchan_buf;
  assign go_7_1L$wnnzsbos_bufchan_r = (! go_7_1L$wnnzsbos_bufchan_buf[0]);
  assign lizzieLet0_1_argbuf_d = (go_7_1L$wnnzsbos_bufchan_buf[0] ? go_7_1L$wnnzsbos_bufchan_buf :
                                  go_7_1L$wnnzsbos_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      go_7_1L$wnnzsbos_bufchan_buf <= {115'd0, 1'd0};
    else
      if ((lizzieLet0_1_argbuf_r && go_7_1L$wnnzsbos_bufchan_buf[0]))
        go_7_1L$wnnzsbos_bufchan_buf <= {115'd0, 1'd0};
      else if (((! lizzieLet0_1_argbuf_r) && (! go_7_1L$wnnzsbos_bufchan_buf[0])))
        go_7_1L$wnnzsbos_bufchan_buf <= go_7_1L$wnnzsbos_bufchan_d;
  
  /* buf (Ty Go) : (go_7_2,Go) > (go_7_2_argbuf,Go) */
  Go_t go_7_2_bufchan_d;
  logic go_7_2_bufchan_r;
  assign go_7_2_r = ((! go_7_2_bufchan_d[0]) || go_7_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_7_2_bufchan_d <= 1'd0;
    else if (go_7_2_r) go_7_2_bufchan_d <= go_7_2_d;
  Go_t go_7_2_bufchan_buf;
  assign go_7_2_bufchan_r = (! go_7_2_bufchan_buf[0]);
  assign go_7_2_argbuf_d = (go_7_2_bufchan_buf[0] ? go_7_2_bufchan_buf :
                            go_7_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_7_2_bufchan_buf <= 1'd0;
    else
      if ((go_7_2_argbuf_r && go_7_2_bufchan_buf[0]))
        go_7_2_bufchan_buf <= 1'd0;
      else if (((! go_7_2_argbuf_r) && (! go_7_2_bufchan_buf[0])))
        go_7_2_bufchan_buf <= go_7_2_bufchan_d;
  
  /* dcon (Ty TupGo___Pointer_QTree_Int___Pointer_CT$wnnz,
      Dcon TupGo___Pointer_QTree_Int___Pointer_CT$wnnz) : [(go_7_2_argbuf,Go),
                                                           (wsiX_1_argbuf,Pointer_QTree_Int),
                                                           (lizzieLet25_1_argbuf,Pointer_CT$wnnz)] > (call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_1,TupGo___Pointer_QTree_Int___Pointer_CT$wnnz) */
  assign call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_1_d = TupGo___Pointer_QTree_Int___Pointer_CT$wnnz_dc((& {go_7_2_argbuf_d[0],
                                                                                                                        wsiX_1_argbuf_d[0],
                                                                                                                        lizzieLet25_1_argbuf_d[0]}), go_7_2_argbuf_d, wsiX_1_argbuf_d, lizzieLet25_1_argbuf_d);
  assign {go_7_2_argbuf_r,
          wsiX_1_argbuf_r,
          lizzieLet25_1_argbuf_r} = {3 {(call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_1_r && call_$wnnzTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_1_d[0])}};
  
  /* buf (Ty MyDTInt_Bool) : (is_z_adda8G_2_2,MyDTInt_Bool) > (is_z_adda8G_2_2_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t is_z_adda8G_2_2_bufchan_d;
  logic is_z_adda8G_2_2_bufchan_r;
  assign is_z_adda8G_2_2_r = ((! is_z_adda8G_2_2_bufchan_d[0]) || is_z_adda8G_2_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) is_z_adda8G_2_2_bufchan_d <= 1'd0;
    else
      if (is_z_adda8G_2_2_r)
        is_z_adda8G_2_2_bufchan_d <= is_z_adda8G_2_2_d;
  MyDTInt_Bool_t is_z_adda8G_2_2_bufchan_buf;
  assign is_z_adda8G_2_2_bufchan_r = (! is_z_adda8G_2_2_bufchan_buf[0]);
  assign is_z_adda8G_2_2_argbuf_d = (is_z_adda8G_2_2_bufchan_buf[0] ? is_z_adda8G_2_2_bufchan_buf :
                                     is_z_adda8G_2_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) is_z_adda8G_2_2_bufchan_buf <= 1'd0;
    else
      if ((is_z_adda8G_2_2_argbuf_r && is_z_adda8G_2_2_bufchan_buf[0]))
        is_z_adda8G_2_2_bufchan_buf <= 1'd0;
      else if (((! is_z_adda8G_2_2_argbuf_r) && (! is_z_adda8G_2_2_bufchan_buf[0])))
        is_z_adda8G_2_2_bufchan_buf <= is_z_adda8G_2_2_bufchan_d;
  
  /* fork (Ty MyDTInt_Bool) : (is_z_adda8G_2_destruct,MyDTInt_Bool) > [(is_z_adda8G_2_1,MyDTInt_Bool),
                                                                  (is_z_adda8G_2_2,MyDTInt_Bool)] */
  logic [1:0] is_z_adda8G_2_destruct_emitted;
  logic [1:0] is_z_adda8G_2_destruct_done;
  assign is_z_adda8G_2_1_d = (is_z_adda8G_2_destruct_d[0] && (! is_z_adda8G_2_destruct_emitted[0]));
  assign is_z_adda8G_2_2_d = (is_z_adda8G_2_destruct_d[0] && (! is_z_adda8G_2_destruct_emitted[1]));
  assign is_z_adda8G_2_destruct_done = (is_z_adda8G_2_destruct_emitted | ({is_z_adda8G_2_2_d[0],
                                                                           is_z_adda8G_2_1_d[0]} & {is_z_adda8G_2_2_r,
                                                                                                    is_z_adda8G_2_1_r}));
  assign is_z_adda8G_2_destruct_r = (& is_z_adda8G_2_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) is_z_adda8G_2_destruct_emitted <= 2'd0;
    else
      is_z_adda8G_2_destruct_emitted <= (is_z_adda8G_2_destruct_r ? 2'd0 :
                                         is_z_adda8G_2_destruct_done);
  
  /* buf (Ty MyDTInt_Bool) : (is_z_adda8G_3_2,MyDTInt_Bool) > (is_z_adda8G_3_2_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t is_z_adda8G_3_2_bufchan_d;
  logic is_z_adda8G_3_2_bufchan_r;
  assign is_z_adda8G_3_2_r = ((! is_z_adda8G_3_2_bufchan_d[0]) || is_z_adda8G_3_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) is_z_adda8G_3_2_bufchan_d <= 1'd0;
    else
      if (is_z_adda8G_3_2_r)
        is_z_adda8G_3_2_bufchan_d <= is_z_adda8G_3_2_d;
  MyDTInt_Bool_t is_z_adda8G_3_2_bufchan_buf;
  assign is_z_adda8G_3_2_bufchan_r = (! is_z_adda8G_3_2_bufchan_buf[0]);
  assign is_z_adda8G_3_2_argbuf_d = (is_z_adda8G_3_2_bufchan_buf[0] ? is_z_adda8G_3_2_bufchan_buf :
                                     is_z_adda8G_3_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) is_z_adda8G_3_2_bufchan_buf <= 1'd0;
    else
      if ((is_z_adda8G_3_2_argbuf_r && is_z_adda8G_3_2_bufchan_buf[0]))
        is_z_adda8G_3_2_bufchan_buf <= 1'd0;
      else if (((! is_z_adda8G_3_2_argbuf_r) && (! is_z_adda8G_3_2_bufchan_buf[0])))
        is_z_adda8G_3_2_bufchan_buf <= is_z_adda8G_3_2_bufchan_d;
  
  /* fork (Ty MyDTInt_Bool) : (is_z_adda8G_3_destruct,MyDTInt_Bool) > [(is_z_adda8G_3_1,MyDTInt_Bool),
                                                                  (is_z_adda8G_3_2,MyDTInt_Bool)] */
  logic [1:0] is_z_adda8G_3_destruct_emitted;
  logic [1:0] is_z_adda8G_3_destruct_done;
  assign is_z_adda8G_3_1_d = (is_z_adda8G_3_destruct_d[0] && (! is_z_adda8G_3_destruct_emitted[0]));
  assign is_z_adda8G_3_2_d = (is_z_adda8G_3_destruct_d[0] && (! is_z_adda8G_3_destruct_emitted[1]));
  assign is_z_adda8G_3_destruct_done = (is_z_adda8G_3_destruct_emitted | ({is_z_adda8G_3_2_d[0],
                                                                           is_z_adda8G_3_1_d[0]} & {is_z_adda8G_3_2_r,
                                                                                                    is_z_adda8G_3_1_r}));
  assign is_z_adda8G_3_destruct_r = (& is_z_adda8G_3_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) is_z_adda8G_3_destruct_emitted <= 2'd0;
    else
      is_z_adda8G_3_destruct_emitted <= (is_z_adda8G_3_destruct_r ? 2'd0 :
                                         is_z_adda8G_3_destruct_done);
  
  /* buf (Ty MyDTInt_Bool) : (is_z_adda8G_4_destruct,MyDTInt_Bool) > (is_z_adda8G_4_1_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t is_z_adda8G_4_destruct_bufchan_d;
  logic is_z_adda8G_4_destruct_bufchan_r;
  assign is_z_adda8G_4_destruct_r = ((! is_z_adda8G_4_destruct_bufchan_d[0]) || is_z_adda8G_4_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) is_z_adda8G_4_destruct_bufchan_d <= 1'd0;
    else
      if (is_z_adda8G_4_destruct_r)
        is_z_adda8G_4_destruct_bufchan_d <= is_z_adda8G_4_destruct_d;
  MyDTInt_Bool_t is_z_adda8G_4_destruct_bufchan_buf;
  assign is_z_adda8G_4_destruct_bufchan_r = (! is_z_adda8G_4_destruct_bufchan_buf[0]);
  assign is_z_adda8G_4_1_argbuf_d = (is_z_adda8G_4_destruct_bufchan_buf[0] ? is_z_adda8G_4_destruct_bufchan_buf :
                                     is_z_adda8G_4_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) is_z_adda8G_4_destruct_bufchan_buf <= 1'd0;
    else
      if ((is_z_adda8G_4_1_argbuf_r && is_z_adda8G_4_destruct_bufchan_buf[0]))
        is_z_adda8G_4_destruct_bufchan_buf <= 1'd0;
      else if (((! is_z_adda8G_4_1_argbuf_r) && (! is_z_adda8G_4_destruct_bufchan_buf[0])))
        is_z_adda8G_4_destruct_bufchan_buf <= is_z_adda8G_4_destruct_bufchan_d;
  
  /* buf (Ty MyDTInt_Bool) : (is_z_mapa8E_2_2,MyDTInt_Bool) > (is_z_mapa8E_2_2_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t is_z_mapa8E_2_2_bufchan_d;
  logic is_z_mapa8E_2_2_bufchan_r;
  assign is_z_mapa8E_2_2_r = ((! is_z_mapa8E_2_2_bufchan_d[0]) || is_z_mapa8E_2_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) is_z_mapa8E_2_2_bufchan_d <= 1'd0;
    else
      if (is_z_mapa8E_2_2_r)
        is_z_mapa8E_2_2_bufchan_d <= is_z_mapa8E_2_2_d;
  MyDTInt_Bool_t is_z_mapa8E_2_2_bufchan_buf;
  assign is_z_mapa8E_2_2_bufchan_r = (! is_z_mapa8E_2_2_bufchan_buf[0]);
  assign is_z_mapa8E_2_2_argbuf_d = (is_z_mapa8E_2_2_bufchan_buf[0] ? is_z_mapa8E_2_2_bufchan_buf :
                                     is_z_mapa8E_2_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) is_z_mapa8E_2_2_bufchan_buf <= 1'd0;
    else
      if ((is_z_mapa8E_2_2_argbuf_r && is_z_mapa8E_2_2_bufchan_buf[0]))
        is_z_mapa8E_2_2_bufchan_buf <= 1'd0;
      else if (((! is_z_mapa8E_2_2_argbuf_r) && (! is_z_mapa8E_2_2_bufchan_buf[0])))
        is_z_mapa8E_2_2_bufchan_buf <= is_z_mapa8E_2_2_bufchan_d;
  
  /* fork (Ty MyDTInt_Bool) : (is_z_mapa8E_2_destruct,MyDTInt_Bool) > [(is_z_mapa8E_2_1,MyDTInt_Bool),
                                                                  (is_z_mapa8E_2_2,MyDTInt_Bool)] */
  logic [1:0] is_z_mapa8E_2_destruct_emitted;
  logic [1:0] is_z_mapa8E_2_destruct_done;
  assign is_z_mapa8E_2_1_d = (is_z_mapa8E_2_destruct_d[0] && (! is_z_mapa8E_2_destruct_emitted[0]));
  assign is_z_mapa8E_2_2_d = (is_z_mapa8E_2_destruct_d[0] && (! is_z_mapa8E_2_destruct_emitted[1]));
  assign is_z_mapa8E_2_destruct_done = (is_z_mapa8E_2_destruct_emitted | ({is_z_mapa8E_2_2_d[0],
                                                                           is_z_mapa8E_2_1_d[0]} & {is_z_mapa8E_2_2_r,
                                                                                                    is_z_mapa8E_2_1_r}));
  assign is_z_mapa8E_2_destruct_r = (& is_z_mapa8E_2_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) is_z_mapa8E_2_destruct_emitted <= 2'd0;
    else
      is_z_mapa8E_2_destruct_emitted <= (is_z_mapa8E_2_destruct_r ? 2'd0 :
                                         is_z_mapa8E_2_destruct_done);
  
  /* buf (Ty MyDTInt_Bool) : (is_z_mapa8E_3_2,MyDTInt_Bool) > (is_z_mapa8E_3_2_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t is_z_mapa8E_3_2_bufchan_d;
  logic is_z_mapa8E_3_2_bufchan_r;
  assign is_z_mapa8E_3_2_r = ((! is_z_mapa8E_3_2_bufchan_d[0]) || is_z_mapa8E_3_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) is_z_mapa8E_3_2_bufchan_d <= 1'd0;
    else
      if (is_z_mapa8E_3_2_r)
        is_z_mapa8E_3_2_bufchan_d <= is_z_mapa8E_3_2_d;
  MyDTInt_Bool_t is_z_mapa8E_3_2_bufchan_buf;
  assign is_z_mapa8E_3_2_bufchan_r = (! is_z_mapa8E_3_2_bufchan_buf[0]);
  assign is_z_mapa8E_3_2_argbuf_d = (is_z_mapa8E_3_2_bufchan_buf[0] ? is_z_mapa8E_3_2_bufchan_buf :
                                     is_z_mapa8E_3_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) is_z_mapa8E_3_2_bufchan_buf <= 1'd0;
    else
      if ((is_z_mapa8E_3_2_argbuf_r && is_z_mapa8E_3_2_bufchan_buf[0]))
        is_z_mapa8E_3_2_bufchan_buf <= 1'd0;
      else if (((! is_z_mapa8E_3_2_argbuf_r) && (! is_z_mapa8E_3_2_bufchan_buf[0])))
        is_z_mapa8E_3_2_bufchan_buf <= is_z_mapa8E_3_2_bufchan_d;
  
  /* fork (Ty MyDTInt_Bool) : (is_z_mapa8E_3_destruct,MyDTInt_Bool) > [(is_z_mapa8E_3_1,MyDTInt_Bool),
                                                                  (is_z_mapa8E_3_2,MyDTInt_Bool)] */
  logic [1:0] is_z_mapa8E_3_destruct_emitted;
  logic [1:0] is_z_mapa8E_3_destruct_done;
  assign is_z_mapa8E_3_1_d = (is_z_mapa8E_3_destruct_d[0] && (! is_z_mapa8E_3_destruct_emitted[0]));
  assign is_z_mapa8E_3_2_d = (is_z_mapa8E_3_destruct_d[0] && (! is_z_mapa8E_3_destruct_emitted[1]));
  assign is_z_mapa8E_3_destruct_done = (is_z_mapa8E_3_destruct_emitted | ({is_z_mapa8E_3_2_d[0],
                                                                           is_z_mapa8E_3_1_d[0]} & {is_z_mapa8E_3_2_r,
                                                                                                    is_z_mapa8E_3_1_r}));
  assign is_z_mapa8E_3_destruct_r = (& is_z_mapa8E_3_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) is_z_mapa8E_3_destruct_emitted <= 2'd0;
    else
      is_z_mapa8E_3_destruct_emitted <= (is_z_mapa8E_3_destruct_r ? 2'd0 :
                                         is_z_mapa8E_3_destruct_done);
  
  /* buf (Ty MyDTInt_Bool) : (is_z_mapa8E_4_destruct,MyDTInt_Bool) > (is_z_mapa8E_4_1_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t is_z_mapa8E_4_destruct_bufchan_d;
  logic is_z_mapa8E_4_destruct_bufchan_r;
  assign is_z_mapa8E_4_destruct_r = ((! is_z_mapa8E_4_destruct_bufchan_d[0]) || is_z_mapa8E_4_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) is_z_mapa8E_4_destruct_bufchan_d <= 1'd0;
    else
      if (is_z_mapa8E_4_destruct_r)
        is_z_mapa8E_4_destruct_bufchan_d <= is_z_mapa8E_4_destruct_d;
  MyDTInt_Bool_t is_z_mapa8E_4_destruct_bufchan_buf;
  assign is_z_mapa8E_4_destruct_bufchan_r = (! is_z_mapa8E_4_destruct_bufchan_buf[0]);
  assign is_z_mapa8E_4_1_argbuf_d = (is_z_mapa8E_4_destruct_bufchan_buf[0] ? is_z_mapa8E_4_destruct_bufchan_buf :
                                     is_z_mapa8E_4_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) is_z_mapa8E_4_destruct_bufchan_buf <= 1'd0;
    else
      if ((is_z_mapa8E_4_1_argbuf_r && is_z_mapa8E_4_destruct_bufchan_buf[0]))
        is_z_mapa8E_4_destruct_bufchan_buf <= 1'd0;
      else if (((! is_z_mapa8E_4_1_argbuf_r) && (! is_z_mapa8E_4_destruct_bufchan_buf[0])))
        is_z_mapa8E_4_destruct_bufchan_buf <= is_z_mapa8E_4_destruct_bufchan_d;
  
  /* buf (Ty MyDTInt_Bool) : (is_z_mapa8v_2_2,MyDTInt_Bool) > (is_z_mapa8v_2_2_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t is_z_mapa8v_2_2_bufchan_d;
  logic is_z_mapa8v_2_2_bufchan_r;
  assign is_z_mapa8v_2_2_r = ((! is_z_mapa8v_2_2_bufchan_d[0]) || is_z_mapa8v_2_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) is_z_mapa8v_2_2_bufchan_d <= 1'd0;
    else
      if (is_z_mapa8v_2_2_r)
        is_z_mapa8v_2_2_bufchan_d <= is_z_mapa8v_2_2_d;
  MyDTInt_Bool_t is_z_mapa8v_2_2_bufchan_buf;
  assign is_z_mapa8v_2_2_bufchan_r = (! is_z_mapa8v_2_2_bufchan_buf[0]);
  assign is_z_mapa8v_2_2_argbuf_d = (is_z_mapa8v_2_2_bufchan_buf[0] ? is_z_mapa8v_2_2_bufchan_buf :
                                     is_z_mapa8v_2_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) is_z_mapa8v_2_2_bufchan_buf <= 1'd0;
    else
      if ((is_z_mapa8v_2_2_argbuf_r && is_z_mapa8v_2_2_bufchan_buf[0]))
        is_z_mapa8v_2_2_bufchan_buf <= 1'd0;
      else if (((! is_z_mapa8v_2_2_argbuf_r) && (! is_z_mapa8v_2_2_bufchan_buf[0])))
        is_z_mapa8v_2_2_bufchan_buf <= is_z_mapa8v_2_2_bufchan_d;
  
  /* fork (Ty MyDTInt_Bool) : (is_z_mapa8v_2_destruct,MyDTInt_Bool) > [(is_z_mapa8v_2_1,MyDTInt_Bool),
                                                                  (is_z_mapa8v_2_2,MyDTInt_Bool)] */
  logic [1:0] is_z_mapa8v_2_destruct_emitted;
  logic [1:0] is_z_mapa8v_2_destruct_done;
  assign is_z_mapa8v_2_1_d = (is_z_mapa8v_2_destruct_d[0] && (! is_z_mapa8v_2_destruct_emitted[0]));
  assign is_z_mapa8v_2_2_d = (is_z_mapa8v_2_destruct_d[0] && (! is_z_mapa8v_2_destruct_emitted[1]));
  assign is_z_mapa8v_2_destruct_done = (is_z_mapa8v_2_destruct_emitted | ({is_z_mapa8v_2_2_d[0],
                                                                           is_z_mapa8v_2_1_d[0]} & {is_z_mapa8v_2_2_r,
                                                                                                    is_z_mapa8v_2_1_r}));
  assign is_z_mapa8v_2_destruct_r = (& is_z_mapa8v_2_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) is_z_mapa8v_2_destruct_emitted <= 2'd0;
    else
      is_z_mapa8v_2_destruct_emitted <= (is_z_mapa8v_2_destruct_r ? 2'd0 :
                                         is_z_mapa8v_2_destruct_done);
  
  /* buf (Ty MyDTInt_Bool) : (is_z_mapa8v_3_2,MyDTInt_Bool) > (is_z_mapa8v_3_2_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t is_z_mapa8v_3_2_bufchan_d;
  logic is_z_mapa8v_3_2_bufchan_r;
  assign is_z_mapa8v_3_2_r = ((! is_z_mapa8v_3_2_bufchan_d[0]) || is_z_mapa8v_3_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) is_z_mapa8v_3_2_bufchan_d <= 1'd0;
    else
      if (is_z_mapa8v_3_2_r)
        is_z_mapa8v_3_2_bufchan_d <= is_z_mapa8v_3_2_d;
  MyDTInt_Bool_t is_z_mapa8v_3_2_bufchan_buf;
  assign is_z_mapa8v_3_2_bufchan_r = (! is_z_mapa8v_3_2_bufchan_buf[0]);
  assign is_z_mapa8v_3_2_argbuf_d = (is_z_mapa8v_3_2_bufchan_buf[0] ? is_z_mapa8v_3_2_bufchan_buf :
                                     is_z_mapa8v_3_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) is_z_mapa8v_3_2_bufchan_buf <= 1'd0;
    else
      if ((is_z_mapa8v_3_2_argbuf_r && is_z_mapa8v_3_2_bufchan_buf[0]))
        is_z_mapa8v_3_2_bufchan_buf <= 1'd0;
      else if (((! is_z_mapa8v_3_2_argbuf_r) && (! is_z_mapa8v_3_2_bufchan_buf[0])))
        is_z_mapa8v_3_2_bufchan_buf <= is_z_mapa8v_3_2_bufchan_d;
  
  /* fork (Ty MyDTInt_Bool) : (is_z_mapa8v_3_destruct,MyDTInt_Bool) > [(is_z_mapa8v_3_1,MyDTInt_Bool),
                                                                  (is_z_mapa8v_3_2,MyDTInt_Bool)] */
  logic [1:0] is_z_mapa8v_3_destruct_emitted;
  logic [1:0] is_z_mapa8v_3_destruct_done;
  assign is_z_mapa8v_3_1_d = (is_z_mapa8v_3_destruct_d[0] && (! is_z_mapa8v_3_destruct_emitted[0]));
  assign is_z_mapa8v_3_2_d = (is_z_mapa8v_3_destruct_d[0] && (! is_z_mapa8v_3_destruct_emitted[1]));
  assign is_z_mapa8v_3_destruct_done = (is_z_mapa8v_3_destruct_emitted | ({is_z_mapa8v_3_2_d[0],
                                                                           is_z_mapa8v_3_1_d[0]} & {is_z_mapa8v_3_2_r,
                                                                                                    is_z_mapa8v_3_1_r}));
  assign is_z_mapa8v_3_destruct_r = (& is_z_mapa8v_3_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) is_z_mapa8v_3_destruct_emitted <= 2'd0;
    else
      is_z_mapa8v_3_destruct_emitted <= (is_z_mapa8v_3_destruct_r ? 2'd0 :
                                         is_z_mapa8v_3_destruct_done);
  
  /* buf (Ty MyDTInt_Bool) : (is_z_mapa8v_4_destruct,MyDTInt_Bool) > (is_z_mapa8v_4_1_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t is_z_mapa8v_4_destruct_bufchan_d;
  logic is_z_mapa8v_4_destruct_bufchan_r;
  assign is_z_mapa8v_4_destruct_r = ((! is_z_mapa8v_4_destruct_bufchan_d[0]) || is_z_mapa8v_4_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) is_z_mapa8v_4_destruct_bufchan_d <= 1'd0;
    else
      if (is_z_mapa8v_4_destruct_r)
        is_z_mapa8v_4_destruct_bufchan_d <= is_z_mapa8v_4_destruct_d;
  MyDTInt_Bool_t is_z_mapa8v_4_destruct_bufchan_buf;
  assign is_z_mapa8v_4_destruct_bufchan_r = (! is_z_mapa8v_4_destruct_bufchan_buf[0]);
  assign is_z_mapa8v_4_1_argbuf_d = (is_z_mapa8v_4_destruct_bufchan_buf[0] ? is_z_mapa8v_4_destruct_bufchan_buf :
                                     is_z_mapa8v_4_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) is_z_mapa8v_4_destruct_bufchan_buf <= 1'd0;
    else
      if ((is_z_mapa8v_4_1_argbuf_r && is_z_mapa8v_4_destruct_bufchan_buf[0]))
        is_z_mapa8v_4_destruct_bufchan_buf <= 1'd0;
      else if (((! is_z_mapa8v_4_1_argbuf_r) && (! is_z_mapa8v_4_destruct_bufchan_buf[0])))
        is_z_mapa8v_4_destruct_bufchan_buf <= is_z_mapa8v_4_destruct_bufchan_d;
  
  /* destruct (Ty QTree_Int,
          Dcon QNode_Int) : (lizzieLet12_1QNode_Int,QTree_Int) > [(q1a8T_destruct,Pointer_QTree_Int),
                                                                  (q2a8U_destruct,Pointer_QTree_Int),
                                                                  (q3a8V_destruct,Pointer_QTree_Int),
                                                                  (q4a8W_destruct,Pointer_QTree_Int)] */
  logic [3:0] lizzieLet12_1QNode_Int_emitted;
  logic [3:0] lizzieLet12_1QNode_Int_done;
  assign q1a8T_destruct_d = {lizzieLet12_1QNode_Int_d[18:3],
                             (lizzieLet12_1QNode_Int_d[0] && (! lizzieLet12_1QNode_Int_emitted[0]))};
  assign q2a8U_destruct_d = {lizzieLet12_1QNode_Int_d[34:19],
                             (lizzieLet12_1QNode_Int_d[0] && (! lizzieLet12_1QNode_Int_emitted[1]))};
  assign q3a8V_destruct_d = {lizzieLet12_1QNode_Int_d[50:35],
                             (lizzieLet12_1QNode_Int_d[0] && (! lizzieLet12_1QNode_Int_emitted[2]))};
  assign q4a8W_destruct_d = {lizzieLet12_1QNode_Int_d[66:51],
                             (lizzieLet12_1QNode_Int_d[0] && (! lizzieLet12_1QNode_Int_emitted[3]))};
  assign lizzieLet12_1QNode_Int_done = (lizzieLet12_1QNode_Int_emitted | ({q4a8W_destruct_d[0],
                                                                           q3a8V_destruct_d[0],
                                                                           q2a8U_destruct_d[0],
                                                                           q1a8T_destruct_d[0]} & {q4a8W_destruct_r,
                                                                                                   q3a8V_destruct_r,
                                                                                                   q2a8U_destruct_r,
                                                                                                   q1a8T_destruct_r}));
  assign lizzieLet12_1QNode_Int_r = (& lizzieLet12_1QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet12_1QNode_Int_emitted <= 4'd0;
    else
      lizzieLet12_1QNode_Int_emitted <= (lizzieLet12_1QNode_Int_r ? 4'd0 :
                                         lizzieLet12_1QNode_Int_done);
  
  /* destruct (Ty QTree_Int,
          Dcon QVal_Int) : (lizzieLet12_1QVal_Int,QTree_Int) > [(v1a8N_destruct,Int)] */
  assign v1a8N_destruct_d = {lizzieLet12_1QVal_Int_d[34:3],
                             lizzieLet12_1QVal_Int_d[0]};
  assign lizzieLet12_1QVal_Int_r = v1a8N_destruct_r;
  
  /* demux (Ty QTree_Int,
       Ty QTree_Int) : (lizzieLet12_2,QTree_Int) (lizzieLet12_1,QTree_Int) > [(_65,QTree_Int),
                                                                              (lizzieLet12_1QVal_Int,QTree_Int),
                                                                              (lizzieLet12_1QNode_Int,QTree_Int),
                                                                              (_64,QTree_Int)] */
  logic [3:0] lizzieLet12_1_onehotd;
  always_comb
    if ((lizzieLet12_2_d[0] && lizzieLet12_1_d[0]))
      unique case (lizzieLet12_2_d[2:1])
        2'd0: lizzieLet12_1_onehotd = 4'd1;
        2'd1: lizzieLet12_1_onehotd = 4'd2;
        2'd2: lizzieLet12_1_onehotd = 4'd4;
        2'd3: lizzieLet12_1_onehotd = 4'd8;
        default: lizzieLet12_1_onehotd = 4'd0;
      endcase
    else lizzieLet12_1_onehotd = 4'd0;
  assign _65_d = {lizzieLet12_1_d[66:1], lizzieLet12_1_onehotd[0]};
  assign lizzieLet12_1QVal_Int_d = {lizzieLet12_1_d[66:1],
                                    lizzieLet12_1_onehotd[1]};
  assign lizzieLet12_1QNode_Int_d = {lizzieLet12_1_d[66:1],
                                     lizzieLet12_1_onehotd[2]};
  assign _64_d = {lizzieLet12_1_d[66:1], lizzieLet12_1_onehotd[3]};
  assign lizzieLet12_1_r = (| (lizzieLet12_1_onehotd & {_64_r,
                                                        lizzieLet12_1QNode_Int_r,
                                                        lizzieLet12_1QVal_Int_r,
                                                        _65_r}));
  assign lizzieLet12_2_r = lizzieLet12_1_r;
  
  /* demux (Ty QTree_Int,
       Ty Go) : (lizzieLet12_3,QTree_Int) (go_12_goMux_data,Go) > [(lizzieLet12_3QNone_Int,Go),
                                                                   (lizzieLet12_3QVal_Int,Go),
                                                                   (lizzieLet12_3QNode_Int,Go),
                                                                   (lizzieLet12_3QError_Int,Go)] */
  logic [3:0] go_12_goMux_data_onehotd;
  always_comb
    if ((lizzieLet12_3_d[0] && go_12_goMux_data_d[0]))
      unique case (lizzieLet12_3_d[2:1])
        2'd0: go_12_goMux_data_onehotd = 4'd1;
        2'd1: go_12_goMux_data_onehotd = 4'd2;
        2'd2: go_12_goMux_data_onehotd = 4'd4;
        2'd3: go_12_goMux_data_onehotd = 4'd8;
        default: go_12_goMux_data_onehotd = 4'd0;
      endcase
    else go_12_goMux_data_onehotd = 4'd0;
  assign lizzieLet12_3QNone_Int_d = go_12_goMux_data_onehotd[0];
  assign lizzieLet12_3QVal_Int_d = go_12_goMux_data_onehotd[1];
  assign lizzieLet12_3QNode_Int_d = go_12_goMux_data_onehotd[2];
  assign lizzieLet12_3QError_Int_d = go_12_goMux_data_onehotd[3];
  assign go_12_goMux_data_r = (| (go_12_goMux_data_onehotd & {lizzieLet12_3QError_Int_r,
                                                              lizzieLet12_3QNode_Int_r,
                                                              lizzieLet12_3QVal_Int_r,
                                                              lizzieLet12_3QNone_Int_r}));
  assign lizzieLet12_3_r = go_12_goMux_data_r;
  
  /* fork (Ty Go) : (lizzieLet12_3QError_Int,Go) > [(lizzieLet12_3QError_Int_1,Go),
                                               (lizzieLet12_3QError_Int_2,Go)] */
  logic [1:0] lizzieLet12_3QError_Int_emitted;
  logic [1:0] lizzieLet12_3QError_Int_done;
  assign lizzieLet12_3QError_Int_1_d = (lizzieLet12_3QError_Int_d[0] && (! lizzieLet12_3QError_Int_emitted[0]));
  assign lizzieLet12_3QError_Int_2_d = (lizzieLet12_3QError_Int_d[0] && (! lizzieLet12_3QError_Int_emitted[1]));
  assign lizzieLet12_3QError_Int_done = (lizzieLet12_3QError_Int_emitted | ({lizzieLet12_3QError_Int_2_d[0],
                                                                             lizzieLet12_3QError_Int_1_d[0]} & {lizzieLet12_3QError_Int_2_r,
                                                                                                                lizzieLet12_3QError_Int_1_r}));
  assign lizzieLet12_3QError_Int_r = (& lizzieLet12_3QError_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet12_3QError_Int_emitted <= 2'd0;
    else
      lizzieLet12_3QError_Int_emitted <= (lizzieLet12_3QError_Int_r ? 2'd0 :
                                          lizzieLet12_3QError_Int_done);
  
  /* dcon (Ty QTree_Int,
      Dcon QError_Int) : [(lizzieLet12_3QError_Int_1,Go)] > (lizzieLet12_3QError_Int_1QError_Int,QTree_Int) */
  assign lizzieLet12_3QError_Int_1QError_Int_d = QError_Int_dc((& {lizzieLet12_3QError_Int_1_d[0]}), lizzieLet12_3QError_Int_1_d);
  assign {lizzieLet12_3QError_Int_1_r} = {1 {(lizzieLet12_3QError_Int_1QError_Int_r && lizzieLet12_3QError_Int_1QError_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (lizzieLet12_3QError_Int_1QError_Int,QTree_Int) > (lizzieLet32_1_argbuf,QTree_Int) */
  QTree_Int_t lizzieLet12_3QError_Int_1QError_Int_bufchan_d;
  logic lizzieLet12_3QError_Int_1QError_Int_bufchan_r;
  assign lizzieLet12_3QError_Int_1QError_Int_r = ((! lizzieLet12_3QError_Int_1QError_Int_bufchan_d[0]) || lizzieLet12_3QError_Int_1QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_3QError_Int_1QError_Int_bufchan_d <= {66'd0, 1'd0};
    else
      if (lizzieLet12_3QError_Int_1QError_Int_r)
        lizzieLet12_3QError_Int_1QError_Int_bufchan_d <= lizzieLet12_3QError_Int_1QError_Int_d;
  QTree_Int_t lizzieLet12_3QError_Int_1QError_Int_bufchan_buf;
  assign lizzieLet12_3QError_Int_1QError_Int_bufchan_r = (! lizzieLet12_3QError_Int_1QError_Int_bufchan_buf[0]);
  assign lizzieLet32_1_argbuf_d = (lizzieLet12_3QError_Int_1QError_Int_bufchan_buf[0] ? lizzieLet12_3QError_Int_1QError_Int_bufchan_buf :
                                   lizzieLet12_3QError_Int_1QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_3QError_Int_1QError_Int_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((lizzieLet32_1_argbuf_r && lizzieLet12_3QError_Int_1QError_Int_bufchan_buf[0]))
        lizzieLet12_3QError_Int_1QError_Int_bufchan_buf <= {66'd0, 1'd0};
      else if (((! lizzieLet32_1_argbuf_r) && (! lizzieLet12_3QError_Int_1QError_Int_bufchan_buf[0])))
        lizzieLet12_3QError_Int_1QError_Int_bufchan_buf <= lizzieLet12_3QError_Int_1QError_Int_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet12_3QError_Int_2,Go) > (lizzieLet12_3QError_Int_2_argbuf,Go) */
  Go_t lizzieLet12_3QError_Int_2_bufchan_d;
  logic lizzieLet12_3QError_Int_2_bufchan_r;
  assign lizzieLet12_3QError_Int_2_r = ((! lizzieLet12_3QError_Int_2_bufchan_d[0]) || lizzieLet12_3QError_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet12_3QError_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet12_3QError_Int_2_r)
        lizzieLet12_3QError_Int_2_bufchan_d <= lizzieLet12_3QError_Int_2_d;
  Go_t lizzieLet12_3QError_Int_2_bufchan_buf;
  assign lizzieLet12_3QError_Int_2_bufchan_r = (! lizzieLet12_3QError_Int_2_bufchan_buf[0]);
  assign lizzieLet12_3QError_Int_2_argbuf_d = (lizzieLet12_3QError_Int_2_bufchan_buf[0] ? lizzieLet12_3QError_Int_2_bufchan_buf :
                                               lizzieLet12_3QError_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet12_3QError_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet12_3QError_Int_2_argbuf_r && lizzieLet12_3QError_Int_2_bufchan_buf[0]))
        lizzieLet12_3QError_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet12_3QError_Int_2_argbuf_r) && (! lizzieLet12_3QError_Int_2_bufchan_buf[0])))
        lizzieLet12_3QError_Int_2_bufchan_buf <= lizzieLet12_3QError_Int_2_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty MyDTInt_Bool) : (lizzieLet12_4,QTree_Int) (is_z_adda8G_goMux_mux,MyDTInt_Bool) > [(_63,MyDTInt_Bool),
                                                                                            (lizzieLet12_4QVal_Int,MyDTInt_Bool),
                                                                                            (lizzieLet12_4QNode_Int,MyDTInt_Bool),
                                                                                            (_62,MyDTInt_Bool)] */
  logic [3:0] is_z_adda8G_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet12_4_d[0] && is_z_adda8G_goMux_mux_d[0]))
      unique case (lizzieLet12_4_d[2:1])
        2'd0: is_z_adda8G_goMux_mux_onehotd = 4'd1;
        2'd1: is_z_adda8G_goMux_mux_onehotd = 4'd2;
        2'd2: is_z_adda8G_goMux_mux_onehotd = 4'd4;
        2'd3: is_z_adda8G_goMux_mux_onehotd = 4'd8;
        default: is_z_adda8G_goMux_mux_onehotd = 4'd0;
      endcase
    else is_z_adda8G_goMux_mux_onehotd = 4'd0;
  assign _63_d = is_z_adda8G_goMux_mux_onehotd[0];
  assign lizzieLet12_4QVal_Int_d = is_z_adda8G_goMux_mux_onehotd[1];
  assign lizzieLet12_4QNode_Int_d = is_z_adda8G_goMux_mux_onehotd[2];
  assign _62_d = is_z_adda8G_goMux_mux_onehotd[3];
  assign is_z_adda8G_goMux_mux_r = (| (is_z_adda8G_goMux_mux_onehotd & {_62_r,
                                                                        lizzieLet12_4QNode_Int_r,
                                                                        lizzieLet12_4QVal_Int_r,
                                                                        _63_r}));
  assign lizzieLet12_4_r = is_z_adda8G_goMux_mux_r;
  
  /* demux (Ty QTree_Int,
       Ty MyDTInt_Bool) : (lizzieLet12_5,QTree_Int) (is_z_mapa8E_goMux_mux,MyDTInt_Bool) > [(lizzieLet12_5QNone_Int,MyDTInt_Bool),
                                                                                            (lizzieLet12_5QVal_Int,MyDTInt_Bool),
                                                                                            (lizzieLet12_5QNode_Int,MyDTInt_Bool),
                                                                                            (_61,MyDTInt_Bool)] */
  logic [3:0] is_z_mapa8E_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet12_5_d[0] && is_z_mapa8E_goMux_mux_d[0]))
      unique case (lizzieLet12_5_d[2:1])
        2'd0: is_z_mapa8E_goMux_mux_onehotd = 4'd1;
        2'd1: is_z_mapa8E_goMux_mux_onehotd = 4'd2;
        2'd2: is_z_mapa8E_goMux_mux_onehotd = 4'd4;
        2'd3: is_z_mapa8E_goMux_mux_onehotd = 4'd8;
        default: is_z_mapa8E_goMux_mux_onehotd = 4'd0;
      endcase
    else is_z_mapa8E_goMux_mux_onehotd = 4'd0;
  assign lizzieLet12_5QNone_Int_d = is_z_mapa8E_goMux_mux_onehotd[0];
  assign lizzieLet12_5QVal_Int_d = is_z_mapa8E_goMux_mux_onehotd[1];
  assign lizzieLet12_5QNode_Int_d = is_z_mapa8E_goMux_mux_onehotd[2];
  assign _61_d = is_z_mapa8E_goMux_mux_onehotd[3];
  assign is_z_mapa8E_goMux_mux_r = (| (is_z_mapa8E_goMux_mux_onehotd & {_61_r,
                                                                        lizzieLet12_5QNode_Int_r,
                                                                        lizzieLet12_5QVal_Int_r,
                                                                        lizzieLet12_5QNone_Int_r}));
  assign lizzieLet12_5_r = is_z_mapa8E_goMux_mux_r;
  
  /* demux (Ty QTree_Int,
       Ty QTree_Int) : (lizzieLet12_6,QTree_Int) (readPointer_QTree_Intm2a8D_1_argbuf_rwb,QTree_Int) > [(lizzieLet12_6QNone_Int,QTree_Int),
                                                                                                        (lizzieLet12_6QVal_Int,QTree_Int),
                                                                                                        (lizzieLet12_6QNode_Int,QTree_Int),
                                                                                                        (_60,QTree_Int)] */
  logic [3:0] readPointer_QTree_Intm2a8D_1_argbuf_rwb_onehotd;
  always_comb
    if ((lizzieLet12_6_d[0] && readPointer_QTree_Intm2a8D_1_argbuf_rwb_d[0]))
      unique case (lizzieLet12_6_d[2:1])
        2'd0: readPointer_QTree_Intm2a8D_1_argbuf_rwb_onehotd = 4'd1;
        2'd1: readPointer_QTree_Intm2a8D_1_argbuf_rwb_onehotd = 4'd2;
        2'd2: readPointer_QTree_Intm2a8D_1_argbuf_rwb_onehotd = 4'd4;
        2'd3: readPointer_QTree_Intm2a8D_1_argbuf_rwb_onehotd = 4'd8;
        default: readPointer_QTree_Intm2a8D_1_argbuf_rwb_onehotd = 4'd0;
      endcase
    else readPointer_QTree_Intm2a8D_1_argbuf_rwb_onehotd = 4'd0;
  assign lizzieLet12_6QNone_Int_d = {readPointer_QTree_Intm2a8D_1_argbuf_rwb_d[66:1],
                                     readPointer_QTree_Intm2a8D_1_argbuf_rwb_onehotd[0]};
  assign lizzieLet12_6QVal_Int_d = {readPointer_QTree_Intm2a8D_1_argbuf_rwb_d[66:1],
                                    readPointer_QTree_Intm2a8D_1_argbuf_rwb_onehotd[1]};
  assign lizzieLet12_6QNode_Int_d = {readPointer_QTree_Intm2a8D_1_argbuf_rwb_d[66:1],
                                     readPointer_QTree_Intm2a8D_1_argbuf_rwb_onehotd[2]};
  assign _60_d = {readPointer_QTree_Intm2a8D_1_argbuf_rwb_d[66:1],
                  readPointer_QTree_Intm2a8D_1_argbuf_rwb_onehotd[3]};
  assign readPointer_QTree_Intm2a8D_1_argbuf_rwb_r = (| (readPointer_QTree_Intm2a8D_1_argbuf_rwb_onehotd & {_60_r,
                                                                                                            lizzieLet12_6QNode_Int_r,
                                                                                                            lizzieLet12_6QVal_Int_r,
                                                                                                            lizzieLet12_6QNone_Int_r}));
  assign lizzieLet12_6_r = readPointer_QTree_Intm2a8D_1_argbuf_rwb_r;
  
  /* fork (Ty QTree_Int) : (lizzieLet12_6QNode_Int,QTree_Int) > [(lizzieLet12_6QNode_Int_1,QTree_Int),
                                                            (lizzieLet12_6QNode_Int_2,QTree_Int),
                                                            (lizzieLet12_6QNode_Int_3,QTree_Int),
                                                            (lizzieLet12_6QNode_Int_4,QTree_Int),
                                                            (lizzieLet12_6QNode_Int_5,QTree_Int),
                                                            (lizzieLet12_6QNode_Int_6,QTree_Int),
                                                            (lizzieLet12_6QNode_Int_7,QTree_Int),
                                                            (lizzieLet12_6QNode_Int_8,QTree_Int),
                                                            (lizzieLet12_6QNode_Int_9,QTree_Int),
                                                            (lizzieLet12_6QNode_Int_10,QTree_Int),
                                                            (lizzieLet12_6QNode_Int_11,QTree_Int),
                                                            (lizzieLet12_6QNode_Int_12,QTree_Int)] */
  logic [11:0] lizzieLet12_6QNode_Int_emitted;
  logic [11:0] lizzieLet12_6QNode_Int_done;
  assign lizzieLet12_6QNode_Int_1_d = {lizzieLet12_6QNode_Int_d[66:1],
                                       (lizzieLet12_6QNode_Int_d[0] && (! lizzieLet12_6QNode_Int_emitted[0]))};
  assign lizzieLet12_6QNode_Int_2_d = {lizzieLet12_6QNode_Int_d[66:1],
                                       (lizzieLet12_6QNode_Int_d[0] && (! lizzieLet12_6QNode_Int_emitted[1]))};
  assign lizzieLet12_6QNode_Int_3_d = {lizzieLet12_6QNode_Int_d[66:1],
                                       (lizzieLet12_6QNode_Int_d[0] && (! lizzieLet12_6QNode_Int_emitted[2]))};
  assign lizzieLet12_6QNode_Int_4_d = {lizzieLet12_6QNode_Int_d[66:1],
                                       (lizzieLet12_6QNode_Int_d[0] && (! lizzieLet12_6QNode_Int_emitted[3]))};
  assign lizzieLet12_6QNode_Int_5_d = {lizzieLet12_6QNode_Int_d[66:1],
                                       (lizzieLet12_6QNode_Int_d[0] && (! lizzieLet12_6QNode_Int_emitted[4]))};
  assign lizzieLet12_6QNode_Int_6_d = {lizzieLet12_6QNode_Int_d[66:1],
                                       (lizzieLet12_6QNode_Int_d[0] && (! lizzieLet12_6QNode_Int_emitted[5]))};
  assign lizzieLet12_6QNode_Int_7_d = {lizzieLet12_6QNode_Int_d[66:1],
                                       (lizzieLet12_6QNode_Int_d[0] && (! lizzieLet12_6QNode_Int_emitted[6]))};
  assign lizzieLet12_6QNode_Int_8_d = {lizzieLet12_6QNode_Int_d[66:1],
                                       (lizzieLet12_6QNode_Int_d[0] && (! lizzieLet12_6QNode_Int_emitted[7]))};
  assign lizzieLet12_6QNode_Int_9_d = {lizzieLet12_6QNode_Int_d[66:1],
                                       (lizzieLet12_6QNode_Int_d[0] && (! lizzieLet12_6QNode_Int_emitted[8]))};
  assign lizzieLet12_6QNode_Int_10_d = {lizzieLet12_6QNode_Int_d[66:1],
                                        (lizzieLet12_6QNode_Int_d[0] && (! lizzieLet12_6QNode_Int_emitted[9]))};
  assign lizzieLet12_6QNode_Int_11_d = {lizzieLet12_6QNode_Int_d[66:1],
                                        (lizzieLet12_6QNode_Int_d[0] && (! lizzieLet12_6QNode_Int_emitted[10]))};
  assign lizzieLet12_6QNode_Int_12_d = {lizzieLet12_6QNode_Int_d[66:1],
                                        (lizzieLet12_6QNode_Int_d[0] && (! lizzieLet12_6QNode_Int_emitted[11]))};
  assign lizzieLet12_6QNode_Int_done = (lizzieLet12_6QNode_Int_emitted | ({lizzieLet12_6QNode_Int_12_d[0],
                                                                           lizzieLet12_6QNode_Int_11_d[0],
                                                                           lizzieLet12_6QNode_Int_10_d[0],
                                                                           lizzieLet12_6QNode_Int_9_d[0],
                                                                           lizzieLet12_6QNode_Int_8_d[0],
                                                                           lizzieLet12_6QNode_Int_7_d[0],
                                                                           lizzieLet12_6QNode_Int_6_d[0],
                                                                           lizzieLet12_6QNode_Int_5_d[0],
                                                                           lizzieLet12_6QNode_Int_4_d[0],
                                                                           lizzieLet12_6QNode_Int_3_d[0],
                                                                           lizzieLet12_6QNode_Int_2_d[0],
                                                                           lizzieLet12_6QNode_Int_1_d[0]} & {lizzieLet12_6QNode_Int_12_r,
                                                                                                             lizzieLet12_6QNode_Int_11_r,
                                                                                                             lizzieLet12_6QNode_Int_10_r,
                                                                                                             lizzieLet12_6QNode_Int_9_r,
                                                                                                             lizzieLet12_6QNode_Int_8_r,
                                                                                                             lizzieLet12_6QNode_Int_7_r,
                                                                                                             lizzieLet12_6QNode_Int_6_r,
                                                                                                             lizzieLet12_6QNode_Int_5_r,
                                                                                                             lizzieLet12_6QNode_Int_4_r,
                                                                                                             lizzieLet12_6QNode_Int_3_r,
                                                                                                             lizzieLet12_6QNode_Int_2_r,
                                                                                                             lizzieLet12_6QNode_Int_1_r}));
  assign lizzieLet12_6QNode_Int_r = (& lizzieLet12_6QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet12_6QNode_Int_emitted <= 12'd0;
    else
      lizzieLet12_6QNode_Int_emitted <= (lizzieLet12_6QNode_Int_r ? 12'd0 :
                                         lizzieLet12_6QNode_Int_done);
  
  /* demux (Ty QTree_Int,
       Ty Pointer_QTree_Int) : (lizzieLet12_6QNode_Int_10,QTree_Int) (q2a8U_destruct,Pointer_QTree_Int) > [(lizzieLet12_6QNode_Int_10QNone_Int,Pointer_QTree_Int),
                                                                                                           (_59,Pointer_QTree_Int),
                                                                                                           (lizzieLet12_6QNode_Int_10QNode_Int,Pointer_QTree_Int),
                                                                                                           (_58,Pointer_QTree_Int)] */
  logic [3:0] q2a8U_destruct_onehotd;
  always_comb
    if ((lizzieLet12_6QNode_Int_10_d[0] && q2a8U_destruct_d[0]))
      unique case (lizzieLet12_6QNode_Int_10_d[2:1])
        2'd0: q2a8U_destruct_onehotd = 4'd1;
        2'd1: q2a8U_destruct_onehotd = 4'd2;
        2'd2: q2a8U_destruct_onehotd = 4'd4;
        2'd3: q2a8U_destruct_onehotd = 4'd8;
        default: q2a8U_destruct_onehotd = 4'd0;
      endcase
    else q2a8U_destruct_onehotd = 4'd0;
  assign lizzieLet12_6QNode_Int_10QNone_Int_d = {q2a8U_destruct_d[16:1],
                                                 q2a8U_destruct_onehotd[0]};
  assign _59_d = {q2a8U_destruct_d[16:1], q2a8U_destruct_onehotd[1]};
  assign lizzieLet12_6QNode_Int_10QNode_Int_d = {q2a8U_destruct_d[16:1],
                                                 q2a8U_destruct_onehotd[2]};
  assign _58_d = {q2a8U_destruct_d[16:1], q2a8U_destruct_onehotd[3]};
  assign q2a8U_destruct_r = (| (q2a8U_destruct_onehotd & {_58_r,
                                                          lizzieLet12_6QNode_Int_10QNode_Int_r,
                                                          _59_r,
                                                          lizzieLet12_6QNode_Int_10QNone_Int_r}));
  assign lizzieLet12_6QNode_Int_10_r = q2a8U_destruct_r;
  
  /* buf (Ty Pointer_QTree_Int) : (lizzieLet12_6QNode_Int_10QNone_Int,Pointer_QTree_Int) > (lizzieLet12_6QNode_Int_10QNone_Int_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t lizzieLet12_6QNode_Int_10QNone_Int_bufchan_d;
  logic lizzieLet12_6QNode_Int_10QNone_Int_bufchan_r;
  assign lizzieLet12_6QNode_Int_10QNone_Int_r = ((! lizzieLet12_6QNode_Int_10QNone_Int_bufchan_d[0]) || lizzieLet12_6QNode_Int_10QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNode_Int_10QNone_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet12_6QNode_Int_10QNone_Int_r)
        lizzieLet12_6QNode_Int_10QNone_Int_bufchan_d <= lizzieLet12_6QNode_Int_10QNone_Int_d;
  Pointer_QTree_Int_t lizzieLet12_6QNode_Int_10QNone_Int_bufchan_buf;
  assign lizzieLet12_6QNode_Int_10QNone_Int_bufchan_r = (! lizzieLet12_6QNode_Int_10QNone_Int_bufchan_buf[0]);
  assign lizzieLet12_6QNode_Int_10QNone_Int_1_argbuf_d = (lizzieLet12_6QNode_Int_10QNone_Int_bufchan_buf[0] ? lizzieLet12_6QNode_Int_10QNone_Int_bufchan_buf :
                                                          lizzieLet12_6QNode_Int_10QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNode_Int_10QNone_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet12_6QNode_Int_10QNone_Int_1_argbuf_r && lizzieLet12_6QNode_Int_10QNone_Int_bufchan_buf[0]))
        lizzieLet12_6QNode_Int_10QNone_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet12_6QNode_Int_10QNone_Int_1_argbuf_r) && (! lizzieLet12_6QNode_Int_10QNone_Int_bufchan_buf[0])))
        lizzieLet12_6QNode_Int_10QNone_Int_bufchan_buf <= lizzieLet12_6QNode_Int_10QNone_Int_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_QTree_Int) : (lizzieLet12_6QNode_Int_11,QTree_Int) (q3a8V_destruct,Pointer_QTree_Int) > [(lizzieLet12_6QNode_Int_11QNone_Int,Pointer_QTree_Int),
                                                                                                           (_57,Pointer_QTree_Int),
                                                                                                           (lizzieLet12_6QNode_Int_11QNode_Int,Pointer_QTree_Int),
                                                                                                           (_56,Pointer_QTree_Int)] */
  logic [3:0] q3a8V_destruct_onehotd;
  always_comb
    if ((lizzieLet12_6QNode_Int_11_d[0] && q3a8V_destruct_d[0]))
      unique case (lizzieLet12_6QNode_Int_11_d[2:1])
        2'd0: q3a8V_destruct_onehotd = 4'd1;
        2'd1: q3a8V_destruct_onehotd = 4'd2;
        2'd2: q3a8V_destruct_onehotd = 4'd4;
        2'd3: q3a8V_destruct_onehotd = 4'd8;
        default: q3a8V_destruct_onehotd = 4'd0;
      endcase
    else q3a8V_destruct_onehotd = 4'd0;
  assign lizzieLet12_6QNode_Int_11QNone_Int_d = {q3a8V_destruct_d[16:1],
                                                 q3a8V_destruct_onehotd[0]};
  assign _57_d = {q3a8V_destruct_d[16:1], q3a8V_destruct_onehotd[1]};
  assign lizzieLet12_6QNode_Int_11QNode_Int_d = {q3a8V_destruct_d[16:1],
                                                 q3a8V_destruct_onehotd[2]};
  assign _56_d = {q3a8V_destruct_d[16:1], q3a8V_destruct_onehotd[3]};
  assign q3a8V_destruct_r = (| (q3a8V_destruct_onehotd & {_56_r,
                                                          lizzieLet12_6QNode_Int_11QNode_Int_r,
                                                          _57_r,
                                                          lizzieLet12_6QNode_Int_11QNone_Int_r}));
  assign lizzieLet12_6QNode_Int_11_r = q3a8V_destruct_r;
  
  /* buf (Ty Pointer_QTree_Int) : (lizzieLet12_6QNode_Int_11QNone_Int,Pointer_QTree_Int) > (lizzieLet12_6QNode_Int_11QNone_Int_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t lizzieLet12_6QNode_Int_11QNone_Int_bufchan_d;
  logic lizzieLet12_6QNode_Int_11QNone_Int_bufchan_r;
  assign lizzieLet12_6QNode_Int_11QNone_Int_r = ((! lizzieLet12_6QNode_Int_11QNone_Int_bufchan_d[0]) || lizzieLet12_6QNode_Int_11QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNode_Int_11QNone_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet12_6QNode_Int_11QNone_Int_r)
        lizzieLet12_6QNode_Int_11QNone_Int_bufchan_d <= lizzieLet12_6QNode_Int_11QNone_Int_d;
  Pointer_QTree_Int_t lizzieLet12_6QNode_Int_11QNone_Int_bufchan_buf;
  assign lizzieLet12_6QNode_Int_11QNone_Int_bufchan_r = (! lizzieLet12_6QNode_Int_11QNone_Int_bufchan_buf[0]);
  assign lizzieLet12_6QNode_Int_11QNone_Int_1_argbuf_d = (lizzieLet12_6QNode_Int_11QNone_Int_bufchan_buf[0] ? lizzieLet12_6QNode_Int_11QNone_Int_bufchan_buf :
                                                          lizzieLet12_6QNode_Int_11QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNode_Int_11QNone_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet12_6QNode_Int_11QNone_Int_1_argbuf_r && lizzieLet12_6QNode_Int_11QNone_Int_bufchan_buf[0]))
        lizzieLet12_6QNode_Int_11QNone_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet12_6QNode_Int_11QNone_Int_1_argbuf_r) && (! lizzieLet12_6QNode_Int_11QNone_Int_bufchan_buf[0])))
        lizzieLet12_6QNode_Int_11QNone_Int_bufchan_buf <= lizzieLet12_6QNode_Int_11QNone_Int_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_QTree_Int) : (lizzieLet12_6QNode_Int_12,QTree_Int) (q4a8W_destruct,Pointer_QTree_Int) > [(lizzieLet12_6QNode_Int_12QNone_Int,Pointer_QTree_Int),
                                                                                                           (_55,Pointer_QTree_Int),
                                                                                                           (lizzieLet12_6QNode_Int_12QNode_Int,Pointer_QTree_Int),
                                                                                                           (_54,Pointer_QTree_Int)] */
  logic [3:0] q4a8W_destruct_onehotd;
  always_comb
    if ((lizzieLet12_6QNode_Int_12_d[0] && q4a8W_destruct_d[0]))
      unique case (lizzieLet12_6QNode_Int_12_d[2:1])
        2'd0: q4a8W_destruct_onehotd = 4'd1;
        2'd1: q4a8W_destruct_onehotd = 4'd2;
        2'd2: q4a8W_destruct_onehotd = 4'd4;
        2'd3: q4a8W_destruct_onehotd = 4'd8;
        default: q4a8W_destruct_onehotd = 4'd0;
      endcase
    else q4a8W_destruct_onehotd = 4'd0;
  assign lizzieLet12_6QNode_Int_12QNone_Int_d = {q4a8W_destruct_d[16:1],
                                                 q4a8W_destruct_onehotd[0]};
  assign _55_d = {q4a8W_destruct_d[16:1], q4a8W_destruct_onehotd[1]};
  assign lizzieLet12_6QNode_Int_12QNode_Int_d = {q4a8W_destruct_d[16:1],
                                                 q4a8W_destruct_onehotd[2]};
  assign _54_d = {q4a8W_destruct_d[16:1], q4a8W_destruct_onehotd[3]};
  assign q4a8W_destruct_r = (| (q4a8W_destruct_onehotd & {_54_r,
                                                          lizzieLet12_6QNode_Int_12QNode_Int_r,
                                                          _55_r,
                                                          lizzieLet12_6QNode_Int_12QNone_Int_r}));
  assign lizzieLet12_6QNode_Int_12_r = q4a8W_destruct_r;
  
  /* buf (Ty Pointer_QTree_Int) : (lizzieLet12_6QNode_Int_12QNode_Int,Pointer_QTree_Int) > (lizzieLet12_6QNode_Int_12QNode_Int_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t lizzieLet12_6QNode_Int_12QNode_Int_bufchan_d;
  logic lizzieLet12_6QNode_Int_12QNode_Int_bufchan_r;
  assign lizzieLet12_6QNode_Int_12QNode_Int_r = ((! lizzieLet12_6QNode_Int_12QNode_Int_bufchan_d[0]) || lizzieLet12_6QNode_Int_12QNode_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNode_Int_12QNode_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet12_6QNode_Int_12QNode_Int_r)
        lizzieLet12_6QNode_Int_12QNode_Int_bufchan_d <= lizzieLet12_6QNode_Int_12QNode_Int_d;
  Pointer_QTree_Int_t lizzieLet12_6QNode_Int_12QNode_Int_bufchan_buf;
  assign lizzieLet12_6QNode_Int_12QNode_Int_bufchan_r = (! lizzieLet12_6QNode_Int_12QNode_Int_bufchan_buf[0]);
  assign lizzieLet12_6QNode_Int_12QNode_Int_1_argbuf_d = (lizzieLet12_6QNode_Int_12QNode_Int_bufchan_buf[0] ? lizzieLet12_6QNode_Int_12QNode_Int_bufchan_buf :
                                                          lizzieLet12_6QNode_Int_12QNode_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNode_Int_12QNode_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet12_6QNode_Int_12QNode_Int_1_argbuf_r && lizzieLet12_6QNode_Int_12QNode_Int_bufchan_buf[0]))
        lizzieLet12_6QNode_Int_12QNode_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet12_6QNode_Int_12QNode_Int_1_argbuf_r) && (! lizzieLet12_6QNode_Int_12QNode_Int_bufchan_buf[0])))
        lizzieLet12_6QNode_Int_12QNode_Int_bufchan_buf <= lizzieLet12_6QNode_Int_12QNode_Int_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (lizzieLet12_6QNode_Int_12QNone_Int,Pointer_QTree_Int) > (lizzieLet12_6QNode_Int_12QNone_Int_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t lizzieLet12_6QNode_Int_12QNone_Int_bufchan_d;
  logic lizzieLet12_6QNode_Int_12QNone_Int_bufchan_r;
  assign lizzieLet12_6QNode_Int_12QNone_Int_r = ((! lizzieLet12_6QNode_Int_12QNone_Int_bufchan_d[0]) || lizzieLet12_6QNode_Int_12QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNode_Int_12QNone_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet12_6QNode_Int_12QNone_Int_r)
        lizzieLet12_6QNode_Int_12QNone_Int_bufchan_d <= lizzieLet12_6QNode_Int_12QNone_Int_d;
  Pointer_QTree_Int_t lizzieLet12_6QNode_Int_12QNone_Int_bufchan_buf;
  assign lizzieLet12_6QNode_Int_12QNone_Int_bufchan_r = (! lizzieLet12_6QNode_Int_12QNone_Int_bufchan_buf[0]);
  assign lizzieLet12_6QNode_Int_12QNone_Int_1_argbuf_d = (lizzieLet12_6QNode_Int_12QNone_Int_bufchan_buf[0] ? lizzieLet12_6QNode_Int_12QNone_Int_bufchan_buf :
                                                          lizzieLet12_6QNode_Int_12QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNode_Int_12QNone_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet12_6QNode_Int_12QNone_Int_1_argbuf_r && lizzieLet12_6QNode_Int_12QNone_Int_bufchan_buf[0]))
        lizzieLet12_6QNode_Int_12QNone_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet12_6QNode_Int_12QNone_Int_1_argbuf_r) && (! lizzieLet12_6QNode_Int_12QNone_Int_bufchan_buf[0])))
        lizzieLet12_6QNode_Int_12QNone_Int_bufchan_buf <= lizzieLet12_6QNode_Int_12QNone_Int_bufchan_d;
  
  /* destruct (Ty QTree_Int,
          Dcon QNode_Int) : (lizzieLet12_6QNode_Int_1QNode_Int,QTree_Int) > [(t1a8Y_destruct,Pointer_QTree_Int),
                                                                             (t2a8Z_destruct,Pointer_QTree_Int),
                                                                             (t3a90_destruct,Pointer_QTree_Int),
                                                                             (t4a91_destruct,Pointer_QTree_Int)] */
  logic [3:0] lizzieLet12_6QNode_Int_1QNode_Int_emitted;
  logic [3:0] lizzieLet12_6QNode_Int_1QNode_Int_done;
  assign t1a8Y_destruct_d = {lizzieLet12_6QNode_Int_1QNode_Int_d[18:3],
                             (lizzieLet12_6QNode_Int_1QNode_Int_d[0] && (! lizzieLet12_6QNode_Int_1QNode_Int_emitted[0]))};
  assign t2a8Z_destruct_d = {lizzieLet12_6QNode_Int_1QNode_Int_d[34:19],
                             (lizzieLet12_6QNode_Int_1QNode_Int_d[0] && (! lizzieLet12_6QNode_Int_1QNode_Int_emitted[1]))};
  assign t3a90_destruct_d = {lizzieLet12_6QNode_Int_1QNode_Int_d[50:35],
                             (lizzieLet12_6QNode_Int_1QNode_Int_d[0] && (! lizzieLet12_6QNode_Int_1QNode_Int_emitted[2]))};
  assign t4a91_destruct_d = {lizzieLet12_6QNode_Int_1QNode_Int_d[66:51],
                             (lizzieLet12_6QNode_Int_1QNode_Int_d[0] && (! lizzieLet12_6QNode_Int_1QNode_Int_emitted[3]))};
  assign lizzieLet12_6QNode_Int_1QNode_Int_done = (lizzieLet12_6QNode_Int_1QNode_Int_emitted | ({t4a91_destruct_d[0],
                                                                                                 t3a90_destruct_d[0],
                                                                                                 t2a8Z_destruct_d[0],
                                                                                                 t1a8Y_destruct_d[0]} & {t4a91_destruct_r,
                                                                                                                         t3a90_destruct_r,
                                                                                                                         t2a8Z_destruct_r,
                                                                                                                         t1a8Y_destruct_r}));
  assign lizzieLet12_6QNode_Int_1QNode_Int_r = (& lizzieLet12_6QNode_Int_1QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNode_Int_1QNode_Int_emitted <= 4'd0;
    else
      lizzieLet12_6QNode_Int_1QNode_Int_emitted <= (lizzieLet12_6QNode_Int_1QNode_Int_r ? 4'd0 :
                                                    lizzieLet12_6QNode_Int_1QNode_Int_done);
  
  /* demux (Ty QTree_Int,
       Ty QTree_Int) : (lizzieLet12_6QNode_Int_2,QTree_Int) (lizzieLet12_6QNode_Int_1,QTree_Int) > [(_53,QTree_Int),
                                                                                                    (_52,QTree_Int),
                                                                                                    (lizzieLet12_6QNode_Int_1QNode_Int,QTree_Int),
                                                                                                    (_51,QTree_Int)] */
  logic [3:0] lizzieLet12_6QNode_Int_1_onehotd;
  always_comb
    if ((lizzieLet12_6QNode_Int_2_d[0] && lizzieLet12_6QNode_Int_1_d[0]))
      unique case (lizzieLet12_6QNode_Int_2_d[2:1])
        2'd0: lizzieLet12_6QNode_Int_1_onehotd = 4'd1;
        2'd1: lizzieLet12_6QNode_Int_1_onehotd = 4'd2;
        2'd2: lizzieLet12_6QNode_Int_1_onehotd = 4'd4;
        2'd3: lizzieLet12_6QNode_Int_1_onehotd = 4'd8;
        default: lizzieLet12_6QNode_Int_1_onehotd = 4'd0;
      endcase
    else lizzieLet12_6QNode_Int_1_onehotd = 4'd0;
  assign _53_d = {lizzieLet12_6QNode_Int_1_d[66:1],
                  lizzieLet12_6QNode_Int_1_onehotd[0]};
  assign _52_d = {lizzieLet12_6QNode_Int_1_d[66:1],
                  lizzieLet12_6QNode_Int_1_onehotd[1]};
  assign lizzieLet12_6QNode_Int_1QNode_Int_d = {lizzieLet12_6QNode_Int_1_d[66:1],
                                                lizzieLet12_6QNode_Int_1_onehotd[2]};
  assign _51_d = {lizzieLet12_6QNode_Int_1_d[66:1],
                  lizzieLet12_6QNode_Int_1_onehotd[3]};
  assign lizzieLet12_6QNode_Int_1_r = (| (lizzieLet12_6QNode_Int_1_onehotd & {_51_r,
                                                                              lizzieLet12_6QNode_Int_1QNode_Int_r,
                                                                              _52_r,
                                                                              _53_r}));
  assign lizzieLet12_6QNode_Int_2_r = lizzieLet12_6QNode_Int_1_r;
  
  /* demux (Ty QTree_Int,
       Ty Go) : (lizzieLet12_6QNode_Int_3,QTree_Int) (lizzieLet12_3QNode_Int,Go) > [(lizzieLet12_6QNode_Int_3QNone_Int,Go),
                                                                                    (lizzieLet12_6QNode_Int_3QVal_Int,Go),
                                                                                    (lizzieLet12_6QNode_Int_3QNode_Int,Go),
                                                                                    (lizzieLet12_6QNode_Int_3QError_Int,Go)] */
  logic [3:0] lizzieLet12_3QNode_Int_onehotd;
  always_comb
    if ((lizzieLet12_6QNode_Int_3_d[0] && lizzieLet12_3QNode_Int_d[0]))
      unique case (lizzieLet12_6QNode_Int_3_d[2:1])
        2'd0: lizzieLet12_3QNode_Int_onehotd = 4'd1;
        2'd1: lizzieLet12_3QNode_Int_onehotd = 4'd2;
        2'd2: lizzieLet12_3QNode_Int_onehotd = 4'd4;
        2'd3: lizzieLet12_3QNode_Int_onehotd = 4'd8;
        default: lizzieLet12_3QNode_Int_onehotd = 4'd0;
      endcase
    else lizzieLet12_3QNode_Int_onehotd = 4'd0;
  assign lizzieLet12_6QNode_Int_3QNone_Int_d = lizzieLet12_3QNode_Int_onehotd[0];
  assign lizzieLet12_6QNode_Int_3QVal_Int_d = lizzieLet12_3QNode_Int_onehotd[1];
  assign lizzieLet12_6QNode_Int_3QNode_Int_d = lizzieLet12_3QNode_Int_onehotd[2];
  assign lizzieLet12_6QNode_Int_3QError_Int_d = lizzieLet12_3QNode_Int_onehotd[3];
  assign lizzieLet12_3QNode_Int_r = (| (lizzieLet12_3QNode_Int_onehotd & {lizzieLet12_6QNode_Int_3QError_Int_r,
                                                                          lizzieLet12_6QNode_Int_3QNode_Int_r,
                                                                          lizzieLet12_6QNode_Int_3QVal_Int_r,
                                                                          lizzieLet12_6QNode_Int_3QNone_Int_r}));
  assign lizzieLet12_6QNode_Int_3_r = lizzieLet12_3QNode_Int_r;
  
  /* fork (Ty Go) : (lizzieLet12_6QNode_Int_3QError_Int,Go) > [(lizzieLet12_6QNode_Int_3QError_Int_1,Go),
                                                          (lizzieLet12_6QNode_Int_3QError_Int_2,Go)] */
  logic [1:0] lizzieLet12_6QNode_Int_3QError_Int_emitted;
  logic [1:0] lizzieLet12_6QNode_Int_3QError_Int_done;
  assign lizzieLet12_6QNode_Int_3QError_Int_1_d = (lizzieLet12_6QNode_Int_3QError_Int_d[0] && (! lizzieLet12_6QNode_Int_3QError_Int_emitted[0]));
  assign lizzieLet12_6QNode_Int_3QError_Int_2_d = (lizzieLet12_6QNode_Int_3QError_Int_d[0] && (! lizzieLet12_6QNode_Int_3QError_Int_emitted[1]));
  assign lizzieLet12_6QNode_Int_3QError_Int_done = (lizzieLet12_6QNode_Int_3QError_Int_emitted | ({lizzieLet12_6QNode_Int_3QError_Int_2_d[0],
                                                                                                   lizzieLet12_6QNode_Int_3QError_Int_1_d[0]} & {lizzieLet12_6QNode_Int_3QError_Int_2_r,
                                                                                                                                                 lizzieLet12_6QNode_Int_3QError_Int_1_r}));
  assign lizzieLet12_6QNode_Int_3QError_Int_r = (& lizzieLet12_6QNode_Int_3QError_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNode_Int_3QError_Int_emitted <= 2'd0;
    else
      lizzieLet12_6QNode_Int_3QError_Int_emitted <= (lizzieLet12_6QNode_Int_3QError_Int_r ? 2'd0 :
                                                     lizzieLet12_6QNode_Int_3QError_Int_done);
  
  /* dcon (Ty QTree_Int,
      Dcon QError_Int) : [(lizzieLet12_6QNode_Int_3QError_Int_1,Go)] > (lizzieLet12_6QNode_Int_3QError_Int_1QError_Int,QTree_Int) */
  assign lizzieLet12_6QNode_Int_3QError_Int_1QError_Int_d = QError_Int_dc((& {lizzieLet12_6QNode_Int_3QError_Int_1_d[0]}), lizzieLet12_6QNode_Int_3QError_Int_1_d);
  assign {lizzieLet12_6QNode_Int_3QError_Int_1_r} = {1 {(lizzieLet12_6QNode_Int_3QError_Int_1QError_Int_r && lizzieLet12_6QNode_Int_3QError_Int_1QError_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (lizzieLet12_6QNode_Int_3QError_Int_1QError_Int,QTree_Int) > (lizzieLet31_1_argbuf,QTree_Int) */
  QTree_Int_t lizzieLet12_6QNode_Int_3QError_Int_1QError_Int_bufchan_d;
  logic lizzieLet12_6QNode_Int_3QError_Int_1QError_Int_bufchan_r;
  assign lizzieLet12_6QNode_Int_3QError_Int_1QError_Int_r = ((! lizzieLet12_6QNode_Int_3QError_Int_1QError_Int_bufchan_d[0]) || lizzieLet12_6QNode_Int_3QError_Int_1QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNode_Int_3QError_Int_1QError_Int_bufchan_d <= {66'd0,
                                                                   1'd0};
    else
      if (lizzieLet12_6QNode_Int_3QError_Int_1QError_Int_r)
        lizzieLet12_6QNode_Int_3QError_Int_1QError_Int_bufchan_d <= lizzieLet12_6QNode_Int_3QError_Int_1QError_Int_d;
  QTree_Int_t lizzieLet12_6QNode_Int_3QError_Int_1QError_Int_bufchan_buf;
  assign lizzieLet12_6QNode_Int_3QError_Int_1QError_Int_bufchan_r = (! lizzieLet12_6QNode_Int_3QError_Int_1QError_Int_bufchan_buf[0]);
  assign lizzieLet31_1_argbuf_d = (lizzieLet12_6QNode_Int_3QError_Int_1QError_Int_bufchan_buf[0] ? lizzieLet12_6QNode_Int_3QError_Int_1QError_Int_bufchan_buf :
                                   lizzieLet12_6QNode_Int_3QError_Int_1QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNode_Int_3QError_Int_1QError_Int_bufchan_buf <= {66'd0,
                                                                     1'd0};
    else
      if ((lizzieLet31_1_argbuf_r && lizzieLet12_6QNode_Int_3QError_Int_1QError_Int_bufchan_buf[0]))
        lizzieLet12_6QNode_Int_3QError_Int_1QError_Int_bufchan_buf <= {66'd0,
                                                                       1'd0};
      else if (((! lizzieLet31_1_argbuf_r) && (! lizzieLet12_6QNode_Int_3QError_Int_1QError_Int_bufchan_buf[0])))
        lizzieLet12_6QNode_Int_3QError_Int_1QError_Int_bufchan_buf <= lizzieLet12_6QNode_Int_3QError_Int_1QError_Int_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet12_6QNode_Int_3QError_Int_2,Go) > (lizzieLet12_6QNode_Int_3QError_Int_2_argbuf,Go) */
  Go_t lizzieLet12_6QNode_Int_3QError_Int_2_bufchan_d;
  logic lizzieLet12_6QNode_Int_3QError_Int_2_bufchan_r;
  assign lizzieLet12_6QNode_Int_3QError_Int_2_r = ((! lizzieLet12_6QNode_Int_3QError_Int_2_bufchan_d[0]) || lizzieLet12_6QNode_Int_3QError_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNode_Int_3QError_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet12_6QNode_Int_3QError_Int_2_r)
        lizzieLet12_6QNode_Int_3QError_Int_2_bufchan_d <= lizzieLet12_6QNode_Int_3QError_Int_2_d;
  Go_t lizzieLet12_6QNode_Int_3QError_Int_2_bufchan_buf;
  assign lizzieLet12_6QNode_Int_3QError_Int_2_bufchan_r = (! lizzieLet12_6QNode_Int_3QError_Int_2_bufchan_buf[0]);
  assign lizzieLet12_6QNode_Int_3QError_Int_2_argbuf_d = (lizzieLet12_6QNode_Int_3QError_Int_2_bufchan_buf[0] ? lizzieLet12_6QNode_Int_3QError_Int_2_bufchan_buf :
                                                          lizzieLet12_6QNode_Int_3QError_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNode_Int_3QError_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet12_6QNode_Int_3QError_Int_2_argbuf_r && lizzieLet12_6QNode_Int_3QError_Int_2_bufchan_buf[0]))
        lizzieLet12_6QNode_Int_3QError_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet12_6QNode_Int_3QError_Int_2_argbuf_r) && (! lizzieLet12_6QNode_Int_3QError_Int_2_bufchan_buf[0])))
        lizzieLet12_6QNode_Int_3QError_Int_2_bufchan_buf <= lizzieLet12_6QNode_Int_3QError_Int_2_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet12_6QNode_Int_3QNode_Int,Go) > (lizzieLet12_6QNode_Int_3QNode_Int_1_argbuf,Go) */
  Go_t lizzieLet12_6QNode_Int_3QNode_Int_bufchan_d;
  logic lizzieLet12_6QNode_Int_3QNode_Int_bufchan_r;
  assign lizzieLet12_6QNode_Int_3QNode_Int_r = ((! lizzieLet12_6QNode_Int_3QNode_Int_bufchan_d[0]) || lizzieLet12_6QNode_Int_3QNode_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNode_Int_3QNode_Int_bufchan_d <= 1'd0;
    else
      if (lizzieLet12_6QNode_Int_3QNode_Int_r)
        lizzieLet12_6QNode_Int_3QNode_Int_bufchan_d <= lizzieLet12_6QNode_Int_3QNode_Int_d;
  Go_t lizzieLet12_6QNode_Int_3QNode_Int_bufchan_buf;
  assign lizzieLet12_6QNode_Int_3QNode_Int_bufchan_r = (! lizzieLet12_6QNode_Int_3QNode_Int_bufchan_buf[0]);
  assign lizzieLet12_6QNode_Int_3QNode_Int_1_argbuf_d = (lizzieLet12_6QNode_Int_3QNode_Int_bufchan_buf[0] ? lizzieLet12_6QNode_Int_3QNode_Int_bufchan_buf :
                                                         lizzieLet12_6QNode_Int_3QNode_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNode_Int_3QNode_Int_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet12_6QNode_Int_3QNode_Int_1_argbuf_r && lizzieLet12_6QNode_Int_3QNode_Int_bufchan_buf[0]))
        lizzieLet12_6QNode_Int_3QNode_Int_bufchan_buf <= 1'd0;
      else if (((! lizzieLet12_6QNode_Int_3QNode_Int_1_argbuf_r) && (! lizzieLet12_6QNode_Int_3QNode_Int_bufchan_buf[0])))
        lizzieLet12_6QNode_Int_3QNode_Int_bufchan_buf <= lizzieLet12_6QNode_Int_3QNode_Int_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet12_6QNode_Int_3QNone_Int,Go) > [(lizzieLet12_6QNode_Int_3QNone_Int_1,Go),
                                                         (lizzieLet12_6QNode_Int_3QNone_Int_2,Go),
                                                         (lizzieLet12_6QNode_Int_3QNone_Int_3,Go),
                                                         (lizzieLet12_6QNode_Int_3QNone_Int_4,Go),
                                                         (lizzieLet12_6QNode_Int_3QNone_Int_5,Go)] */
  logic [4:0] lizzieLet12_6QNode_Int_3QNone_Int_emitted;
  logic [4:0] lizzieLet12_6QNode_Int_3QNone_Int_done;
  assign lizzieLet12_6QNode_Int_3QNone_Int_1_d = (lizzieLet12_6QNode_Int_3QNone_Int_d[0] && (! lizzieLet12_6QNode_Int_3QNone_Int_emitted[0]));
  assign lizzieLet12_6QNode_Int_3QNone_Int_2_d = (lizzieLet12_6QNode_Int_3QNone_Int_d[0] && (! lizzieLet12_6QNode_Int_3QNone_Int_emitted[1]));
  assign lizzieLet12_6QNode_Int_3QNone_Int_3_d = (lizzieLet12_6QNode_Int_3QNone_Int_d[0] && (! lizzieLet12_6QNode_Int_3QNone_Int_emitted[2]));
  assign lizzieLet12_6QNode_Int_3QNone_Int_4_d = (lizzieLet12_6QNode_Int_3QNone_Int_d[0] && (! lizzieLet12_6QNode_Int_3QNone_Int_emitted[3]));
  assign lizzieLet12_6QNode_Int_3QNone_Int_5_d = (lizzieLet12_6QNode_Int_3QNone_Int_d[0] && (! lizzieLet12_6QNode_Int_3QNone_Int_emitted[4]));
  assign lizzieLet12_6QNode_Int_3QNone_Int_done = (lizzieLet12_6QNode_Int_3QNone_Int_emitted | ({lizzieLet12_6QNode_Int_3QNone_Int_5_d[0],
                                                                                                 lizzieLet12_6QNode_Int_3QNone_Int_4_d[0],
                                                                                                 lizzieLet12_6QNode_Int_3QNone_Int_3_d[0],
                                                                                                 lizzieLet12_6QNode_Int_3QNone_Int_2_d[0],
                                                                                                 lizzieLet12_6QNode_Int_3QNone_Int_1_d[0]} & {lizzieLet12_6QNode_Int_3QNone_Int_5_r,
                                                                                                                                              lizzieLet12_6QNode_Int_3QNone_Int_4_r,
                                                                                                                                              lizzieLet12_6QNode_Int_3QNone_Int_3_r,
                                                                                                                                              lizzieLet12_6QNode_Int_3QNone_Int_2_r,
                                                                                                                                              lizzieLet12_6QNode_Int_3QNone_Int_1_r}));
  assign lizzieLet12_6QNode_Int_3QNone_Int_r = (& lizzieLet12_6QNode_Int_3QNone_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNode_Int_3QNone_Int_emitted <= 5'd0;
    else
      lizzieLet12_6QNode_Int_3QNone_Int_emitted <= (lizzieLet12_6QNode_Int_3QNone_Int_r ? 5'd0 :
                                                    lizzieLet12_6QNode_Int_3QNone_Int_done);
  
  /* buf (Ty Go) : (lizzieLet12_6QNode_Int_3QNone_Int_1,Go) > (lizzieLet12_6QNode_Int_3QNone_Int_1_argbuf,Go) */
  Go_t lizzieLet12_6QNode_Int_3QNone_Int_1_bufchan_d;
  logic lizzieLet12_6QNode_Int_3QNone_Int_1_bufchan_r;
  assign lizzieLet12_6QNode_Int_3QNone_Int_1_r = ((! lizzieLet12_6QNode_Int_3QNone_Int_1_bufchan_d[0]) || lizzieLet12_6QNode_Int_3QNone_Int_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNode_Int_3QNone_Int_1_bufchan_d <= 1'd0;
    else
      if (lizzieLet12_6QNode_Int_3QNone_Int_1_r)
        lizzieLet12_6QNode_Int_3QNone_Int_1_bufchan_d <= lizzieLet12_6QNode_Int_3QNone_Int_1_d;
  Go_t lizzieLet12_6QNode_Int_3QNone_Int_1_bufchan_buf;
  assign lizzieLet12_6QNode_Int_3QNone_Int_1_bufchan_r = (! lizzieLet12_6QNode_Int_3QNone_Int_1_bufchan_buf[0]);
  assign lizzieLet12_6QNode_Int_3QNone_Int_1_argbuf_d = (lizzieLet12_6QNode_Int_3QNone_Int_1_bufchan_buf[0] ? lizzieLet12_6QNode_Int_3QNone_Int_1_bufchan_buf :
                                                         lizzieLet12_6QNode_Int_3QNone_Int_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNode_Int_3QNone_Int_1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet12_6QNode_Int_3QNone_Int_1_argbuf_r && lizzieLet12_6QNode_Int_3QNone_Int_1_bufchan_buf[0]))
        lizzieLet12_6QNode_Int_3QNone_Int_1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet12_6QNode_Int_3QNone_Int_1_argbuf_r) && (! lizzieLet12_6QNode_Int_3QNone_Int_1_bufchan_buf[0])))
        lizzieLet12_6QNode_Int_3QNone_Int_1_bufchan_buf <= lizzieLet12_6QNode_Int_3QNone_Int_1_bufchan_d;
  
  /* dcon (Ty TupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int,
      Dcon TupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int) : [(lizzieLet12_6QNode_Int_3QNone_Int_1_argbuf,Go),
                                                                      (lizzieLet12_6QNode_Int_12QNone_Int_1_argbuf,Pointer_QTree_Int),
                                                                      (lizzieLet12_6QNode_Int_5QNone_Int_1_argbuf,MyDTInt_Bool),
                                                                      (lizzieLet12_6QNode_Int_7QNone_Int_1_argbuf,MyDTInt_Int)] > (f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int5,TupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int) */
  assign \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int5_d  = TupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_dc((& {lizzieLet12_6QNode_Int_3QNone_Int_1_argbuf_d[0],
                                                                                                                                                                lizzieLet12_6QNode_Int_12QNone_Int_1_argbuf_d[0],
                                                                                                                                                                lizzieLet12_6QNode_Int_5QNone_Int_1_argbuf_d[0],
                                                                                                                                                                lizzieLet12_6QNode_Int_7QNone_Int_1_argbuf_d[0]}), lizzieLet12_6QNode_Int_3QNone_Int_1_argbuf_d, lizzieLet12_6QNode_Int_12QNone_Int_1_argbuf_d, lizzieLet12_6QNode_Int_5QNone_Int_1_argbuf_d, lizzieLet12_6QNode_Int_7QNone_Int_1_argbuf_d);
  assign {lizzieLet12_6QNode_Int_3QNone_Int_1_argbuf_r,
          lizzieLet12_6QNode_Int_12QNone_Int_1_argbuf_r,
          lizzieLet12_6QNode_Int_5QNone_Int_1_argbuf_r,
          lizzieLet12_6QNode_Int_7QNone_Int_1_argbuf_r} = {4 {(\f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int5_r  && \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int5_d [0])}};
  
  /* buf (Ty Go) : (lizzieLet12_6QNode_Int_3QNone_Int_2,Go) > (lizzieLet12_6QNode_Int_3QNone_Int_2_argbuf,Go) */
  Go_t lizzieLet12_6QNode_Int_3QNone_Int_2_bufchan_d;
  logic lizzieLet12_6QNode_Int_3QNone_Int_2_bufchan_r;
  assign lizzieLet12_6QNode_Int_3QNone_Int_2_r = ((! lizzieLet12_6QNode_Int_3QNone_Int_2_bufchan_d[0]) || lizzieLet12_6QNode_Int_3QNone_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNode_Int_3QNone_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet12_6QNode_Int_3QNone_Int_2_r)
        lizzieLet12_6QNode_Int_3QNone_Int_2_bufchan_d <= lizzieLet12_6QNode_Int_3QNone_Int_2_d;
  Go_t lizzieLet12_6QNode_Int_3QNone_Int_2_bufchan_buf;
  assign lizzieLet12_6QNode_Int_3QNone_Int_2_bufchan_r = (! lizzieLet12_6QNode_Int_3QNone_Int_2_bufchan_buf[0]);
  assign lizzieLet12_6QNode_Int_3QNone_Int_2_argbuf_d = (lizzieLet12_6QNode_Int_3QNone_Int_2_bufchan_buf[0] ? lizzieLet12_6QNode_Int_3QNone_Int_2_bufchan_buf :
                                                         lizzieLet12_6QNode_Int_3QNone_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNode_Int_3QNone_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet12_6QNode_Int_3QNone_Int_2_argbuf_r && lizzieLet12_6QNode_Int_3QNone_Int_2_bufchan_buf[0]))
        lizzieLet12_6QNode_Int_3QNone_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet12_6QNode_Int_3QNone_Int_2_argbuf_r) && (! lizzieLet12_6QNode_Int_3QNone_Int_2_bufchan_buf[0])))
        lizzieLet12_6QNode_Int_3QNone_Int_2_bufchan_buf <= lizzieLet12_6QNode_Int_3QNone_Int_2_bufchan_d;
  
  /* dcon (Ty TupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int,
      Dcon TupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int) : [(lizzieLet12_6QNode_Int_3QNone_Int_2_argbuf,Go),
                                                                      (lizzieLet12_6QNode_Int_11QNone_Int_1_argbuf,Pointer_QTree_Int),
                                                                      (lizzieLet12_6QNode_Int_5QNone_Int_2_argbuf,MyDTInt_Bool),
                                                                      (lizzieLet12_6QNode_Int_7QNone_Int_2_argbuf,MyDTInt_Int)] > (f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int6,TupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int) */
  assign \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int6_d  = TupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_dc((& {lizzieLet12_6QNode_Int_3QNone_Int_2_argbuf_d[0],
                                                                                                                                                                lizzieLet12_6QNode_Int_11QNone_Int_1_argbuf_d[0],
                                                                                                                                                                lizzieLet12_6QNode_Int_5QNone_Int_2_argbuf_d[0],
                                                                                                                                                                lizzieLet12_6QNode_Int_7QNone_Int_2_argbuf_d[0]}), lizzieLet12_6QNode_Int_3QNone_Int_2_argbuf_d, lizzieLet12_6QNode_Int_11QNone_Int_1_argbuf_d, lizzieLet12_6QNode_Int_5QNone_Int_2_argbuf_d, lizzieLet12_6QNode_Int_7QNone_Int_2_argbuf_d);
  assign {lizzieLet12_6QNode_Int_3QNone_Int_2_argbuf_r,
          lizzieLet12_6QNode_Int_11QNone_Int_1_argbuf_r,
          lizzieLet12_6QNode_Int_5QNone_Int_2_argbuf_r,
          lizzieLet12_6QNode_Int_7QNone_Int_2_argbuf_r} = {4 {(\f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int6_r  && \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int6_d [0])}};
  
  /* buf (Ty Go) : (lizzieLet12_6QNode_Int_3QNone_Int_3,Go) > (lizzieLet12_6QNode_Int_3QNone_Int_3_argbuf,Go) */
  Go_t lizzieLet12_6QNode_Int_3QNone_Int_3_bufchan_d;
  logic lizzieLet12_6QNode_Int_3QNone_Int_3_bufchan_r;
  assign lizzieLet12_6QNode_Int_3QNone_Int_3_r = ((! lizzieLet12_6QNode_Int_3QNone_Int_3_bufchan_d[0]) || lizzieLet12_6QNode_Int_3QNone_Int_3_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNode_Int_3QNone_Int_3_bufchan_d <= 1'd0;
    else
      if (lizzieLet12_6QNode_Int_3QNone_Int_3_r)
        lizzieLet12_6QNode_Int_3QNone_Int_3_bufchan_d <= lizzieLet12_6QNode_Int_3QNone_Int_3_d;
  Go_t lizzieLet12_6QNode_Int_3QNone_Int_3_bufchan_buf;
  assign lizzieLet12_6QNode_Int_3QNone_Int_3_bufchan_r = (! lizzieLet12_6QNode_Int_3QNone_Int_3_bufchan_buf[0]);
  assign lizzieLet12_6QNode_Int_3QNone_Int_3_argbuf_d = (lizzieLet12_6QNode_Int_3QNone_Int_3_bufchan_buf[0] ? lizzieLet12_6QNode_Int_3QNone_Int_3_bufchan_buf :
                                                         lizzieLet12_6QNode_Int_3QNone_Int_3_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNode_Int_3QNone_Int_3_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet12_6QNode_Int_3QNone_Int_3_argbuf_r && lizzieLet12_6QNode_Int_3QNone_Int_3_bufchan_buf[0]))
        lizzieLet12_6QNode_Int_3QNone_Int_3_bufchan_buf <= 1'd0;
      else if (((! lizzieLet12_6QNode_Int_3QNone_Int_3_argbuf_r) && (! lizzieLet12_6QNode_Int_3QNone_Int_3_bufchan_buf[0])))
        lizzieLet12_6QNode_Int_3QNone_Int_3_bufchan_buf <= lizzieLet12_6QNode_Int_3QNone_Int_3_bufchan_d;
  
  /* dcon (Ty TupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int,
      Dcon TupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int) : [(lizzieLet12_6QNode_Int_3QNone_Int_3_argbuf,Go),
                                                                      (lizzieLet12_6QNode_Int_10QNone_Int_1_argbuf,Pointer_QTree_Int),
                                                                      (lizzieLet12_6QNode_Int_5QNone_Int_3_argbuf,MyDTInt_Bool),
                                                                      (lizzieLet12_6QNode_Int_7QNone_Int_3_argbuf,MyDTInt_Int)] > (f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int7,TupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int) */
  assign \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int7_d  = TupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_dc((& {lizzieLet12_6QNode_Int_3QNone_Int_3_argbuf_d[0],
                                                                                                                                                                lizzieLet12_6QNode_Int_10QNone_Int_1_argbuf_d[0],
                                                                                                                                                                lizzieLet12_6QNode_Int_5QNone_Int_3_argbuf_d[0],
                                                                                                                                                                lizzieLet12_6QNode_Int_7QNone_Int_3_argbuf_d[0]}), lizzieLet12_6QNode_Int_3QNone_Int_3_argbuf_d, lizzieLet12_6QNode_Int_10QNone_Int_1_argbuf_d, lizzieLet12_6QNode_Int_5QNone_Int_3_argbuf_d, lizzieLet12_6QNode_Int_7QNone_Int_3_argbuf_d);
  assign {lizzieLet12_6QNode_Int_3QNone_Int_3_argbuf_r,
          lizzieLet12_6QNode_Int_10QNone_Int_1_argbuf_r,
          lizzieLet12_6QNode_Int_5QNone_Int_3_argbuf_r,
          lizzieLet12_6QNode_Int_7QNone_Int_3_argbuf_r} = {4 {(\f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int7_r  && \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int7_d [0])}};
  
  /* buf (Ty Go) : (lizzieLet12_6QNode_Int_3QNone_Int_4,Go) > (lizzieLet12_6QNode_Int_3QNone_Int_4_argbuf,Go) */
  Go_t lizzieLet12_6QNode_Int_3QNone_Int_4_bufchan_d;
  logic lizzieLet12_6QNode_Int_3QNone_Int_4_bufchan_r;
  assign lizzieLet12_6QNode_Int_3QNone_Int_4_r = ((! lizzieLet12_6QNode_Int_3QNone_Int_4_bufchan_d[0]) || lizzieLet12_6QNode_Int_3QNone_Int_4_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNode_Int_3QNone_Int_4_bufchan_d <= 1'd0;
    else
      if (lizzieLet12_6QNode_Int_3QNone_Int_4_r)
        lizzieLet12_6QNode_Int_3QNone_Int_4_bufchan_d <= lizzieLet12_6QNode_Int_3QNone_Int_4_d;
  Go_t lizzieLet12_6QNode_Int_3QNone_Int_4_bufchan_buf;
  assign lizzieLet12_6QNode_Int_3QNone_Int_4_bufchan_r = (! lizzieLet12_6QNode_Int_3QNone_Int_4_bufchan_buf[0]);
  assign lizzieLet12_6QNode_Int_3QNone_Int_4_argbuf_d = (lizzieLet12_6QNode_Int_3QNone_Int_4_bufchan_buf[0] ? lizzieLet12_6QNode_Int_3QNone_Int_4_bufchan_buf :
                                                         lizzieLet12_6QNode_Int_3QNone_Int_4_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNode_Int_3QNone_Int_4_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet12_6QNode_Int_3QNone_Int_4_argbuf_r && lizzieLet12_6QNode_Int_3QNone_Int_4_bufchan_buf[0]))
        lizzieLet12_6QNode_Int_3QNone_Int_4_bufchan_buf <= 1'd0;
      else if (((! lizzieLet12_6QNode_Int_3QNone_Int_4_argbuf_r) && (! lizzieLet12_6QNode_Int_3QNone_Int_4_bufchan_buf[0])))
        lizzieLet12_6QNode_Int_3QNone_Int_4_bufchan_buf <= lizzieLet12_6QNode_Int_3QNone_Int_4_bufchan_d;
  
  /* dcon (Ty TupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int,
      Dcon TupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int) : [(lizzieLet12_6QNode_Int_3QNone_Int_4_argbuf,Go),
                                                                      (lizzieLet12_6QNode_Int_9QNone_Int_1_argbuf,Pointer_QTree_Int),
                                                                      (lizzieLet12_6QNode_Int_5QNone_Int_4_argbuf,MyDTInt_Bool),
                                                                      (lizzieLet12_6QNode_Int_7QNone_Int_4_argbuf,MyDTInt_Int)] > (f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int8,TupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int) */
  assign \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int8_d  = TupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_dc((& {lizzieLet12_6QNode_Int_3QNone_Int_4_argbuf_d[0],
                                                                                                                                                                lizzieLet12_6QNode_Int_9QNone_Int_1_argbuf_d[0],
                                                                                                                                                                lizzieLet12_6QNode_Int_5QNone_Int_4_argbuf_d[0],
                                                                                                                                                                lizzieLet12_6QNode_Int_7QNone_Int_4_argbuf_d[0]}), lizzieLet12_6QNode_Int_3QNone_Int_4_argbuf_d, lizzieLet12_6QNode_Int_9QNone_Int_1_argbuf_d, lizzieLet12_6QNode_Int_5QNone_Int_4_argbuf_d, lizzieLet12_6QNode_Int_7QNone_Int_4_argbuf_d);
  assign {lizzieLet12_6QNode_Int_3QNone_Int_4_argbuf_r,
          lizzieLet12_6QNode_Int_9QNone_Int_1_argbuf_r,
          lizzieLet12_6QNode_Int_5QNone_Int_4_argbuf_r,
          lizzieLet12_6QNode_Int_7QNone_Int_4_argbuf_r} = {4 {(\f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int8_r  && \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int8_d [0])}};
  
  /* buf (Ty Go) : (lizzieLet12_6QNode_Int_3QNone_Int_5,Go) > (lizzieLet12_6QNode_Int_3QNone_Int_5_argbuf,Go) */
  Go_t lizzieLet12_6QNode_Int_3QNone_Int_5_bufchan_d;
  logic lizzieLet12_6QNode_Int_3QNone_Int_5_bufchan_r;
  assign lizzieLet12_6QNode_Int_3QNone_Int_5_r = ((! lizzieLet12_6QNode_Int_3QNone_Int_5_bufchan_d[0]) || lizzieLet12_6QNode_Int_3QNone_Int_5_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNode_Int_3QNone_Int_5_bufchan_d <= 1'd0;
    else
      if (lizzieLet12_6QNode_Int_3QNone_Int_5_r)
        lizzieLet12_6QNode_Int_3QNone_Int_5_bufchan_d <= lizzieLet12_6QNode_Int_3QNone_Int_5_d;
  Go_t lizzieLet12_6QNode_Int_3QNone_Int_5_bufchan_buf;
  assign lizzieLet12_6QNode_Int_3QNone_Int_5_bufchan_r = (! lizzieLet12_6QNode_Int_3QNone_Int_5_bufchan_buf[0]);
  assign lizzieLet12_6QNode_Int_3QNone_Int_5_argbuf_d = (lizzieLet12_6QNode_Int_3QNone_Int_5_bufchan_buf[0] ? lizzieLet12_6QNode_Int_3QNone_Int_5_bufchan_buf :
                                                         lizzieLet12_6QNode_Int_3QNone_Int_5_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNode_Int_3QNone_Int_5_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet12_6QNode_Int_3QNone_Int_5_argbuf_r && lizzieLet12_6QNode_Int_3QNone_Int_5_bufchan_buf[0]))
        lizzieLet12_6QNode_Int_3QNone_Int_5_bufchan_buf <= 1'd0;
      else if (((! lizzieLet12_6QNode_Int_3QNone_Int_5_argbuf_r) && (! lizzieLet12_6QNode_Int_3QNone_Int_5_bufchan_buf[0])))
        lizzieLet12_6QNode_Int_3QNone_Int_5_bufchan_buf <= lizzieLet12_6QNode_Int_3QNone_Int_5_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet12_6QNode_Int_3QVal_Int,Go) > [(lizzieLet12_6QNode_Int_3QVal_Int_1,Go),
                                                        (lizzieLet12_6QNode_Int_3QVal_Int_2,Go)] */
  logic [1:0] lizzieLet12_6QNode_Int_3QVal_Int_emitted;
  logic [1:0] lizzieLet12_6QNode_Int_3QVal_Int_done;
  assign lizzieLet12_6QNode_Int_3QVal_Int_1_d = (lizzieLet12_6QNode_Int_3QVal_Int_d[0] && (! lizzieLet12_6QNode_Int_3QVal_Int_emitted[0]));
  assign lizzieLet12_6QNode_Int_3QVal_Int_2_d = (lizzieLet12_6QNode_Int_3QVal_Int_d[0] && (! lizzieLet12_6QNode_Int_3QVal_Int_emitted[1]));
  assign lizzieLet12_6QNode_Int_3QVal_Int_done = (lizzieLet12_6QNode_Int_3QVal_Int_emitted | ({lizzieLet12_6QNode_Int_3QVal_Int_2_d[0],
                                                                                               lizzieLet12_6QNode_Int_3QVal_Int_1_d[0]} & {lizzieLet12_6QNode_Int_3QVal_Int_2_r,
                                                                                                                                           lizzieLet12_6QNode_Int_3QVal_Int_1_r}));
  assign lizzieLet12_6QNode_Int_3QVal_Int_r = (& lizzieLet12_6QNode_Int_3QVal_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNode_Int_3QVal_Int_emitted <= 2'd0;
    else
      lizzieLet12_6QNode_Int_3QVal_Int_emitted <= (lizzieLet12_6QNode_Int_3QVal_Int_r ? 2'd0 :
                                                   lizzieLet12_6QNode_Int_3QVal_Int_done);
  
  /* dcon (Ty QTree_Int,
      Dcon QError_Int) : [(lizzieLet12_6QNode_Int_3QVal_Int_1,Go)] > (lizzieLet12_6QNode_Int_3QVal_Int_1QError_Int,QTree_Int) */
  assign lizzieLet12_6QNode_Int_3QVal_Int_1QError_Int_d = QError_Int_dc((& {lizzieLet12_6QNode_Int_3QVal_Int_1_d[0]}), lizzieLet12_6QNode_Int_3QVal_Int_1_d);
  assign {lizzieLet12_6QNode_Int_3QVal_Int_1_r} = {1 {(lizzieLet12_6QNode_Int_3QVal_Int_1QError_Int_r && lizzieLet12_6QNode_Int_3QVal_Int_1QError_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (lizzieLet12_6QNode_Int_3QVal_Int_1QError_Int,QTree_Int) > (lizzieLet29_1_argbuf,QTree_Int) */
  QTree_Int_t lizzieLet12_6QNode_Int_3QVal_Int_1QError_Int_bufchan_d;
  logic lizzieLet12_6QNode_Int_3QVal_Int_1QError_Int_bufchan_r;
  assign lizzieLet12_6QNode_Int_3QVal_Int_1QError_Int_r = ((! lizzieLet12_6QNode_Int_3QVal_Int_1QError_Int_bufchan_d[0]) || lizzieLet12_6QNode_Int_3QVal_Int_1QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNode_Int_3QVal_Int_1QError_Int_bufchan_d <= {66'd0,
                                                                 1'd0};
    else
      if (lizzieLet12_6QNode_Int_3QVal_Int_1QError_Int_r)
        lizzieLet12_6QNode_Int_3QVal_Int_1QError_Int_bufchan_d <= lizzieLet12_6QNode_Int_3QVal_Int_1QError_Int_d;
  QTree_Int_t lizzieLet12_6QNode_Int_3QVal_Int_1QError_Int_bufchan_buf;
  assign lizzieLet12_6QNode_Int_3QVal_Int_1QError_Int_bufchan_r = (! lizzieLet12_6QNode_Int_3QVal_Int_1QError_Int_bufchan_buf[0]);
  assign lizzieLet29_1_argbuf_d = (lizzieLet12_6QNode_Int_3QVal_Int_1QError_Int_bufchan_buf[0] ? lizzieLet12_6QNode_Int_3QVal_Int_1QError_Int_bufchan_buf :
                                   lizzieLet12_6QNode_Int_3QVal_Int_1QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNode_Int_3QVal_Int_1QError_Int_bufchan_buf <= {66'd0,
                                                                   1'd0};
    else
      if ((lizzieLet29_1_argbuf_r && lizzieLet12_6QNode_Int_3QVal_Int_1QError_Int_bufchan_buf[0]))
        lizzieLet12_6QNode_Int_3QVal_Int_1QError_Int_bufchan_buf <= {66'd0,
                                                                     1'd0};
      else if (((! lizzieLet29_1_argbuf_r) && (! lizzieLet12_6QNode_Int_3QVal_Int_1QError_Int_bufchan_buf[0])))
        lizzieLet12_6QNode_Int_3QVal_Int_1QError_Int_bufchan_buf <= lizzieLet12_6QNode_Int_3QVal_Int_1QError_Int_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet12_6QNode_Int_3QVal_Int_2,Go) > (lizzieLet12_6QNode_Int_3QVal_Int_2_argbuf,Go) */
  Go_t lizzieLet12_6QNode_Int_3QVal_Int_2_bufchan_d;
  logic lizzieLet12_6QNode_Int_3QVal_Int_2_bufchan_r;
  assign lizzieLet12_6QNode_Int_3QVal_Int_2_r = ((! lizzieLet12_6QNode_Int_3QVal_Int_2_bufchan_d[0]) || lizzieLet12_6QNode_Int_3QVal_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNode_Int_3QVal_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet12_6QNode_Int_3QVal_Int_2_r)
        lizzieLet12_6QNode_Int_3QVal_Int_2_bufchan_d <= lizzieLet12_6QNode_Int_3QVal_Int_2_d;
  Go_t lizzieLet12_6QNode_Int_3QVal_Int_2_bufchan_buf;
  assign lizzieLet12_6QNode_Int_3QVal_Int_2_bufchan_r = (! lizzieLet12_6QNode_Int_3QVal_Int_2_bufchan_buf[0]);
  assign lizzieLet12_6QNode_Int_3QVal_Int_2_argbuf_d = (lizzieLet12_6QNode_Int_3QVal_Int_2_bufchan_buf[0] ? lizzieLet12_6QNode_Int_3QVal_Int_2_bufchan_buf :
                                                        lizzieLet12_6QNode_Int_3QVal_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNode_Int_3QVal_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet12_6QNode_Int_3QVal_Int_2_argbuf_r && lizzieLet12_6QNode_Int_3QVal_Int_2_bufchan_buf[0]))
        lizzieLet12_6QNode_Int_3QVal_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet12_6QNode_Int_3QVal_Int_2_argbuf_r) && (! lizzieLet12_6QNode_Int_3QVal_Int_2_bufchan_buf[0])))
        lizzieLet12_6QNode_Int_3QVal_Int_2_bufchan_buf <= lizzieLet12_6QNode_Int_3QVal_Int_2_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty MyDTInt_Bool) : (lizzieLet12_6QNode_Int_4,QTree_Int) (lizzieLet12_4QNode_Int,MyDTInt_Bool) > [(_50,MyDTInt_Bool),
                                                                                                        (_49,MyDTInt_Bool),
                                                                                                        (lizzieLet12_6QNode_Int_4QNode_Int,MyDTInt_Bool),
                                                                                                        (_48,MyDTInt_Bool)] */
  logic [3:0] lizzieLet12_4QNode_Int_onehotd;
  always_comb
    if ((lizzieLet12_6QNode_Int_4_d[0] && lizzieLet12_4QNode_Int_d[0]))
      unique case (lizzieLet12_6QNode_Int_4_d[2:1])
        2'd0: lizzieLet12_4QNode_Int_onehotd = 4'd1;
        2'd1: lizzieLet12_4QNode_Int_onehotd = 4'd2;
        2'd2: lizzieLet12_4QNode_Int_onehotd = 4'd4;
        2'd3: lizzieLet12_4QNode_Int_onehotd = 4'd8;
        default: lizzieLet12_4QNode_Int_onehotd = 4'd0;
      endcase
    else lizzieLet12_4QNode_Int_onehotd = 4'd0;
  assign _50_d = lizzieLet12_4QNode_Int_onehotd[0];
  assign _49_d = lizzieLet12_4QNode_Int_onehotd[1];
  assign lizzieLet12_6QNode_Int_4QNode_Int_d = lizzieLet12_4QNode_Int_onehotd[2];
  assign _48_d = lizzieLet12_4QNode_Int_onehotd[3];
  assign lizzieLet12_4QNode_Int_r = (| (lizzieLet12_4QNode_Int_onehotd & {_48_r,
                                                                          lizzieLet12_6QNode_Int_4QNode_Int_r,
                                                                          _49_r,
                                                                          _50_r}));
  assign lizzieLet12_6QNode_Int_4_r = lizzieLet12_4QNode_Int_r;
  
  /* fork (Ty MyDTInt_Bool) : (lizzieLet12_6QNode_Int_4QNode_Int,MyDTInt_Bool) > [(lizzieLet12_6QNode_Int_4QNode_Int_1,MyDTInt_Bool),
                                                                             (lizzieLet12_6QNode_Int_4QNode_Int_2,MyDTInt_Bool)] */
  logic [1:0] lizzieLet12_6QNode_Int_4QNode_Int_emitted;
  logic [1:0] lizzieLet12_6QNode_Int_4QNode_Int_done;
  assign lizzieLet12_6QNode_Int_4QNode_Int_1_d = (lizzieLet12_6QNode_Int_4QNode_Int_d[0] && (! lizzieLet12_6QNode_Int_4QNode_Int_emitted[0]));
  assign lizzieLet12_6QNode_Int_4QNode_Int_2_d = (lizzieLet12_6QNode_Int_4QNode_Int_d[0] && (! lizzieLet12_6QNode_Int_4QNode_Int_emitted[1]));
  assign lizzieLet12_6QNode_Int_4QNode_Int_done = (lizzieLet12_6QNode_Int_4QNode_Int_emitted | ({lizzieLet12_6QNode_Int_4QNode_Int_2_d[0],
                                                                                                 lizzieLet12_6QNode_Int_4QNode_Int_1_d[0]} & {lizzieLet12_6QNode_Int_4QNode_Int_2_r,
                                                                                                                                              lizzieLet12_6QNode_Int_4QNode_Int_1_r}));
  assign lizzieLet12_6QNode_Int_4QNode_Int_r = (& lizzieLet12_6QNode_Int_4QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNode_Int_4QNode_Int_emitted <= 2'd0;
    else
      lizzieLet12_6QNode_Int_4QNode_Int_emitted <= (lizzieLet12_6QNode_Int_4QNode_Int_r ? 2'd0 :
                                                    lizzieLet12_6QNode_Int_4QNode_Int_done);
  
  /* buf (Ty MyDTInt_Bool) : (lizzieLet12_6QNode_Int_4QNode_Int_2,MyDTInt_Bool) > (lizzieLet12_6QNode_Int_4QNode_Int_2_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t lizzieLet12_6QNode_Int_4QNode_Int_2_bufchan_d;
  logic lizzieLet12_6QNode_Int_4QNode_Int_2_bufchan_r;
  assign lizzieLet12_6QNode_Int_4QNode_Int_2_r = ((! lizzieLet12_6QNode_Int_4QNode_Int_2_bufchan_d[0]) || lizzieLet12_6QNode_Int_4QNode_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNode_Int_4QNode_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet12_6QNode_Int_4QNode_Int_2_r)
        lizzieLet12_6QNode_Int_4QNode_Int_2_bufchan_d <= lizzieLet12_6QNode_Int_4QNode_Int_2_d;
  MyDTInt_Bool_t lizzieLet12_6QNode_Int_4QNode_Int_2_bufchan_buf;
  assign lizzieLet12_6QNode_Int_4QNode_Int_2_bufchan_r = (! lizzieLet12_6QNode_Int_4QNode_Int_2_bufchan_buf[0]);
  assign lizzieLet12_6QNode_Int_4QNode_Int_2_argbuf_d = (lizzieLet12_6QNode_Int_4QNode_Int_2_bufchan_buf[0] ? lizzieLet12_6QNode_Int_4QNode_Int_2_bufchan_buf :
                                                         lizzieLet12_6QNode_Int_4QNode_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNode_Int_4QNode_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet12_6QNode_Int_4QNode_Int_2_argbuf_r && lizzieLet12_6QNode_Int_4QNode_Int_2_bufchan_buf[0]))
        lizzieLet12_6QNode_Int_4QNode_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet12_6QNode_Int_4QNode_Int_2_argbuf_r) && (! lizzieLet12_6QNode_Int_4QNode_Int_2_bufchan_buf[0])))
        lizzieLet12_6QNode_Int_4QNode_Int_2_bufchan_buf <= lizzieLet12_6QNode_Int_4QNode_Int_2_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty MyDTInt_Bool) : (lizzieLet12_6QNode_Int_5,QTree_Int) (lizzieLet12_5QNode_Int,MyDTInt_Bool) > [(lizzieLet12_6QNode_Int_5QNone_Int,MyDTInt_Bool),
                                                                                                        (_47,MyDTInt_Bool),
                                                                                                        (lizzieLet12_6QNode_Int_5QNode_Int,MyDTInt_Bool),
                                                                                                        (_46,MyDTInt_Bool)] */
  logic [3:0] lizzieLet12_5QNode_Int_onehotd;
  always_comb
    if ((lizzieLet12_6QNode_Int_5_d[0] && lizzieLet12_5QNode_Int_d[0]))
      unique case (lizzieLet12_6QNode_Int_5_d[2:1])
        2'd0: lizzieLet12_5QNode_Int_onehotd = 4'd1;
        2'd1: lizzieLet12_5QNode_Int_onehotd = 4'd2;
        2'd2: lizzieLet12_5QNode_Int_onehotd = 4'd4;
        2'd3: lizzieLet12_5QNode_Int_onehotd = 4'd8;
        default: lizzieLet12_5QNode_Int_onehotd = 4'd0;
      endcase
    else lizzieLet12_5QNode_Int_onehotd = 4'd0;
  assign lizzieLet12_6QNode_Int_5QNone_Int_d = lizzieLet12_5QNode_Int_onehotd[0];
  assign _47_d = lizzieLet12_5QNode_Int_onehotd[1];
  assign lizzieLet12_6QNode_Int_5QNode_Int_d = lizzieLet12_5QNode_Int_onehotd[2];
  assign _46_d = lizzieLet12_5QNode_Int_onehotd[3];
  assign lizzieLet12_5QNode_Int_r = (| (lizzieLet12_5QNode_Int_onehotd & {_46_r,
                                                                          lizzieLet12_6QNode_Int_5QNode_Int_r,
                                                                          _47_r,
                                                                          lizzieLet12_6QNode_Int_5QNone_Int_r}));
  assign lizzieLet12_6QNode_Int_5_r = lizzieLet12_5QNode_Int_r;
  
  /* fork (Ty MyDTInt_Bool) : (lizzieLet12_6QNode_Int_5QNode_Int,MyDTInt_Bool) > [(lizzieLet12_6QNode_Int_5QNode_Int_1,MyDTInt_Bool),
                                                                             (lizzieLet12_6QNode_Int_5QNode_Int_2,MyDTInt_Bool)] */
  logic [1:0] lizzieLet12_6QNode_Int_5QNode_Int_emitted;
  logic [1:0] lizzieLet12_6QNode_Int_5QNode_Int_done;
  assign lizzieLet12_6QNode_Int_5QNode_Int_1_d = (lizzieLet12_6QNode_Int_5QNode_Int_d[0] && (! lizzieLet12_6QNode_Int_5QNode_Int_emitted[0]));
  assign lizzieLet12_6QNode_Int_5QNode_Int_2_d = (lizzieLet12_6QNode_Int_5QNode_Int_d[0] && (! lizzieLet12_6QNode_Int_5QNode_Int_emitted[1]));
  assign lizzieLet12_6QNode_Int_5QNode_Int_done = (lizzieLet12_6QNode_Int_5QNode_Int_emitted | ({lizzieLet12_6QNode_Int_5QNode_Int_2_d[0],
                                                                                                 lizzieLet12_6QNode_Int_5QNode_Int_1_d[0]} & {lizzieLet12_6QNode_Int_5QNode_Int_2_r,
                                                                                                                                              lizzieLet12_6QNode_Int_5QNode_Int_1_r}));
  assign lizzieLet12_6QNode_Int_5QNode_Int_r = (& lizzieLet12_6QNode_Int_5QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNode_Int_5QNode_Int_emitted <= 2'd0;
    else
      lizzieLet12_6QNode_Int_5QNode_Int_emitted <= (lizzieLet12_6QNode_Int_5QNode_Int_r ? 2'd0 :
                                                    lizzieLet12_6QNode_Int_5QNode_Int_done);
  
  /* buf (Ty MyDTInt_Bool) : (lizzieLet12_6QNode_Int_5QNode_Int_2,MyDTInt_Bool) > (lizzieLet12_6QNode_Int_5QNode_Int_2_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t lizzieLet12_6QNode_Int_5QNode_Int_2_bufchan_d;
  logic lizzieLet12_6QNode_Int_5QNode_Int_2_bufchan_r;
  assign lizzieLet12_6QNode_Int_5QNode_Int_2_r = ((! lizzieLet12_6QNode_Int_5QNode_Int_2_bufchan_d[0]) || lizzieLet12_6QNode_Int_5QNode_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNode_Int_5QNode_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet12_6QNode_Int_5QNode_Int_2_r)
        lizzieLet12_6QNode_Int_5QNode_Int_2_bufchan_d <= lizzieLet12_6QNode_Int_5QNode_Int_2_d;
  MyDTInt_Bool_t lizzieLet12_6QNode_Int_5QNode_Int_2_bufchan_buf;
  assign lizzieLet12_6QNode_Int_5QNode_Int_2_bufchan_r = (! lizzieLet12_6QNode_Int_5QNode_Int_2_bufchan_buf[0]);
  assign lizzieLet12_6QNode_Int_5QNode_Int_2_argbuf_d = (lizzieLet12_6QNode_Int_5QNode_Int_2_bufchan_buf[0] ? lizzieLet12_6QNode_Int_5QNode_Int_2_bufchan_buf :
                                                         lizzieLet12_6QNode_Int_5QNode_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNode_Int_5QNode_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet12_6QNode_Int_5QNode_Int_2_argbuf_r && lizzieLet12_6QNode_Int_5QNode_Int_2_bufchan_buf[0]))
        lizzieLet12_6QNode_Int_5QNode_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet12_6QNode_Int_5QNode_Int_2_argbuf_r) && (! lizzieLet12_6QNode_Int_5QNode_Int_2_bufchan_buf[0])))
        lizzieLet12_6QNode_Int_5QNode_Int_2_bufchan_buf <= lizzieLet12_6QNode_Int_5QNode_Int_2_bufchan_d;
  
  /* fork (Ty MyDTInt_Bool) : (lizzieLet12_6QNode_Int_5QNone_Int,MyDTInt_Bool) > [(lizzieLet12_6QNode_Int_5QNone_Int_1,MyDTInt_Bool),
                                                                             (lizzieLet12_6QNode_Int_5QNone_Int_2,MyDTInt_Bool),
                                                                             (lizzieLet12_6QNode_Int_5QNone_Int_3,MyDTInt_Bool),
                                                                             (lizzieLet12_6QNode_Int_5QNone_Int_4,MyDTInt_Bool)] */
  logic [3:0] lizzieLet12_6QNode_Int_5QNone_Int_emitted;
  logic [3:0] lizzieLet12_6QNode_Int_5QNone_Int_done;
  assign lizzieLet12_6QNode_Int_5QNone_Int_1_d = (lizzieLet12_6QNode_Int_5QNone_Int_d[0] && (! lizzieLet12_6QNode_Int_5QNone_Int_emitted[0]));
  assign lizzieLet12_6QNode_Int_5QNone_Int_2_d = (lizzieLet12_6QNode_Int_5QNone_Int_d[0] && (! lizzieLet12_6QNode_Int_5QNone_Int_emitted[1]));
  assign lizzieLet12_6QNode_Int_5QNone_Int_3_d = (lizzieLet12_6QNode_Int_5QNone_Int_d[0] && (! lizzieLet12_6QNode_Int_5QNone_Int_emitted[2]));
  assign lizzieLet12_6QNode_Int_5QNone_Int_4_d = (lizzieLet12_6QNode_Int_5QNone_Int_d[0] && (! lizzieLet12_6QNode_Int_5QNone_Int_emitted[3]));
  assign lizzieLet12_6QNode_Int_5QNone_Int_done = (lizzieLet12_6QNode_Int_5QNone_Int_emitted | ({lizzieLet12_6QNode_Int_5QNone_Int_4_d[0],
                                                                                                 lizzieLet12_6QNode_Int_5QNone_Int_3_d[0],
                                                                                                 lizzieLet12_6QNode_Int_5QNone_Int_2_d[0],
                                                                                                 lizzieLet12_6QNode_Int_5QNone_Int_1_d[0]} & {lizzieLet12_6QNode_Int_5QNone_Int_4_r,
                                                                                                                                              lizzieLet12_6QNode_Int_5QNone_Int_3_r,
                                                                                                                                              lizzieLet12_6QNode_Int_5QNone_Int_2_r,
                                                                                                                                              lizzieLet12_6QNode_Int_5QNone_Int_1_r}));
  assign lizzieLet12_6QNode_Int_5QNone_Int_r = (& lizzieLet12_6QNode_Int_5QNone_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNode_Int_5QNone_Int_emitted <= 4'd0;
    else
      lizzieLet12_6QNode_Int_5QNone_Int_emitted <= (lizzieLet12_6QNode_Int_5QNone_Int_r ? 4'd0 :
                                                    lizzieLet12_6QNode_Int_5QNone_Int_done);
  
  /* buf (Ty MyDTInt_Bool) : (lizzieLet12_6QNode_Int_5QNone_Int_1,MyDTInt_Bool) > (lizzieLet12_6QNode_Int_5QNone_Int_1_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t lizzieLet12_6QNode_Int_5QNone_Int_1_bufchan_d;
  logic lizzieLet12_6QNode_Int_5QNone_Int_1_bufchan_r;
  assign lizzieLet12_6QNode_Int_5QNone_Int_1_r = ((! lizzieLet12_6QNode_Int_5QNone_Int_1_bufchan_d[0]) || lizzieLet12_6QNode_Int_5QNone_Int_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNode_Int_5QNone_Int_1_bufchan_d <= 1'd0;
    else
      if (lizzieLet12_6QNode_Int_5QNone_Int_1_r)
        lizzieLet12_6QNode_Int_5QNone_Int_1_bufchan_d <= lizzieLet12_6QNode_Int_5QNone_Int_1_d;
  MyDTInt_Bool_t lizzieLet12_6QNode_Int_5QNone_Int_1_bufchan_buf;
  assign lizzieLet12_6QNode_Int_5QNone_Int_1_bufchan_r = (! lizzieLet12_6QNode_Int_5QNone_Int_1_bufchan_buf[0]);
  assign lizzieLet12_6QNode_Int_5QNone_Int_1_argbuf_d = (lizzieLet12_6QNode_Int_5QNone_Int_1_bufchan_buf[0] ? lizzieLet12_6QNode_Int_5QNone_Int_1_bufchan_buf :
                                                         lizzieLet12_6QNode_Int_5QNone_Int_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNode_Int_5QNone_Int_1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet12_6QNode_Int_5QNone_Int_1_argbuf_r && lizzieLet12_6QNode_Int_5QNone_Int_1_bufchan_buf[0]))
        lizzieLet12_6QNode_Int_5QNone_Int_1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet12_6QNode_Int_5QNone_Int_1_argbuf_r) && (! lizzieLet12_6QNode_Int_5QNone_Int_1_bufchan_buf[0])))
        lizzieLet12_6QNode_Int_5QNone_Int_1_bufchan_buf <= lizzieLet12_6QNode_Int_5QNone_Int_1_bufchan_d;
  
  /* buf (Ty MyDTInt_Bool) : (lizzieLet12_6QNode_Int_5QNone_Int_2,MyDTInt_Bool) > (lizzieLet12_6QNode_Int_5QNone_Int_2_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t lizzieLet12_6QNode_Int_5QNone_Int_2_bufchan_d;
  logic lizzieLet12_6QNode_Int_5QNone_Int_2_bufchan_r;
  assign lizzieLet12_6QNode_Int_5QNone_Int_2_r = ((! lizzieLet12_6QNode_Int_5QNone_Int_2_bufchan_d[0]) || lizzieLet12_6QNode_Int_5QNone_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNode_Int_5QNone_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet12_6QNode_Int_5QNone_Int_2_r)
        lizzieLet12_6QNode_Int_5QNone_Int_2_bufchan_d <= lizzieLet12_6QNode_Int_5QNone_Int_2_d;
  MyDTInt_Bool_t lizzieLet12_6QNode_Int_5QNone_Int_2_bufchan_buf;
  assign lizzieLet12_6QNode_Int_5QNone_Int_2_bufchan_r = (! lizzieLet12_6QNode_Int_5QNone_Int_2_bufchan_buf[0]);
  assign lizzieLet12_6QNode_Int_5QNone_Int_2_argbuf_d = (lizzieLet12_6QNode_Int_5QNone_Int_2_bufchan_buf[0] ? lizzieLet12_6QNode_Int_5QNone_Int_2_bufchan_buf :
                                                         lizzieLet12_6QNode_Int_5QNone_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNode_Int_5QNone_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet12_6QNode_Int_5QNone_Int_2_argbuf_r && lizzieLet12_6QNode_Int_5QNone_Int_2_bufchan_buf[0]))
        lizzieLet12_6QNode_Int_5QNone_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet12_6QNode_Int_5QNone_Int_2_argbuf_r) && (! lizzieLet12_6QNode_Int_5QNone_Int_2_bufchan_buf[0])))
        lizzieLet12_6QNode_Int_5QNone_Int_2_bufchan_buf <= lizzieLet12_6QNode_Int_5QNone_Int_2_bufchan_d;
  
  /* buf (Ty MyDTInt_Bool) : (lizzieLet12_6QNode_Int_5QNone_Int_3,MyDTInt_Bool) > (lizzieLet12_6QNode_Int_5QNone_Int_3_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t lizzieLet12_6QNode_Int_5QNone_Int_3_bufchan_d;
  logic lizzieLet12_6QNode_Int_5QNone_Int_3_bufchan_r;
  assign lizzieLet12_6QNode_Int_5QNone_Int_3_r = ((! lizzieLet12_6QNode_Int_5QNone_Int_3_bufchan_d[0]) || lizzieLet12_6QNode_Int_5QNone_Int_3_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNode_Int_5QNone_Int_3_bufchan_d <= 1'd0;
    else
      if (lizzieLet12_6QNode_Int_5QNone_Int_3_r)
        lizzieLet12_6QNode_Int_5QNone_Int_3_bufchan_d <= lizzieLet12_6QNode_Int_5QNone_Int_3_d;
  MyDTInt_Bool_t lizzieLet12_6QNode_Int_5QNone_Int_3_bufchan_buf;
  assign lizzieLet12_6QNode_Int_5QNone_Int_3_bufchan_r = (! lizzieLet12_6QNode_Int_5QNone_Int_3_bufchan_buf[0]);
  assign lizzieLet12_6QNode_Int_5QNone_Int_3_argbuf_d = (lizzieLet12_6QNode_Int_5QNone_Int_3_bufchan_buf[0] ? lizzieLet12_6QNode_Int_5QNone_Int_3_bufchan_buf :
                                                         lizzieLet12_6QNode_Int_5QNone_Int_3_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNode_Int_5QNone_Int_3_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet12_6QNode_Int_5QNone_Int_3_argbuf_r && lizzieLet12_6QNode_Int_5QNone_Int_3_bufchan_buf[0]))
        lizzieLet12_6QNode_Int_5QNone_Int_3_bufchan_buf <= 1'd0;
      else if (((! lizzieLet12_6QNode_Int_5QNone_Int_3_argbuf_r) && (! lizzieLet12_6QNode_Int_5QNone_Int_3_bufchan_buf[0])))
        lizzieLet12_6QNode_Int_5QNone_Int_3_bufchan_buf <= lizzieLet12_6QNode_Int_5QNone_Int_3_bufchan_d;
  
  /* buf (Ty MyDTInt_Bool) : (lizzieLet12_6QNode_Int_5QNone_Int_4,MyDTInt_Bool) > (lizzieLet12_6QNode_Int_5QNone_Int_4_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t lizzieLet12_6QNode_Int_5QNone_Int_4_bufchan_d;
  logic lizzieLet12_6QNode_Int_5QNone_Int_4_bufchan_r;
  assign lizzieLet12_6QNode_Int_5QNone_Int_4_r = ((! lizzieLet12_6QNode_Int_5QNone_Int_4_bufchan_d[0]) || lizzieLet12_6QNode_Int_5QNone_Int_4_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNode_Int_5QNone_Int_4_bufchan_d <= 1'd0;
    else
      if (lizzieLet12_6QNode_Int_5QNone_Int_4_r)
        lizzieLet12_6QNode_Int_5QNone_Int_4_bufchan_d <= lizzieLet12_6QNode_Int_5QNone_Int_4_d;
  MyDTInt_Bool_t lizzieLet12_6QNode_Int_5QNone_Int_4_bufchan_buf;
  assign lizzieLet12_6QNode_Int_5QNone_Int_4_bufchan_r = (! lizzieLet12_6QNode_Int_5QNone_Int_4_bufchan_buf[0]);
  assign lizzieLet12_6QNode_Int_5QNone_Int_4_argbuf_d = (lizzieLet12_6QNode_Int_5QNone_Int_4_bufchan_buf[0] ? lizzieLet12_6QNode_Int_5QNone_Int_4_bufchan_buf :
                                                         lizzieLet12_6QNode_Int_5QNone_Int_4_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNode_Int_5QNone_Int_4_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet12_6QNode_Int_5QNone_Int_4_argbuf_r && lizzieLet12_6QNode_Int_5QNone_Int_4_bufchan_buf[0]))
        lizzieLet12_6QNode_Int_5QNone_Int_4_bufchan_buf <= 1'd0;
      else if (((! lizzieLet12_6QNode_Int_5QNone_Int_4_argbuf_r) && (! lizzieLet12_6QNode_Int_5QNone_Int_4_bufchan_buf[0])))
        lizzieLet12_6QNode_Int_5QNone_Int_4_bufchan_buf <= lizzieLet12_6QNode_Int_5QNone_Int_4_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty MyDTInt_Int_Int) : (lizzieLet12_6QNode_Int_6,QTree_Int) (lizzieLet12_7QNode_Int,MyDTInt_Int_Int) > [(_45,MyDTInt_Int_Int),
                                                                                                              (_44,MyDTInt_Int_Int),
                                                                                                              (lizzieLet12_6QNode_Int_6QNode_Int,MyDTInt_Int_Int),
                                                                                                              (_43,MyDTInt_Int_Int)] */
  logic [3:0] lizzieLet12_7QNode_Int_onehotd;
  always_comb
    if ((lizzieLet12_6QNode_Int_6_d[0] && lizzieLet12_7QNode_Int_d[0]))
      unique case (lizzieLet12_6QNode_Int_6_d[2:1])
        2'd0: lizzieLet12_7QNode_Int_onehotd = 4'd1;
        2'd1: lizzieLet12_7QNode_Int_onehotd = 4'd2;
        2'd2: lizzieLet12_7QNode_Int_onehotd = 4'd4;
        2'd3: lizzieLet12_7QNode_Int_onehotd = 4'd8;
        default: lizzieLet12_7QNode_Int_onehotd = 4'd0;
      endcase
    else lizzieLet12_7QNode_Int_onehotd = 4'd0;
  assign _45_d = lizzieLet12_7QNode_Int_onehotd[0];
  assign _44_d = lizzieLet12_7QNode_Int_onehotd[1];
  assign lizzieLet12_6QNode_Int_6QNode_Int_d = lizzieLet12_7QNode_Int_onehotd[2];
  assign _43_d = lizzieLet12_7QNode_Int_onehotd[3];
  assign lizzieLet12_7QNode_Int_r = (| (lizzieLet12_7QNode_Int_onehotd & {_43_r,
                                                                          lizzieLet12_6QNode_Int_6QNode_Int_r,
                                                                          _44_r,
                                                                          _45_r}));
  assign lizzieLet12_6QNode_Int_6_r = lizzieLet12_7QNode_Int_r;
  
  /* fork (Ty MyDTInt_Int_Int) : (lizzieLet12_6QNode_Int_6QNode_Int,MyDTInt_Int_Int) > [(lizzieLet12_6QNode_Int_6QNode_Int_1,MyDTInt_Int_Int),
                                                                                   (lizzieLet12_6QNode_Int_6QNode_Int_2,MyDTInt_Int_Int)] */
  logic [1:0] lizzieLet12_6QNode_Int_6QNode_Int_emitted;
  logic [1:0] lizzieLet12_6QNode_Int_6QNode_Int_done;
  assign lizzieLet12_6QNode_Int_6QNode_Int_1_d = (lizzieLet12_6QNode_Int_6QNode_Int_d[0] && (! lizzieLet12_6QNode_Int_6QNode_Int_emitted[0]));
  assign lizzieLet12_6QNode_Int_6QNode_Int_2_d = (lizzieLet12_6QNode_Int_6QNode_Int_d[0] && (! lizzieLet12_6QNode_Int_6QNode_Int_emitted[1]));
  assign lizzieLet12_6QNode_Int_6QNode_Int_done = (lizzieLet12_6QNode_Int_6QNode_Int_emitted | ({lizzieLet12_6QNode_Int_6QNode_Int_2_d[0],
                                                                                                 lizzieLet12_6QNode_Int_6QNode_Int_1_d[0]} & {lizzieLet12_6QNode_Int_6QNode_Int_2_r,
                                                                                                                                              lizzieLet12_6QNode_Int_6QNode_Int_1_r}));
  assign lizzieLet12_6QNode_Int_6QNode_Int_r = (& lizzieLet12_6QNode_Int_6QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNode_Int_6QNode_Int_emitted <= 2'd0;
    else
      lizzieLet12_6QNode_Int_6QNode_Int_emitted <= (lizzieLet12_6QNode_Int_6QNode_Int_r ? 2'd0 :
                                                    lizzieLet12_6QNode_Int_6QNode_Int_done);
  
  /* buf (Ty MyDTInt_Int_Int) : (lizzieLet12_6QNode_Int_6QNode_Int_2,MyDTInt_Int_Int) > (lizzieLet12_6QNode_Int_6QNode_Int_2_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t lizzieLet12_6QNode_Int_6QNode_Int_2_bufchan_d;
  logic lizzieLet12_6QNode_Int_6QNode_Int_2_bufchan_r;
  assign lizzieLet12_6QNode_Int_6QNode_Int_2_r = ((! lizzieLet12_6QNode_Int_6QNode_Int_2_bufchan_d[0]) || lizzieLet12_6QNode_Int_6QNode_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNode_Int_6QNode_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet12_6QNode_Int_6QNode_Int_2_r)
        lizzieLet12_6QNode_Int_6QNode_Int_2_bufchan_d <= lizzieLet12_6QNode_Int_6QNode_Int_2_d;
  MyDTInt_Int_Int_t lizzieLet12_6QNode_Int_6QNode_Int_2_bufchan_buf;
  assign lizzieLet12_6QNode_Int_6QNode_Int_2_bufchan_r = (! lizzieLet12_6QNode_Int_6QNode_Int_2_bufchan_buf[0]);
  assign lizzieLet12_6QNode_Int_6QNode_Int_2_argbuf_d = (lizzieLet12_6QNode_Int_6QNode_Int_2_bufchan_buf[0] ? lizzieLet12_6QNode_Int_6QNode_Int_2_bufchan_buf :
                                                         lizzieLet12_6QNode_Int_6QNode_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNode_Int_6QNode_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet12_6QNode_Int_6QNode_Int_2_argbuf_r && lizzieLet12_6QNode_Int_6QNode_Int_2_bufchan_buf[0]))
        lizzieLet12_6QNode_Int_6QNode_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet12_6QNode_Int_6QNode_Int_2_argbuf_r) && (! lizzieLet12_6QNode_Int_6QNode_Int_2_bufchan_buf[0])))
        lizzieLet12_6QNode_Int_6QNode_Int_2_bufchan_buf <= lizzieLet12_6QNode_Int_6QNode_Int_2_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty MyDTInt_Int) : (lizzieLet12_6QNode_Int_7,QTree_Int) (lizzieLet12_8QNode_Int,MyDTInt_Int) > [(lizzieLet12_6QNode_Int_7QNone_Int,MyDTInt_Int),
                                                                                                      (_42,MyDTInt_Int),
                                                                                                      (lizzieLet12_6QNode_Int_7QNode_Int,MyDTInt_Int),
                                                                                                      (_41,MyDTInt_Int)] */
  logic [3:0] lizzieLet12_8QNode_Int_onehotd;
  always_comb
    if ((lizzieLet12_6QNode_Int_7_d[0] && lizzieLet12_8QNode_Int_d[0]))
      unique case (lizzieLet12_6QNode_Int_7_d[2:1])
        2'd0: lizzieLet12_8QNode_Int_onehotd = 4'd1;
        2'd1: lizzieLet12_8QNode_Int_onehotd = 4'd2;
        2'd2: lizzieLet12_8QNode_Int_onehotd = 4'd4;
        2'd3: lizzieLet12_8QNode_Int_onehotd = 4'd8;
        default: lizzieLet12_8QNode_Int_onehotd = 4'd0;
      endcase
    else lizzieLet12_8QNode_Int_onehotd = 4'd0;
  assign lizzieLet12_6QNode_Int_7QNone_Int_d = lizzieLet12_8QNode_Int_onehotd[0];
  assign _42_d = lizzieLet12_8QNode_Int_onehotd[1];
  assign lizzieLet12_6QNode_Int_7QNode_Int_d = lizzieLet12_8QNode_Int_onehotd[2];
  assign _41_d = lizzieLet12_8QNode_Int_onehotd[3];
  assign lizzieLet12_8QNode_Int_r = (| (lizzieLet12_8QNode_Int_onehotd & {_41_r,
                                                                          lizzieLet12_6QNode_Int_7QNode_Int_r,
                                                                          _42_r,
                                                                          lizzieLet12_6QNode_Int_7QNone_Int_r}));
  assign lizzieLet12_6QNode_Int_7_r = lizzieLet12_8QNode_Int_r;
  
  /* fork (Ty MyDTInt_Int) : (lizzieLet12_6QNode_Int_7QNode_Int,MyDTInt_Int) > [(lizzieLet12_6QNode_Int_7QNode_Int_1,MyDTInt_Int),
                                                                           (lizzieLet12_6QNode_Int_7QNode_Int_2,MyDTInt_Int)] */
  logic [1:0] lizzieLet12_6QNode_Int_7QNode_Int_emitted;
  logic [1:0] lizzieLet12_6QNode_Int_7QNode_Int_done;
  assign lizzieLet12_6QNode_Int_7QNode_Int_1_d = (lizzieLet12_6QNode_Int_7QNode_Int_d[0] && (! lizzieLet12_6QNode_Int_7QNode_Int_emitted[0]));
  assign lizzieLet12_6QNode_Int_7QNode_Int_2_d = (lizzieLet12_6QNode_Int_7QNode_Int_d[0] && (! lizzieLet12_6QNode_Int_7QNode_Int_emitted[1]));
  assign lizzieLet12_6QNode_Int_7QNode_Int_done = (lizzieLet12_6QNode_Int_7QNode_Int_emitted | ({lizzieLet12_6QNode_Int_7QNode_Int_2_d[0],
                                                                                                 lizzieLet12_6QNode_Int_7QNode_Int_1_d[0]} & {lizzieLet12_6QNode_Int_7QNode_Int_2_r,
                                                                                                                                              lizzieLet12_6QNode_Int_7QNode_Int_1_r}));
  assign lizzieLet12_6QNode_Int_7QNode_Int_r = (& lizzieLet12_6QNode_Int_7QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNode_Int_7QNode_Int_emitted <= 2'd0;
    else
      lizzieLet12_6QNode_Int_7QNode_Int_emitted <= (lizzieLet12_6QNode_Int_7QNode_Int_r ? 2'd0 :
                                                    lizzieLet12_6QNode_Int_7QNode_Int_done);
  
  /* buf (Ty MyDTInt_Int) : (lizzieLet12_6QNode_Int_7QNode_Int_2,MyDTInt_Int) > (lizzieLet12_6QNode_Int_7QNode_Int_2_argbuf,MyDTInt_Int) */
  MyDTInt_Int_t lizzieLet12_6QNode_Int_7QNode_Int_2_bufchan_d;
  logic lizzieLet12_6QNode_Int_7QNode_Int_2_bufchan_r;
  assign lizzieLet12_6QNode_Int_7QNode_Int_2_r = ((! lizzieLet12_6QNode_Int_7QNode_Int_2_bufchan_d[0]) || lizzieLet12_6QNode_Int_7QNode_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNode_Int_7QNode_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet12_6QNode_Int_7QNode_Int_2_r)
        lizzieLet12_6QNode_Int_7QNode_Int_2_bufchan_d <= lizzieLet12_6QNode_Int_7QNode_Int_2_d;
  MyDTInt_Int_t lizzieLet12_6QNode_Int_7QNode_Int_2_bufchan_buf;
  assign lizzieLet12_6QNode_Int_7QNode_Int_2_bufchan_r = (! lizzieLet12_6QNode_Int_7QNode_Int_2_bufchan_buf[0]);
  assign lizzieLet12_6QNode_Int_7QNode_Int_2_argbuf_d = (lizzieLet12_6QNode_Int_7QNode_Int_2_bufchan_buf[0] ? lizzieLet12_6QNode_Int_7QNode_Int_2_bufchan_buf :
                                                         lizzieLet12_6QNode_Int_7QNode_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNode_Int_7QNode_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet12_6QNode_Int_7QNode_Int_2_argbuf_r && lizzieLet12_6QNode_Int_7QNode_Int_2_bufchan_buf[0]))
        lizzieLet12_6QNode_Int_7QNode_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet12_6QNode_Int_7QNode_Int_2_argbuf_r) && (! lizzieLet12_6QNode_Int_7QNode_Int_2_bufchan_buf[0])))
        lizzieLet12_6QNode_Int_7QNode_Int_2_bufchan_buf <= lizzieLet12_6QNode_Int_7QNode_Int_2_bufchan_d;
  
  /* fork (Ty MyDTInt_Int) : (lizzieLet12_6QNode_Int_7QNone_Int,MyDTInt_Int) > [(lizzieLet12_6QNode_Int_7QNone_Int_1,MyDTInt_Int),
                                                                           (lizzieLet12_6QNode_Int_7QNone_Int_2,MyDTInt_Int),
                                                                           (lizzieLet12_6QNode_Int_7QNone_Int_3,MyDTInt_Int),
                                                                           (lizzieLet12_6QNode_Int_7QNone_Int_4,MyDTInt_Int)] */
  logic [3:0] lizzieLet12_6QNode_Int_7QNone_Int_emitted;
  logic [3:0] lizzieLet12_6QNode_Int_7QNone_Int_done;
  assign lizzieLet12_6QNode_Int_7QNone_Int_1_d = (lizzieLet12_6QNode_Int_7QNone_Int_d[0] && (! lizzieLet12_6QNode_Int_7QNone_Int_emitted[0]));
  assign lizzieLet12_6QNode_Int_7QNone_Int_2_d = (lizzieLet12_6QNode_Int_7QNone_Int_d[0] && (! lizzieLet12_6QNode_Int_7QNone_Int_emitted[1]));
  assign lizzieLet12_6QNode_Int_7QNone_Int_3_d = (lizzieLet12_6QNode_Int_7QNone_Int_d[0] && (! lizzieLet12_6QNode_Int_7QNone_Int_emitted[2]));
  assign lizzieLet12_6QNode_Int_7QNone_Int_4_d = (lizzieLet12_6QNode_Int_7QNone_Int_d[0] && (! lizzieLet12_6QNode_Int_7QNone_Int_emitted[3]));
  assign lizzieLet12_6QNode_Int_7QNone_Int_done = (lizzieLet12_6QNode_Int_7QNone_Int_emitted | ({lizzieLet12_6QNode_Int_7QNone_Int_4_d[0],
                                                                                                 lizzieLet12_6QNode_Int_7QNone_Int_3_d[0],
                                                                                                 lizzieLet12_6QNode_Int_7QNone_Int_2_d[0],
                                                                                                 lizzieLet12_6QNode_Int_7QNone_Int_1_d[0]} & {lizzieLet12_6QNode_Int_7QNone_Int_4_r,
                                                                                                                                              lizzieLet12_6QNode_Int_7QNone_Int_3_r,
                                                                                                                                              lizzieLet12_6QNode_Int_7QNone_Int_2_r,
                                                                                                                                              lizzieLet12_6QNode_Int_7QNone_Int_1_r}));
  assign lizzieLet12_6QNode_Int_7QNone_Int_r = (& lizzieLet12_6QNode_Int_7QNone_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNode_Int_7QNone_Int_emitted <= 4'd0;
    else
      lizzieLet12_6QNode_Int_7QNone_Int_emitted <= (lizzieLet12_6QNode_Int_7QNone_Int_r ? 4'd0 :
                                                    lizzieLet12_6QNode_Int_7QNone_Int_done);
  
  /* buf (Ty MyDTInt_Int) : (lizzieLet12_6QNode_Int_7QNone_Int_1,MyDTInt_Int) > (lizzieLet12_6QNode_Int_7QNone_Int_1_argbuf,MyDTInt_Int) */
  MyDTInt_Int_t lizzieLet12_6QNode_Int_7QNone_Int_1_bufchan_d;
  logic lizzieLet12_6QNode_Int_7QNone_Int_1_bufchan_r;
  assign lizzieLet12_6QNode_Int_7QNone_Int_1_r = ((! lizzieLet12_6QNode_Int_7QNone_Int_1_bufchan_d[0]) || lizzieLet12_6QNode_Int_7QNone_Int_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNode_Int_7QNone_Int_1_bufchan_d <= 1'd0;
    else
      if (lizzieLet12_6QNode_Int_7QNone_Int_1_r)
        lizzieLet12_6QNode_Int_7QNone_Int_1_bufchan_d <= lizzieLet12_6QNode_Int_7QNone_Int_1_d;
  MyDTInt_Int_t lizzieLet12_6QNode_Int_7QNone_Int_1_bufchan_buf;
  assign lizzieLet12_6QNode_Int_7QNone_Int_1_bufchan_r = (! lizzieLet12_6QNode_Int_7QNone_Int_1_bufchan_buf[0]);
  assign lizzieLet12_6QNode_Int_7QNone_Int_1_argbuf_d = (lizzieLet12_6QNode_Int_7QNone_Int_1_bufchan_buf[0] ? lizzieLet12_6QNode_Int_7QNone_Int_1_bufchan_buf :
                                                         lizzieLet12_6QNode_Int_7QNone_Int_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNode_Int_7QNone_Int_1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet12_6QNode_Int_7QNone_Int_1_argbuf_r && lizzieLet12_6QNode_Int_7QNone_Int_1_bufchan_buf[0]))
        lizzieLet12_6QNode_Int_7QNone_Int_1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet12_6QNode_Int_7QNone_Int_1_argbuf_r) && (! lizzieLet12_6QNode_Int_7QNone_Int_1_bufchan_buf[0])))
        lizzieLet12_6QNode_Int_7QNone_Int_1_bufchan_buf <= lizzieLet12_6QNode_Int_7QNone_Int_1_bufchan_d;
  
  /* buf (Ty MyDTInt_Int) : (lizzieLet12_6QNode_Int_7QNone_Int_2,MyDTInt_Int) > (lizzieLet12_6QNode_Int_7QNone_Int_2_argbuf,MyDTInt_Int) */
  MyDTInt_Int_t lizzieLet12_6QNode_Int_7QNone_Int_2_bufchan_d;
  logic lizzieLet12_6QNode_Int_7QNone_Int_2_bufchan_r;
  assign lizzieLet12_6QNode_Int_7QNone_Int_2_r = ((! lizzieLet12_6QNode_Int_7QNone_Int_2_bufchan_d[0]) || lizzieLet12_6QNode_Int_7QNone_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNode_Int_7QNone_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet12_6QNode_Int_7QNone_Int_2_r)
        lizzieLet12_6QNode_Int_7QNone_Int_2_bufchan_d <= lizzieLet12_6QNode_Int_7QNone_Int_2_d;
  MyDTInt_Int_t lizzieLet12_6QNode_Int_7QNone_Int_2_bufchan_buf;
  assign lizzieLet12_6QNode_Int_7QNone_Int_2_bufchan_r = (! lizzieLet12_6QNode_Int_7QNone_Int_2_bufchan_buf[0]);
  assign lizzieLet12_6QNode_Int_7QNone_Int_2_argbuf_d = (lizzieLet12_6QNode_Int_7QNone_Int_2_bufchan_buf[0] ? lizzieLet12_6QNode_Int_7QNone_Int_2_bufchan_buf :
                                                         lizzieLet12_6QNode_Int_7QNone_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNode_Int_7QNone_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet12_6QNode_Int_7QNone_Int_2_argbuf_r && lizzieLet12_6QNode_Int_7QNone_Int_2_bufchan_buf[0]))
        lizzieLet12_6QNode_Int_7QNone_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet12_6QNode_Int_7QNone_Int_2_argbuf_r) && (! lizzieLet12_6QNode_Int_7QNone_Int_2_bufchan_buf[0])))
        lizzieLet12_6QNode_Int_7QNone_Int_2_bufchan_buf <= lizzieLet12_6QNode_Int_7QNone_Int_2_bufchan_d;
  
  /* buf (Ty MyDTInt_Int) : (lizzieLet12_6QNode_Int_7QNone_Int_3,MyDTInt_Int) > (lizzieLet12_6QNode_Int_7QNone_Int_3_argbuf,MyDTInt_Int) */
  MyDTInt_Int_t lizzieLet12_6QNode_Int_7QNone_Int_3_bufchan_d;
  logic lizzieLet12_6QNode_Int_7QNone_Int_3_bufchan_r;
  assign lizzieLet12_6QNode_Int_7QNone_Int_3_r = ((! lizzieLet12_6QNode_Int_7QNone_Int_3_bufchan_d[0]) || lizzieLet12_6QNode_Int_7QNone_Int_3_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNode_Int_7QNone_Int_3_bufchan_d <= 1'd0;
    else
      if (lizzieLet12_6QNode_Int_7QNone_Int_3_r)
        lizzieLet12_6QNode_Int_7QNone_Int_3_bufchan_d <= lizzieLet12_6QNode_Int_7QNone_Int_3_d;
  MyDTInt_Int_t lizzieLet12_6QNode_Int_7QNone_Int_3_bufchan_buf;
  assign lizzieLet12_6QNode_Int_7QNone_Int_3_bufchan_r = (! lizzieLet12_6QNode_Int_7QNone_Int_3_bufchan_buf[0]);
  assign lizzieLet12_6QNode_Int_7QNone_Int_3_argbuf_d = (lizzieLet12_6QNode_Int_7QNone_Int_3_bufchan_buf[0] ? lizzieLet12_6QNode_Int_7QNone_Int_3_bufchan_buf :
                                                         lizzieLet12_6QNode_Int_7QNone_Int_3_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNode_Int_7QNone_Int_3_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet12_6QNode_Int_7QNone_Int_3_argbuf_r && lizzieLet12_6QNode_Int_7QNone_Int_3_bufchan_buf[0]))
        lizzieLet12_6QNode_Int_7QNone_Int_3_bufchan_buf <= 1'd0;
      else if (((! lizzieLet12_6QNode_Int_7QNone_Int_3_argbuf_r) && (! lizzieLet12_6QNode_Int_7QNone_Int_3_bufchan_buf[0])))
        lizzieLet12_6QNode_Int_7QNone_Int_3_bufchan_buf <= lizzieLet12_6QNode_Int_7QNone_Int_3_bufchan_d;
  
  /* buf (Ty MyDTInt_Int) : (lizzieLet12_6QNode_Int_7QNone_Int_4,MyDTInt_Int) > (lizzieLet12_6QNode_Int_7QNone_Int_4_argbuf,MyDTInt_Int) */
  MyDTInt_Int_t lizzieLet12_6QNode_Int_7QNone_Int_4_bufchan_d;
  logic lizzieLet12_6QNode_Int_7QNone_Int_4_bufchan_r;
  assign lizzieLet12_6QNode_Int_7QNone_Int_4_r = ((! lizzieLet12_6QNode_Int_7QNone_Int_4_bufchan_d[0]) || lizzieLet12_6QNode_Int_7QNone_Int_4_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNode_Int_7QNone_Int_4_bufchan_d <= 1'd0;
    else
      if (lizzieLet12_6QNode_Int_7QNone_Int_4_r)
        lizzieLet12_6QNode_Int_7QNone_Int_4_bufchan_d <= lizzieLet12_6QNode_Int_7QNone_Int_4_d;
  MyDTInt_Int_t lizzieLet12_6QNode_Int_7QNone_Int_4_bufchan_buf;
  assign lizzieLet12_6QNode_Int_7QNone_Int_4_bufchan_r = (! lizzieLet12_6QNode_Int_7QNone_Int_4_bufchan_buf[0]);
  assign lizzieLet12_6QNode_Int_7QNone_Int_4_argbuf_d = (lizzieLet12_6QNode_Int_7QNone_Int_4_bufchan_buf[0] ? lizzieLet12_6QNode_Int_7QNone_Int_4_bufchan_buf :
                                                         lizzieLet12_6QNode_Int_7QNone_Int_4_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNode_Int_7QNone_Int_4_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet12_6QNode_Int_7QNone_Int_4_argbuf_r && lizzieLet12_6QNode_Int_7QNone_Int_4_bufchan_buf[0]))
        lizzieLet12_6QNode_Int_7QNone_Int_4_bufchan_buf <= 1'd0;
      else if (((! lizzieLet12_6QNode_Int_7QNone_Int_4_argbuf_r) && (! lizzieLet12_6QNode_Int_7QNone_Int_4_bufchan_buf[0])))
        lizzieLet12_6QNode_Int_7QNone_Int_4_bufchan_buf <= lizzieLet12_6QNode_Int_7QNone_Int_4_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_CTf_f_Int_Int) : (lizzieLet12_6QNode_Int_8,QTree_Int) (lizzieLet12_9QNode_Int,Pointer_CTf_f_Int_Int) > [(lizzieLet12_6QNode_Int_8QNone_Int,Pointer_CTf_f_Int_Int),
                                                                                                                          (lizzieLet12_6QNode_Int_8QVal_Int,Pointer_CTf_f_Int_Int),
                                                                                                                          (lizzieLet12_6QNode_Int_8QNode_Int,Pointer_CTf_f_Int_Int),
                                                                                                                          (lizzieLet12_6QNode_Int_8QError_Int,Pointer_CTf_f_Int_Int)] */
  logic [3:0] lizzieLet12_9QNode_Int_onehotd;
  always_comb
    if ((lizzieLet12_6QNode_Int_8_d[0] && lizzieLet12_9QNode_Int_d[0]))
      unique case (lizzieLet12_6QNode_Int_8_d[2:1])
        2'd0: lizzieLet12_9QNode_Int_onehotd = 4'd1;
        2'd1: lizzieLet12_9QNode_Int_onehotd = 4'd2;
        2'd2: lizzieLet12_9QNode_Int_onehotd = 4'd4;
        2'd3: lizzieLet12_9QNode_Int_onehotd = 4'd8;
        default: lizzieLet12_9QNode_Int_onehotd = 4'd0;
      endcase
    else lizzieLet12_9QNode_Int_onehotd = 4'd0;
  assign lizzieLet12_6QNode_Int_8QNone_Int_d = {lizzieLet12_9QNode_Int_d[16:1],
                                                lizzieLet12_9QNode_Int_onehotd[0]};
  assign lizzieLet12_6QNode_Int_8QVal_Int_d = {lizzieLet12_9QNode_Int_d[16:1],
                                               lizzieLet12_9QNode_Int_onehotd[1]};
  assign lizzieLet12_6QNode_Int_8QNode_Int_d = {lizzieLet12_9QNode_Int_d[16:1],
                                                lizzieLet12_9QNode_Int_onehotd[2]};
  assign lizzieLet12_6QNode_Int_8QError_Int_d = {lizzieLet12_9QNode_Int_d[16:1],
                                                 lizzieLet12_9QNode_Int_onehotd[3]};
  assign lizzieLet12_9QNode_Int_r = (| (lizzieLet12_9QNode_Int_onehotd & {lizzieLet12_6QNode_Int_8QError_Int_r,
                                                                          lizzieLet12_6QNode_Int_8QNode_Int_r,
                                                                          lizzieLet12_6QNode_Int_8QVal_Int_r,
                                                                          lizzieLet12_6QNode_Int_8QNone_Int_r}));
  assign lizzieLet12_6QNode_Int_8_r = lizzieLet12_9QNode_Int_r;
  
  /* buf (Ty Pointer_CTf_f_Int_Int) : (lizzieLet12_6QNode_Int_8QError_Int,Pointer_CTf_f_Int_Int) > (lizzieLet12_6QNode_Int_8QError_Int_1_argbuf,Pointer_CTf_f_Int_Int) */
  Pointer_CTf_f_Int_Int_t lizzieLet12_6QNode_Int_8QError_Int_bufchan_d;
  logic lizzieLet12_6QNode_Int_8QError_Int_bufchan_r;
  assign lizzieLet12_6QNode_Int_8QError_Int_r = ((! lizzieLet12_6QNode_Int_8QError_Int_bufchan_d[0]) || lizzieLet12_6QNode_Int_8QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNode_Int_8QError_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet12_6QNode_Int_8QError_Int_r)
        lizzieLet12_6QNode_Int_8QError_Int_bufchan_d <= lizzieLet12_6QNode_Int_8QError_Int_d;
  Pointer_CTf_f_Int_Int_t lizzieLet12_6QNode_Int_8QError_Int_bufchan_buf;
  assign lizzieLet12_6QNode_Int_8QError_Int_bufchan_r = (! lizzieLet12_6QNode_Int_8QError_Int_bufchan_buf[0]);
  assign lizzieLet12_6QNode_Int_8QError_Int_1_argbuf_d = (lizzieLet12_6QNode_Int_8QError_Int_bufchan_buf[0] ? lizzieLet12_6QNode_Int_8QError_Int_bufchan_buf :
                                                          lizzieLet12_6QNode_Int_8QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNode_Int_8QError_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet12_6QNode_Int_8QError_Int_1_argbuf_r && lizzieLet12_6QNode_Int_8QError_Int_bufchan_buf[0]))
        lizzieLet12_6QNode_Int_8QError_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet12_6QNode_Int_8QError_Int_1_argbuf_r) && (! lizzieLet12_6QNode_Int_8QError_Int_bufchan_buf[0])))
        lizzieLet12_6QNode_Int_8QError_Int_bufchan_buf <= lizzieLet12_6QNode_Int_8QError_Int_bufchan_d;
  
  /* dcon (Ty CTf_f_Int_Int,
      Dcon Lcall_f_f_Int_Int3) : [(lizzieLet12_6QNode_Int_8QNode_Int,Pointer_CTf_f_Int_Int),
                                  (lizzieLet12_6QNode_Int_9QNode_Int,Pointer_QTree_Int),
                                  (t1a8Y_destruct,Pointer_QTree_Int),
                                  (lizzieLet12_6QNode_Int_5QNode_Int_1,MyDTInt_Bool),
                                  (lizzieLet12_6QNode_Int_7QNode_Int_1,MyDTInt_Int),
                                  (lizzieLet12_6QNode_Int_4QNode_Int_1,MyDTInt_Bool),
                                  (lizzieLet12_6QNode_Int_6QNode_Int_1,MyDTInt_Int_Int),
                                  (lizzieLet12_6QNode_Int_10QNode_Int,Pointer_QTree_Int),
                                  (t2a8Z_destruct,Pointer_QTree_Int),
                                  (lizzieLet12_6QNode_Int_11QNode_Int,Pointer_QTree_Int),
                                  (t3a90_destruct,Pointer_QTree_Int)] > (lizzieLet12_6QNode_Int_8QNode_Int_1lizzieLet12_6QNode_Int_9QNode_Int_1t1a8Y_1lizzieLet12_6QNode_Int_5QNode_Int_1lizzieLet12_6QNode_Int_7QNode_Int_1lizzieLet12_6QNode_Int_4QNode_Int_1lizzieLet12_6QNode_Int_6QNode_Int_1lizzieLet12_6QNode_Int_10QNode_Int_1t2a8Z_1lizzieLet12_6QNode_Int_11QNode_Int_1t3a90_1Lcall_f_f_Int_Int3,CTf_f_Int_Int) */
  assign lizzieLet12_6QNode_Int_8QNode_Int_1lizzieLet12_6QNode_Int_9QNode_Int_1t1a8Y_1lizzieLet12_6QNode_Int_5QNode_Int_1lizzieLet12_6QNode_Int_7QNode_Int_1lizzieLet12_6QNode_Int_4QNode_Int_1lizzieLet12_6QNode_Int_6QNode_Int_1lizzieLet12_6QNode_Int_10QNode_Int_1t2a8Z_1lizzieLet12_6QNode_Int_11QNode_Int_1t3a90_1Lcall_f_f_Int_Int3_d = Lcall_f_f_Int_Int3_dc((& {lizzieLet12_6QNode_Int_8QNode_Int_d[0],
                                                                                                                                                                                                                                                                                                                                                                         lizzieLet12_6QNode_Int_9QNode_Int_d[0],
                                                                                                                                                                                                                                                                                                                                                                         t1a8Y_destruct_d[0],
                                                                                                                                                                                                                                                                                                                                                                         lizzieLet12_6QNode_Int_5QNode_Int_1_d[0],
                                                                                                                                                                                                                                                                                                                                                                         lizzieLet12_6QNode_Int_7QNode_Int_1_d[0],
                                                                                                                                                                                                                                                                                                                                                                         lizzieLet12_6QNode_Int_4QNode_Int_1_d[0],
                                                                                                                                                                                                                                                                                                                                                                         lizzieLet12_6QNode_Int_6QNode_Int_1_d[0],
                                                                                                                                                                                                                                                                                                                                                                         lizzieLet12_6QNode_Int_10QNode_Int_d[0],
                                                                                                                                                                                                                                                                                                                                                                         t2a8Z_destruct_d[0],
                                                                                                                                                                                                                                                                                                                                                                         lizzieLet12_6QNode_Int_11QNode_Int_d[0],
                                                                                                                                                                                                                                                                                                                                                                         t3a90_destruct_d[0]}), lizzieLet12_6QNode_Int_8QNode_Int_d, lizzieLet12_6QNode_Int_9QNode_Int_d, t1a8Y_destruct_d, lizzieLet12_6QNode_Int_5QNode_Int_1_d, lizzieLet12_6QNode_Int_7QNode_Int_1_d, lizzieLet12_6QNode_Int_4QNode_Int_1_d, lizzieLet12_6QNode_Int_6QNode_Int_1_d, lizzieLet12_6QNode_Int_10QNode_Int_d, t2a8Z_destruct_d, lizzieLet12_6QNode_Int_11QNode_Int_d, t3a90_destruct_d);
  assign {lizzieLet12_6QNode_Int_8QNode_Int_r,
          lizzieLet12_6QNode_Int_9QNode_Int_r,
          t1a8Y_destruct_r,
          lizzieLet12_6QNode_Int_5QNode_Int_1_r,
          lizzieLet12_6QNode_Int_7QNode_Int_1_r,
          lizzieLet12_6QNode_Int_4QNode_Int_1_r,
          lizzieLet12_6QNode_Int_6QNode_Int_1_r,
          lizzieLet12_6QNode_Int_10QNode_Int_r,
          t2a8Z_destruct_r,
          lizzieLet12_6QNode_Int_11QNode_Int_r,
          t3a90_destruct_r} = {11 {(lizzieLet12_6QNode_Int_8QNode_Int_1lizzieLet12_6QNode_Int_9QNode_Int_1t1a8Y_1lizzieLet12_6QNode_Int_5QNode_Int_1lizzieLet12_6QNode_Int_7QNode_Int_1lizzieLet12_6QNode_Int_4QNode_Int_1lizzieLet12_6QNode_Int_6QNode_Int_1lizzieLet12_6QNode_Int_10QNode_Int_1t2a8Z_1lizzieLet12_6QNode_Int_11QNode_Int_1t3a90_1Lcall_f_f_Int_Int3_r && lizzieLet12_6QNode_Int_8QNode_Int_1lizzieLet12_6QNode_Int_9QNode_Int_1t1a8Y_1lizzieLet12_6QNode_Int_5QNode_Int_1lizzieLet12_6QNode_Int_7QNode_Int_1lizzieLet12_6QNode_Int_4QNode_Int_1lizzieLet12_6QNode_Int_6QNode_Int_1lizzieLet12_6QNode_Int_10QNode_Int_1t2a8Z_1lizzieLet12_6QNode_Int_11QNode_Int_1t3a90_1Lcall_f_f_Int_Int3_d[0])}};
  
  /* buf (Ty CTf_f_Int_Int) : (lizzieLet12_6QNode_Int_8QNode_Int_1lizzieLet12_6QNode_Int_9QNode_Int_1t1a8Y_1lizzieLet12_6QNode_Int_5QNode_Int_1lizzieLet12_6QNode_Int_7QNode_Int_1lizzieLet12_6QNode_Int_4QNode_Int_1lizzieLet12_6QNode_Int_6QNode_Int_1lizzieLet12_6QNode_Int_10QNode_Int_1t2a8Z_1lizzieLet12_6QNode_Int_11QNode_Int_1t3a90_1Lcall_f_f_Int_Int3,CTf_f_Int_Int) > (lizzieLet30_1_argbuf,CTf_f_Int_Int) */
  CTf_f_Int_Int_t lizzieLet12_6QNode_Int_8QNode_Int_1lizzieLet12_6QNode_Int_9QNode_Int_1t1a8Y_1lizzieLet12_6QNode_Int_5QNode_Int_1lizzieLet12_6QNode_Int_7QNode_Int_1lizzieLet12_6QNode_Int_4QNode_Int_1lizzieLet12_6QNode_Int_6QNode_Int_1lizzieLet12_6QNode_Int_10QNode_Int_1t2a8Z_1lizzieLet12_6QNode_Int_11QNode_Int_1t3a90_1Lcall_f_f_Int_Int3_bufchan_d;
  logic lizzieLet12_6QNode_Int_8QNode_Int_1lizzieLet12_6QNode_Int_9QNode_Int_1t1a8Y_1lizzieLet12_6QNode_Int_5QNode_Int_1lizzieLet12_6QNode_Int_7QNode_Int_1lizzieLet12_6QNode_Int_4QNode_Int_1lizzieLet12_6QNode_Int_6QNode_Int_1lizzieLet12_6QNode_Int_10QNode_Int_1t2a8Z_1lizzieLet12_6QNode_Int_11QNode_Int_1t3a90_1Lcall_f_f_Int_Int3_bufchan_r;
  assign lizzieLet12_6QNode_Int_8QNode_Int_1lizzieLet12_6QNode_Int_9QNode_Int_1t1a8Y_1lizzieLet12_6QNode_Int_5QNode_Int_1lizzieLet12_6QNode_Int_7QNode_Int_1lizzieLet12_6QNode_Int_4QNode_Int_1lizzieLet12_6QNode_Int_6QNode_Int_1lizzieLet12_6QNode_Int_10QNode_Int_1t2a8Z_1lizzieLet12_6QNode_Int_11QNode_Int_1t3a90_1Lcall_f_f_Int_Int3_r = ((! lizzieLet12_6QNode_Int_8QNode_Int_1lizzieLet12_6QNode_Int_9QNode_Int_1t1a8Y_1lizzieLet12_6QNode_Int_5QNode_Int_1lizzieLet12_6QNode_Int_7QNode_Int_1lizzieLet12_6QNode_Int_4QNode_Int_1lizzieLet12_6QNode_Int_6QNode_Int_1lizzieLet12_6QNode_Int_10QNode_Int_1t2a8Z_1lizzieLet12_6QNode_Int_11QNode_Int_1t3a90_1Lcall_f_f_Int_Int3_bufchan_d[0]) || lizzieLet12_6QNode_Int_8QNode_Int_1lizzieLet12_6QNode_Int_9QNode_Int_1t1a8Y_1lizzieLet12_6QNode_Int_5QNode_Int_1lizzieLet12_6QNode_Int_7QNode_Int_1lizzieLet12_6QNode_Int_4QNode_Int_1lizzieLet12_6QNode_Int_6QNode_Int_1lizzieLet12_6QNode_Int_10QNode_Int_1t2a8Z_1lizzieLet12_6QNode_Int_11QNode_Int_1t3a90_1Lcall_f_f_Int_Int3_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNode_Int_8QNode_Int_1lizzieLet12_6QNode_Int_9QNode_Int_1t1a8Y_1lizzieLet12_6QNode_Int_5QNode_Int_1lizzieLet12_6QNode_Int_7QNode_Int_1lizzieLet12_6QNode_Int_4QNode_Int_1lizzieLet12_6QNode_Int_6QNode_Int_1lizzieLet12_6QNode_Int_10QNode_Int_1t2a8Z_1lizzieLet12_6QNode_Int_11QNode_Int_1t3a90_1Lcall_f_f_Int_Int3_bufchan_d <= {115'd0,
                                                                                                                                                                                                                                                                                                                                                      1'd0};
    else
      if (lizzieLet12_6QNode_Int_8QNode_Int_1lizzieLet12_6QNode_Int_9QNode_Int_1t1a8Y_1lizzieLet12_6QNode_Int_5QNode_Int_1lizzieLet12_6QNode_Int_7QNode_Int_1lizzieLet12_6QNode_Int_4QNode_Int_1lizzieLet12_6QNode_Int_6QNode_Int_1lizzieLet12_6QNode_Int_10QNode_Int_1t2a8Z_1lizzieLet12_6QNode_Int_11QNode_Int_1t3a90_1Lcall_f_f_Int_Int3_r)
        lizzieLet12_6QNode_Int_8QNode_Int_1lizzieLet12_6QNode_Int_9QNode_Int_1t1a8Y_1lizzieLet12_6QNode_Int_5QNode_Int_1lizzieLet12_6QNode_Int_7QNode_Int_1lizzieLet12_6QNode_Int_4QNode_Int_1lizzieLet12_6QNode_Int_6QNode_Int_1lizzieLet12_6QNode_Int_10QNode_Int_1t2a8Z_1lizzieLet12_6QNode_Int_11QNode_Int_1t3a90_1Lcall_f_f_Int_Int3_bufchan_d <= lizzieLet12_6QNode_Int_8QNode_Int_1lizzieLet12_6QNode_Int_9QNode_Int_1t1a8Y_1lizzieLet12_6QNode_Int_5QNode_Int_1lizzieLet12_6QNode_Int_7QNode_Int_1lizzieLet12_6QNode_Int_4QNode_Int_1lizzieLet12_6QNode_Int_6QNode_Int_1lizzieLet12_6QNode_Int_10QNode_Int_1t2a8Z_1lizzieLet12_6QNode_Int_11QNode_Int_1t3a90_1Lcall_f_f_Int_Int3_d;
  CTf_f_Int_Int_t lizzieLet12_6QNode_Int_8QNode_Int_1lizzieLet12_6QNode_Int_9QNode_Int_1t1a8Y_1lizzieLet12_6QNode_Int_5QNode_Int_1lizzieLet12_6QNode_Int_7QNode_Int_1lizzieLet12_6QNode_Int_4QNode_Int_1lizzieLet12_6QNode_Int_6QNode_Int_1lizzieLet12_6QNode_Int_10QNode_Int_1t2a8Z_1lizzieLet12_6QNode_Int_11QNode_Int_1t3a90_1Lcall_f_f_Int_Int3_bufchan_buf;
  assign lizzieLet12_6QNode_Int_8QNode_Int_1lizzieLet12_6QNode_Int_9QNode_Int_1t1a8Y_1lizzieLet12_6QNode_Int_5QNode_Int_1lizzieLet12_6QNode_Int_7QNode_Int_1lizzieLet12_6QNode_Int_4QNode_Int_1lizzieLet12_6QNode_Int_6QNode_Int_1lizzieLet12_6QNode_Int_10QNode_Int_1t2a8Z_1lizzieLet12_6QNode_Int_11QNode_Int_1t3a90_1Lcall_f_f_Int_Int3_bufchan_r = (! lizzieLet12_6QNode_Int_8QNode_Int_1lizzieLet12_6QNode_Int_9QNode_Int_1t1a8Y_1lizzieLet12_6QNode_Int_5QNode_Int_1lizzieLet12_6QNode_Int_7QNode_Int_1lizzieLet12_6QNode_Int_4QNode_Int_1lizzieLet12_6QNode_Int_6QNode_Int_1lizzieLet12_6QNode_Int_10QNode_Int_1t2a8Z_1lizzieLet12_6QNode_Int_11QNode_Int_1t3a90_1Lcall_f_f_Int_Int3_bufchan_buf[0]);
  assign lizzieLet30_1_argbuf_d = (lizzieLet12_6QNode_Int_8QNode_Int_1lizzieLet12_6QNode_Int_9QNode_Int_1t1a8Y_1lizzieLet12_6QNode_Int_5QNode_Int_1lizzieLet12_6QNode_Int_7QNode_Int_1lizzieLet12_6QNode_Int_4QNode_Int_1lizzieLet12_6QNode_Int_6QNode_Int_1lizzieLet12_6QNode_Int_10QNode_Int_1t2a8Z_1lizzieLet12_6QNode_Int_11QNode_Int_1t3a90_1Lcall_f_f_Int_Int3_bufchan_buf[0] ? lizzieLet12_6QNode_Int_8QNode_Int_1lizzieLet12_6QNode_Int_9QNode_Int_1t1a8Y_1lizzieLet12_6QNode_Int_5QNode_Int_1lizzieLet12_6QNode_Int_7QNode_Int_1lizzieLet12_6QNode_Int_4QNode_Int_1lizzieLet12_6QNode_Int_6QNode_Int_1lizzieLet12_6QNode_Int_10QNode_Int_1t2a8Z_1lizzieLet12_6QNode_Int_11QNode_Int_1t3a90_1Lcall_f_f_Int_Int3_bufchan_buf :
                                   lizzieLet12_6QNode_Int_8QNode_Int_1lizzieLet12_6QNode_Int_9QNode_Int_1t1a8Y_1lizzieLet12_6QNode_Int_5QNode_Int_1lizzieLet12_6QNode_Int_7QNode_Int_1lizzieLet12_6QNode_Int_4QNode_Int_1lizzieLet12_6QNode_Int_6QNode_Int_1lizzieLet12_6QNode_Int_10QNode_Int_1t2a8Z_1lizzieLet12_6QNode_Int_11QNode_Int_1t3a90_1Lcall_f_f_Int_Int3_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNode_Int_8QNode_Int_1lizzieLet12_6QNode_Int_9QNode_Int_1t1a8Y_1lizzieLet12_6QNode_Int_5QNode_Int_1lizzieLet12_6QNode_Int_7QNode_Int_1lizzieLet12_6QNode_Int_4QNode_Int_1lizzieLet12_6QNode_Int_6QNode_Int_1lizzieLet12_6QNode_Int_10QNode_Int_1t2a8Z_1lizzieLet12_6QNode_Int_11QNode_Int_1t3a90_1Lcall_f_f_Int_Int3_bufchan_buf <= {115'd0,
                                                                                                                                                                                                                                                                                                                                                        1'd0};
    else
      if ((lizzieLet30_1_argbuf_r && lizzieLet12_6QNode_Int_8QNode_Int_1lizzieLet12_6QNode_Int_9QNode_Int_1t1a8Y_1lizzieLet12_6QNode_Int_5QNode_Int_1lizzieLet12_6QNode_Int_7QNode_Int_1lizzieLet12_6QNode_Int_4QNode_Int_1lizzieLet12_6QNode_Int_6QNode_Int_1lizzieLet12_6QNode_Int_10QNode_Int_1t2a8Z_1lizzieLet12_6QNode_Int_11QNode_Int_1t3a90_1Lcall_f_f_Int_Int3_bufchan_buf[0]))
        lizzieLet12_6QNode_Int_8QNode_Int_1lizzieLet12_6QNode_Int_9QNode_Int_1t1a8Y_1lizzieLet12_6QNode_Int_5QNode_Int_1lizzieLet12_6QNode_Int_7QNode_Int_1lizzieLet12_6QNode_Int_4QNode_Int_1lizzieLet12_6QNode_Int_6QNode_Int_1lizzieLet12_6QNode_Int_10QNode_Int_1t2a8Z_1lizzieLet12_6QNode_Int_11QNode_Int_1t3a90_1Lcall_f_f_Int_Int3_bufchan_buf <= {115'd0,
                                                                                                                                                                                                                                                                                                                                                          1'd0};
      else if (((! lizzieLet30_1_argbuf_r) && (! lizzieLet12_6QNode_Int_8QNode_Int_1lizzieLet12_6QNode_Int_9QNode_Int_1t1a8Y_1lizzieLet12_6QNode_Int_5QNode_Int_1lizzieLet12_6QNode_Int_7QNode_Int_1lizzieLet12_6QNode_Int_4QNode_Int_1lizzieLet12_6QNode_Int_6QNode_Int_1lizzieLet12_6QNode_Int_10QNode_Int_1t2a8Z_1lizzieLet12_6QNode_Int_11QNode_Int_1t3a90_1Lcall_f_f_Int_Int3_bufchan_buf[0])))
        lizzieLet12_6QNode_Int_8QNode_Int_1lizzieLet12_6QNode_Int_9QNode_Int_1t1a8Y_1lizzieLet12_6QNode_Int_5QNode_Int_1lizzieLet12_6QNode_Int_7QNode_Int_1lizzieLet12_6QNode_Int_4QNode_Int_1lizzieLet12_6QNode_Int_6QNode_Int_1lizzieLet12_6QNode_Int_10QNode_Int_1t2a8Z_1lizzieLet12_6QNode_Int_11QNode_Int_1t3a90_1Lcall_f_f_Int_Int3_bufchan_buf <= lizzieLet12_6QNode_Int_8QNode_Int_1lizzieLet12_6QNode_Int_9QNode_Int_1t1a8Y_1lizzieLet12_6QNode_Int_5QNode_Int_1lizzieLet12_6QNode_Int_7QNode_Int_1lizzieLet12_6QNode_Int_4QNode_Int_1lizzieLet12_6QNode_Int_6QNode_Int_1lizzieLet12_6QNode_Int_10QNode_Int_1t2a8Z_1lizzieLet12_6QNode_Int_11QNode_Int_1t3a90_1Lcall_f_f_Int_Int3_bufchan_d;
  
  /* buf (Ty Pointer_CTf_f_Int_Int) : (lizzieLet12_6QNode_Int_8QNone_Int,Pointer_CTf_f_Int_Int) > (lizzieLet12_6QNode_Int_8QNone_Int_1_argbuf,Pointer_CTf_f_Int_Int) */
  Pointer_CTf_f_Int_Int_t lizzieLet12_6QNode_Int_8QNone_Int_bufchan_d;
  logic lizzieLet12_6QNode_Int_8QNone_Int_bufchan_r;
  assign lizzieLet12_6QNode_Int_8QNone_Int_r = ((! lizzieLet12_6QNode_Int_8QNone_Int_bufchan_d[0]) || lizzieLet12_6QNode_Int_8QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNode_Int_8QNone_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet12_6QNode_Int_8QNone_Int_r)
        lizzieLet12_6QNode_Int_8QNone_Int_bufchan_d <= lizzieLet12_6QNode_Int_8QNone_Int_d;
  Pointer_CTf_f_Int_Int_t lizzieLet12_6QNode_Int_8QNone_Int_bufchan_buf;
  assign lizzieLet12_6QNode_Int_8QNone_Int_bufchan_r = (! lizzieLet12_6QNode_Int_8QNone_Int_bufchan_buf[0]);
  assign lizzieLet12_6QNode_Int_8QNone_Int_1_argbuf_d = (lizzieLet12_6QNode_Int_8QNone_Int_bufchan_buf[0] ? lizzieLet12_6QNode_Int_8QNone_Int_bufchan_buf :
                                                         lizzieLet12_6QNode_Int_8QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNode_Int_8QNone_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet12_6QNode_Int_8QNone_Int_1_argbuf_r && lizzieLet12_6QNode_Int_8QNone_Int_bufchan_buf[0]))
        lizzieLet12_6QNode_Int_8QNone_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet12_6QNode_Int_8QNone_Int_1_argbuf_r) && (! lizzieLet12_6QNode_Int_8QNone_Int_bufchan_buf[0])))
        lizzieLet12_6QNode_Int_8QNone_Int_bufchan_buf <= lizzieLet12_6QNode_Int_8QNone_Int_bufchan_d;
  
  /* buf (Ty Pointer_CTf_f_Int_Int) : (lizzieLet12_6QNode_Int_8QVal_Int,Pointer_CTf_f_Int_Int) > (lizzieLet12_6QNode_Int_8QVal_Int_1_argbuf,Pointer_CTf_f_Int_Int) */
  Pointer_CTf_f_Int_Int_t lizzieLet12_6QNode_Int_8QVal_Int_bufchan_d;
  logic lizzieLet12_6QNode_Int_8QVal_Int_bufchan_r;
  assign lizzieLet12_6QNode_Int_8QVal_Int_r = ((! lizzieLet12_6QNode_Int_8QVal_Int_bufchan_d[0]) || lizzieLet12_6QNode_Int_8QVal_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNode_Int_8QVal_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet12_6QNode_Int_8QVal_Int_r)
        lizzieLet12_6QNode_Int_8QVal_Int_bufchan_d <= lizzieLet12_6QNode_Int_8QVal_Int_d;
  Pointer_CTf_f_Int_Int_t lizzieLet12_6QNode_Int_8QVal_Int_bufchan_buf;
  assign lizzieLet12_6QNode_Int_8QVal_Int_bufchan_r = (! lizzieLet12_6QNode_Int_8QVal_Int_bufchan_buf[0]);
  assign lizzieLet12_6QNode_Int_8QVal_Int_1_argbuf_d = (lizzieLet12_6QNode_Int_8QVal_Int_bufchan_buf[0] ? lizzieLet12_6QNode_Int_8QVal_Int_bufchan_buf :
                                                        lizzieLet12_6QNode_Int_8QVal_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNode_Int_8QVal_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet12_6QNode_Int_8QVal_Int_1_argbuf_r && lizzieLet12_6QNode_Int_8QVal_Int_bufchan_buf[0]))
        lizzieLet12_6QNode_Int_8QVal_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet12_6QNode_Int_8QVal_Int_1_argbuf_r) && (! lizzieLet12_6QNode_Int_8QVal_Int_bufchan_buf[0])))
        lizzieLet12_6QNode_Int_8QVal_Int_bufchan_buf <= lizzieLet12_6QNode_Int_8QVal_Int_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_QTree_Int) : (lizzieLet12_6QNode_Int_9,QTree_Int) (q1a8T_destruct,Pointer_QTree_Int) > [(lizzieLet12_6QNode_Int_9QNone_Int,Pointer_QTree_Int),
                                                                                                          (_40,Pointer_QTree_Int),
                                                                                                          (lizzieLet12_6QNode_Int_9QNode_Int,Pointer_QTree_Int),
                                                                                                          (_39,Pointer_QTree_Int)] */
  logic [3:0] q1a8T_destruct_onehotd;
  always_comb
    if ((lizzieLet12_6QNode_Int_9_d[0] && q1a8T_destruct_d[0]))
      unique case (lizzieLet12_6QNode_Int_9_d[2:1])
        2'd0: q1a8T_destruct_onehotd = 4'd1;
        2'd1: q1a8T_destruct_onehotd = 4'd2;
        2'd2: q1a8T_destruct_onehotd = 4'd4;
        2'd3: q1a8T_destruct_onehotd = 4'd8;
        default: q1a8T_destruct_onehotd = 4'd0;
      endcase
    else q1a8T_destruct_onehotd = 4'd0;
  assign lizzieLet12_6QNode_Int_9QNone_Int_d = {q1a8T_destruct_d[16:1],
                                                q1a8T_destruct_onehotd[0]};
  assign _40_d = {q1a8T_destruct_d[16:1], q1a8T_destruct_onehotd[1]};
  assign lizzieLet12_6QNode_Int_9QNode_Int_d = {q1a8T_destruct_d[16:1],
                                                q1a8T_destruct_onehotd[2]};
  assign _39_d = {q1a8T_destruct_d[16:1], q1a8T_destruct_onehotd[3]};
  assign q1a8T_destruct_r = (| (q1a8T_destruct_onehotd & {_39_r,
                                                          lizzieLet12_6QNode_Int_9QNode_Int_r,
                                                          _40_r,
                                                          lizzieLet12_6QNode_Int_9QNone_Int_r}));
  assign lizzieLet12_6QNode_Int_9_r = q1a8T_destruct_r;
  
  /* buf (Ty Pointer_QTree_Int) : (lizzieLet12_6QNode_Int_9QNone_Int,Pointer_QTree_Int) > (lizzieLet12_6QNode_Int_9QNone_Int_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t lizzieLet12_6QNode_Int_9QNone_Int_bufchan_d;
  logic lizzieLet12_6QNode_Int_9QNone_Int_bufchan_r;
  assign lizzieLet12_6QNode_Int_9QNone_Int_r = ((! lizzieLet12_6QNode_Int_9QNone_Int_bufchan_d[0]) || lizzieLet12_6QNode_Int_9QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNode_Int_9QNone_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet12_6QNode_Int_9QNone_Int_r)
        lizzieLet12_6QNode_Int_9QNone_Int_bufchan_d <= lizzieLet12_6QNode_Int_9QNone_Int_d;
  Pointer_QTree_Int_t lizzieLet12_6QNode_Int_9QNone_Int_bufchan_buf;
  assign lizzieLet12_6QNode_Int_9QNone_Int_bufchan_r = (! lizzieLet12_6QNode_Int_9QNone_Int_bufchan_buf[0]);
  assign lizzieLet12_6QNode_Int_9QNone_Int_1_argbuf_d = (lizzieLet12_6QNode_Int_9QNone_Int_bufchan_buf[0] ? lizzieLet12_6QNode_Int_9QNone_Int_bufchan_buf :
                                                         lizzieLet12_6QNode_Int_9QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNode_Int_9QNone_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet12_6QNode_Int_9QNone_Int_1_argbuf_r && lizzieLet12_6QNode_Int_9QNone_Int_bufchan_buf[0]))
        lizzieLet12_6QNode_Int_9QNone_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet12_6QNode_Int_9QNone_Int_1_argbuf_r) && (! lizzieLet12_6QNode_Int_9QNone_Int_bufchan_buf[0])))
        lizzieLet12_6QNode_Int_9QNone_Int_bufchan_buf <= lizzieLet12_6QNode_Int_9QNone_Int_bufchan_d;
  
  /* fork (Ty QTree_Int) : (lizzieLet12_6QNone_Int,QTree_Int) > [(lizzieLet12_6QNone_Int_1,QTree_Int),
                                                            (lizzieLet12_6QNone_Int_2,QTree_Int),
                                                            (lizzieLet12_6QNone_Int_3,QTree_Int),
                                                            (lizzieLet12_6QNone_Int_4,QTree_Int),
                                                            (lizzieLet12_6QNone_Int_5,QTree_Int),
                                                            (lizzieLet12_6QNone_Int_6,QTree_Int)] */
  logic [5:0] lizzieLet12_6QNone_Int_emitted;
  logic [5:0] lizzieLet12_6QNone_Int_done;
  assign lizzieLet12_6QNone_Int_1_d = {lizzieLet12_6QNone_Int_d[66:1],
                                       (lizzieLet12_6QNone_Int_d[0] && (! lizzieLet12_6QNone_Int_emitted[0]))};
  assign lizzieLet12_6QNone_Int_2_d = {lizzieLet12_6QNone_Int_d[66:1],
                                       (lizzieLet12_6QNone_Int_d[0] && (! lizzieLet12_6QNone_Int_emitted[1]))};
  assign lizzieLet12_6QNone_Int_3_d = {lizzieLet12_6QNone_Int_d[66:1],
                                       (lizzieLet12_6QNone_Int_d[0] && (! lizzieLet12_6QNone_Int_emitted[2]))};
  assign lizzieLet12_6QNone_Int_4_d = {lizzieLet12_6QNone_Int_d[66:1],
                                       (lizzieLet12_6QNone_Int_d[0] && (! lizzieLet12_6QNone_Int_emitted[3]))};
  assign lizzieLet12_6QNone_Int_5_d = {lizzieLet12_6QNone_Int_d[66:1],
                                       (lizzieLet12_6QNone_Int_d[0] && (! lizzieLet12_6QNone_Int_emitted[4]))};
  assign lizzieLet12_6QNone_Int_6_d = {lizzieLet12_6QNone_Int_d[66:1],
                                       (lizzieLet12_6QNone_Int_d[0] && (! lizzieLet12_6QNone_Int_emitted[5]))};
  assign lizzieLet12_6QNone_Int_done = (lizzieLet12_6QNone_Int_emitted | ({lizzieLet12_6QNone_Int_6_d[0],
                                                                           lizzieLet12_6QNone_Int_5_d[0],
                                                                           lizzieLet12_6QNone_Int_4_d[0],
                                                                           lizzieLet12_6QNone_Int_3_d[0],
                                                                           lizzieLet12_6QNone_Int_2_d[0],
                                                                           lizzieLet12_6QNone_Int_1_d[0]} & {lizzieLet12_6QNone_Int_6_r,
                                                                                                             lizzieLet12_6QNone_Int_5_r,
                                                                                                             lizzieLet12_6QNone_Int_4_r,
                                                                                                             lizzieLet12_6QNone_Int_3_r,
                                                                                                             lizzieLet12_6QNone_Int_2_r,
                                                                                                             lizzieLet12_6QNone_Int_1_r}));
  assign lizzieLet12_6QNone_Int_r = (& lizzieLet12_6QNone_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet12_6QNone_Int_emitted <= 6'd0;
    else
      lizzieLet12_6QNone_Int_emitted <= (lizzieLet12_6QNone_Int_r ? 6'd0 :
                                         lizzieLet12_6QNone_Int_done);
  
  /* destruct (Ty QTree_Int,
          Dcon QNode_Int) : (lizzieLet12_6QNone_Int_1QNode_Int,QTree_Int) > [(tla8J_destruct,Pointer_QTree_Int),
                                                                             (tra8K_destruct,Pointer_QTree_Int),
                                                                             (bla8L_destruct,Pointer_QTree_Int),
                                                                             (bra8M_destruct,Pointer_QTree_Int)] */
  logic [3:0] lizzieLet12_6QNone_Int_1QNode_Int_emitted;
  logic [3:0] lizzieLet12_6QNone_Int_1QNode_Int_done;
  assign tla8J_destruct_d = {lizzieLet12_6QNone_Int_1QNode_Int_d[18:3],
                             (lizzieLet12_6QNone_Int_1QNode_Int_d[0] && (! lizzieLet12_6QNone_Int_1QNode_Int_emitted[0]))};
  assign tra8K_destruct_d = {lizzieLet12_6QNone_Int_1QNode_Int_d[34:19],
                             (lizzieLet12_6QNone_Int_1QNode_Int_d[0] && (! lizzieLet12_6QNone_Int_1QNode_Int_emitted[1]))};
  assign bla8L_destruct_d = {lizzieLet12_6QNone_Int_1QNode_Int_d[50:35],
                             (lizzieLet12_6QNone_Int_1QNode_Int_d[0] && (! lizzieLet12_6QNone_Int_1QNode_Int_emitted[2]))};
  assign bra8M_destruct_d = {lizzieLet12_6QNone_Int_1QNode_Int_d[66:51],
                             (lizzieLet12_6QNone_Int_1QNode_Int_d[0] && (! lizzieLet12_6QNone_Int_1QNode_Int_emitted[3]))};
  assign lizzieLet12_6QNone_Int_1QNode_Int_done = (lizzieLet12_6QNone_Int_1QNode_Int_emitted | ({bra8M_destruct_d[0],
                                                                                                 bla8L_destruct_d[0],
                                                                                                 tra8K_destruct_d[0],
                                                                                                 tla8J_destruct_d[0]} & {bra8M_destruct_r,
                                                                                                                         bla8L_destruct_r,
                                                                                                                         tra8K_destruct_r,
                                                                                                                         tla8J_destruct_r}));
  assign lizzieLet12_6QNone_Int_1QNode_Int_r = (& lizzieLet12_6QNone_Int_1QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNone_Int_1QNode_Int_emitted <= 4'd0;
    else
      lizzieLet12_6QNone_Int_1QNode_Int_emitted <= (lizzieLet12_6QNone_Int_1QNode_Int_r ? 4'd0 :
                                                    lizzieLet12_6QNone_Int_1QNode_Int_done);
  
  /* destruct (Ty QTree_Int,
          Dcon QVal_Int) : (lizzieLet12_6QNone_Int_1QVal_Int,QTree_Int) > [(va8I_destruct,Int)] */
  assign va8I_destruct_d = {lizzieLet12_6QNone_Int_1QVal_Int_d[34:3],
                            lizzieLet12_6QNone_Int_1QVal_Int_d[0]};
  assign lizzieLet12_6QNone_Int_1QVal_Int_r = va8I_destruct_r;
  
  /* demux (Ty QTree_Int,
       Ty QTree_Int) : (lizzieLet12_6QNone_Int_2,QTree_Int) (lizzieLet12_6QNone_Int_1,QTree_Int) > [(_38,QTree_Int),
                                                                                                    (lizzieLet12_6QNone_Int_1QVal_Int,QTree_Int),
                                                                                                    (lizzieLet12_6QNone_Int_1QNode_Int,QTree_Int),
                                                                                                    (_37,QTree_Int)] */
  logic [3:0] lizzieLet12_6QNone_Int_1_onehotd;
  always_comb
    if ((lizzieLet12_6QNone_Int_2_d[0] && lizzieLet12_6QNone_Int_1_d[0]))
      unique case (lizzieLet12_6QNone_Int_2_d[2:1])
        2'd0: lizzieLet12_6QNone_Int_1_onehotd = 4'd1;
        2'd1: lizzieLet12_6QNone_Int_1_onehotd = 4'd2;
        2'd2: lizzieLet12_6QNone_Int_1_onehotd = 4'd4;
        2'd3: lizzieLet12_6QNone_Int_1_onehotd = 4'd8;
        default: lizzieLet12_6QNone_Int_1_onehotd = 4'd0;
      endcase
    else lizzieLet12_6QNone_Int_1_onehotd = 4'd0;
  assign _38_d = {lizzieLet12_6QNone_Int_1_d[66:1],
                  lizzieLet12_6QNone_Int_1_onehotd[0]};
  assign lizzieLet12_6QNone_Int_1QVal_Int_d = {lizzieLet12_6QNone_Int_1_d[66:1],
                                               lizzieLet12_6QNone_Int_1_onehotd[1]};
  assign lizzieLet12_6QNone_Int_1QNode_Int_d = {lizzieLet12_6QNone_Int_1_d[66:1],
                                                lizzieLet12_6QNone_Int_1_onehotd[2]};
  assign _37_d = {lizzieLet12_6QNone_Int_1_d[66:1],
                  lizzieLet12_6QNone_Int_1_onehotd[3]};
  assign lizzieLet12_6QNone_Int_1_r = (| (lizzieLet12_6QNone_Int_1_onehotd & {_37_r,
                                                                              lizzieLet12_6QNone_Int_1QNode_Int_r,
                                                                              lizzieLet12_6QNone_Int_1QVal_Int_r,
                                                                              _38_r}));
  assign lizzieLet12_6QNone_Int_2_r = lizzieLet12_6QNone_Int_1_r;
  
  /* demux (Ty QTree_Int,
       Ty Go) : (lizzieLet12_6QNone_Int_3,QTree_Int) (lizzieLet12_3QNone_Int,Go) > [(lizzieLet12_6QNone_Int_3QNone_Int,Go),
                                                                                    (lizzieLet12_6QNone_Int_3QVal_Int,Go),
                                                                                    (lizzieLet12_6QNone_Int_3QNode_Int,Go),
                                                                                    (lizzieLet12_6QNone_Int_3QError_Int,Go)] */
  logic [3:0] lizzieLet12_3QNone_Int_onehotd;
  always_comb
    if ((lizzieLet12_6QNone_Int_3_d[0] && lizzieLet12_3QNone_Int_d[0]))
      unique case (lizzieLet12_6QNone_Int_3_d[2:1])
        2'd0: lizzieLet12_3QNone_Int_onehotd = 4'd1;
        2'd1: lizzieLet12_3QNone_Int_onehotd = 4'd2;
        2'd2: lizzieLet12_3QNone_Int_onehotd = 4'd4;
        2'd3: lizzieLet12_3QNone_Int_onehotd = 4'd8;
        default: lizzieLet12_3QNone_Int_onehotd = 4'd0;
      endcase
    else lizzieLet12_3QNone_Int_onehotd = 4'd0;
  assign lizzieLet12_6QNone_Int_3QNone_Int_d = lizzieLet12_3QNone_Int_onehotd[0];
  assign lizzieLet12_6QNone_Int_3QVal_Int_d = lizzieLet12_3QNone_Int_onehotd[1];
  assign lizzieLet12_6QNone_Int_3QNode_Int_d = lizzieLet12_3QNone_Int_onehotd[2];
  assign lizzieLet12_6QNone_Int_3QError_Int_d = lizzieLet12_3QNone_Int_onehotd[3];
  assign lizzieLet12_3QNone_Int_r = (| (lizzieLet12_3QNone_Int_onehotd & {lizzieLet12_6QNone_Int_3QError_Int_r,
                                                                          lizzieLet12_6QNone_Int_3QNode_Int_r,
                                                                          lizzieLet12_6QNone_Int_3QVal_Int_r,
                                                                          lizzieLet12_6QNone_Int_3QNone_Int_r}));
  assign lizzieLet12_6QNone_Int_3_r = lizzieLet12_3QNone_Int_r;
  
  /* fork (Ty Go) : (lizzieLet12_6QNone_Int_3QError_Int,Go) > [(lizzieLet12_6QNone_Int_3QError_Int_1,Go),
                                                          (lizzieLet12_6QNone_Int_3QError_Int_2,Go)] */
  logic [1:0] lizzieLet12_6QNone_Int_3QError_Int_emitted;
  logic [1:0] lizzieLet12_6QNone_Int_3QError_Int_done;
  assign lizzieLet12_6QNone_Int_3QError_Int_1_d = (lizzieLet12_6QNone_Int_3QError_Int_d[0] && (! lizzieLet12_6QNone_Int_3QError_Int_emitted[0]));
  assign lizzieLet12_6QNone_Int_3QError_Int_2_d = (lizzieLet12_6QNone_Int_3QError_Int_d[0] && (! lizzieLet12_6QNone_Int_3QError_Int_emitted[1]));
  assign lizzieLet12_6QNone_Int_3QError_Int_done = (lizzieLet12_6QNone_Int_3QError_Int_emitted | ({lizzieLet12_6QNone_Int_3QError_Int_2_d[0],
                                                                                                   lizzieLet12_6QNone_Int_3QError_Int_1_d[0]} & {lizzieLet12_6QNone_Int_3QError_Int_2_r,
                                                                                                                                                 lizzieLet12_6QNone_Int_3QError_Int_1_r}));
  assign lizzieLet12_6QNone_Int_3QError_Int_r = (& lizzieLet12_6QNone_Int_3QError_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNone_Int_3QError_Int_emitted <= 2'd0;
    else
      lizzieLet12_6QNone_Int_3QError_Int_emitted <= (lizzieLet12_6QNone_Int_3QError_Int_r ? 2'd0 :
                                                     lizzieLet12_6QNone_Int_3QError_Int_done);
  
  /* dcon (Ty QTree_Int,
      Dcon QError_Int) : [(lizzieLet12_6QNone_Int_3QError_Int_1,Go)] > (lizzieLet12_6QNone_Int_3QError_Int_1QError_Int,QTree_Int) */
  assign lizzieLet12_6QNone_Int_3QError_Int_1QError_Int_d = QError_Int_dc((& {lizzieLet12_6QNone_Int_3QError_Int_1_d[0]}), lizzieLet12_6QNone_Int_3QError_Int_1_d);
  assign {lizzieLet12_6QNone_Int_3QError_Int_1_r} = {1 {(lizzieLet12_6QNone_Int_3QError_Int_1QError_Int_r && lizzieLet12_6QNone_Int_3QError_Int_1QError_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (lizzieLet12_6QNone_Int_3QError_Int_1QError_Int,QTree_Int) > (lizzieLet18_1_argbuf,QTree_Int) */
  QTree_Int_t lizzieLet12_6QNone_Int_3QError_Int_1QError_Int_bufchan_d;
  logic lizzieLet12_6QNone_Int_3QError_Int_1QError_Int_bufchan_r;
  assign lizzieLet12_6QNone_Int_3QError_Int_1QError_Int_r = ((! lizzieLet12_6QNone_Int_3QError_Int_1QError_Int_bufchan_d[0]) || lizzieLet12_6QNone_Int_3QError_Int_1QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNone_Int_3QError_Int_1QError_Int_bufchan_d <= {66'd0,
                                                                   1'd0};
    else
      if (lizzieLet12_6QNone_Int_3QError_Int_1QError_Int_r)
        lizzieLet12_6QNone_Int_3QError_Int_1QError_Int_bufchan_d <= lizzieLet12_6QNone_Int_3QError_Int_1QError_Int_d;
  QTree_Int_t lizzieLet12_6QNone_Int_3QError_Int_1QError_Int_bufchan_buf;
  assign lizzieLet12_6QNone_Int_3QError_Int_1QError_Int_bufchan_r = (! lizzieLet12_6QNone_Int_3QError_Int_1QError_Int_bufchan_buf[0]);
  assign lizzieLet18_1_argbuf_d = (lizzieLet12_6QNone_Int_3QError_Int_1QError_Int_bufchan_buf[0] ? lizzieLet12_6QNone_Int_3QError_Int_1QError_Int_bufchan_buf :
                                   lizzieLet12_6QNone_Int_3QError_Int_1QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNone_Int_3QError_Int_1QError_Int_bufchan_buf <= {66'd0,
                                                                     1'd0};
    else
      if ((lizzieLet18_1_argbuf_r && lizzieLet12_6QNone_Int_3QError_Int_1QError_Int_bufchan_buf[0]))
        lizzieLet12_6QNone_Int_3QError_Int_1QError_Int_bufchan_buf <= {66'd0,
                                                                       1'd0};
      else if (((! lizzieLet18_1_argbuf_r) && (! lizzieLet12_6QNone_Int_3QError_Int_1QError_Int_bufchan_buf[0])))
        lizzieLet12_6QNone_Int_3QError_Int_1QError_Int_bufchan_buf <= lizzieLet12_6QNone_Int_3QError_Int_1QError_Int_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet12_6QNone_Int_3QError_Int_2,Go) > (lizzieLet12_6QNone_Int_3QError_Int_2_argbuf,Go) */
  Go_t lizzieLet12_6QNone_Int_3QError_Int_2_bufchan_d;
  logic lizzieLet12_6QNone_Int_3QError_Int_2_bufchan_r;
  assign lizzieLet12_6QNone_Int_3QError_Int_2_r = ((! lizzieLet12_6QNone_Int_3QError_Int_2_bufchan_d[0]) || lizzieLet12_6QNone_Int_3QError_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNone_Int_3QError_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet12_6QNone_Int_3QError_Int_2_r)
        lizzieLet12_6QNone_Int_3QError_Int_2_bufchan_d <= lizzieLet12_6QNone_Int_3QError_Int_2_d;
  Go_t lizzieLet12_6QNone_Int_3QError_Int_2_bufchan_buf;
  assign lizzieLet12_6QNone_Int_3QError_Int_2_bufchan_r = (! lizzieLet12_6QNone_Int_3QError_Int_2_bufchan_buf[0]);
  assign lizzieLet12_6QNone_Int_3QError_Int_2_argbuf_d = (lizzieLet12_6QNone_Int_3QError_Int_2_bufchan_buf[0] ? lizzieLet12_6QNone_Int_3QError_Int_2_bufchan_buf :
                                                          lizzieLet12_6QNone_Int_3QError_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNone_Int_3QError_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet12_6QNone_Int_3QError_Int_2_argbuf_r && lizzieLet12_6QNone_Int_3QError_Int_2_bufchan_buf[0]))
        lizzieLet12_6QNone_Int_3QError_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet12_6QNone_Int_3QError_Int_2_argbuf_r) && (! lizzieLet12_6QNone_Int_3QError_Int_2_bufchan_buf[0])))
        lizzieLet12_6QNone_Int_3QError_Int_2_bufchan_buf <= lizzieLet12_6QNone_Int_3QError_Int_2_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet12_6QNone_Int_3QNode_Int,Go) > [(lizzieLet12_6QNone_Int_3QNode_Int_1,Go),
                                                         (lizzieLet12_6QNone_Int_3QNode_Int_2,Go),
                                                         (lizzieLet12_6QNone_Int_3QNode_Int_3,Go),
                                                         (lizzieLet12_6QNone_Int_3QNode_Int_4,Go),
                                                         (lizzieLet12_6QNone_Int_3QNode_Int_5,Go)] */
  logic [4:0] lizzieLet12_6QNone_Int_3QNode_Int_emitted;
  logic [4:0] lizzieLet12_6QNone_Int_3QNode_Int_done;
  assign lizzieLet12_6QNone_Int_3QNode_Int_1_d = (lizzieLet12_6QNone_Int_3QNode_Int_d[0] && (! lizzieLet12_6QNone_Int_3QNode_Int_emitted[0]));
  assign lizzieLet12_6QNone_Int_3QNode_Int_2_d = (lizzieLet12_6QNone_Int_3QNode_Int_d[0] && (! lizzieLet12_6QNone_Int_3QNode_Int_emitted[1]));
  assign lizzieLet12_6QNone_Int_3QNode_Int_3_d = (lizzieLet12_6QNone_Int_3QNode_Int_d[0] && (! lizzieLet12_6QNone_Int_3QNode_Int_emitted[2]));
  assign lizzieLet12_6QNone_Int_3QNode_Int_4_d = (lizzieLet12_6QNone_Int_3QNode_Int_d[0] && (! lizzieLet12_6QNone_Int_3QNode_Int_emitted[3]));
  assign lizzieLet12_6QNone_Int_3QNode_Int_5_d = (lizzieLet12_6QNone_Int_3QNode_Int_d[0] && (! lizzieLet12_6QNone_Int_3QNode_Int_emitted[4]));
  assign lizzieLet12_6QNone_Int_3QNode_Int_done = (lizzieLet12_6QNone_Int_3QNode_Int_emitted | ({lizzieLet12_6QNone_Int_3QNode_Int_5_d[0],
                                                                                                 lizzieLet12_6QNone_Int_3QNode_Int_4_d[0],
                                                                                                 lizzieLet12_6QNone_Int_3QNode_Int_3_d[0],
                                                                                                 lizzieLet12_6QNone_Int_3QNode_Int_2_d[0],
                                                                                                 lizzieLet12_6QNone_Int_3QNode_Int_1_d[0]} & {lizzieLet12_6QNone_Int_3QNode_Int_5_r,
                                                                                                                                              lizzieLet12_6QNone_Int_3QNode_Int_4_r,
                                                                                                                                              lizzieLet12_6QNone_Int_3QNode_Int_3_r,
                                                                                                                                              lizzieLet12_6QNone_Int_3QNode_Int_2_r,
                                                                                                                                              lizzieLet12_6QNone_Int_3QNode_Int_1_r}));
  assign lizzieLet12_6QNone_Int_3QNode_Int_r = (& lizzieLet12_6QNone_Int_3QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNone_Int_3QNode_Int_emitted <= 5'd0;
    else
      lizzieLet12_6QNone_Int_3QNode_Int_emitted <= (lizzieLet12_6QNone_Int_3QNode_Int_r ? 5'd0 :
                                                    lizzieLet12_6QNone_Int_3QNode_Int_done);
  
  /* buf (Ty Go) : (lizzieLet12_6QNone_Int_3QNode_Int_1,Go) > (lizzieLet12_6QNone_Int_3QNode_Int_1_argbuf,Go) */
  Go_t lizzieLet12_6QNone_Int_3QNode_Int_1_bufchan_d;
  logic lizzieLet12_6QNone_Int_3QNode_Int_1_bufchan_r;
  assign lizzieLet12_6QNone_Int_3QNode_Int_1_r = ((! lizzieLet12_6QNone_Int_3QNode_Int_1_bufchan_d[0]) || lizzieLet12_6QNone_Int_3QNode_Int_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNone_Int_3QNode_Int_1_bufchan_d <= 1'd0;
    else
      if (lizzieLet12_6QNone_Int_3QNode_Int_1_r)
        lizzieLet12_6QNone_Int_3QNode_Int_1_bufchan_d <= lizzieLet12_6QNone_Int_3QNode_Int_1_d;
  Go_t lizzieLet12_6QNone_Int_3QNode_Int_1_bufchan_buf;
  assign lizzieLet12_6QNone_Int_3QNode_Int_1_bufchan_r = (! lizzieLet12_6QNone_Int_3QNode_Int_1_bufchan_buf[0]);
  assign lizzieLet12_6QNone_Int_3QNode_Int_1_argbuf_d = (lizzieLet12_6QNone_Int_3QNode_Int_1_bufchan_buf[0] ? lizzieLet12_6QNone_Int_3QNode_Int_1_bufchan_buf :
                                                         lizzieLet12_6QNone_Int_3QNode_Int_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNone_Int_3QNode_Int_1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet12_6QNone_Int_3QNode_Int_1_argbuf_r && lizzieLet12_6QNone_Int_3QNode_Int_1_bufchan_buf[0]))
        lizzieLet12_6QNone_Int_3QNode_Int_1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet12_6QNone_Int_3QNode_Int_1_argbuf_r) && (! lizzieLet12_6QNone_Int_3QNode_Int_1_bufchan_buf[0])))
        lizzieLet12_6QNone_Int_3QNode_Int_1_bufchan_buf <= lizzieLet12_6QNone_Int_3QNode_Int_1_bufchan_d;
  
  /* dcon (Ty TupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int,
      Dcon TupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int) : [(lizzieLet12_6QNone_Int_3QNode_Int_1_argbuf,Go),
                                                                      (bra8M_1_argbuf,Pointer_QTree_Int),
                                                                      (lizzieLet12_6QNone_Int_4QNode_Int_1_argbuf,MyDTInt_Bool),
                                                                      (lizzieLet12_6QNone_Int_5QNode_Int_1_argbuf,MyDTInt_Int)] > (f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_1,TupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int) */
  assign \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_1_d  = TupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_dc((& {lizzieLet12_6QNone_Int_3QNode_Int_1_argbuf_d[0],
                                                                                                                                                                 bra8M_1_argbuf_d[0],
                                                                                                                                                                 lizzieLet12_6QNone_Int_4QNode_Int_1_argbuf_d[0],
                                                                                                                                                                 lizzieLet12_6QNone_Int_5QNode_Int_1_argbuf_d[0]}), lizzieLet12_6QNone_Int_3QNode_Int_1_argbuf_d, bra8M_1_argbuf_d, lizzieLet12_6QNone_Int_4QNode_Int_1_argbuf_d, lizzieLet12_6QNone_Int_5QNode_Int_1_argbuf_d);
  assign {lizzieLet12_6QNone_Int_3QNode_Int_1_argbuf_r,
          bra8M_1_argbuf_r,
          lizzieLet12_6QNone_Int_4QNode_Int_1_argbuf_r,
          lizzieLet12_6QNone_Int_5QNode_Int_1_argbuf_r} = {4 {(\f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_1_r  && \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_1_d [0])}};
  
  /* buf (Ty Go) : (lizzieLet12_6QNone_Int_3QNode_Int_2,Go) > (lizzieLet12_6QNone_Int_3QNode_Int_2_argbuf,Go) */
  Go_t lizzieLet12_6QNone_Int_3QNode_Int_2_bufchan_d;
  logic lizzieLet12_6QNone_Int_3QNode_Int_2_bufchan_r;
  assign lizzieLet12_6QNone_Int_3QNode_Int_2_r = ((! lizzieLet12_6QNone_Int_3QNode_Int_2_bufchan_d[0]) || lizzieLet12_6QNone_Int_3QNode_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNone_Int_3QNode_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet12_6QNone_Int_3QNode_Int_2_r)
        lizzieLet12_6QNone_Int_3QNode_Int_2_bufchan_d <= lizzieLet12_6QNone_Int_3QNode_Int_2_d;
  Go_t lizzieLet12_6QNone_Int_3QNode_Int_2_bufchan_buf;
  assign lizzieLet12_6QNone_Int_3QNode_Int_2_bufchan_r = (! lizzieLet12_6QNone_Int_3QNode_Int_2_bufchan_buf[0]);
  assign lizzieLet12_6QNone_Int_3QNode_Int_2_argbuf_d = (lizzieLet12_6QNone_Int_3QNode_Int_2_bufchan_buf[0] ? lizzieLet12_6QNone_Int_3QNode_Int_2_bufchan_buf :
                                                         lizzieLet12_6QNone_Int_3QNode_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNone_Int_3QNode_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet12_6QNone_Int_3QNode_Int_2_argbuf_r && lizzieLet12_6QNone_Int_3QNode_Int_2_bufchan_buf[0]))
        lizzieLet12_6QNone_Int_3QNode_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet12_6QNone_Int_3QNode_Int_2_argbuf_r) && (! lizzieLet12_6QNone_Int_3QNode_Int_2_bufchan_buf[0])))
        lizzieLet12_6QNone_Int_3QNode_Int_2_bufchan_buf <= lizzieLet12_6QNone_Int_3QNode_Int_2_bufchan_d;
  
  /* dcon (Ty TupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int,
      Dcon TupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int) : [(lizzieLet12_6QNone_Int_3QNode_Int_2_argbuf,Go),
                                                                      (bla8L_1_argbuf,Pointer_QTree_Int),
                                                                      (lizzieLet12_6QNone_Int_4QNode_Int_2_argbuf,MyDTInt_Bool),
                                                                      (lizzieLet12_6QNone_Int_5QNode_Int_2_argbuf,MyDTInt_Int)] > (f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int2,TupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int) */
  assign \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int2_d  = TupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_dc((& {lizzieLet12_6QNone_Int_3QNode_Int_2_argbuf_d[0],
                                                                                                                                                                bla8L_1_argbuf_d[0],
                                                                                                                                                                lizzieLet12_6QNone_Int_4QNode_Int_2_argbuf_d[0],
                                                                                                                                                                lizzieLet12_6QNone_Int_5QNode_Int_2_argbuf_d[0]}), lizzieLet12_6QNone_Int_3QNode_Int_2_argbuf_d, bla8L_1_argbuf_d, lizzieLet12_6QNone_Int_4QNode_Int_2_argbuf_d, lizzieLet12_6QNone_Int_5QNode_Int_2_argbuf_d);
  assign {lizzieLet12_6QNone_Int_3QNode_Int_2_argbuf_r,
          bla8L_1_argbuf_r,
          lizzieLet12_6QNone_Int_4QNode_Int_2_argbuf_r,
          lizzieLet12_6QNone_Int_5QNode_Int_2_argbuf_r} = {4 {(\f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int2_r  && \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int2_d [0])}};
  
  /* buf (Ty Go) : (lizzieLet12_6QNone_Int_3QNode_Int_3,Go) > (lizzieLet12_6QNone_Int_3QNode_Int_3_argbuf,Go) */
  Go_t lizzieLet12_6QNone_Int_3QNode_Int_3_bufchan_d;
  logic lizzieLet12_6QNone_Int_3QNode_Int_3_bufchan_r;
  assign lizzieLet12_6QNone_Int_3QNode_Int_3_r = ((! lizzieLet12_6QNone_Int_3QNode_Int_3_bufchan_d[0]) || lizzieLet12_6QNone_Int_3QNode_Int_3_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNone_Int_3QNode_Int_3_bufchan_d <= 1'd0;
    else
      if (lizzieLet12_6QNone_Int_3QNode_Int_3_r)
        lizzieLet12_6QNone_Int_3QNode_Int_3_bufchan_d <= lizzieLet12_6QNone_Int_3QNode_Int_3_d;
  Go_t lizzieLet12_6QNone_Int_3QNode_Int_3_bufchan_buf;
  assign lizzieLet12_6QNone_Int_3QNode_Int_3_bufchan_r = (! lizzieLet12_6QNone_Int_3QNode_Int_3_bufchan_buf[0]);
  assign lizzieLet12_6QNone_Int_3QNode_Int_3_argbuf_d = (lizzieLet12_6QNone_Int_3QNode_Int_3_bufchan_buf[0] ? lizzieLet12_6QNone_Int_3QNode_Int_3_bufchan_buf :
                                                         lizzieLet12_6QNone_Int_3QNode_Int_3_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNone_Int_3QNode_Int_3_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet12_6QNone_Int_3QNode_Int_3_argbuf_r && lizzieLet12_6QNone_Int_3QNode_Int_3_bufchan_buf[0]))
        lizzieLet12_6QNone_Int_3QNode_Int_3_bufchan_buf <= 1'd0;
      else if (((! lizzieLet12_6QNone_Int_3QNode_Int_3_argbuf_r) && (! lizzieLet12_6QNone_Int_3QNode_Int_3_bufchan_buf[0])))
        lizzieLet12_6QNone_Int_3QNode_Int_3_bufchan_buf <= lizzieLet12_6QNone_Int_3QNode_Int_3_bufchan_d;
  
  /* dcon (Ty TupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int,
      Dcon TupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int) : [(lizzieLet12_6QNone_Int_3QNode_Int_3_argbuf,Go),
                                                                      (tra8K_1_argbuf,Pointer_QTree_Int),
                                                                      (lizzieLet12_6QNone_Int_4QNode_Int_3_argbuf,MyDTInt_Bool),
                                                                      (lizzieLet12_6QNone_Int_5QNode_Int_3_argbuf,MyDTInt_Int)] > (f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int3,TupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int) */
  assign \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int3_d  = TupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_dc((& {lizzieLet12_6QNone_Int_3QNode_Int_3_argbuf_d[0],
                                                                                                                                                                tra8K_1_argbuf_d[0],
                                                                                                                                                                lizzieLet12_6QNone_Int_4QNode_Int_3_argbuf_d[0],
                                                                                                                                                                lizzieLet12_6QNone_Int_5QNode_Int_3_argbuf_d[0]}), lizzieLet12_6QNone_Int_3QNode_Int_3_argbuf_d, tra8K_1_argbuf_d, lizzieLet12_6QNone_Int_4QNode_Int_3_argbuf_d, lizzieLet12_6QNone_Int_5QNode_Int_3_argbuf_d);
  assign {lizzieLet12_6QNone_Int_3QNode_Int_3_argbuf_r,
          tra8K_1_argbuf_r,
          lizzieLet12_6QNone_Int_4QNode_Int_3_argbuf_r,
          lizzieLet12_6QNone_Int_5QNode_Int_3_argbuf_r} = {4 {(\f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int3_r  && \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int3_d [0])}};
  
  /* buf (Ty Go) : (lizzieLet12_6QNone_Int_3QNode_Int_4,Go) > (lizzieLet12_6QNone_Int_3QNode_Int_4_argbuf,Go) */
  Go_t lizzieLet12_6QNone_Int_3QNode_Int_4_bufchan_d;
  logic lizzieLet12_6QNone_Int_3QNode_Int_4_bufchan_r;
  assign lizzieLet12_6QNone_Int_3QNode_Int_4_r = ((! lizzieLet12_6QNone_Int_3QNode_Int_4_bufchan_d[0]) || lizzieLet12_6QNone_Int_3QNode_Int_4_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNone_Int_3QNode_Int_4_bufchan_d <= 1'd0;
    else
      if (lizzieLet12_6QNone_Int_3QNode_Int_4_r)
        lizzieLet12_6QNone_Int_3QNode_Int_4_bufchan_d <= lizzieLet12_6QNone_Int_3QNode_Int_4_d;
  Go_t lizzieLet12_6QNone_Int_3QNode_Int_4_bufchan_buf;
  assign lizzieLet12_6QNone_Int_3QNode_Int_4_bufchan_r = (! lizzieLet12_6QNone_Int_3QNode_Int_4_bufchan_buf[0]);
  assign lizzieLet12_6QNone_Int_3QNode_Int_4_argbuf_d = (lizzieLet12_6QNone_Int_3QNode_Int_4_bufchan_buf[0] ? lizzieLet12_6QNone_Int_3QNode_Int_4_bufchan_buf :
                                                         lizzieLet12_6QNone_Int_3QNode_Int_4_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNone_Int_3QNode_Int_4_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet12_6QNone_Int_3QNode_Int_4_argbuf_r && lizzieLet12_6QNone_Int_3QNode_Int_4_bufchan_buf[0]))
        lizzieLet12_6QNone_Int_3QNode_Int_4_bufchan_buf <= 1'd0;
      else if (((! lizzieLet12_6QNone_Int_3QNode_Int_4_argbuf_r) && (! lizzieLet12_6QNone_Int_3QNode_Int_4_bufchan_buf[0])))
        lizzieLet12_6QNone_Int_3QNode_Int_4_bufchan_buf <= lizzieLet12_6QNone_Int_3QNode_Int_4_bufchan_d;
  
  /* dcon (Ty TupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int,
      Dcon TupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int) : [(lizzieLet12_6QNone_Int_3QNode_Int_4_argbuf,Go),
                                                                      (tla8J_1_argbuf,Pointer_QTree_Int),
                                                                      (lizzieLet12_6QNone_Int_4QNode_Int_4_argbuf,MyDTInt_Bool),
                                                                      (lizzieLet12_6QNone_Int_5QNode_Int_4_argbuf,MyDTInt_Int)] > (f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int4,TupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int) */
  assign \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int4_d  = TupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_dc((& {lizzieLet12_6QNone_Int_3QNode_Int_4_argbuf_d[0],
                                                                                                                                                                tla8J_1_argbuf_d[0],
                                                                                                                                                                lizzieLet12_6QNone_Int_4QNode_Int_4_argbuf_d[0],
                                                                                                                                                                lizzieLet12_6QNone_Int_5QNode_Int_4_argbuf_d[0]}), lizzieLet12_6QNone_Int_3QNode_Int_4_argbuf_d, tla8J_1_argbuf_d, lizzieLet12_6QNone_Int_4QNode_Int_4_argbuf_d, lizzieLet12_6QNone_Int_5QNode_Int_4_argbuf_d);
  assign {lizzieLet12_6QNone_Int_3QNode_Int_4_argbuf_r,
          tla8J_1_argbuf_r,
          lizzieLet12_6QNone_Int_4QNode_Int_4_argbuf_r,
          lizzieLet12_6QNone_Int_5QNode_Int_4_argbuf_r} = {4 {(\f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int4_r  && \f''''''''_f''''''''_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int4_d [0])}};
  
  /* buf (Ty Go) : (lizzieLet12_6QNone_Int_3QNode_Int_5,Go) > (lizzieLet12_6QNone_Int_3QNode_Int_5_argbuf,Go) */
  Go_t lizzieLet12_6QNone_Int_3QNode_Int_5_bufchan_d;
  logic lizzieLet12_6QNone_Int_3QNode_Int_5_bufchan_r;
  assign lizzieLet12_6QNone_Int_3QNode_Int_5_r = ((! lizzieLet12_6QNone_Int_3QNode_Int_5_bufchan_d[0]) || lizzieLet12_6QNone_Int_3QNode_Int_5_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNone_Int_3QNode_Int_5_bufchan_d <= 1'd0;
    else
      if (lizzieLet12_6QNone_Int_3QNode_Int_5_r)
        lizzieLet12_6QNone_Int_3QNode_Int_5_bufchan_d <= lizzieLet12_6QNone_Int_3QNode_Int_5_d;
  Go_t lizzieLet12_6QNone_Int_3QNode_Int_5_bufchan_buf;
  assign lizzieLet12_6QNone_Int_3QNode_Int_5_bufchan_r = (! lizzieLet12_6QNone_Int_3QNode_Int_5_bufchan_buf[0]);
  assign lizzieLet12_6QNone_Int_3QNode_Int_5_argbuf_d = (lizzieLet12_6QNone_Int_3QNode_Int_5_bufchan_buf[0] ? lizzieLet12_6QNone_Int_3QNode_Int_5_bufchan_buf :
                                                         lizzieLet12_6QNone_Int_3QNode_Int_5_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNone_Int_3QNode_Int_5_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet12_6QNone_Int_3QNode_Int_5_argbuf_r && lizzieLet12_6QNone_Int_3QNode_Int_5_bufchan_buf[0]))
        lizzieLet12_6QNone_Int_3QNode_Int_5_bufchan_buf <= 1'd0;
      else if (((! lizzieLet12_6QNone_Int_3QNode_Int_5_argbuf_r) && (! lizzieLet12_6QNone_Int_3QNode_Int_5_bufchan_buf[0])))
        lizzieLet12_6QNone_Int_3QNode_Int_5_bufchan_buf <= lizzieLet12_6QNone_Int_3QNode_Int_5_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet12_6QNone_Int_3QNone_Int,Go) > [(lizzieLet12_6QNone_Int_3QNone_Int_1,Go),
                                                         (lizzieLet12_6QNone_Int_3QNone_Int_2,Go)] */
  logic [1:0] lizzieLet12_6QNone_Int_3QNone_Int_emitted;
  logic [1:0] lizzieLet12_6QNone_Int_3QNone_Int_done;
  assign lizzieLet12_6QNone_Int_3QNone_Int_1_d = (lizzieLet12_6QNone_Int_3QNone_Int_d[0] && (! lizzieLet12_6QNone_Int_3QNone_Int_emitted[0]));
  assign lizzieLet12_6QNone_Int_3QNone_Int_2_d = (lizzieLet12_6QNone_Int_3QNone_Int_d[0] && (! lizzieLet12_6QNone_Int_3QNone_Int_emitted[1]));
  assign lizzieLet12_6QNone_Int_3QNone_Int_done = (lizzieLet12_6QNone_Int_3QNone_Int_emitted | ({lizzieLet12_6QNone_Int_3QNone_Int_2_d[0],
                                                                                                 lizzieLet12_6QNone_Int_3QNone_Int_1_d[0]} & {lizzieLet12_6QNone_Int_3QNone_Int_2_r,
                                                                                                                                              lizzieLet12_6QNone_Int_3QNone_Int_1_r}));
  assign lizzieLet12_6QNone_Int_3QNone_Int_r = (& lizzieLet12_6QNone_Int_3QNone_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNone_Int_3QNone_Int_emitted <= 2'd0;
    else
      lizzieLet12_6QNone_Int_3QNone_Int_emitted <= (lizzieLet12_6QNone_Int_3QNone_Int_r ? 2'd0 :
                                                    lizzieLet12_6QNone_Int_3QNone_Int_done);
  
  /* dcon (Ty QTree_Int,
      Dcon QNone_Int) : [(lizzieLet12_6QNone_Int_3QNone_Int_1,Go)] > (lizzieLet12_6QNone_Int_3QNone_Int_1QNone_Int,QTree_Int) */
  assign lizzieLet12_6QNone_Int_3QNone_Int_1QNone_Int_d = QNone_Int_dc((& {lizzieLet12_6QNone_Int_3QNone_Int_1_d[0]}), lizzieLet12_6QNone_Int_3QNone_Int_1_d);
  assign {lizzieLet12_6QNone_Int_3QNone_Int_1_r} = {1 {(lizzieLet12_6QNone_Int_3QNone_Int_1QNone_Int_r && lizzieLet12_6QNone_Int_3QNone_Int_1QNone_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (lizzieLet12_6QNone_Int_3QNone_Int_1QNone_Int,QTree_Int) > (lizzieLet14_1_argbuf,QTree_Int) */
  QTree_Int_t lizzieLet12_6QNone_Int_3QNone_Int_1QNone_Int_bufchan_d;
  logic lizzieLet12_6QNone_Int_3QNone_Int_1QNone_Int_bufchan_r;
  assign lizzieLet12_6QNone_Int_3QNone_Int_1QNone_Int_r = ((! lizzieLet12_6QNone_Int_3QNone_Int_1QNone_Int_bufchan_d[0]) || lizzieLet12_6QNone_Int_3QNone_Int_1QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNone_Int_3QNone_Int_1QNone_Int_bufchan_d <= {66'd0,
                                                                 1'd0};
    else
      if (lizzieLet12_6QNone_Int_3QNone_Int_1QNone_Int_r)
        lizzieLet12_6QNone_Int_3QNone_Int_1QNone_Int_bufchan_d <= lizzieLet12_6QNone_Int_3QNone_Int_1QNone_Int_d;
  QTree_Int_t lizzieLet12_6QNone_Int_3QNone_Int_1QNone_Int_bufchan_buf;
  assign lizzieLet12_6QNone_Int_3QNone_Int_1QNone_Int_bufchan_r = (! lizzieLet12_6QNone_Int_3QNone_Int_1QNone_Int_bufchan_buf[0]);
  assign lizzieLet14_1_argbuf_d = (lizzieLet12_6QNone_Int_3QNone_Int_1QNone_Int_bufchan_buf[0] ? lizzieLet12_6QNone_Int_3QNone_Int_1QNone_Int_bufchan_buf :
                                   lizzieLet12_6QNone_Int_3QNone_Int_1QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNone_Int_3QNone_Int_1QNone_Int_bufchan_buf <= {66'd0,
                                                                   1'd0};
    else
      if ((lizzieLet14_1_argbuf_r && lizzieLet12_6QNone_Int_3QNone_Int_1QNone_Int_bufchan_buf[0]))
        lizzieLet12_6QNone_Int_3QNone_Int_1QNone_Int_bufchan_buf <= {66'd0,
                                                                     1'd0};
      else if (((! lizzieLet14_1_argbuf_r) && (! lizzieLet12_6QNone_Int_3QNone_Int_1QNone_Int_bufchan_buf[0])))
        lizzieLet12_6QNone_Int_3QNone_Int_1QNone_Int_bufchan_buf <= lizzieLet12_6QNone_Int_3QNone_Int_1QNone_Int_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet12_6QNone_Int_3QNone_Int_2,Go) > (lizzieLet12_6QNone_Int_3QNone_Int_2_argbuf,Go) */
  Go_t lizzieLet12_6QNone_Int_3QNone_Int_2_bufchan_d;
  logic lizzieLet12_6QNone_Int_3QNone_Int_2_bufchan_r;
  assign lizzieLet12_6QNone_Int_3QNone_Int_2_r = ((! lizzieLet12_6QNone_Int_3QNone_Int_2_bufchan_d[0]) || lizzieLet12_6QNone_Int_3QNone_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNone_Int_3QNone_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet12_6QNone_Int_3QNone_Int_2_r)
        lizzieLet12_6QNone_Int_3QNone_Int_2_bufchan_d <= lizzieLet12_6QNone_Int_3QNone_Int_2_d;
  Go_t lizzieLet12_6QNone_Int_3QNone_Int_2_bufchan_buf;
  assign lizzieLet12_6QNone_Int_3QNone_Int_2_bufchan_r = (! lizzieLet12_6QNone_Int_3QNone_Int_2_bufchan_buf[0]);
  assign lizzieLet12_6QNone_Int_3QNone_Int_2_argbuf_d = (lizzieLet12_6QNone_Int_3QNone_Int_2_bufchan_buf[0] ? lizzieLet12_6QNone_Int_3QNone_Int_2_bufchan_buf :
                                                         lizzieLet12_6QNone_Int_3QNone_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNone_Int_3QNone_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet12_6QNone_Int_3QNone_Int_2_argbuf_r && lizzieLet12_6QNone_Int_3QNone_Int_2_bufchan_buf[0]))
        lizzieLet12_6QNone_Int_3QNone_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet12_6QNone_Int_3QNone_Int_2_argbuf_r) && (! lizzieLet12_6QNone_Int_3QNone_Int_2_bufchan_buf[0])))
        lizzieLet12_6QNone_Int_3QNone_Int_2_bufchan_buf <= lizzieLet12_6QNone_Int_3QNone_Int_2_bufchan_d;
  
  /* mergectrl (Ty C17,
           Ty Go) : [(lizzieLet12_6QNone_Int_3QNone_Int_2_argbuf,Go),
                     (lizzieLet44_3Lcall_f_f_Int_Int0_1_argbuf,Go),
                     (es_2_1_1MyFalse_2_argbuf,Go),
                     (es_2_1_1MyTrue_2_argbuf,Go),
                     (lizzieLet12_6QNone_Int_3QNode_Int_5_argbuf,Go),
                     (lizzieLet12_6QNone_Int_3QError_Int_2_argbuf,Go),
                     (es_10_1MyFalse_2_argbuf,Go),
                     (es_10_1MyTrue_2_argbuf,Go),
                     (es_19_1MyFalse_2_argbuf,Go),
                     (es_19_1MyTrue_2_argbuf,Go),
                     (es_14_1MyTrue_2_argbuf,Go),
                     (lizzieLet12_6QVal_Int_3QNode_Int_2_argbuf,Go),
                     (lizzieLet12_6QVal_Int_3QError_Int_2_argbuf,Go),
                     (lizzieLet12_6QNode_Int_3QNone_Int_5_argbuf,Go),
                     (lizzieLet12_6QNode_Int_3QVal_Int_2_argbuf,Go),
                     (lizzieLet12_6QNode_Int_3QError_Int_2_argbuf,Go),
                     (lizzieLet12_3QError_Int_2_argbuf,Go)] > (go_17_goMux_choice,C17) (go_17_goMux_data,Go) */
  logic [16:0] lizzieLet12_6QNone_Int_3QNone_Int_2_argbuf_select_d;
  assign lizzieLet12_6QNone_Int_3QNone_Int_2_argbuf_select_d = ((| lizzieLet12_6QNone_Int_3QNone_Int_2_argbuf_select_q) ? lizzieLet12_6QNone_Int_3QNone_Int_2_argbuf_select_q :
                                                                (lizzieLet12_6QNone_Int_3QNone_Int_2_argbuf_d[0] ? 17'd1 :
                                                                 (lizzieLet44_3Lcall_f_f_Int_Int0_1_argbuf_d[0] ? 17'd2 :
                                                                  (es_2_1_1MyFalse_2_argbuf_d[0] ? 17'd4 :
                                                                   (es_2_1_1MyTrue_2_argbuf_d[0] ? 17'd8 :
                                                                    (lizzieLet12_6QNone_Int_3QNode_Int_5_argbuf_d[0] ? 17'd16 :
                                                                     (lizzieLet12_6QNone_Int_3QError_Int_2_argbuf_d[0] ? 17'd32 :
                                                                      (es_10_1MyFalse_2_argbuf_d[0] ? 17'd64 :
                                                                       (es_10_1MyTrue_2_argbuf_d[0] ? 17'd128 :
                                                                        (es_19_1MyFalse_2_argbuf_d[0] ? 17'd256 :
                                                                         (es_19_1MyTrue_2_argbuf_d[0] ? 17'd512 :
                                                                          (es_14_1MyTrue_2_argbuf_d[0] ? 17'd1024 :
                                                                           (lizzieLet12_6QVal_Int_3QNode_Int_2_argbuf_d[0] ? 17'd2048 :
                                                                            (lizzieLet12_6QVal_Int_3QError_Int_2_argbuf_d[0] ? 17'd4096 :
                                                                             (lizzieLet12_6QNode_Int_3QNone_Int_5_argbuf_d[0] ? 17'd8192 :
                                                                              (lizzieLet12_6QNode_Int_3QVal_Int_2_argbuf_d[0] ? 17'd16384 :
                                                                               (lizzieLet12_6QNode_Int_3QError_Int_2_argbuf_d[0] ? 17'd32768 :
                                                                                (lizzieLet12_3QError_Int_2_argbuf_d[0] ? 17'd65536 :
                                                                                 17'd0))))))))))))))))));
  logic [16:0] lizzieLet12_6QNone_Int_3QNone_Int_2_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNone_Int_3QNone_Int_2_argbuf_select_q <= 17'd0;
    else
      lizzieLet12_6QNone_Int_3QNone_Int_2_argbuf_select_q <= (lizzieLet12_6QNone_Int_3QNone_Int_2_argbuf_done ? 17'd0 :
                                                              lizzieLet12_6QNone_Int_3QNone_Int_2_argbuf_select_d);
  logic [1:0] lizzieLet12_6QNone_Int_3QNone_Int_2_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNone_Int_3QNone_Int_2_argbuf_emit_q <= 2'd0;
    else
      lizzieLet12_6QNone_Int_3QNone_Int_2_argbuf_emit_q <= (lizzieLet12_6QNone_Int_3QNone_Int_2_argbuf_done ? 2'd0 :
                                                            lizzieLet12_6QNone_Int_3QNone_Int_2_argbuf_emit_d);
  logic [1:0] lizzieLet12_6QNone_Int_3QNone_Int_2_argbuf_emit_d;
  assign lizzieLet12_6QNone_Int_3QNone_Int_2_argbuf_emit_d = (lizzieLet12_6QNone_Int_3QNone_Int_2_argbuf_emit_q | ({go_17_goMux_choice_d[0],
                                                                                                                    go_17_goMux_data_d[0]} & {go_17_goMux_choice_r,
                                                                                                                                              go_17_goMux_data_r}));
  logic lizzieLet12_6QNone_Int_3QNone_Int_2_argbuf_done;
  assign lizzieLet12_6QNone_Int_3QNone_Int_2_argbuf_done = (& lizzieLet12_6QNone_Int_3QNone_Int_2_argbuf_emit_d);
  assign {lizzieLet12_3QError_Int_2_argbuf_r,
          lizzieLet12_6QNode_Int_3QError_Int_2_argbuf_r,
          lizzieLet12_6QNode_Int_3QVal_Int_2_argbuf_r,
          lizzieLet12_6QNode_Int_3QNone_Int_5_argbuf_r,
          lizzieLet12_6QVal_Int_3QError_Int_2_argbuf_r,
          lizzieLet12_6QVal_Int_3QNode_Int_2_argbuf_r,
          es_14_1MyTrue_2_argbuf_r,
          es_19_1MyTrue_2_argbuf_r,
          es_19_1MyFalse_2_argbuf_r,
          es_10_1MyTrue_2_argbuf_r,
          es_10_1MyFalse_2_argbuf_r,
          lizzieLet12_6QNone_Int_3QError_Int_2_argbuf_r,
          lizzieLet12_6QNone_Int_3QNode_Int_5_argbuf_r,
          es_2_1_1MyTrue_2_argbuf_r,
          es_2_1_1MyFalse_2_argbuf_r,
          lizzieLet44_3Lcall_f_f_Int_Int0_1_argbuf_r,
          lizzieLet12_6QNone_Int_3QNone_Int_2_argbuf_r} = (lizzieLet12_6QNone_Int_3QNone_Int_2_argbuf_done ? lizzieLet12_6QNone_Int_3QNone_Int_2_argbuf_select_d :
                                                           17'd0);
  assign go_17_goMux_data_d = ((lizzieLet12_6QNone_Int_3QNone_Int_2_argbuf_select_d[0] && (! lizzieLet12_6QNone_Int_3QNone_Int_2_argbuf_emit_q[0])) ? lizzieLet12_6QNone_Int_3QNone_Int_2_argbuf_d :
                               ((lizzieLet12_6QNone_Int_3QNone_Int_2_argbuf_select_d[1] && (! lizzieLet12_6QNone_Int_3QNone_Int_2_argbuf_emit_q[0])) ? lizzieLet44_3Lcall_f_f_Int_Int0_1_argbuf_d :
                                ((lizzieLet12_6QNone_Int_3QNone_Int_2_argbuf_select_d[2] && (! lizzieLet12_6QNone_Int_3QNone_Int_2_argbuf_emit_q[0])) ? es_2_1_1MyFalse_2_argbuf_d :
                                 ((lizzieLet12_6QNone_Int_3QNone_Int_2_argbuf_select_d[3] && (! lizzieLet12_6QNone_Int_3QNone_Int_2_argbuf_emit_q[0])) ? es_2_1_1MyTrue_2_argbuf_d :
                                  ((lizzieLet12_6QNone_Int_3QNone_Int_2_argbuf_select_d[4] && (! lizzieLet12_6QNone_Int_3QNone_Int_2_argbuf_emit_q[0])) ? lizzieLet12_6QNone_Int_3QNode_Int_5_argbuf_d :
                                   ((lizzieLet12_6QNone_Int_3QNone_Int_2_argbuf_select_d[5] && (! lizzieLet12_6QNone_Int_3QNone_Int_2_argbuf_emit_q[0])) ? lizzieLet12_6QNone_Int_3QError_Int_2_argbuf_d :
                                    ((lizzieLet12_6QNone_Int_3QNone_Int_2_argbuf_select_d[6] && (! lizzieLet12_6QNone_Int_3QNone_Int_2_argbuf_emit_q[0])) ? es_10_1MyFalse_2_argbuf_d :
                                     ((lizzieLet12_6QNone_Int_3QNone_Int_2_argbuf_select_d[7] && (! lizzieLet12_6QNone_Int_3QNone_Int_2_argbuf_emit_q[0])) ? es_10_1MyTrue_2_argbuf_d :
                                      ((lizzieLet12_6QNone_Int_3QNone_Int_2_argbuf_select_d[8] && (! lizzieLet12_6QNone_Int_3QNone_Int_2_argbuf_emit_q[0])) ? es_19_1MyFalse_2_argbuf_d :
                                       ((lizzieLet12_6QNone_Int_3QNone_Int_2_argbuf_select_d[9] && (! lizzieLet12_6QNone_Int_3QNone_Int_2_argbuf_emit_q[0])) ? es_19_1MyTrue_2_argbuf_d :
                                        ((lizzieLet12_6QNone_Int_3QNone_Int_2_argbuf_select_d[10] && (! lizzieLet12_6QNone_Int_3QNone_Int_2_argbuf_emit_q[0])) ? es_14_1MyTrue_2_argbuf_d :
                                         ((lizzieLet12_6QNone_Int_3QNone_Int_2_argbuf_select_d[11] && (! lizzieLet12_6QNone_Int_3QNone_Int_2_argbuf_emit_q[0])) ? lizzieLet12_6QVal_Int_3QNode_Int_2_argbuf_d :
                                          ((lizzieLet12_6QNone_Int_3QNone_Int_2_argbuf_select_d[12] && (! lizzieLet12_6QNone_Int_3QNone_Int_2_argbuf_emit_q[0])) ? lizzieLet12_6QVal_Int_3QError_Int_2_argbuf_d :
                                           ((lizzieLet12_6QNone_Int_3QNone_Int_2_argbuf_select_d[13] && (! lizzieLet12_6QNone_Int_3QNone_Int_2_argbuf_emit_q[0])) ? lizzieLet12_6QNode_Int_3QNone_Int_5_argbuf_d :
                                            ((lizzieLet12_6QNone_Int_3QNone_Int_2_argbuf_select_d[14] && (! lizzieLet12_6QNone_Int_3QNone_Int_2_argbuf_emit_q[0])) ? lizzieLet12_6QNode_Int_3QVal_Int_2_argbuf_d :
                                             ((lizzieLet12_6QNone_Int_3QNone_Int_2_argbuf_select_d[15] && (! lizzieLet12_6QNone_Int_3QNone_Int_2_argbuf_emit_q[0])) ? lizzieLet12_6QNode_Int_3QError_Int_2_argbuf_d :
                                              ((lizzieLet12_6QNone_Int_3QNone_Int_2_argbuf_select_d[16] && (! lizzieLet12_6QNone_Int_3QNone_Int_2_argbuf_emit_q[0])) ? lizzieLet12_3QError_Int_2_argbuf_d :
                                               1'd0)))))))))))))))));
  assign go_17_goMux_choice_d = ((lizzieLet12_6QNone_Int_3QNone_Int_2_argbuf_select_d[0] && (! lizzieLet12_6QNone_Int_3QNone_Int_2_argbuf_emit_q[1])) ? C1_17_dc(1'd1) :
                                 ((lizzieLet12_6QNone_Int_3QNone_Int_2_argbuf_select_d[1] && (! lizzieLet12_6QNone_Int_3QNone_Int_2_argbuf_emit_q[1])) ? C2_17_dc(1'd1) :
                                  ((lizzieLet12_6QNone_Int_3QNone_Int_2_argbuf_select_d[2] && (! lizzieLet12_6QNone_Int_3QNone_Int_2_argbuf_emit_q[1])) ? C3_17_dc(1'd1) :
                                   ((lizzieLet12_6QNone_Int_3QNone_Int_2_argbuf_select_d[3] && (! lizzieLet12_6QNone_Int_3QNone_Int_2_argbuf_emit_q[1])) ? C4_17_dc(1'd1) :
                                    ((lizzieLet12_6QNone_Int_3QNone_Int_2_argbuf_select_d[4] && (! lizzieLet12_6QNone_Int_3QNone_Int_2_argbuf_emit_q[1])) ? C5_17_dc(1'd1) :
                                     ((lizzieLet12_6QNone_Int_3QNone_Int_2_argbuf_select_d[5] && (! lizzieLet12_6QNone_Int_3QNone_Int_2_argbuf_emit_q[1])) ? C6_17_dc(1'd1) :
                                      ((lizzieLet12_6QNone_Int_3QNone_Int_2_argbuf_select_d[6] && (! lizzieLet12_6QNone_Int_3QNone_Int_2_argbuf_emit_q[1])) ? C7_17_dc(1'd1) :
                                       ((lizzieLet12_6QNone_Int_3QNone_Int_2_argbuf_select_d[7] && (! lizzieLet12_6QNone_Int_3QNone_Int_2_argbuf_emit_q[1])) ? C8_17_dc(1'd1) :
                                        ((lizzieLet12_6QNone_Int_3QNone_Int_2_argbuf_select_d[8] && (! lizzieLet12_6QNone_Int_3QNone_Int_2_argbuf_emit_q[1])) ? C9_17_dc(1'd1) :
                                         ((lizzieLet12_6QNone_Int_3QNone_Int_2_argbuf_select_d[9] && (! lizzieLet12_6QNone_Int_3QNone_Int_2_argbuf_emit_q[1])) ? C10_17_dc(1'd1) :
                                          ((lizzieLet12_6QNone_Int_3QNone_Int_2_argbuf_select_d[10] && (! lizzieLet12_6QNone_Int_3QNone_Int_2_argbuf_emit_q[1])) ? C11_17_dc(1'd1) :
                                           ((lizzieLet12_6QNone_Int_3QNone_Int_2_argbuf_select_d[11] && (! lizzieLet12_6QNone_Int_3QNone_Int_2_argbuf_emit_q[1])) ? C12_17_dc(1'd1) :
                                            ((lizzieLet12_6QNone_Int_3QNone_Int_2_argbuf_select_d[12] && (! lizzieLet12_6QNone_Int_3QNone_Int_2_argbuf_emit_q[1])) ? C13_17_dc(1'd1) :
                                             ((lizzieLet12_6QNone_Int_3QNone_Int_2_argbuf_select_d[13] && (! lizzieLet12_6QNone_Int_3QNone_Int_2_argbuf_emit_q[1])) ? C14_17_dc(1'd1) :
                                              ((lizzieLet12_6QNone_Int_3QNone_Int_2_argbuf_select_d[14] && (! lizzieLet12_6QNone_Int_3QNone_Int_2_argbuf_emit_q[1])) ? C15_17_dc(1'd1) :
                                               ((lizzieLet12_6QNone_Int_3QNone_Int_2_argbuf_select_d[15] && (! lizzieLet12_6QNone_Int_3QNone_Int_2_argbuf_emit_q[1])) ? C16_17_dc(1'd1) :
                                                ((lizzieLet12_6QNone_Int_3QNone_Int_2_argbuf_select_d[16] && (! lizzieLet12_6QNone_Int_3QNone_Int_2_argbuf_emit_q[1])) ? C17_17_dc(1'd1) :
                                                 {5'd0, 1'd0})))))))))))))))));
  
  /* fork (Ty Go) : (lizzieLet12_6QNone_Int_3QVal_Int,Go) > [(lizzieLet12_6QNone_Int_3QVal_Int_1,Go),
                                                        (lizzieLet12_6QNone_Int_3QVal_Int_2,Go),
                                                        (lizzieLet12_6QNone_Int_3QVal_Int_3,Go)] */
  logic [2:0] lizzieLet12_6QNone_Int_3QVal_Int_emitted;
  logic [2:0] lizzieLet12_6QNone_Int_3QVal_Int_done;
  assign lizzieLet12_6QNone_Int_3QVal_Int_1_d = (lizzieLet12_6QNone_Int_3QVal_Int_d[0] && (! lizzieLet12_6QNone_Int_3QVal_Int_emitted[0]));
  assign lizzieLet12_6QNone_Int_3QVal_Int_2_d = (lizzieLet12_6QNone_Int_3QVal_Int_d[0] && (! lizzieLet12_6QNone_Int_3QVal_Int_emitted[1]));
  assign lizzieLet12_6QNone_Int_3QVal_Int_3_d = (lizzieLet12_6QNone_Int_3QVal_Int_d[0] && (! lizzieLet12_6QNone_Int_3QVal_Int_emitted[2]));
  assign lizzieLet12_6QNone_Int_3QVal_Int_done = (lizzieLet12_6QNone_Int_3QVal_Int_emitted | ({lizzieLet12_6QNone_Int_3QVal_Int_3_d[0],
                                                                                               lizzieLet12_6QNone_Int_3QVal_Int_2_d[0],
                                                                                               lizzieLet12_6QNone_Int_3QVal_Int_1_d[0]} & {lizzieLet12_6QNone_Int_3QVal_Int_3_r,
                                                                                                                                           lizzieLet12_6QNone_Int_3QVal_Int_2_r,
                                                                                                                                           lizzieLet12_6QNone_Int_3QVal_Int_1_r}));
  assign lizzieLet12_6QNone_Int_3QVal_Int_r = (& lizzieLet12_6QNone_Int_3QVal_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNone_Int_3QVal_Int_emitted <= 3'd0;
    else
      lizzieLet12_6QNone_Int_3QVal_Int_emitted <= (lizzieLet12_6QNone_Int_3QVal_Int_r ? 3'd0 :
                                                   lizzieLet12_6QNone_Int_3QVal_Int_done);
  
  /* buf (Ty Go) : (lizzieLet12_6QNone_Int_3QVal_Int_1,Go) > (lizzieLet12_6QNone_Int_3QVal_Int_1_argbuf,Go) */
  Go_t lizzieLet12_6QNone_Int_3QVal_Int_1_bufchan_d;
  logic lizzieLet12_6QNone_Int_3QVal_Int_1_bufchan_r;
  assign lizzieLet12_6QNone_Int_3QVal_Int_1_r = ((! lizzieLet12_6QNone_Int_3QVal_Int_1_bufchan_d[0]) || lizzieLet12_6QNone_Int_3QVal_Int_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNone_Int_3QVal_Int_1_bufchan_d <= 1'd0;
    else
      if (lizzieLet12_6QNone_Int_3QVal_Int_1_r)
        lizzieLet12_6QNone_Int_3QVal_Int_1_bufchan_d <= lizzieLet12_6QNone_Int_3QVal_Int_1_d;
  Go_t lizzieLet12_6QNone_Int_3QVal_Int_1_bufchan_buf;
  assign lizzieLet12_6QNone_Int_3QVal_Int_1_bufchan_r = (! lizzieLet12_6QNone_Int_3QVal_Int_1_bufchan_buf[0]);
  assign lizzieLet12_6QNone_Int_3QVal_Int_1_argbuf_d = (lizzieLet12_6QNone_Int_3QVal_Int_1_bufchan_buf[0] ? lizzieLet12_6QNone_Int_3QVal_Int_1_bufchan_buf :
                                                        lizzieLet12_6QNone_Int_3QVal_Int_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNone_Int_3QVal_Int_1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet12_6QNone_Int_3QVal_Int_1_argbuf_r && lizzieLet12_6QNone_Int_3QVal_Int_1_bufchan_buf[0]))
        lizzieLet12_6QNone_Int_3QVal_Int_1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet12_6QNone_Int_3QVal_Int_1_argbuf_r) && (! lizzieLet12_6QNone_Int_3QVal_Int_1_bufchan_buf[0])))
        lizzieLet12_6QNone_Int_3QVal_Int_1_bufchan_buf <= lizzieLet12_6QNone_Int_3QVal_Int_1_bufchan_d;
  
  /* dcon (Ty TupGo___MyDTInt_Int___Int,
      Dcon TupGo___MyDTInt_Int___Int) : [(lizzieLet12_6QNone_Int_3QVal_Int_1_argbuf,Go),
                                         (lizzieLet12_6QNone_Int_5QVal_Int_1_argbuf,MyDTInt_Int),
                                         (va8I_1_argbuf,Int)] > (applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1,TupGo___MyDTInt_Int___Int) */
  assign applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_d = TupGo___MyDTInt_Int___Int_dc((& {lizzieLet12_6QNone_Int_3QVal_Int_1_argbuf_d[0],
                                                                                          lizzieLet12_6QNone_Int_5QVal_Int_1_argbuf_d[0],
                                                                                          va8I_1_argbuf_d[0]}), lizzieLet12_6QNone_Int_3QVal_Int_1_argbuf_d, lizzieLet12_6QNone_Int_5QVal_Int_1_argbuf_d, va8I_1_argbuf_d);
  assign {lizzieLet12_6QNone_Int_3QVal_Int_1_argbuf_r,
          lizzieLet12_6QNone_Int_5QVal_Int_1_argbuf_r,
          va8I_1_argbuf_r} = {3 {(applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_r && applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_d[0])}};
  
  /* buf (Ty Go) : (lizzieLet12_6QNone_Int_3QVal_Int_2,Go) > (lizzieLet12_6QNone_Int_3QVal_Int_2_argbuf,Go) */
  Go_t lizzieLet12_6QNone_Int_3QVal_Int_2_bufchan_d;
  logic lizzieLet12_6QNone_Int_3QVal_Int_2_bufchan_r;
  assign lizzieLet12_6QNone_Int_3QVal_Int_2_r = ((! lizzieLet12_6QNone_Int_3QVal_Int_2_bufchan_d[0]) || lizzieLet12_6QNone_Int_3QVal_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNone_Int_3QVal_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet12_6QNone_Int_3QVal_Int_2_r)
        lizzieLet12_6QNone_Int_3QVal_Int_2_bufchan_d <= lizzieLet12_6QNone_Int_3QVal_Int_2_d;
  Go_t lizzieLet12_6QNone_Int_3QVal_Int_2_bufchan_buf;
  assign lizzieLet12_6QNone_Int_3QVal_Int_2_bufchan_r = (! lizzieLet12_6QNone_Int_3QVal_Int_2_bufchan_buf[0]);
  assign lizzieLet12_6QNone_Int_3QVal_Int_2_argbuf_d = (lizzieLet12_6QNone_Int_3QVal_Int_2_bufchan_buf[0] ? lizzieLet12_6QNone_Int_3QVal_Int_2_bufchan_buf :
                                                        lizzieLet12_6QNone_Int_3QVal_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNone_Int_3QVal_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet12_6QNone_Int_3QVal_Int_2_argbuf_r && lizzieLet12_6QNone_Int_3QVal_Int_2_bufchan_buf[0]))
        lizzieLet12_6QNone_Int_3QVal_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet12_6QNone_Int_3QVal_Int_2_argbuf_r) && (! lizzieLet12_6QNone_Int_3QVal_Int_2_bufchan_buf[0])))
        lizzieLet12_6QNone_Int_3QVal_Int_2_bufchan_buf <= lizzieLet12_6QNone_Int_3QVal_Int_2_bufchan_d;
  
  /* dcon (Ty TupGo___MyDTInt_Bool___Int,
      Dcon TupGo___MyDTInt_Bool___Int) : [(lizzieLet12_6QNone_Int_3QVal_Int_2_argbuf,Go),
                                          (lizzieLet12_6QNone_Int_4QVal_Int_1_argbuf,MyDTInt_Bool),
                                          (es_1_1_1_argbuf,Int)] > (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1,TupGo___MyDTInt_Bool___Int) */
  assign applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_d = TupGo___MyDTInt_Bool___Int_dc((& {lizzieLet12_6QNone_Int_3QVal_Int_2_argbuf_d[0],
                                                                                             lizzieLet12_6QNone_Int_4QVal_Int_1_argbuf_d[0],
                                                                                             es_1_1_1_argbuf_d[0]}), lizzieLet12_6QNone_Int_3QVal_Int_2_argbuf_d, lizzieLet12_6QNone_Int_4QVal_Int_1_argbuf_d, es_1_1_1_argbuf_d);
  assign {lizzieLet12_6QNone_Int_3QVal_Int_2_argbuf_r,
          lizzieLet12_6QNone_Int_4QVal_Int_1_argbuf_r,
          es_1_1_1_argbuf_r} = {3 {(applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_r && applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_d[0])}};
  
  /* demux (Ty QTree_Int,
       Ty MyDTInt_Bool) : (lizzieLet12_6QNone_Int_4,QTree_Int) (lizzieLet12_5QNone_Int,MyDTInt_Bool) > [(_36,MyDTInt_Bool),
                                                                                                        (lizzieLet12_6QNone_Int_4QVal_Int,MyDTInt_Bool),
                                                                                                        (lizzieLet12_6QNone_Int_4QNode_Int,MyDTInt_Bool),
                                                                                                        (_35,MyDTInt_Bool)] */
  logic [3:0] lizzieLet12_5QNone_Int_onehotd;
  always_comb
    if ((lizzieLet12_6QNone_Int_4_d[0] && lizzieLet12_5QNone_Int_d[0]))
      unique case (lizzieLet12_6QNone_Int_4_d[2:1])
        2'd0: lizzieLet12_5QNone_Int_onehotd = 4'd1;
        2'd1: lizzieLet12_5QNone_Int_onehotd = 4'd2;
        2'd2: lizzieLet12_5QNone_Int_onehotd = 4'd4;
        2'd3: lizzieLet12_5QNone_Int_onehotd = 4'd8;
        default: lizzieLet12_5QNone_Int_onehotd = 4'd0;
      endcase
    else lizzieLet12_5QNone_Int_onehotd = 4'd0;
  assign _36_d = lizzieLet12_5QNone_Int_onehotd[0];
  assign lizzieLet12_6QNone_Int_4QVal_Int_d = lizzieLet12_5QNone_Int_onehotd[1];
  assign lizzieLet12_6QNone_Int_4QNode_Int_d = lizzieLet12_5QNone_Int_onehotd[2];
  assign _35_d = lizzieLet12_5QNone_Int_onehotd[3];
  assign lizzieLet12_5QNone_Int_r = (| (lizzieLet12_5QNone_Int_onehotd & {_35_r,
                                                                          lizzieLet12_6QNone_Int_4QNode_Int_r,
                                                                          lizzieLet12_6QNone_Int_4QVal_Int_r,
                                                                          _36_r}));
  assign lizzieLet12_6QNone_Int_4_r = lizzieLet12_5QNone_Int_r;
  
  /* fork (Ty MyDTInt_Bool) : (lizzieLet12_6QNone_Int_4QNode_Int,MyDTInt_Bool) > [(lizzieLet12_6QNone_Int_4QNode_Int_1,MyDTInt_Bool),
                                                                             (lizzieLet12_6QNone_Int_4QNode_Int_2,MyDTInt_Bool),
                                                                             (lizzieLet12_6QNone_Int_4QNode_Int_3,MyDTInt_Bool),
                                                                             (lizzieLet12_6QNone_Int_4QNode_Int_4,MyDTInt_Bool)] */
  logic [3:0] lizzieLet12_6QNone_Int_4QNode_Int_emitted;
  logic [3:0] lizzieLet12_6QNone_Int_4QNode_Int_done;
  assign lizzieLet12_6QNone_Int_4QNode_Int_1_d = (lizzieLet12_6QNone_Int_4QNode_Int_d[0] && (! lizzieLet12_6QNone_Int_4QNode_Int_emitted[0]));
  assign lizzieLet12_6QNone_Int_4QNode_Int_2_d = (lizzieLet12_6QNone_Int_4QNode_Int_d[0] && (! lizzieLet12_6QNone_Int_4QNode_Int_emitted[1]));
  assign lizzieLet12_6QNone_Int_4QNode_Int_3_d = (lizzieLet12_6QNone_Int_4QNode_Int_d[0] && (! lizzieLet12_6QNone_Int_4QNode_Int_emitted[2]));
  assign lizzieLet12_6QNone_Int_4QNode_Int_4_d = (lizzieLet12_6QNone_Int_4QNode_Int_d[0] && (! lizzieLet12_6QNone_Int_4QNode_Int_emitted[3]));
  assign lizzieLet12_6QNone_Int_4QNode_Int_done = (lizzieLet12_6QNone_Int_4QNode_Int_emitted | ({lizzieLet12_6QNone_Int_4QNode_Int_4_d[0],
                                                                                                 lizzieLet12_6QNone_Int_4QNode_Int_3_d[0],
                                                                                                 lizzieLet12_6QNone_Int_4QNode_Int_2_d[0],
                                                                                                 lizzieLet12_6QNone_Int_4QNode_Int_1_d[0]} & {lizzieLet12_6QNone_Int_4QNode_Int_4_r,
                                                                                                                                              lizzieLet12_6QNone_Int_4QNode_Int_3_r,
                                                                                                                                              lizzieLet12_6QNone_Int_4QNode_Int_2_r,
                                                                                                                                              lizzieLet12_6QNone_Int_4QNode_Int_1_r}));
  assign lizzieLet12_6QNone_Int_4QNode_Int_r = (& lizzieLet12_6QNone_Int_4QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNone_Int_4QNode_Int_emitted <= 4'd0;
    else
      lizzieLet12_6QNone_Int_4QNode_Int_emitted <= (lizzieLet12_6QNone_Int_4QNode_Int_r ? 4'd0 :
                                                    lizzieLet12_6QNone_Int_4QNode_Int_done);
  
  /* buf (Ty MyDTInt_Bool) : (lizzieLet12_6QNone_Int_4QNode_Int_1,MyDTInt_Bool) > (lizzieLet12_6QNone_Int_4QNode_Int_1_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t lizzieLet12_6QNone_Int_4QNode_Int_1_bufchan_d;
  logic lizzieLet12_6QNone_Int_4QNode_Int_1_bufchan_r;
  assign lizzieLet12_6QNone_Int_4QNode_Int_1_r = ((! lizzieLet12_6QNone_Int_4QNode_Int_1_bufchan_d[0]) || lizzieLet12_6QNone_Int_4QNode_Int_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNone_Int_4QNode_Int_1_bufchan_d <= 1'd0;
    else
      if (lizzieLet12_6QNone_Int_4QNode_Int_1_r)
        lizzieLet12_6QNone_Int_4QNode_Int_1_bufchan_d <= lizzieLet12_6QNone_Int_4QNode_Int_1_d;
  MyDTInt_Bool_t lizzieLet12_6QNone_Int_4QNode_Int_1_bufchan_buf;
  assign lizzieLet12_6QNone_Int_4QNode_Int_1_bufchan_r = (! lizzieLet12_6QNone_Int_4QNode_Int_1_bufchan_buf[0]);
  assign lizzieLet12_6QNone_Int_4QNode_Int_1_argbuf_d = (lizzieLet12_6QNone_Int_4QNode_Int_1_bufchan_buf[0] ? lizzieLet12_6QNone_Int_4QNode_Int_1_bufchan_buf :
                                                         lizzieLet12_6QNone_Int_4QNode_Int_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNone_Int_4QNode_Int_1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet12_6QNone_Int_4QNode_Int_1_argbuf_r && lizzieLet12_6QNone_Int_4QNode_Int_1_bufchan_buf[0]))
        lizzieLet12_6QNone_Int_4QNode_Int_1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet12_6QNone_Int_4QNode_Int_1_argbuf_r) && (! lizzieLet12_6QNone_Int_4QNode_Int_1_bufchan_buf[0])))
        lizzieLet12_6QNone_Int_4QNode_Int_1_bufchan_buf <= lizzieLet12_6QNone_Int_4QNode_Int_1_bufchan_d;
  
  /* buf (Ty MyDTInt_Bool) : (lizzieLet12_6QNone_Int_4QNode_Int_2,MyDTInt_Bool) > (lizzieLet12_6QNone_Int_4QNode_Int_2_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t lizzieLet12_6QNone_Int_4QNode_Int_2_bufchan_d;
  logic lizzieLet12_6QNone_Int_4QNode_Int_2_bufchan_r;
  assign lizzieLet12_6QNone_Int_4QNode_Int_2_r = ((! lizzieLet12_6QNone_Int_4QNode_Int_2_bufchan_d[0]) || lizzieLet12_6QNone_Int_4QNode_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNone_Int_4QNode_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet12_6QNone_Int_4QNode_Int_2_r)
        lizzieLet12_6QNone_Int_4QNode_Int_2_bufchan_d <= lizzieLet12_6QNone_Int_4QNode_Int_2_d;
  MyDTInt_Bool_t lizzieLet12_6QNone_Int_4QNode_Int_2_bufchan_buf;
  assign lizzieLet12_6QNone_Int_4QNode_Int_2_bufchan_r = (! lizzieLet12_6QNone_Int_4QNode_Int_2_bufchan_buf[0]);
  assign lizzieLet12_6QNone_Int_4QNode_Int_2_argbuf_d = (lizzieLet12_6QNone_Int_4QNode_Int_2_bufchan_buf[0] ? lizzieLet12_6QNone_Int_4QNode_Int_2_bufchan_buf :
                                                         lizzieLet12_6QNone_Int_4QNode_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNone_Int_4QNode_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet12_6QNone_Int_4QNode_Int_2_argbuf_r && lizzieLet12_6QNone_Int_4QNode_Int_2_bufchan_buf[0]))
        lizzieLet12_6QNone_Int_4QNode_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet12_6QNone_Int_4QNode_Int_2_argbuf_r) && (! lizzieLet12_6QNone_Int_4QNode_Int_2_bufchan_buf[0])))
        lizzieLet12_6QNone_Int_4QNode_Int_2_bufchan_buf <= lizzieLet12_6QNone_Int_4QNode_Int_2_bufchan_d;
  
  /* buf (Ty MyDTInt_Bool) : (lizzieLet12_6QNone_Int_4QNode_Int_3,MyDTInt_Bool) > (lizzieLet12_6QNone_Int_4QNode_Int_3_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t lizzieLet12_6QNone_Int_4QNode_Int_3_bufchan_d;
  logic lizzieLet12_6QNone_Int_4QNode_Int_3_bufchan_r;
  assign lizzieLet12_6QNone_Int_4QNode_Int_3_r = ((! lizzieLet12_6QNone_Int_4QNode_Int_3_bufchan_d[0]) || lizzieLet12_6QNone_Int_4QNode_Int_3_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNone_Int_4QNode_Int_3_bufchan_d <= 1'd0;
    else
      if (lizzieLet12_6QNone_Int_4QNode_Int_3_r)
        lizzieLet12_6QNone_Int_4QNode_Int_3_bufchan_d <= lizzieLet12_6QNone_Int_4QNode_Int_3_d;
  MyDTInt_Bool_t lizzieLet12_6QNone_Int_4QNode_Int_3_bufchan_buf;
  assign lizzieLet12_6QNone_Int_4QNode_Int_3_bufchan_r = (! lizzieLet12_6QNone_Int_4QNode_Int_3_bufchan_buf[0]);
  assign lizzieLet12_6QNone_Int_4QNode_Int_3_argbuf_d = (lizzieLet12_6QNone_Int_4QNode_Int_3_bufchan_buf[0] ? lizzieLet12_6QNone_Int_4QNode_Int_3_bufchan_buf :
                                                         lizzieLet12_6QNone_Int_4QNode_Int_3_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNone_Int_4QNode_Int_3_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet12_6QNone_Int_4QNode_Int_3_argbuf_r && lizzieLet12_6QNone_Int_4QNode_Int_3_bufchan_buf[0]))
        lizzieLet12_6QNone_Int_4QNode_Int_3_bufchan_buf <= 1'd0;
      else if (((! lizzieLet12_6QNone_Int_4QNode_Int_3_argbuf_r) && (! lizzieLet12_6QNone_Int_4QNode_Int_3_bufchan_buf[0])))
        lizzieLet12_6QNone_Int_4QNode_Int_3_bufchan_buf <= lizzieLet12_6QNone_Int_4QNode_Int_3_bufchan_d;
  
  /* buf (Ty MyDTInt_Bool) : (lizzieLet12_6QNone_Int_4QNode_Int_4,MyDTInt_Bool) > (lizzieLet12_6QNone_Int_4QNode_Int_4_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t lizzieLet12_6QNone_Int_4QNode_Int_4_bufchan_d;
  logic lizzieLet12_6QNone_Int_4QNode_Int_4_bufchan_r;
  assign lizzieLet12_6QNone_Int_4QNode_Int_4_r = ((! lizzieLet12_6QNone_Int_4QNode_Int_4_bufchan_d[0]) || lizzieLet12_6QNone_Int_4QNode_Int_4_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNone_Int_4QNode_Int_4_bufchan_d <= 1'd0;
    else
      if (lizzieLet12_6QNone_Int_4QNode_Int_4_r)
        lizzieLet12_6QNone_Int_4QNode_Int_4_bufchan_d <= lizzieLet12_6QNone_Int_4QNode_Int_4_d;
  MyDTInt_Bool_t lizzieLet12_6QNone_Int_4QNode_Int_4_bufchan_buf;
  assign lizzieLet12_6QNone_Int_4QNode_Int_4_bufchan_r = (! lizzieLet12_6QNone_Int_4QNode_Int_4_bufchan_buf[0]);
  assign lizzieLet12_6QNone_Int_4QNode_Int_4_argbuf_d = (lizzieLet12_6QNone_Int_4QNode_Int_4_bufchan_buf[0] ? lizzieLet12_6QNone_Int_4QNode_Int_4_bufchan_buf :
                                                         lizzieLet12_6QNone_Int_4QNode_Int_4_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNone_Int_4QNode_Int_4_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet12_6QNone_Int_4QNode_Int_4_argbuf_r && lizzieLet12_6QNone_Int_4QNode_Int_4_bufchan_buf[0]))
        lizzieLet12_6QNone_Int_4QNode_Int_4_bufchan_buf <= 1'd0;
      else if (((! lizzieLet12_6QNone_Int_4QNode_Int_4_argbuf_r) && (! lizzieLet12_6QNone_Int_4QNode_Int_4_bufchan_buf[0])))
        lizzieLet12_6QNone_Int_4QNode_Int_4_bufchan_buf <= lizzieLet12_6QNone_Int_4QNode_Int_4_bufchan_d;
  
  /* buf (Ty MyDTInt_Bool) : (lizzieLet12_6QNone_Int_4QVal_Int,MyDTInt_Bool) > (lizzieLet12_6QNone_Int_4QVal_Int_1_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t lizzieLet12_6QNone_Int_4QVal_Int_bufchan_d;
  logic lizzieLet12_6QNone_Int_4QVal_Int_bufchan_r;
  assign lizzieLet12_6QNone_Int_4QVal_Int_r = ((! lizzieLet12_6QNone_Int_4QVal_Int_bufchan_d[0]) || lizzieLet12_6QNone_Int_4QVal_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNone_Int_4QVal_Int_bufchan_d <= 1'd0;
    else
      if (lizzieLet12_6QNone_Int_4QVal_Int_r)
        lizzieLet12_6QNone_Int_4QVal_Int_bufchan_d <= lizzieLet12_6QNone_Int_4QVal_Int_d;
  MyDTInt_Bool_t lizzieLet12_6QNone_Int_4QVal_Int_bufchan_buf;
  assign lizzieLet12_6QNone_Int_4QVal_Int_bufchan_r = (! lizzieLet12_6QNone_Int_4QVal_Int_bufchan_buf[0]);
  assign lizzieLet12_6QNone_Int_4QVal_Int_1_argbuf_d = (lizzieLet12_6QNone_Int_4QVal_Int_bufchan_buf[0] ? lizzieLet12_6QNone_Int_4QVal_Int_bufchan_buf :
                                                        lizzieLet12_6QNone_Int_4QVal_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNone_Int_4QVal_Int_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet12_6QNone_Int_4QVal_Int_1_argbuf_r && lizzieLet12_6QNone_Int_4QVal_Int_bufchan_buf[0]))
        lizzieLet12_6QNone_Int_4QVal_Int_bufchan_buf <= 1'd0;
      else if (((! lizzieLet12_6QNone_Int_4QVal_Int_1_argbuf_r) && (! lizzieLet12_6QNone_Int_4QVal_Int_bufchan_buf[0])))
        lizzieLet12_6QNone_Int_4QVal_Int_bufchan_buf <= lizzieLet12_6QNone_Int_4QVal_Int_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty MyDTInt_Int) : (lizzieLet12_6QNone_Int_5,QTree_Int) (lizzieLet12_8QNone_Int,MyDTInt_Int) > [(_34,MyDTInt_Int),
                                                                                                      (lizzieLet12_6QNone_Int_5QVal_Int,MyDTInt_Int),
                                                                                                      (lizzieLet12_6QNone_Int_5QNode_Int,MyDTInt_Int),
                                                                                                      (_33,MyDTInt_Int)] */
  logic [3:0] lizzieLet12_8QNone_Int_onehotd;
  always_comb
    if ((lizzieLet12_6QNone_Int_5_d[0] && lizzieLet12_8QNone_Int_d[0]))
      unique case (lizzieLet12_6QNone_Int_5_d[2:1])
        2'd0: lizzieLet12_8QNone_Int_onehotd = 4'd1;
        2'd1: lizzieLet12_8QNone_Int_onehotd = 4'd2;
        2'd2: lizzieLet12_8QNone_Int_onehotd = 4'd4;
        2'd3: lizzieLet12_8QNone_Int_onehotd = 4'd8;
        default: lizzieLet12_8QNone_Int_onehotd = 4'd0;
      endcase
    else lizzieLet12_8QNone_Int_onehotd = 4'd0;
  assign _34_d = lizzieLet12_8QNone_Int_onehotd[0];
  assign lizzieLet12_6QNone_Int_5QVal_Int_d = lizzieLet12_8QNone_Int_onehotd[1];
  assign lizzieLet12_6QNone_Int_5QNode_Int_d = lizzieLet12_8QNone_Int_onehotd[2];
  assign _33_d = lizzieLet12_8QNone_Int_onehotd[3];
  assign lizzieLet12_8QNone_Int_r = (| (lizzieLet12_8QNone_Int_onehotd & {_33_r,
                                                                          lizzieLet12_6QNone_Int_5QNode_Int_r,
                                                                          lizzieLet12_6QNone_Int_5QVal_Int_r,
                                                                          _34_r}));
  assign lizzieLet12_6QNone_Int_5_r = lizzieLet12_8QNone_Int_r;
  
  /* fork (Ty MyDTInt_Int) : (lizzieLet12_6QNone_Int_5QNode_Int,MyDTInt_Int) > [(lizzieLet12_6QNone_Int_5QNode_Int_1,MyDTInt_Int),
                                                                           (lizzieLet12_6QNone_Int_5QNode_Int_2,MyDTInt_Int),
                                                                           (lizzieLet12_6QNone_Int_5QNode_Int_3,MyDTInt_Int),
                                                                           (lizzieLet12_6QNone_Int_5QNode_Int_4,MyDTInt_Int)] */
  logic [3:0] lizzieLet12_6QNone_Int_5QNode_Int_emitted;
  logic [3:0] lizzieLet12_6QNone_Int_5QNode_Int_done;
  assign lizzieLet12_6QNone_Int_5QNode_Int_1_d = (lizzieLet12_6QNone_Int_5QNode_Int_d[0] && (! lizzieLet12_6QNone_Int_5QNode_Int_emitted[0]));
  assign lizzieLet12_6QNone_Int_5QNode_Int_2_d = (lizzieLet12_6QNone_Int_5QNode_Int_d[0] && (! lizzieLet12_6QNone_Int_5QNode_Int_emitted[1]));
  assign lizzieLet12_6QNone_Int_5QNode_Int_3_d = (lizzieLet12_6QNone_Int_5QNode_Int_d[0] && (! lizzieLet12_6QNone_Int_5QNode_Int_emitted[2]));
  assign lizzieLet12_6QNone_Int_5QNode_Int_4_d = (lizzieLet12_6QNone_Int_5QNode_Int_d[0] && (! lizzieLet12_6QNone_Int_5QNode_Int_emitted[3]));
  assign lizzieLet12_6QNone_Int_5QNode_Int_done = (lizzieLet12_6QNone_Int_5QNode_Int_emitted | ({lizzieLet12_6QNone_Int_5QNode_Int_4_d[0],
                                                                                                 lizzieLet12_6QNone_Int_5QNode_Int_3_d[0],
                                                                                                 lizzieLet12_6QNone_Int_5QNode_Int_2_d[0],
                                                                                                 lizzieLet12_6QNone_Int_5QNode_Int_1_d[0]} & {lizzieLet12_6QNone_Int_5QNode_Int_4_r,
                                                                                                                                              lizzieLet12_6QNone_Int_5QNode_Int_3_r,
                                                                                                                                              lizzieLet12_6QNone_Int_5QNode_Int_2_r,
                                                                                                                                              lizzieLet12_6QNone_Int_5QNode_Int_1_r}));
  assign lizzieLet12_6QNone_Int_5QNode_Int_r = (& lizzieLet12_6QNone_Int_5QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNone_Int_5QNode_Int_emitted <= 4'd0;
    else
      lizzieLet12_6QNone_Int_5QNode_Int_emitted <= (lizzieLet12_6QNone_Int_5QNode_Int_r ? 4'd0 :
                                                    lizzieLet12_6QNone_Int_5QNode_Int_done);
  
  /* buf (Ty MyDTInt_Int) : (lizzieLet12_6QNone_Int_5QNode_Int_1,MyDTInt_Int) > (lizzieLet12_6QNone_Int_5QNode_Int_1_argbuf,MyDTInt_Int) */
  MyDTInt_Int_t lizzieLet12_6QNone_Int_5QNode_Int_1_bufchan_d;
  logic lizzieLet12_6QNone_Int_5QNode_Int_1_bufchan_r;
  assign lizzieLet12_6QNone_Int_5QNode_Int_1_r = ((! lizzieLet12_6QNone_Int_5QNode_Int_1_bufchan_d[0]) || lizzieLet12_6QNone_Int_5QNode_Int_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNone_Int_5QNode_Int_1_bufchan_d <= 1'd0;
    else
      if (lizzieLet12_6QNone_Int_5QNode_Int_1_r)
        lizzieLet12_6QNone_Int_5QNode_Int_1_bufchan_d <= lizzieLet12_6QNone_Int_5QNode_Int_1_d;
  MyDTInt_Int_t lizzieLet12_6QNone_Int_5QNode_Int_1_bufchan_buf;
  assign lizzieLet12_6QNone_Int_5QNode_Int_1_bufchan_r = (! lizzieLet12_6QNone_Int_5QNode_Int_1_bufchan_buf[0]);
  assign lizzieLet12_6QNone_Int_5QNode_Int_1_argbuf_d = (lizzieLet12_6QNone_Int_5QNode_Int_1_bufchan_buf[0] ? lizzieLet12_6QNone_Int_5QNode_Int_1_bufchan_buf :
                                                         lizzieLet12_6QNone_Int_5QNode_Int_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNone_Int_5QNode_Int_1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet12_6QNone_Int_5QNode_Int_1_argbuf_r && lizzieLet12_6QNone_Int_5QNode_Int_1_bufchan_buf[0]))
        lizzieLet12_6QNone_Int_5QNode_Int_1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet12_6QNone_Int_5QNode_Int_1_argbuf_r) && (! lizzieLet12_6QNone_Int_5QNode_Int_1_bufchan_buf[0])))
        lizzieLet12_6QNone_Int_5QNode_Int_1_bufchan_buf <= lizzieLet12_6QNone_Int_5QNode_Int_1_bufchan_d;
  
  /* buf (Ty MyDTInt_Int) : (lizzieLet12_6QNone_Int_5QNode_Int_2,MyDTInt_Int) > (lizzieLet12_6QNone_Int_5QNode_Int_2_argbuf,MyDTInt_Int) */
  MyDTInt_Int_t lizzieLet12_6QNone_Int_5QNode_Int_2_bufchan_d;
  logic lizzieLet12_6QNone_Int_5QNode_Int_2_bufchan_r;
  assign lizzieLet12_6QNone_Int_5QNode_Int_2_r = ((! lizzieLet12_6QNone_Int_5QNode_Int_2_bufchan_d[0]) || lizzieLet12_6QNone_Int_5QNode_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNone_Int_5QNode_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet12_6QNone_Int_5QNode_Int_2_r)
        lizzieLet12_6QNone_Int_5QNode_Int_2_bufchan_d <= lizzieLet12_6QNone_Int_5QNode_Int_2_d;
  MyDTInt_Int_t lizzieLet12_6QNone_Int_5QNode_Int_2_bufchan_buf;
  assign lizzieLet12_6QNone_Int_5QNode_Int_2_bufchan_r = (! lizzieLet12_6QNone_Int_5QNode_Int_2_bufchan_buf[0]);
  assign lizzieLet12_6QNone_Int_5QNode_Int_2_argbuf_d = (lizzieLet12_6QNone_Int_5QNode_Int_2_bufchan_buf[0] ? lizzieLet12_6QNone_Int_5QNode_Int_2_bufchan_buf :
                                                         lizzieLet12_6QNone_Int_5QNode_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNone_Int_5QNode_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet12_6QNone_Int_5QNode_Int_2_argbuf_r && lizzieLet12_6QNone_Int_5QNode_Int_2_bufchan_buf[0]))
        lizzieLet12_6QNone_Int_5QNode_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet12_6QNone_Int_5QNode_Int_2_argbuf_r) && (! lizzieLet12_6QNone_Int_5QNode_Int_2_bufchan_buf[0])))
        lizzieLet12_6QNone_Int_5QNode_Int_2_bufchan_buf <= lizzieLet12_6QNone_Int_5QNode_Int_2_bufchan_d;
  
  /* buf (Ty MyDTInt_Int) : (lizzieLet12_6QNone_Int_5QNode_Int_3,MyDTInt_Int) > (lizzieLet12_6QNone_Int_5QNode_Int_3_argbuf,MyDTInt_Int) */
  MyDTInt_Int_t lizzieLet12_6QNone_Int_5QNode_Int_3_bufchan_d;
  logic lizzieLet12_6QNone_Int_5QNode_Int_3_bufchan_r;
  assign lizzieLet12_6QNone_Int_5QNode_Int_3_r = ((! lizzieLet12_6QNone_Int_5QNode_Int_3_bufchan_d[0]) || lizzieLet12_6QNone_Int_5QNode_Int_3_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNone_Int_5QNode_Int_3_bufchan_d <= 1'd0;
    else
      if (lizzieLet12_6QNone_Int_5QNode_Int_3_r)
        lizzieLet12_6QNone_Int_5QNode_Int_3_bufchan_d <= lizzieLet12_6QNone_Int_5QNode_Int_3_d;
  MyDTInt_Int_t lizzieLet12_6QNone_Int_5QNode_Int_3_bufchan_buf;
  assign lizzieLet12_6QNone_Int_5QNode_Int_3_bufchan_r = (! lizzieLet12_6QNone_Int_5QNode_Int_3_bufchan_buf[0]);
  assign lizzieLet12_6QNone_Int_5QNode_Int_3_argbuf_d = (lizzieLet12_6QNone_Int_5QNode_Int_3_bufchan_buf[0] ? lizzieLet12_6QNone_Int_5QNode_Int_3_bufchan_buf :
                                                         lizzieLet12_6QNone_Int_5QNode_Int_3_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNone_Int_5QNode_Int_3_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet12_6QNone_Int_5QNode_Int_3_argbuf_r && lizzieLet12_6QNone_Int_5QNode_Int_3_bufchan_buf[0]))
        lizzieLet12_6QNone_Int_5QNode_Int_3_bufchan_buf <= 1'd0;
      else if (((! lizzieLet12_6QNone_Int_5QNode_Int_3_argbuf_r) && (! lizzieLet12_6QNone_Int_5QNode_Int_3_bufchan_buf[0])))
        lizzieLet12_6QNone_Int_5QNode_Int_3_bufchan_buf <= lizzieLet12_6QNone_Int_5QNode_Int_3_bufchan_d;
  
  /* buf (Ty MyDTInt_Int) : (lizzieLet12_6QNone_Int_5QNode_Int_4,MyDTInt_Int) > (lizzieLet12_6QNone_Int_5QNode_Int_4_argbuf,MyDTInt_Int) */
  MyDTInt_Int_t lizzieLet12_6QNone_Int_5QNode_Int_4_bufchan_d;
  logic lizzieLet12_6QNone_Int_5QNode_Int_4_bufchan_r;
  assign lizzieLet12_6QNone_Int_5QNode_Int_4_r = ((! lizzieLet12_6QNone_Int_5QNode_Int_4_bufchan_d[0]) || lizzieLet12_6QNone_Int_5QNode_Int_4_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNone_Int_5QNode_Int_4_bufchan_d <= 1'd0;
    else
      if (lizzieLet12_6QNone_Int_5QNode_Int_4_r)
        lizzieLet12_6QNone_Int_5QNode_Int_4_bufchan_d <= lizzieLet12_6QNone_Int_5QNode_Int_4_d;
  MyDTInt_Int_t lizzieLet12_6QNone_Int_5QNode_Int_4_bufchan_buf;
  assign lizzieLet12_6QNone_Int_5QNode_Int_4_bufchan_r = (! lizzieLet12_6QNone_Int_5QNode_Int_4_bufchan_buf[0]);
  assign lizzieLet12_6QNone_Int_5QNode_Int_4_argbuf_d = (lizzieLet12_6QNone_Int_5QNode_Int_4_bufchan_buf[0] ? lizzieLet12_6QNone_Int_5QNode_Int_4_bufchan_buf :
                                                         lizzieLet12_6QNone_Int_5QNode_Int_4_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNone_Int_5QNode_Int_4_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet12_6QNone_Int_5QNode_Int_4_argbuf_r && lizzieLet12_6QNone_Int_5QNode_Int_4_bufchan_buf[0]))
        lizzieLet12_6QNone_Int_5QNode_Int_4_bufchan_buf <= 1'd0;
      else if (((! lizzieLet12_6QNone_Int_5QNode_Int_4_argbuf_r) && (! lizzieLet12_6QNone_Int_5QNode_Int_4_bufchan_buf[0])))
        lizzieLet12_6QNone_Int_5QNode_Int_4_bufchan_buf <= lizzieLet12_6QNone_Int_5QNode_Int_4_bufchan_d;
  
  /* fork (Ty MyDTInt_Int) : (lizzieLet12_6QNone_Int_5QVal_Int,MyDTInt_Int) > [(lizzieLet12_6QNone_Int_5QVal_Int_1,MyDTInt_Int),
                                                                          (lizzieLet12_6QNone_Int_5QVal_Int_2,MyDTInt_Int)] */
  logic [1:0] lizzieLet12_6QNone_Int_5QVal_Int_emitted;
  logic [1:0] lizzieLet12_6QNone_Int_5QVal_Int_done;
  assign lizzieLet12_6QNone_Int_5QVal_Int_1_d = (lizzieLet12_6QNone_Int_5QVal_Int_d[0] && (! lizzieLet12_6QNone_Int_5QVal_Int_emitted[0]));
  assign lizzieLet12_6QNone_Int_5QVal_Int_2_d = (lizzieLet12_6QNone_Int_5QVal_Int_d[0] && (! lizzieLet12_6QNone_Int_5QVal_Int_emitted[1]));
  assign lizzieLet12_6QNone_Int_5QVal_Int_done = (lizzieLet12_6QNone_Int_5QVal_Int_emitted | ({lizzieLet12_6QNone_Int_5QVal_Int_2_d[0],
                                                                                               lizzieLet12_6QNone_Int_5QVal_Int_1_d[0]} & {lizzieLet12_6QNone_Int_5QVal_Int_2_r,
                                                                                                                                           lizzieLet12_6QNone_Int_5QVal_Int_1_r}));
  assign lizzieLet12_6QNone_Int_5QVal_Int_r = (& lizzieLet12_6QNone_Int_5QVal_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNone_Int_5QVal_Int_emitted <= 2'd0;
    else
      lizzieLet12_6QNone_Int_5QVal_Int_emitted <= (lizzieLet12_6QNone_Int_5QVal_Int_r ? 2'd0 :
                                                   lizzieLet12_6QNone_Int_5QVal_Int_done);
  
  /* buf (Ty MyDTInt_Int) : (lizzieLet12_6QNone_Int_5QVal_Int_1,MyDTInt_Int) > (lizzieLet12_6QNone_Int_5QVal_Int_1_argbuf,MyDTInt_Int) */
  MyDTInt_Int_t lizzieLet12_6QNone_Int_5QVal_Int_1_bufchan_d;
  logic lizzieLet12_6QNone_Int_5QVal_Int_1_bufchan_r;
  assign lizzieLet12_6QNone_Int_5QVal_Int_1_r = ((! lizzieLet12_6QNone_Int_5QVal_Int_1_bufchan_d[0]) || lizzieLet12_6QNone_Int_5QVal_Int_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNone_Int_5QVal_Int_1_bufchan_d <= 1'd0;
    else
      if (lizzieLet12_6QNone_Int_5QVal_Int_1_r)
        lizzieLet12_6QNone_Int_5QVal_Int_1_bufchan_d <= lizzieLet12_6QNone_Int_5QVal_Int_1_d;
  MyDTInt_Int_t lizzieLet12_6QNone_Int_5QVal_Int_1_bufchan_buf;
  assign lizzieLet12_6QNone_Int_5QVal_Int_1_bufchan_r = (! lizzieLet12_6QNone_Int_5QVal_Int_1_bufchan_buf[0]);
  assign lizzieLet12_6QNone_Int_5QVal_Int_1_argbuf_d = (lizzieLet12_6QNone_Int_5QVal_Int_1_bufchan_buf[0] ? lizzieLet12_6QNone_Int_5QVal_Int_1_bufchan_buf :
                                                        lizzieLet12_6QNone_Int_5QVal_Int_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNone_Int_5QVal_Int_1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet12_6QNone_Int_5QVal_Int_1_argbuf_r && lizzieLet12_6QNone_Int_5QVal_Int_1_bufchan_buf[0]))
        lizzieLet12_6QNone_Int_5QVal_Int_1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet12_6QNone_Int_5QVal_Int_1_argbuf_r) && (! lizzieLet12_6QNone_Int_5QVal_Int_1_bufchan_buf[0])))
        lizzieLet12_6QNone_Int_5QVal_Int_1_bufchan_buf <= lizzieLet12_6QNone_Int_5QVal_Int_1_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_CTf_f_Int_Int) : (lizzieLet12_6QNone_Int_6,QTree_Int) (lizzieLet12_9QNone_Int,Pointer_CTf_f_Int_Int) > [(lizzieLet12_6QNone_Int_6QNone_Int,Pointer_CTf_f_Int_Int),
                                                                                                                          (lizzieLet12_6QNone_Int_6QVal_Int,Pointer_CTf_f_Int_Int),
                                                                                                                          (lizzieLet12_6QNone_Int_6QNode_Int,Pointer_CTf_f_Int_Int),
                                                                                                                          (lizzieLet12_6QNone_Int_6QError_Int,Pointer_CTf_f_Int_Int)] */
  logic [3:0] lizzieLet12_9QNone_Int_onehotd;
  always_comb
    if ((lizzieLet12_6QNone_Int_6_d[0] && lizzieLet12_9QNone_Int_d[0]))
      unique case (lizzieLet12_6QNone_Int_6_d[2:1])
        2'd0: lizzieLet12_9QNone_Int_onehotd = 4'd1;
        2'd1: lizzieLet12_9QNone_Int_onehotd = 4'd2;
        2'd2: lizzieLet12_9QNone_Int_onehotd = 4'd4;
        2'd3: lizzieLet12_9QNone_Int_onehotd = 4'd8;
        default: lizzieLet12_9QNone_Int_onehotd = 4'd0;
      endcase
    else lizzieLet12_9QNone_Int_onehotd = 4'd0;
  assign lizzieLet12_6QNone_Int_6QNone_Int_d = {lizzieLet12_9QNone_Int_d[16:1],
                                                lizzieLet12_9QNone_Int_onehotd[0]};
  assign lizzieLet12_6QNone_Int_6QVal_Int_d = {lizzieLet12_9QNone_Int_d[16:1],
                                               lizzieLet12_9QNone_Int_onehotd[1]};
  assign lizzieLet12_6QNone_Int_6QNode_Int_d = {lizzieLet12_9QNone_Int_d[16:1],
                                                lizzieLet12_9QNone_Int_onehotd[2]};
  assign lizzieLet12_6QNone_Int_6QError_Int_d = {lizzieLet12_9QNone_Int_d[16:1],
                                                 lizzieLet12_9QNone_Int_onehotd[3]};
  assign lizzieLet12_9QNone_Int_r = (| (lizzieLet12_9QNone_Int_onehotd & {lizzieLet12_6QNone_Int_6QError_Int_r,
                                                                          lizzieLet12_6QNone_Int_6QNode_Int_r,
                                                                          lizzieLet12_6QNone_Int_6QVal_Int_r,
                                                                          lizzieLet12_6QNone_Int_6QNone_Int_r}));
  assign lizzieLet12_6QNone_Int_6_r = lizzieLet12_9QNone_Int_r;
  
  /* buf (Ty Pointer_CTf_f_Int_Int) : (lizzieLet12_6QNone_Int_6QError_Int,Pointer_CTf_f_Int_Int) > (lizzieLet12_6QNone_Int_6QError_Int_1_argbuf,Pointer_CTf_f_Int_Int) */
  Pointer_CTf_f_Int_Int_t lizzieLet12_6QNone_Int_6QError_Int_bufchan_d;
  logic lizzieLet12_6QNone_Int_6QError_Int_bufchan_r;
  assign lizzieLet12_6QNone_Int_6QError_Int_r = ((! lizzieLet12_6QNone_Int_6QError_Int_bufchan_d[0]) || lizzieLet12_6QNone_Int_6QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNone_Int_6QError_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet12_6QNone_Int_6QError_Int_r)
        lizzieLet12_6QNone_Int_6QError_Int_bufchan_d <= lizzieLet12_6QNone_Int_6QError_Int_d;
  Pointer_CTf_f_Int_Int_t lizzieLet12_6QNone_Int_6QError_Int_bufchan_buf;
  assign lizzieLet12_6QNone_Int_6QError_Int_bufchan_r = (! lizzieLet12_6QNone_Int_6QError_Int_bufchan_buf[0]);
  assign lizzieLet12_6QNone_Int_6QError_Int_1_argbuf_d = (lizzieLet12_6QNone_Int_6QError_Int_bufchan_buf[0] ? lizzieLet12_6QNone_Int_6QError_Int_bufchan_buf :
                                                          lizzieLet12_6QNone_Int_6QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNone_Int_6QError_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet12_6QNone_Int_6QError_Int_1_argbuf_r && lizzieLet12_6QNone_Int_6QError_Int_bufchan_buf[0]))
        lizzieLet12_6QNone_Int_6QError_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet12_6QNone_Int_6QError_Int_1_argbuf_r) && (! lizzieLet12_6QNone_Int_6QError_Int_bufchan_buf[0])))
        lizzieLet12_6QNone_Int_6QError_Int_bufchan_buf <= lizzieLet12_6QNone_Int_6QError_Int_bufchan_d;
  
  /* buf (Ty Pointer_CTf_f_Int_Int) : (lizzieLet12_6QNone_Int_6QNode_Int,Pointer_CTf_f_Int_Int) > (lizzieLet12_6QNone_Int_6QNode_Int_1_argbuf,Pointer_CTf_f_Int_Int) */
  Pointer_CTf_f_Int_Int_t lizzieLet12_6QNone_Int_6QNode_Int_bufchan_d;
  logic lizzieLet12_6QNone_Int_6QNode_Int_bufchan_r;
  assign lizzieLet12_6QNone_Int_6QNode_Int_r = ((! lizzieLet12_6QNone_Int_6QNode_Int_bufchan_d[0]) || lizzieLet12_6QNone_Int_6QNode_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNone_Int_6QNode_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet12_6QNone_Int_6QNode_Int_r)
        lizzieLet12_6QNone_Int_6QNode_Int_bufchan_d <= lizzieLet12_6QNone_Int_6QNode_Int_d;
  Pointer_CTf_f_Int_Int_t lizzieLet12_6QNone_Int_6QNode_Int_bufchan_buf;
  assign lizzieLet12_6QNone_Int_6QNode_Int_bufchan_r = (! lizzieLet12_6QNone_Int_6QNode_Int_bufchan_buf[0]);
  assign lizzieLet12_6QNone_Int_6QNode_Int_1_argbuf_d = (lizzieLet12_6QNone_Int_6QNode_Int_bufchan_buf[0] ? lizzieLet12_6QNone_Int_6QNode_Int_bufchan_buf :
                                                         lizzieLet12_6QNone_Int_6QNode_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNone_Int_6QNode_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet12_6QNone_Int_6QNode_Int_1_argbuf_r && lizzieLet12_6QNone_Int_6QNode_Int_bufchan_buf[0]))
        lizzieLet12_6QNone_Int_6QNode_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet12_6QNone_Int_6QNode_Int_1_argbuf_r) && (! lizzieLet12_6QNone_Int_6QNode_Int_bufchan_buf[0])))
        lizzieLet12_6QNone_Int_6QNode_Int_bufchan_buf <= lizzieLet12_6QNone_Int_6QNode_Int_bufchan_d;
  
  /* buf (Ty Pointer_CTf_f_Int_Int) : (lizzieLet12_6QNone_Int_6QNone_Int,Pointer_CTf_f_Int_Int) > (lizzieLet12_6QNone_Int_6QNone_Int_1_argbuf,Pointer_CTf_f_Int_Int) */
  Pointer_CTf_f_Int_Int_t lizzieLet12_6QNone_Int_6QNone_Int_bufchan_d;
  logic lizzieLet12_6QNone_Int_6QNone_Int_bufchan_r;
  assign lizzieLet12_6QNone_Int_6QNone_Int_r = ((! lizzieLet12_6QNone_Int_6QNone_Int_bufchan_d[0]) || lizzieLet12_6QNone_Int_6QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNone_Int_6QNone_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet12_6QNone_Int_6QNone_Int_r)
        lizzieLet12_6QNone_Int_6QNone_Int_bufchan_d <= lizzieLet12_6QNone_Int_6QNone_Int_d;
  Pointer_CTf_f_Int_Int_t lizzieLet12_6QNone_Int_6QNone_Int_bufchan_buf;
  assign lizzieLet12_6QNone_Int_6QNone_Int_bufchan_r = (! lizzieLet12_6QNone_Int_6QNone_Int_bufchan_buf[0]);
  assign lizzieLet12_6QNone_Int_6QNone_Int_1_argbuf_d = (lizzieLet12_6QNone_Int_6QNone_Int_bufchan_buf[0] ? lizzieLet12_6QNone_Int_6QNone_Int_bufchan_buf :
                                                         lizzieLet12_6QNone_Int_6QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QNone_Int_6QNone_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet12_6QNone_Int_6QNone_Int_1_argbuf_r && lizzieLet12_6QNone_Int_6QNone_Int_bufchan_buf[0]))
        lizzieLet12_6QNone_Int_6QNone_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet12_6QNone_Int_6QNone_Int_1_argbuf_r) && (! lizzieLet12_6QNone_Int_6QNone_Int_bufchan_buf[0])))
        lizzieLet12_6QNone_Int_6QNone_Int_bufchan_buf <= lizzieLet12_6QNone_Int_6QNone_Int_bufchan_d;
  
  /* fork (Ty QTree_Int) : (lizzieLet12_6QVal_Int,QTree_Int) > [(lizzieLet12_6QVal_Int_1,QTree_Int),
                                                           (lizzieLet12_6QVal_Int_2,QTree_Int),
                                                           (lizzieLet12_6QVal_Int_3,QTree_Int),
                                                           (lizzieLet12_6QVal_Int_4,QTree_Int),
                                                           (lizzieLet12_6QVal_Int_5,QTree_Int),
                                                           (lizzieLet12_6QVal_Int_6,QTree_Int),
                                                           (lizzieLet12_6QVal_Int_7,QTree_Int),
                                                           (lizzieLet12_6QVal_Int_8,QTree_Int),
                                                           (lizzieLet12_6QVal_Int_9,QTree_Int)] */
  logic [8:0] lizzieLet12_6QVal_Int_emitted;
  logic [8:0] lizzieLet12_6QVal_Int_done;
  assign lizzieLet12_6QVal_Int_1_d = {lizzieLet12_6QVal_Int_d[66:1],
                                      (lizzieLet12_6QVal_Int_d[0] && (! lizzieLet12_6QVal_Int_emitted[0]))};
  assign lizzieLet12_6QVal_Int_2_d = {lizzieLet12_6QVal_Int_d[66:1],
                                      (lizzieLet12_6QVal_Int_d[0] && (! lizzieLet12_6QVal_Int_emitted[1]))};
  assign lizzieLet12_6QVal_Int_3_d = {lizzieLet12_6QVal_Int_d[66:1],
                                      (lizzieLet12_6QVal_Int_d[0] && (! lizzieLet12_6QVal_Int_emitted[2]))};
  assign lizzieLet12_6QVal_Int_4_d = {lizzieLet12_6QVal_Int_d[66:1],
                                      (lizzieLet12_6QVal_Int_d[0] && (! lizzieLet12_6QVal_Int_emitted[3]))};
  assign lizzieLet12_6QVal_Int_5_d = {lizzieLet12_6QVal_Int_d[66:1],
                                      (lizzieLet12_6QVal_Int_d[0] && (! lizzieLet12_6QVal_Int_emitted[4]))};
  assign lizzieLet12_6QVal_Int_6_d = {lizzieLet12_6QVal_Int_d[66:1],
                                      (lizzieLet12_6QVal_Int_d[0] && (! lizzieLet12_6QVal_Int_emitted[5]))};
  assign lizzieLet12_6QVal_Int_7_d = {lizzieLet12_6QVal_Int_d[66:1],
                                      (lizzieLet12_6QVal_Int_d[0] && (! lizzieLet12_6QVal_Int_emitted[6]))};
  assign lizzieLet12_6QVal_Int_8_d = {lizzieLet12_6QVal_Int_d[66:1],
                                      (lizzieLet12_6QVal_Int_d[0] && (! lizzieLet12_6QVal_Int_emitted[7]))};
  assign lizzieLet12_6QVal_Int_9_d = {lizzieLet12_6QVal_Int_d[66:1],
                                      (lizzieLet12_6QVal_Int_d[0] && (! lizzieLet12_6QVal_Int_emitted[8]))};
  assign lizzieLet12_6QVal_Int_done = (lizzieLet12_6QVal_Int_emitted | ({lizzieLet12_6QVal_Int_9_d[0],
                                                                         lizzieLet12_6QVal_Int_8_d[0],
                                                                         lizzieLet12_6QVal_Int_7_d[0],
                                                                         lizzieLet12_6QVal_Int_6_d[0],
                                                                         lizzieLet12_6QVal_Int_5_d[0],
                                                                         lizzieLet12_6QVal_Int_4_d[0],
                                                                         lizzieLet12_6QVal_Int_3_d[0],
                                                                         lizzieLet12_6QVal_Int_2_d[0],
                                                                         lizzieLet12_6QVal_Int_1_d[0]} & {lizzieLet12_6QVal_Int_9_r,
                                                                                                          lizzieLet12_6QVal_Int_8_r,
                                                                                                          lizzieLet12_6QVal_Int_7_r,
                                                                                                          lizzieLet12_6QVal_Int_6_r,
                                                                                                          lizzieLet12_6QVal_Int_5_r,
                                                                                                          lizzieLet12_6QVal_Int_4_r,
                                                                                                          lizzieLet12_6QVal_Int_3_r,
                                                                                                          lizzieLet12_6QVal_Int_2_r,
                                                                                                          lizzieLet12_6QVal_Int_1_r}));
  assign lizzieLet12_6QVal_Int_r = (& lizzieLet12_6QVal_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet12_6QVal_Int_emitted <= 9'd0;
    else
      lizzieLet12_6QVal_Int_emitted <= (lizzieLet12_6QVal_Int_r ? 9'd0 :
                                        lizzieLet12_6QVal_Int_done);
  
  /* destruct (Ty QTree_Int,
          Dcon QVal_Int) : (lizzieLet12_6QVal_Int_1QVal_Int,QTree_Int) > [(va8O_destruct,Int)] */
  assign va8O_destruct_d = {lizzieLet12_6QVal_Int_1QVal_Int_d[34:3],
                            lizzieLet12_6QVal_Int_1QVal_Int_d[0]};
  assign lizzieLet12_6QVal_Int_1QVal_Int_r = va8O_destruct_r;
  
  /* demux (Ty QTree_Int,
       Ty QTree_Int) : (lizzieLet12_6QVal_Int_2,QTree_Int) (lizzieLet12_6QVal_Int_1,QTree_Int) > [(_32,QTree_Int),
                                                                                                  (lizzieLet12_6QVal_Int_1QVal_Int,QTree_Int),
                                                                                                  (_31,QTree_Int),
                                                                                                  (_30,QTree_Int)] */
  logic [3:0] lizzieLet12_6QVal_Int_1_onehotd;
  always_comb
    if ((lizzieLet12_6QVal_Int_2_d[0] && lizzieLet12_6QVal_Int_1_d[0]))
      unique case (lizzieLet12_6QVal_Int_2_d[2:1])
        2'd0: lizzieLet12_6QVal_Int_1_onehotd = 4'd1;
        2'd1: lizzieLet12_6QVal_Int_1_onehotd = 4'd2;
        2'd2: lizzieLet12_6QVal_Int_1_onehotd = 4'd4;
        2'd3: lizzieLet12_6QVal_Int_1_onehotd = 4'd8;
        default: lizzieLet12_6QVal_Int_1_onehotd = 4'd0;
      endcase
    else lizzieLet12_6QVal_Int_1_onehotd = 4'd0;
  assign _32_d = {lizzieLet12_6QVal_Int_1_d[66:1],
                  lizzieLet12_6QVal_Int_1_onehotd[0]};
  assign lizzieLet12_6QVal_Int_1QVal_Int_d = {lizzieLet12_6QVal_Int_1_d[66:1],
                                              lizzieLet12_6QVal_Int_1_onehotd[1]};
  assign _31_d = {lizzieLet12_6QVal_Int_1_d[66:1],
                  lizzieLet12_6QVal_Int_1_onehotd[2]};
  assign _30_d = {lizzieLet12_6QVal_Int_1_d[66:1],
                  lizzieLet12_6QVal_Int_1_onehotd[3]};
  assign lizzieLet12_6QVal_Int_1_r = (| (lizzieLet12_6QVal_Int_1_onehotd & {_30_r,
                                                                            _31_r,
                                                                            lizzieLet12_6QVal_Int_1QVal_Int_r,
                                                                            _32_r}));
  assign lizzieLet12_6QVal_Int_2_r = lizzieLet12_6QVal_Int_1_r;
  
  /* demux (Ty QTree_Int,
       Ty Go) : (lizzieLet12_6QVal_Int_3,QTree_Int) (lizzieLet12_3QVal_Int,Go) > [(lizzieLet12_6QVal_Int_3QNone_Int,Go),
                                                                                  (lizzieLet12_6QVal_Int_3QVal_Int,Go),
                                                                                  (lizzieLet12_6QVal_Int_3QNode_Int,Go),
                                                                                  (lizzieLet12_6QVal_Int_3QError_Int,Go)] */
  logic [3:0] lizzieLet12_3QVal_Int_onehotd;
  always_comb
    if ((lizzieLet12_6QVal_Int_3_d[0] && lizzieLet12_3QVal_Int_d[0]))
      unique case (lizzieLet12_6QVal_Int_3_d[2:1])
        2'd0: lizzieLet12_3QVal_Int_onehotd = 4'd1;
        2'd1: lizzieLet12_3QVal_Int_onehotd = 4'd2;
        2'd2: lizzieLet12_3QVal_Int_onehotd = 4'd4;
        2'd3: lizzieLet12_3QVal_Int_onehotd = 4'd8;
        default: lizzieLet12_3QVal_Int_onehotd = 4'd0;
      endcase
    else lizzieLet12_3QVal_Int_onehotd = 4'd0;
  assign lizzieLet12_6QVal_Int_3QNone_Int_d = lizzieLet12_3QVal_Int_onehotd[0];
  assign lizzieLet12_6QVal_Int_3QVal_Int_d = lizzieLet12_3QVal_Int_onehotd[1];
  assign lizzieLet12_6QVal_Int_3QNode_Int_d = lizzieLet12_3QVal_Int_onehotd[2];
  assign lizzieLet12_6QVal_Int_3QError_Int_d = lizzieLet12_3QVal_Int_onehotd[3];
  assign lizzieLet12_3QVal_Int_r = (| (lizzieLet12_3QVal_Int_onehotd & {lizzieLet12_6QVal_Int_3QError_Int_r,
                                                                        lizzieLet12_6QVal_Int_3QNode_Int_r,
                                                                        lizzieLet12_6QVal_Int_3QVal_Int_r,
                                                                        lizzieLet12_6QVal_Int_3QNone_Int_r}));
  assign lizzieLet12_6QVal_Int_3_r = lizzieLet12_3QVal_Int_r;
  
  /* fork (Ty Go) : (lizzieLet12_6QVal_Int_3QError_Int,Go) > [(lizzieLet12_6QVal_Int_3QError_Int_1,Go),
                                                         (lizzieLet12_6QVal_Int_3QError_Int_2,Go)] */
  logic [1:0] lizzieLet12_6QVal_Int_3QError_Int_emitted;
  logic [1:0] lizzieLet12_6QVal_Int_3QError_Int_done;
  assign lizzieLet12_6QVal_Int_3QError_Int_1_d = (lizzieLet12_6QVal_Int_3QError_Int_d[0] && (! lizzieLet12_6QVal_Int_3QError_Int_emitted[0]));
  assign lizzieLet12_6QVal_Int_3QError_Int_2_d = (lizzieLet12_6QVal_Int_3QError_Int_d[0] && (! lizzieLet12_6QVal_Int_3QError_Int_emitted[1]));
  assign lizzieLet12_6QVal_Int_3QError_Int_done = (lizzieLet12_6QVal_Int_3QError_Int_emitted | ({lizzieLet12_6QVal_Int_3QError_Int_2_d[0],
                                                                                                 lizzieLet12_6QVal_Int_3QError_Int_1_d[0]} & {lizzieLet12_6QVal_Int_3QError_Int_2_r,
                                                                                                                                              lizzieLet12_6QVal_Int_3QError_Int_1_r}));
  assign lizzieLet12_6QVal_Int_3QError_Int_r = (& lizzieLet12_6QVal_Int_3QError_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QVal_Int_3QError_Int_emitted <= 2'd0;
    else
      lizzieLet12_6QVal_Int_3QError_Int_emitted <= (lizzieLet12_6QVal_Int_3QError_Int_r ? 2'd0 :
                                                    lizzieLet12_6QVal_Int_3QError_Int_done);
  
  /* dcon (Ty QTree_Int,
      Dcon QError_Int) : [(lizzieLet12_6QVal_Int_3QError_Int_1,Go)] > (lizzieLet12_6QVal_Int_3QError_Int_1QError_Int,QTree_Int) */
  assign lizzieLet12_6QVal_Int_3QError_Int_1QError_Int_d = QError_Int_dc((& {lizzieLet12_6QVal_Int_3QError_Int_1_d[0]}), lizzieLet12_6QVal_Int_3QError_Int_1_d);
  assign {lizzieLet12_6QVal_Int_3QError_Int_1_r} = {1 {(lizzieLet12_6QVal_Int_3QError_Int_1QError_Int_r && lizzieLet12_6QVal_Int_3QError_Int_1QError_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (lizzieLet12_6QVal_Int_3QError_Int_1QError_Int,QTree_Int) > (lizzieLet26_1_argbuf,QTree_Int) */
  QTree_Int_t lizzieLet12_6QVal_Int_3QError_Int_1QError_Int_bufchan_d;
  logic lizzieLet12_6QVal_Int_3QError_Int_1QError_Int_bufchan_r;
  assign lizzieLet12_6QVal_Int_3QError_Int_1QError_Int_r = ((! lizzieLet12_6QVal_Int_3QError_Int_1QError_Int_bufchan_d[0]) || lizzieLet12_6QVal_Int_3QError_Int_1QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QVal_Int_3QError_Int_1QError_Int_bufchan_d <= {66'd0,
                                                                  1'd0};
    else
      if (lizzieLet12_6QVal_Int_3QError_Int_1QError_Int_r)
        lizzieLet12_6QVal_Int_3QError_Int_1QError_Int_bufchan_d <= lizzieLet12_6QVal_Int_3QError_Int_1QError_Int_d;
  QTree_Int_t lizzieLet12_6QVal_Int_3QError_Int_1QError_Int_bufchan_buf;
  assign lizzieLet12_6QVal_Int_3QError_Int_1QError_Int_bufchan_r = (! lizzieLet12_6QVal_Int_3QError_Int_1QError_Int_bufchan_buf[0]);
  assign lizzieLet26_1_argbuf_d = (lizzieLet12_6QVal_Int_3QError_Int_1QError_Int_bufchan_buf[0] ? lizzieLet12_6QVal_Int_3QError_Int_1QError_Int_bufchan_buf :
                                   lizzieLet12_6QVal_Int_3QError_Int_1QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QVal_Int_3QError_Int_1QError_Int_bufchan_buf <= {66'd0,
                                                                    1'd0};
    else
      if ((lizzieLet26_1_argbuf_r && lizzieLet12_6QVal_Int_3QError_Int_1QError_Int_bufchan_buf[0]))
        lizzieLet12_6QVal_Int_3QError_Int_1QError_Int_bufchan_buf <= {66'd0,
                                                                      1'd0};
      else if (((! lizzieLet26_1_argbuf_r) && (! lizzieLet12_6QVal_Int_3QError_Int_1QError_Int_bufchan_buf[0])))
        lizzieLet12_6QVal_Int_3QError_Int_1QError_Int_bufchan_buf <= lizzieLet12_6QVal_Int_3QError_Int_1QError_Int_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet12_6QVal_Int_3QError_Int_2,Go) > (lizzieLet12_6QVal_Int_3QError_Int_2_argbuf,Go) */
  Go_t lizzieLet12_6QVal_Int_3QError_Int_2_bufchan_d;
  logic lizzieLet12_6QVal_Int_3QError_Int_2_bufchan_r;
  assign lizzieLet12_6QVal_Int_3QError_Int_2_r = ((! lizzieLet12_6QVal_Int_3QError_Int_2_bufchan_d[0]) || lizzieLet12_6QVal_Int_3QError_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QVal_Int_3QError_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet12_6QVal_Int_3QError_Int_2_r)
        lizzieLet12_6QVal_Int_3QError_Int_2_bufchan_d <= lizzieLet12_6QVal_Int_3QError_Int_2_d;
  Go_t lizzieLet12_6QVal_Int_3QError_Int_2_bufchan_buf;
  assign lizzieLet12_6QVal_Int_3QError_Int_2_bufchan_r = (! lizzieLet12_6QVal_Int_3QError_Int_2_bufchan_buf[0]);
  assign lizzieLet12_6QVal_Int_3QError_Int_2_argbuf_d = (lizzieLet12_6QVal_Int_3QError_Int_2_bufchan_buf[0] ? lizzieLet12_6QVal_Int_3QError_Int_2_bufchan_buf :
                                                         lizzieLet12_6QVal_Int_3QError_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QVal_Int_3QError_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet12_6QVal_Int_3QError_Int_2_argbuf_r && lizzieLet12_6QVal_Int_3QError_Int_2_bufchan_buf[0]))
        lizzieLet12_6QVal_Int_3QError_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet12_6QVal_Int_3QError_Int_2_argbuf_r) && (! lizzieLet12_6QVal_Int_3QError_Int_2_bufchan_buf[0])))
        lizzieLet12_6QVal_Int_3QError_Int_2_bufchan_buf <= lizzieLet12_6QVal_Int_3QError_Int_2_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet12_6QVal_Int_3QNode_Int,Go) > [(lizzieLet12_6QVal_Int_3QNode_Int_1,Go),
                                                        (lizzieLet12_6QVal_Int_3QNode_Int_2,Go)] */
  logic [1:0] lizzieLet12_6QVal_Int_3QNode_Int_emitted;
  logic [1:0] lizzieLet12_6QVal_Int_3QNode_Int_done;
  assign lizzieLet12_6QVal_Int_3QNode_Int_1_d = (lizzieLet12_6QVal_Int_3QNode_Int_d[0] && (! lizzieLet12_6QVal_Int_3QNode_Int_emitted[0]));
  assign lizzieLet12_6QVal_Int_3QNode_Int_2_d = (lizzieLet12_6QVal_Int_3QNode_Int_d[0] && (! lizzieLet12_6QVal_Int_3QNode_Int_emitted[1]));
  assign lizzieLet12_6QVal_Int_3QNode_Int_done = (lizzieLet12_6QVal_Int_3QNode_Int_emitted | ({lizzieLet12_6QVal_Int_3QNode_Int_2_d[0],
                                                                                               lizzieLet12_6QVal_Int_3QNode_Int_1_d[0]} & {lizzieLet12_6QVal_Int_3QNode_Int_2_r,
                                                                                                                                           lizzieLet12_6QVal_Int_3QNode_Int_1_r}));
  assign lizzieLet12_6QVal_Int_3QNode_Int_r = (& lizzieLet12_6QVal_Int_3QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QVal_Int_3QNode_Int_emitted <= 2'd0;
    else
      lizzieLet12_6QVal_Int_3QNode_Int_emitted <= (lizzieLet12_6QVal_Int_3QNode_Int_r ? 2'd0 :
                                                   lizzieLet12_6QVal_Int_3QNode_Int_done);
  
  /* dcon (Ty QTree_Int,
      Dcon QError_Int) : [(lizzieLet12_6QVal_Int_3QNode_Int_1,Go)] > (lizzieLet12_6QVal_Int_3QNode_Int_1QError_Int,QTree_Int) */
  assign lizzieLet12_6QVal_Int_3QNode_Int_1QError_Int_d = QError_Int_dc((& {lizzieLet12_6QVal_Int_3QNode_Int_1_d[0]}), lizzieLet12_6QVal_Int_3QNode_Int_1_d);
  assign {lizzieLet12_6QVal_Int_3QNode_Int_1_r} = {1 {(lizzieLet12_6QVal_Int_3QNode_Int_1QError_Int_r && lizzieLet12_6QVal_Int_3QNode_Int_1QError_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (lizzieLet12_6QVal_Int_3QNode_Int_1QError_Int,QTree_Int) > (lizzieLet25_1_1_argbuf,QTree_Int) */
  QTree_Int_t lizzieLet12_6QVal_Int_3QNode_Int_1QError_Int_bufchan_d;
  logic lizzieLet12_6QVal_Int_3QNode_Int_1QError_Int_bufchan_r;
  assign lizzieLet12_6QVal_Int_3QNode_Int_1QError_Int_r = ((! lizzieLet12_6QVal_Int_3QNode_Int_1QError_Int_bufchan_d[0]) || lizzieLet12_6QVal_Int_3QNode_Int_1QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QVal_Int_3QNode_Int_1QError_Int_bufchan_d <= {66'd0,
                                                                 1'd0};
    else
      if (lizzieLet12_6QVal_Int_3QNode_Int_1QError_Int_r)
        lizzieLet12_6QVal_Int_3QNode_Int_1QError_Int_bufchan_d <= lizzieLet12_6QVal_Int_3QNode_Int_1QError_Int_d;
  QTree_Int_t lizzieLet12_6QVal_Int_3QNode_Int_1QError_Int_bufchan_buf;
  assign lizzieLet12_6QVal_Int_3QNode_Int_1QError_Int_bufchan_r = (! lizzieLet12_6QVal_Int_3QNode_Int_1QError_Int_bufchan_buf[0]);
  assign lizzieLet25_1_1_argbuf_d = (lizzieLet12_6QVal_Int_3QNode_Int_1QError_Int_bufchan_buf[0] ? lizzieLet12_6QVal_Int_3QNode_Int_1QError_Int_bufchan_buf :
                                     lizzieLet12_6QVal_Int_3QNode_Int_1QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QVal_Int_3QNode_Int_1QError_Int_bufchan_buf <= {66'd0,
                                                                   1'd0};
    else
      if ((lizzieLet25_1_1_argbuf_r && lizzieLet12_6QVal_Int_3QNode_Int_1QError_Int_bufchan_buf[0]))
        lizzieLet12_6QVal_Int_3QNode_Int_1QError_Int_bufchan_buf <= {66'd0,
                                                                     1'd0};
      else if (((! lizzieLet25_1_1_argbuf_r) && (! lizzieLet12_6QVal_Int_3QNode_Int_1QError_Int_bufchan_buf[0])))
        lizzieLet12_6QVal_Int_3QNode_Int_1QError_Int_bufchan_buf <= lizzieLet12_6QVal_Int_3QNode_Int_1QError_Int_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet12_6QVal_Int_3QNode_Int_2,Go) > (lizzieLet12_6QVal_Int_3QNode_Int_2_argbuf,Go) */
  Go_t lizzieLet12_6QVal_Int_3QNode_Int_2_bufchan_d;
  logic lizzieLet12_6QVal_Int_3QNode_Int_2_bufchan_r;
  assign lizzieLet12_6QVal_Int_3QNode_Int_2_r = ((! lizzieLet12_6QVal_Int_3QNode_Int_2_bufchan_d[0]) || lizzieLet12_6QVal_Int_3QNode_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QVal_Int_3QNode_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet12_6QVal_Int_3QNode_Int_2_r)
        lizzieLet12_6QVal_Int_3QNode_Int_2_bufchan_d <= lizzieLet12_6QVal_Int_3QNode_Int_2_d;
  Go_t lizzieLet12_6QVal_Int_3QNode_Int_2_bufchan_buf;
  assign lizzieLet12_6QVal_Int_3QNode_Int_2_bufchan_r = (! lizzieLet12_6QVal_Int_3QNode_Int_2_bufchan_buf[0]);
  assign lizzieLet12_6QVal_Int_3QNode_Int_2_argbuf_d = (lizzieLet12_6QVal_Int_3QNode_Int_2_bufchan_buf[0] ? lizzieLet12_6QVal_Int_3QNode_Int_2_bufchan_buf :
                                                        lizzieLet12_6QVal_Int_3QNode_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QVal_Int_3QNode_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet12_6QVal_Int_3QNode_Int_2_argbuf_r && lizzieLet12_6QVal_Int_3QNode_Int_2_bufchan_buf[0]))
        lizzieLet12_6QVal_Int_3QNode_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet12_6QVal_Int_3QNode_Int_2_argbuf_r) && (! lizzieLet12_6QVal_Int_3QNode_Int_2_bufchan_buf[0])))
        lizzieLet12_6QVal_Int_3QNode_Int_2_bufchan_buf <= lizzieLet12_6QVal_Int_3QNode_Int_2_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet12_6QVal_Int_3QNone_Int,Go) > [(lizzieLet12_6QVal_Int_3QNone_Int_1,Go),
                                                        (lizzieLet12_6QVal_Int_3QNone_Int_2,Go),
                                                        (lizzieLet12_6QVal_Int_3QNone_Int_3,Go)] */
  logic [2:0] lizzieLet12_6QVal_Int_3QNone_Int_emitted;
  logic [2:0] lizzieLet12_6QVal_Int_3QNone_Int_done;
  assign lizzieLet12_6QVal_Int_3QNone_Int_1_d = (lizzieLet12_6QVal_Int_3QNone_Int_d[0] && (! lizzieLet12_6QVal_Int_3QNone_Int_emitted[0]));
  assign lizzieLet12_6QVal_Int_3QNone_Int_2_d = (lizzieLet12_6QVal_Int_3QNone_Int_d[0] && (! lizzieLet12_6QVal_Int_3QNone_Int_emitted[1]));
  assign lizzieLet12_6QVal_Int_3QNone_Int_3_d = (lizzieLet12_6QVal_Int_3QNone_Int_d[0] && (! lizzieLet12_6QVal_Int_3QNone_Int_emitted[2]));
  assign lizzieLet12_6QVal_Int_3QNone_Int_done = (lizzieLet12_6QVal_Int_3QNone_Int_emitted | ({lizzieLet12_6QVal_Int_3QNone_Int_3_d[0],
                                                                                               lizzieLet12_6QVal_Int_3QNone_Int_2_d[0],
                                                                                               lizzieLet12_6QVal_Int_3QNone_Int_1_d[0]} & {lizzieLet12_6QVal_Int_3QNone_Int_3_r,
                                                                                                                                           lizzieLet12_6QVal_Int_3QNone_Int_2_r,
                                                                                                                                           lizzieLet12_6QVal_Int_3QNone_Int_1_r}));
  assign lizzieLet12_6QVal_Int_3QNone_Int_r = (& lizzieLet12_6QVal_Int_3QNone_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QVal_Int_3QNone_Int_emitted <= 3'd0;
    else
      lizzieLet12_6QVal_Int_3QNone_Int_emitted <= (lizzieLet12_6QVal_Int_3QNone_Int_r ? 3'd0 :
                                                   lizzieLet12_6QVal_Int_3QNone_Int_done);
  
  /* buf (Ty Go) : (lizzieLet12_6QVal_Int_3QNone_Int_1,Go) > (lizzieLet12_6QVal_Int_3QNone_Int_1_argbuf,Go) */
  Go_t lizzieLet12_6QVal_Int_3QNone_Int_1_bufchan_d;
  logic lizzieLet12_6QVal_Int_3QNone_Int_1_bufchan_r;
  assign lizzieLet12_6QVal_Int_3QNone_Int_1_r = ((! lizzieLet12_6QVal_Int_3QNone_Int_1_bufchan_d[0]) || lizzieLet12_6QVal_Int_3QNone_Int_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QVal_Int_3QNone_Int_1_bufchan_d <= 1'd0;
    else
      if (lizzieLet12_6QVal_Int_3QNone_Int_1_r)
        lizzieLet12_6QVal_Int_3QNone_Int_1_bufchan_d <= lizzieLet12_6QVal_Int_3QNone_Int_1_d;
  Go_t lizzieLet12_6QVal_Int_3QNone_Int_1_bufchan_buf;
  assign lizzieLet12_6QVal_Int_3QNone_Int_1_bufchan_r = (! lizzieLet12_6QVal_Int_3QNone_Int_1_bufchan_buf[0]);
  assign lizzieLet12_6QVal_Int_3QNone_Int_1_argbuf_d = (lizzieLet12_6QVal_Int_3QNone_Int_1_bufchan_buf[0] ? lizzieLet12_6QVal_Int_3QNone_Int_1_bufchan_buf :
                                                        lizzieLet12_6QVal_Int_3QNone_Int_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QVal_Int_3QNone_Int_1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet12_6QVal_Int_3QNone_Int_1_argbuf_r && lizzieLet12_6QVal_Int_3QNone_Int_1_bufchan_buf[0]))
        lizzieLet12_6QVal_Int_3QNone_Int_1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet12_6QVal_Int_3QNone_Int_1_argbuf_r) && (! lizzieLet12_6QVal_Int_3QNone_Int_1_bufchan_buf[0])))
        lizzieLet12_6QVal_Int_3QNone_Int_1_bufchan_buf <= lizzieLet12_6QVal_Int_3QNone_Int_1_bufchan_d;
  
  /* dcon (Ty TupGo___MyDTInt_Int___Int,
      Dcon TupGo___MyDTInt_Int___Int) : [(lizzieLet12_6QVal_Int_3QNone_Int_1_argbuf,Go),
                                         (lizzieLet12_6QVal_Int_7QNone_Int_1_argbuf,MyDTInt_Int),
                                         (lizzieLet12_6QVal_Int_9QNone_Int_1_argbuf,Int)] > (applyfnInt_Int_5TupGo___MyDTInt_Int___Int5,TupGo___MyDTInt_Int___Int) */
  assign applyfnInt_Int_5TupGo___MyDTInt_Int___Int5_d = TupGo___MyDTInt_Int___Int_dc((& {lizzieLet12_6QVal_Int_3QNone_Int_1_argbuf_d[0],
                                                                                         lizzieLet12_6QVal_Int_7QNone_Int_1_argbuf_d[0],
                                                                                         lizzieLet12_6QVal_Int_9QNone_Int_1_argbuf_d[0]}), lizzieLet12_6QVal_Int_3QNone_Int_1_argbuf_d, lizzieLet12_6QVal_Int_7QNone_Int_1_argbuf_d, lizzieLet12_6QVal_Int_9QNone_Int_1_argbuf_d);
  assign {lizzieLet12_6QVal_Int_3QNone_Int_1_argbuf_r,
          lizzieLet12_6QVal_Int_7QNone_Int_1_argbuf_r,
          lizzieLet12_6QVal_Int_9QNone_Int_1_argbuf_r} = {3 {(applyfnInt_Int_5TupGo___MyDTInt_Int___Int5_r && applyfnInt_Int_5TupGo___MyDTInt_Int___Int5_d[0])}};
  
  /* buf (Ty Go) : (lizzieLet12_6QVal_Int_3QNone_Int_2,Go) > (lizzieLet12_6QVal_Int_3QNone_Int_2_argbuf,Go) */
  Go_t lizzieLet12_6QVal_Int_3QNone_Int_2_bufchan_d;
  logic lizzieLet12_6QVal_Int_3QNone_Int_2_bufchan_r;
  assign lizzieLet12_6QVal_Int_3QNone_Int_2_r = ((! lizzieLet12_6QVal_Int_3QNone_Int_2_bufchan_d[0]) || lizzieLet12_6QVal_Int_3QNone_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QVal_Int_3QNone_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet12_6QVal_Int_3QNone_Int_2_r)
        lizzieLet12_6QVal_Int_3QNone_Int_2_bufchan_d <= lizzieLet12_6QVal_Int_3QNone_Int_2_d;
  Go_t lizzieLet12_6QVal_Int_3QNone_Int_2_bufchan_buf;
  assign lizzieLet12_6QVal_Int_3QNone_Int_2_bufchan_r = (! lizzieLet12_6QVal_Int_3QNone_Int_2_bufchan_buf[0]);
  assign lizzieLet12_6QVal_Int_3QNone_Int_2_argbuf_d = (lizzieLet12_6QVal_Int_3QNone_Int_2_bufchan_buf[0] ? lizzieLet12_6QVal_Int_3QNone_Int_2_bufchan_buf :
                                                        lizzieLet12_6QVal_Int_3QNone_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QVal_Int_3QNone_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet12_6QVal_Int_3QNone_Int_2_argbuf_r && lizzieLet12_6QVal_Int_3QNone_Int_2_bufchan_buf[0]))
        lizzieLet12_6QVal_Int_3QNone_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet12_6QVal_Int_3QNone_Int_2_argbuf_r) && (! lizzieLet12_6QVal_Int_3QNone_Int_2_bufchan_buf[0])))
        lizzieLet12_6QVal_Int_3QNone_Int_2_bufchan_buf <= lizzieLet12_6QVal_Int_3QNone_Int_2_bufchan_d;
  
  /* dcon (Ty TupGo___MyDTInt_Bool___Int,
      Dcon TupGo___MyDTInt_Bool___Int) : [(lizzieLet12_6QVal_Int_3QNone_Int_2_argbuf,Go),
                                          (lizzieLet12_6QVal_Int_5QNone_Int_1_argbuf,MyDTInt_Bool),
                                          (es_9_1_argbuf,Int)] > (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int3,TupGo___MyDTInt_Bool___Int) */
  assign applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int3_d = TupGo___MyDTInt_Bool___Int_dc((& {lizzieLet12_6QVal_Int_3QNone_Int_2_argbuf_d[0],
                                                                                            lizzieLet12_6QVal_Int_5QNone_Int_1_argbuf_d[0],
                                                                                            es_9_1_argbuf_d[0]}), lizzieLet12_6QVal_Int_3QNone_Int_2_argbuf_d, lizzieLet12_6QVal_Int_5QNone_Int_1_argbuf_d, es_9_1_argbuf_d);
  assign {lizzieLet12_6QVal_Int_3QNone_Int_2_argbuf_r,
          lizzieLet12_6QVal_Int_5QNone_Int_1_argbuf_r,
          es_9_1_argbuf_r} = {3 {(applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int3_r && applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int3_d[0])}};
  
  /* fork (Ty Go) : (lizzieLet12_6QVal_Int_3QVal_Int,Go) > [(lizzieLet12_6QVal_Int_3QVal_Int_1,Go),
                                                       (lizzieLet12_6QVal_Int_3QVal_Int_2,Go)] */
  logic [1:0] lizzieLet12_6QVal_Int_3QVal_Int_emitted;
  logic [1:0] lizzieLet12_6QVal_Int_3QVal_Int_done;
  assign lizzieLet12_6QVal_Int_3QVal_Int_1_d = (lizzieLet12_6QVal_Int_3QVal_Int_d[0] && (! lizzieLet12_6QVal_Int_3QVal_Int_emitted[0]));
  assign lizzieLet12_6QVal_Int_3QVal_Int_2_d = (lizzieLet12_6QVal_Int_3QVal_Int_d[0] && (! lizzieLet12_6QVal_Int_3QVal_Int_emitted[1]));
  assign lizzieLet12_6QVal_Int_3QVal_Int_done = (lizzieLet12_6QVal_Int_3QVal_Int_emitted | ({lizzieLet12_6QVal_Int_3QVal_Int_2_d[0],
                                                                                             lizzieLet12_6QVal_Int_3QVal_Int_1_d[0]} & {lizzieLet12_6QVal_Int_3QVal_Int_2_r,
                                                                                                                                        lizzieLet12_6QVal_Int_3QVal_Int_1_r}));
  assign lizzieLet12_6QVal_Int_3QVal_Int_r = (& lizzieLet12_6QVal_Int_3QVal_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QVal_Int_3QVal_Int_emitted <= 2'd0;
    else
      lizzieLet12_6QVal_Int_3QVal_Int_emitted <= (lizzieLet12_6QVal_Int_3QVal_Int_r ? 2'd0 :
                                                  lizzieLet12_6QVal_Int_3QVal_Int_done);
  
  /* buf (Ty Go) : (lizzieLet12_6QVal_Int_3QVal_Int_1,Go) > (lizzieLet12_6QVal_Int_3QVal_Int_1_argbuf,Go) */
  Go_t lizzieLet12_6QVal_Int_3QVal_Int_1_bufchan_d;
  logic lizzieLet12_6QVal_Int_3QVal_Int_1_bufchan_r;
  assign lizzieLet12_6QVal_Int_3QVal_Int_1_r = ((! lizzieLet12_6QVal_Int_3QVal_Int_1_bufchan_d[0]) || lizzieLet12_6QVal_Int_3QVal_Int_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QVal_Int_3QVal_Int_1_bufchan_d <= 1'd0;
    else
      if (lizzieLet12_6QVal_Int_3QVal_Int_1_r)
        lizzieLet12_6QVal_Int_3QVal_Int_1_bufchan_d <= lizzieLet12_6QVal_Int_3QVal_Int_1_d;
  Go_t lizzieLet12_6QVal_Int_3QVal_Int_1_bufchan_buf;
  assign lizzieLet12_6QVal_Int_3QVal_Int_1_bufchan_r = (! lizzieLet12_6QVal_Int_3QVal_Int_1_bufchan_buf[0]);
  assign lizzieLet12_6QVal_Int_3QVal_Int_1_argbuf_d = (lizzieLet12_6QVal_Int_3QVal_Int_1_bufchan_buf[0] ? lizzieLet12_6QVal_Int_3QVal_Int_1_bufchan_buf :
                                                       lizzieLet12_6QVal_Int_3QVal_Int_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QVal_Int_3QVal_Int_1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet12_6QVal_Int_3QVal_Int_1_argbuf_r && lizzieLet12_6QVal_Int_3QVal_Int_1_bufchan_buf[0]))
        lizzieLet12_6QVal_Int_3QVal_Int_1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet12_6QVal_Int_3QVal_Int_1_argbuf_r) && (! lizzieLet12_6QVal_Int_3QVal_Int_1_bufchan_buf[0])))
        lizzieLet12_6QVal_Int_3QVal_Int_1_bufchan_buf <= lizzieLet12_6QVal_Int_3QVal_Int_1_bufchan_d;
  
  /* dcon (Ty TupGo___MyDTInt_Bool___Int,
      Dcon TupGo___MyDTInt_Bool___Int) : [(lizzieLet12_6QVal_Int_3QVal_Int_1_argbuf,Go),
                                          (lizzieLet12_6QVal_Int_4QVal_Int_1_argbuf,MyDTInt_Bool),
                                          (es_13_1_argbuf,Int)] > (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int4,TupGo___MyDTInt_Bool___Int) */
  assign applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int4_d = TupGo___MyDTInt_Bool___Int_dc((& {lizzieLet12_6QVal_Int_3QVal_Int_1_argbuf_d[0],
                                                                                            lizzieLet12_6QVal_Int_4QVal_Int_1_argbuf_d[0],
                                                                                            es_13_1_argbuf_d[0]}), lizzieLet12_6QVal_Int_3QVal_Int_1_argbuf_d, lizzieLet12_6QVal_Int_4QVal_Int_1_argbuf_d, es_13_1_argbuf_d);
  assign {lizzieLet12_6QVal_Int_3QVal_Int_1_argbuf_r,
          lizzieLet12_6QVal_Int_4QVal_Int_1_argbuf_r,
          es_13_1_argbuf_r} = {3 {(applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int4_r && applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int4_d[0])}};
  
  /* demux (Ty QTree_Int,
       Ty MyDTInt_Bool) : (lizzieLet12_6QVal_Int_4,QTree_Int) (lizzieLet12_4QVal_Int,MyDTInt_Bool) > [(_29,MyDTInt_Bool),
                                                                                                      (lizzieLet12_6QVal_Int_4QVal_Int,MyDTInt_Bool),
                                                                                                      (_28,MyDTInt_Bool),
                                                                                                      (_27,MyDTInt_Bool)] */
  logic [3:0] lizzieLet12_4QVal_Int_onehotd;
  always_comb
    if ((lizzieLet12_6QVal_Int_4_d[0] && lizzieLet12_4QVal_Int_d[0]))
      unique case (lizzieLet12_6QVal_Int_4_d[2:1])
        2'd0: lizzieLet12_4QVal_Int_onehotd = 4'd1;
        2'd1: lizzieLet12_4QVal_Int_onehotd = 4'd2;
        2'd2: lizzieLet12_4QVal_Int_onehotd = 4'd4;
        2'd3: lizzieLet12_4QVal_Int_onehotd = 4'd8;
        default: lizzieLet12_4QVal_Int_onehotd = 4'd0;
      endcase
    else lizzieLet12_4QVal_Int_onehotd = 4'd0;
  assign _29_d = lizzieLet12_4QVal_Int_onehotd[0];
  assign lizzieLet12_6QVal_Int_4QVal_Int_d = lizzieLet12_4QVal_Int_onehotd[1];
  assign _28_d = lizzieLet12_4QVal_Int_onehotd[2];
  assign _27_d = lizzieLet12_4QVal_Int_onehotd[3];
  assign lizzieLet12_4QVal_Int_r = (| (lizzieLet12_4QVal_Int_onehotd & {_27_r,
                                                                        _28_r,
                                                                        lizzieLet12_6QVal_Int_4QVal_Int_r,
                                                                        _29_r}));
  assign lizzieLet12_6QVal_Int_4_r = lizzieLet12_4QVal_Int_r;
  
  /* buf (Ty MyDTInt_Bool) : (lizzieLet12_6QVal_Int_4QVal_Int,MyDTInt_Bool) > (lizzieLet12_6QVal_Int_4QVal_Int_1_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t lizzieLet12_6QVal_Int_4QVal_Int_bufchan_d;
  logic lizzieLet12_6QVal_Int_4QVal_Int_bufchan_r;
  assign lizzieLet12_6QVal_Int_4QVal_Int_r = ((! lizzieLet12_6QVal_Int_4QVal_Int_bufchan_d[0]) || lizzieLet12_6QVal_Int_4QVal_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QVal_Int_4QVal_Int_bufchan_d <= 1'd0;
    else
      if (lizzieLet12_6QVal_Int_4QVal_Int_r)
        lizzieLet12_6QVal_Int_4QVal_Int_bufchan_d <= lizzieLet12_6QVal_Int_4QVal_Int_d;
  MyDTInt_Bool_t lizzieLet12_6QVal_Int_4QVal_Int_bufchan_buf;
  assign lizzieLet12_6QVal_Int_4QVal_Int_bufchan_r = (! lizzieLet12_6QVal_Int_4QVal_Int_bufchan_buf[0]);
  assign lizzieLet12_6QVal_Int_4QVal_Int_1_argbuf_d = (lizzieLet12_6QVal_Int_4QVal_Int_bufchan_buf[0] ? lizzieLet12_6QVal_Int_4QVal_Int_bufchan_buf :
                                                       lizzieLet12_6QVal_Int_4QVal_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QVal_Int_4QVal_Int_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet12_6QVal_Int_4QVal_Int_1_argbuf_r && lizzieLet12_6QVal_Int_4QVal_Int_bufchan_buf[0]))
        lizzieLet12_6QVal_Int_4QVal_Int_bufchan_buf <= 1'd0;
      else if (((! lizzieLet12_6QVal_Int_4QVal_Int_1_argbuf_r) && (! lizzieLet12_6QVal_Int_4QVal_Int_bufchan_buf[0])))
        lizzieLet12_6QVal_Int_4QVal_Int_bufchan_buf <= lizzieLet12_6QVal_Int_4QVal_Int_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty MyDTInt_Bool) : (lizzieLet12_6QVal_Int_5,QTree_Int) (lizzieLet12_5QVal_Int,MyDTInt_Bool) > [(lizzieLet12_6QVal_Int_5QNone_Int,MyDTInt_Bool),
                                                                                                      (lizzieLet12_6QVal_Int_5QVal_Int,MyDTInt_Bool),
                                                                                                      (_26,MyDTInt_Bool),
                                                                                                      (_25,MyDTInt_Bool)] */
  logic [3:0] lizzieLet12_5QVal_Int_onehotd;
  always_comb
    if ((lizzieLet12_6QVal_Int_5_d[0] && lizzieLet12_5QVal_Int_d[0]))
      unique case (lizzieLet12_6QVal_Int_5_d[2:1])
        2'd0: lizzieLet12_5QVal_Int_onehotd = 4'd1;
        2'd1: lizzieLet12_5QVal_Int_onehotd = 4'd2;
        2'd2: lizzieLet12_5QVal_Int_onehotd = 4'd4;
        2'd3: lizzieLet12_5QVal_Int_onehotd = 4'd8;
        default: lizzieLet12_5QVal_Int_onehotd = 4'd0;
      endcase
    else lizzieLet12_5QVal_Int_onehotd = 4'd0;
  assign lizzieLet12_6QVal_Int_5QNone_Int_d = lizzieLet12_5QVal_Int_onehotd[0];
  assign lizzieLet12_6QVal_Int_5QVal_Int_d = lizzieLet12_5QVal_Int_onehotd[1];
  assign _26_d = lizzieLet12_5QVal_Int_onehotd[2];
  assign _25_d = lizzieLet12_5QVal_Int_onehotd[3];
  assign lizzieLet12_5QVal_Int_r = (| (lizzieLet12_5QVal_Int_onehotd & {_25_r,
                                                                        _26_r,
                                                                        lizzieLet12_6QVal_Int_5QVal_Int_r,
                                                                        lizzieLet12_6QVal_Int_5QNone_Int_r}));
  assign lizzieLet12_6QVal_Int_5_r = lizzieLet12_5QVal_Int_r;
  
  /* buf (Ty MyDTInt_Bool) : (lizzieLet12_6QVal_Int_5QNone_Int,MyDTInt_Bool) > (lizzieLet12_6QVal_Int_5QNone_Int_1_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t lizzieLet12_6QVal_Int_5QNone_Int_bufchan_d;
  logic lizzieLet12_6QVal_Int_5QNone_Int_bufchan_r;
  assign lizzieLet12_6QVal_Int_5QNone_Int_r = ((! lizzieLet12_6QVal_Int_5QNone_Int_bufchan_d[0]) || lizzieLet12_6QVal_Int_5QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QVal_Int_5QNone_Int_bufchan_d <= 1'd0;
    else
      if (lizzieLet12_6QVal_Int_5QNone_Int_r)
        lizzieLet12_6QVal_Int_5QNone_Int_bufchan_d <= lizzieLet12_6QVal_Int_5QNone_Int_d;
  MyDTInt_Bool_t lizzieLet12_6QVal_Int_5QNone_Int_bufchan_buf;
  assign lizzieLet12_6QVal_Int_5QNone_Int_bufchan_r = (! lizzieLet12_6QVal_Int_5QNone_Int_bufchan_buf[0]);
  assign lizzieLet12_6QVal_Int_5QNone_Int_1_argbuf_d = (lizzieLet12_6QVal_Int_5QNone_Int_bufchan_buf[0] ? lizzieLet12_6QVal_Int_5QNone_Int_bufchan_buf :
                                                        lizzieLet12_6QVal_Int_5QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QVal_Int_5QNone_Int_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet12_6QVal_Int_5QNone_Int_1_argbuf_r && lizzieLet12_6QVal_Int_5QNone_Int_bufchan_buf[0]))
        lizzieLet12_6QVal_Int_5QNone_Int_bufchan_buf <= 1'd0;
      else if (((! lizzieLet12_6QVal_Int_5QNone_Int_1_argbuf_r) && (! lizzieLet12_6QVal_Int_5QNone_Int_bufchan_buf[0])))
        lizzieLet12_6QVal_Int_5QNone_Int_bufchan_buf <= lizzieLet12_6QVal_Int_5QNone_Int_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty MyDTInt_Int_Int) : (lizzieLet12_6QVal_Int_6,QTree_Int) (lizzieLet12_7QVal_Int,MyDTInt_Int_Int) > [(_24,MyDTInt_Int_Int),
                                                                                                            (lizzieLet12_6QVal_Int_6QVal_Int,MyDTInt_Int_Int),
                                                                                                            (_23,MyDTInt_Int_Int),
                                                                                                            (_22,MyDTInt_Int_Int)] */
  logic [3:0] lizzieLet12_7QVal_Int_onehotd;
  always_comb
    if ((lizzieLet12_6QVal_Int_6_d[0] && lizzieLet12_7QVal_Int_d[0]))
      unique case (lizzieLet12_6QVal_Int_6_d[2:1])
        2'd0: lizzieLet12_7QVal_Int_onehotd = 4'd1;
        2'd1: lizzieLet12_7QVal_Int_onehotd = 4'd2;
        2'd2: lizzieLet12_7QVal_Int_onehotd = 4'd4;
        2'd3: lizzieLet12_7QVal_Int_onehotd = 4'd8;
        default: lizzieLet12_7QVal_Int_onehotd = 4'd0;
      endcase
    else lizzieLet12_7QVal_Int_onehotd = 4'd0;
  assign _24_d = lizzieLet12_7QVal_Int_onehotd[0];
  assign lizzieLet12_6QVal_Int_6QVal_Int_d = lizzieLet12_7QVal_Int_onehotd[1];
  assign _23_d = lizzieLet12_7QVal_Int_onehotd[2];
  assign _22_d = lizzieLet12_7QVal_Int_onehotd[3];
  assign lizzieLet12_7QVal_Int_r = (| (lizzieLet12_7QVal_Int_onehotd & {_22_r,
                                                                        _23_r,
                                                                        lizzieLet12_6QVal_Int_6QVal_Int_r,
                                                                        _24_r}));
  assign lizzieLet12_6QVal_Int_6_r = lizzieLet12_7QVal_Int_r;
  
  /* fork (Ty MyDTInt_Int_Int) : (lizzieLet12_6QVal_Int_6QVal_Int,MyDTInt_Int_Int) > [(lizzieLet12_6QVal_Int_6QVal_Int_1,MyDTInt_Int_Int),
                                                                                 (lizzieLet12_6QVal_Int_6QVal_Int_2,MyDTInt_Int_Int)] */
  logic [1:0] lizzieLet12_6QVal_Int_6QVal_Int_emitted;
  logic [1:0] lizzieLet12_6QVal_Int_6QVal_Int_done;
  assign lizzieLet12_6QVal_Int_6QVal_Int_1_d = (lizzieLet12_6QVal_Int_6QVal_Int_d[0] && (! lizzieLet12_6QVal_Int_6QVal_Int_emitted[0]));
  assign lizzieLet12_6QVal_Int_6QVal_Int_2_d = (lizzieLet12_6QVal_Int_6QVal_Int_d[0] && (! lizzieLet12_6QVal_Int_6QVal_Int_emitted[1]));
  assign lizzieLet12_6QVal_Int_6QVal_Int_done = (lizzieLet12_6QVal_Int_6QVal_Int_emitted | ({lizzieLet12_6QVal_Int_6QVal_Int_2_d[0],
                                                                                             lizzieLet12_6QVal_Int_6QVal_Int_1_d[0]} & {lizzieLet12_6QVal_Int_6QVal_Int_2_r,
                                                                                                                                        lizzieLet12_6QVal_Int_6QVal_Int_1_r}));
  assign lizzieLet12_6QVal_Int_6QVal_Int_r = (& lizzieLet12_6QVal_Int_6QVal_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QVal_Int_6QVal_Int_emitted <= 2'd0;
    else
      lizzieLet12_6QVal_Int_6QVal_Int_emitted <= (lizzieLet12_6QVal_Int_6QVal_Int_r ? 2'd0 :
                                                  lizzieLet12_6QVal_Int_6QVal_Int_done);
  
  /* buf (Ty MyDTInt_Int_Int) : (lizzieLet12_6QVal_Int_6QVal_Int_1,MyDTInt_Int_Int) > (lizzieLet12_6QVal_Int_6QVal_Int_1_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t lizzieLet12_6QVal_Int_6QVal_Int_1_bufchan_d;
  logic lizzieLet12_6QVal_Int_6QVal_Int_1_bufchan_r;
  assign lizzieLet12_6QVal_Int_6QVal_Int_1_r = ((! lizzieLet12_6QVal_Int_6QVal_Int_1_bufchan_d[0]) || lizzieLet12_6QVal_Int_6QVal_Int_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QVal_Int_6QVal_Int_1_bufchan_d <= 1'd0;
    else
      if (lizzieLet12_6QVal_Int_6QVal_Int_1_r)
        lizzieLet12_6QVal_Int_6QVal_Int_1_bufchan_d <= lizzieLet12_6QVal_Int_6QVal_Int_1_d;
  MyDTInt_Int_Int_t lizzieLet12_6QVal_Int_6QVal_Int_1_bufchan_buf;
  assign lizzieLet12_6QVal_Int_6QVal_Int_1_bufchan_r = (! lizzieLet12_6QVal_Int_6QVal_Int_1_bufchan_buf[0]);
  assign lizzieLet12_6QVal_Int_6QVal_Int_1_argbuf_d = (lizzieLet12_6QVal_Int_6QVal_Int_1_bufchan_buf[0] ? lizzieLet12_6QVal_Int_6QVal_Int_1_bufchan_buf :
                                                       lizzieLet12_6QVal_Int_6QVal_Int_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QVal_Int_6QVal_Int_1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet12_6QVal_Int_6QVal_Int_1_argbuf_r && lizzieLet12_6QVal_Int_6QVal_Int_1_bufchan_buf[0]))
        lizzieLet12_6QVal_Int_6QVal_Int_1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet12_6QVal_Int_6QVal_Int_1_argbuf_r) && (! lizzieLet12_6QVal_Int_6QVal_Int_1_bufchan_buf[0])))
        lizzieLet12_6QVal_Int_6QVal_Int_1_bufchan_buf <= lizzieLet12_6QVal_Int_6QVal_Int_1_bufchan_d;
  
  /* dcon (Ty TupMyDTInt_Int_Int___Int___Int,
      Dcon TupMyDTInt_Int_Int___Int___Int) : [(lizzieLet12_6QVal_Int_6QVal_Int_1_argbuf,MyDTInt_Int_Int),
                                              (lizzieLet12_6QVal_Int_9QVal_Int_1_argbuf,Int),
                                              (va8O_1_argbuf,Int)] > (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1,TupMyDTInt_Int_Int___Int___Int) */
  assign applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_d = TupMyDTInt_Int_Int___Int___Int_dc((& {lizzieLet12_6QVal_Int_6QVal_Int_1_argbuf_d[0],
                                                                                                        lizzieLet12_6QVal_Int_9QVal_Int_1_argbuf_d[0],
                                                                                                        va8O_1_argbuf_d[0]}), lizzieLet12_6QVal_Int_6QVal_Int_1_argbuf_d, lizzieLet12_6QVal_Int_9QVal_Int_1_argbuf_d, va8O_1_argbuf_d);
  assign {lizzieLet12_6QVal_Int_6QVal_Int_1_argbuf_r,
          lizzieLet12_6QVal_Int_9QVal_Int_1_argbuf_r,
          va8O_1_argbuf_r} = {3 {(applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_r && applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_d[0])}};
  
  /* demux (Ty QTree_Int,
       Ty MyDTInt_Int) : (lizzieLet12_6QVal_Int_7,QTree_Int) (lizzieLet12_8QVal_Int,MyDTInt_Int) > [(lizzieLet12_6QVal_Int_7QNone_Int,MyDTInt_Int),
                                                                                                    (lizzieLet12_6QVal_Int_7QVal_Int,MyDTInt_Int),
                                                                                                    (_21,MyDTInt_Int),
                                                                                                    (_20,MyDTInt_Int)] */
  logic [3:0] lizzieLet12_8QVal_Int_onehotd;
  always_comb
    if ((lizzieLet12_6QVal_Int_7_d[0] && lizzieLet12_8QVal_Int_d[0]))
      unique case (lizzieLet12_6QVal_Int_7_d[2:1])
        2'd0: lizzieLet12_8QVal_Int_onehotd = 4'd1;
        2'd1: lizzieLet12_8QVal_Int_onehotd = 4'd2;
        2'd2: lizzieLet12_8QVal_Int_onehotd = 4'd4;
        2'd3: lizzieLet12_8QVal_Int_onehotd = 4'd8;
        default: lizzieLet12_8QVal_Int_onehotd = 4'd0;
      endcase
    else lizzieLet12_8QVal_Int_onehotd = 4'd0;
  assign lizzieLet12_6QVal_Int_7QNone_Int_d = lizzieLet12_8QVal_Int_onehotd[0];
  assign lizzieLet12_6QVal_Int_7QVal_Int_d = lizzieLet12_8QVal_Int_onehotd[1];
  assign _21_d = lizzieLet12_8QVal_Int_onehotd[2];
  assign _20_d = lizzieLet12_8QVal_Int_onehotd[3];
  assign lizzieLet12_8QVal_Int_r = (| (lizzieLet12_8QVal_Int_onehotd & {_20_r,
                                                                        _21_r,
                                                                        lizzieLet12_6QVal_Int_7QVal_Int_r,
                                                                        lizzieLet12_6QVal_Int_7QNone_Int_r}));
  assign lizzieLet12_6QVal_Int_7_r = lizzieLet12_8QVal_Int_r;
  
  /* fork (Ty MyDTInt_Int) : (lizzieLet12_6QVal_Int_7QNone_Int,MyDTInt_Int) > [(lizzieLet12_6QVal_Int_7QNone_Int_1,MyDTInt_Int),
                                                                          (lizzieLet12_6QVal_Int_7QNone_Int_2,MyDTInt_Int)] */
  logic [1:0] lizzieLet12_6QVal_Int_7QNone_Int_emitted;
  logic [1:0] lizzieLet12_6QVal_Int_7QNone_Int_done;
  assign lizzieLet12_6QVal_Int_7QNone_Int_1_d = (lizzieLet12_6QVal_Int_7QNone_Int_d[0] && (! lizzieLet12_6QVal_Int_7QNone_Int_emitted[0]));
  assign lizzieLet12_6QVal_Int_7QNone_Int_2_d = (lizzieLet12_6QVal_Int_7QNone_Int_d[0] && (! lizzieLet12_6QVal_Int_7QNone_Int_emitted[1]));
  assign lizzieLet12_6QVal_Int_7QNone_Int_done = (lizzieLet12_6QVal_Int_7QNone_Int_emitted | ({lizzieLet12_6QVal_Int_7QNone_Int_2_d[0],
                                                                                               lizzieLet12_6QVal_Int_7QNone_Int_1_d[0]} & {lizzieLet12_6QVal_Int_7QNone_Int_2_r,
                                                                                                                                           lizzieLet12_6QVal_Int_7QNone_Int_1_r}));
  assign lizzieLet12_6QVal_Int_7QNone_Int_r = (& lizzieLet12_6QVal_Int_7QNone_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QVal_Int_7QNone_Int_emitted <= 2'd0;
    else
      lizzieLet12_6QVal_Int_7QNone_Int_emitted <= (lizzieLet12_6QVal_Int_7QNone_Int_r ? 2'd0 :
                                                   lizzieLet12_6QVal_Int_7QNone_Int_done);
  
  /* buf (Ty MyDTInt_Int) : (lizzieLet12_6QVal_Int_7QNone_Int_1,MyDTInt_Int) > (lizzieLet12_6QVal_Int_7QNone_Int_1_argbuf,MyDTInt_Int) */
  MyDTInt_Int_t lizzieLet12_6QVal_Int_7QNone_Int_1_bufchan_d;
  logic lizzieLet12_6QVal_Int_7QNone_Int_1_bufchan_r;
  assign lizzieLet12_6QVal_Int_7QNone_Int_1_r = ((! lizzieLet12_6QVal_Int_7QNone_Int_1_bufchan_d[0]) || lizzieLet12_6QVal_Int_7QNone_Int_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QVal_Int_7QNone_Int_1_bufchan_d <= 1'd0;
    else
      if (lizzieLet12_6QVal_Int_7QNone_Int_1_r)
        lizzieLet12_6QVal_Int_7QNone_Int_1_bufchan_d <= lizzieLet12_6QVal_Int_7QNone_Int_1_d;
  MyDTInt_Int_t lizzieLet12_6QVal_Int_7QNone_Int_1_bufchan_buf;
  assign lizzieLet12_6QVal_Int_7QNone_Int_1_bufchan_r = (! lizzieLet12_6QVal_Int_7QNone_Int_1_bufchan_buf[0]);
  assign lizzieLet12_6QVal_Int_7QNone_Int_1_argbuf_d = (lizzieLet12_6QVal_Int_7QNone_Int_1_bufchan_buf[0] ? lizzieLet12_6QVal_Int_7QNone_Int_1_bufchan_buf :
                                                        lizzieLet12_6QVal_Int_7QNone_Int_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QVal_Int_7QNone_Int_1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet12_6QVal_Int_7QNone_Int_1_argbuf_r && lizzieLet12_6QVal_Int_7QNone_Int_1_bufchan_buf[0]))
        lizzieLet12_6QVal_Int_7QNone_Int_1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet12_6QVal_Int_7QNone_Int_1_argbuf_r) && (! lizzieLet12_6QVal_Int_7QNone_Int_1_bufchan_buf[0])))
        lizzieLet12_6QVal_Int_7QNone_Int_1_bufchan_buf <= lizzieLet12_6QVal_Int_7QNone_Int_1_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_CTf_f_Int_Int) : (lizzieLet12_6QVal_Int_8,QTree_Int) (lizzieLet12_9QVal_Int,Pointer_CTf_f_Int_Int) > [(lizzieLet12_6QVal_Int_8QNone_Int,Pointer_CTf_f_Int_Int),
                                                                                                                        (lizzieLet12_6QVal_Int_8QVal_Int,Pointer_CTf_f_Int_Int),
                                                                                                                        (lizzieLet12_6QVal_Int_8QNode_Int,Pointer_CTf_f_Int_Int),
                                                                                                                        (lizzieLet12_6QVal_Int_8QError_Int,Pointer_CTf_f_Int_Int)] */
  logic [3:0] lizzieLet12_9QVal_Int_onehotd;
  always_comb
    if ((lizzieLet12_6QVal_Int_8_d[0] && lizzieLet12_9QVal_Int_d[0]))
      unique case (lizzieLet12_6QVal_Int_8_d[2:1])
        2'd0: lizzieLet12_9QVal_Int_onehotd = 4'd1;
        2'd1: lizzieLet12_9QVal_Int_onehotd = 4'd2;
        2'd2: lizzieLet12_9QVal_Int_onehotd = 4'd4;
        2'd3: lizzieLet12_9QVal_Int_onehotd = 4'd8;
        default: lizzieLet12_9QVal_Int_onehotd = 4'd0;
      endcase
    else lizzieLet12_9QVal_Int_onehotd = 4'd0;
  assign lizzieLet12_6QVal_Int_8QNone_Int_d = {lizzieLet12_9QVal_Int_d[16:1],
                                               lizzieLet12_9QVal_Int_onehotd[0]};
  assign lizzieLet12_6QVal_Int_8QVal_Int_d = {lizzieLet12_9QVal_Int_d[16:1],
                                              lizzieLet12_9QVal_Int_onehotd[1]};
  assign lizzieLet12_6QVal_Int_8QNode_Int_d = {lizzieLet12_9QVal_Int_d[16:1],
                                               lizzieLet12_9QVal_Int_onehotd[2]};
  assign lizzieLet12_6QVal_Int_8QError_Int_d = {lizzieLet12_9QVal_Int_d[16:1],
                                                lizzieLet12_9QVal_Int_onehotd[3]};
  assign lizzieLet12_9QVal_Int_r = (| (lizzieLet12_9QVal_Int_onehotd & {lizzieLet12_6QVal_Int_8QError_Int_r,
                                                                        lizzieLet12_6QVal_Int_8QNode_Int_r,
                                                                        lizzieLet12_6QVal_Int_8QVal_Int_r,
                                                                        lizzieLet12_6QVal_Int_8QNone_Int_r}));
  assign lizzieLet12_6QVal_Int_8_r = lizzieLet12_9QVal_Int_r;
  
  /* buf (Ty Pointer_CTf_f_Int_Int) : (lizzieLet12_6QVal_Int_8QError_Int,Pointer_CTf_f_Int_Int) > (lizzieLet12_6QVal_Int_8QError_Int_1_argbuf,Pointer_CTf_f_Int_Int) */
  Pointer_CTf_f_Int_Int_t lizzieLet12_6QVal_Int_8QError_Int_bufchan_d;
  logic lizzieLet12_6QVal_Int_8QError_Int_bufchan_r;
  assign lizzieLet12_6QVal_Int_8QError_Int_r = ((! lizzieLet12_6QVal_Int_8QError_Int_bufchan_d[0]) || lizzieLet12_6QVal_Int_8QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QVal_Int_8QError_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet12_6QVal_Int_8QError_Int_r)
        lizzieLet12_6QVal_Int_8QError_Int_bufchan_d <= lizzieLet12_6QVal_Int_8QError_Int_d;
  Pointer_CTf_f_Int_Int_t lizzieLet12_6QVal_Int_8QError_Int_bufchan_buf;
  assign lizzieLet12_6QVal_Int_8QError_Int_bufchan_r = (! lizzieLet12_6QVal_Int_8QError_Int_bufchan_buf[0]);
  assign lizzieLet12_6QVal_Int_8QError_Int_1_argbuf_d = (lizzieLet12_6QVal_Int_8QError_Int_bufchan_buf[0] ? lizzieLet12_6QVal_Int_8QError_Int_bufchan_buf :
                                                         lizzieLet12_6QVal_Int_8QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QVal_Int_8QError_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet12_6QVal_Int_8QError_Int_1_argbuf_r && lizzieLet12_6QVal_Int_8QError_Int_bufchan_buf[0]))
        lizzieLet12_6QVal_Int_8QError_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet12_6QVal_Int_8QError_Int_1_argbuf_r) && (! lizzieLet12_6QVal_Int_8QError_Int_bufchan_buf[0])))
        lizzieLet12_6QVal_Int_8QError_Int_bufchan_buf <= lizzieLet12_6QVal_Int_8QError_Int_bufchan_d;
  
  /* buf (Ty Pointer_CTf_f_Int_Int) : (lizzieLet12_6QVal_Int_8QNode_Int,Pointer_CTf_f_Int_Int) > (lizzieLet12_6QVal_Int_8QNode_Int_1_argbuf,Pointer_CTf_f_Int_Int) */
  Pointer_CTf_f_Int_Int_t lizzieLet12_6QVal_Int_8QNode_Int_bufchan_d;
  logic lizzieLet12_6QVal_Int_8QNode_Int_bufchan_r;
  assign lizzieLet12_6QVal_Int_8QNode_Int_r = ((! lizzieLet12_6QVal_Int_8QNode_Int_bufchan_d[0]) || lizzieLet12_6QVal_Int_8QNode_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QVal_Int_8QNode_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet12_6QVal_Int_8QNode_Int_r)
        lizzieLet12_6QVal_Int_8QNode_Int_bufchan_d <= lizzieLet12_6QVal_Int_8QNode_Int_d;
  Pointer_CTf_f_Int_Int_t lizzieLet12_6QVal_Int_8QNode_Int_bufchan_buf;
  assign lizzieLet12_6QVal_Int_8QNode_Int_bufchan_r = (! lizzieLet12_6QVal_Int_8QNode_Int_bufchan_buf[0]);
  assign lizzieLet12_6QVal_Int_8QNode_Int_1_argbuf_d = (lizzieLet12_6QVal_Int_8QNode_Int_bufchan_buf[0] ? lizzieLet12_6QVal_Int_8QNode_Int_bufchan_buf :
                                                        lizzieLet12_6QVal_Int_8QNode_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QVal_Int_8QNode_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet12_6QVal_Int_8QNode_Int_1_argbuf_r && lizzieLet12_6QVal_Int_8QNode_Int_bufchan_buf[0]))
        lizzieLet12_6QVal_Int_8QNode_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet12_6QVal_Int_8QNode_Int_1_argbuf_r) && (! lizzieLet12_6QVal_Int_8QNode_Int_bufchan_buf[0])))
        lizzieLet12_6QVal_Int_8QNode_Int_bufchan_buf <= lizzieLet12_6QVal_Int_8QNode_Int_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Int) : (lizzieLet12_6QVal_Int_9,QTree_Int) (v1a8N_destruct,Int) > [(lizzieLet12_6QVal_Int_9QNone_Int,Int),
                                                                             (lizzieLet12_6QVal_Int_9QVal_Int,Int),
                                                                             (_19,Int),
                                                                             (_18,Int)] */
  logic [3:0] v1a8N_destruct_onehotd;
  always_comb
    if ((lizzieLet12_6QVal_Int_9_d[0] && v1a8N_destruct_d[0]))
      unique case (lizzieLet12_6QVal_Int_9_d[2:1])
        2'd0: v1a8N_destruct_onehotd = 4'd1;
        2'd1: v1a8N_destruct_onehotd = 4'd2;
        2'd2: v1a8N_destruct_onehotd = 4'd4;
        2'd3: v1a8N_destruct_onehotd = 4'd8;
        default: v1a8N_destruct_onehotd = 4'd0;
      endcase
    else v1a8N_destruct_onehotd = 4'd0;
  assign lizzieLet12_6QVal_Int_9QNone_Int_d = {v1a8N_destruct_d[32:1],
                                               v1a8N_destruct_onehotd[0]};
  assign lizzieLet12_6QVal_Int_9QVal_Int_d = {v1a8N_destruct_d[32:1],
                                              v1a8N_destruct_onehotd[1]};
  assign _19_d = {v1a8N_destruct_d[32:1], v1a8N_destruct_onehotd[2]};
  assign _18_d = {v1a8N_destruct_d[32:1], v1a8N_destruct_onehotd[3]};
  assign v1a8N_destruct_r = (| (v1a8N_destruct_onehotd & {_18_r,
                                                          _19_r,
                                                          lizzieLet12_6QVal_Int_9QVal_Int_r,
                                                          lizzieLet12_6QVal_Int_9QNone_Int_r}));
  assign lizzieLet12_6QVal_Int_9_r = v1a8N_destruct_r;
  
  /* fork (Ty Int) : (lizzieLet12_6QVal_Int_9QNone_Int,Int) > [(lizzieLet12_6QVal_Int_9QNone_Int_1,Int),
                                                          (lizzieLet12_6QVal_Int_9QNone_Int_2,Int)] */
  logic [1:0] lizzieLet12_6QVal_Int_9QNone_Int_emitted;
  logic [1:0] lizzieLet12_6QVal_Int_9QNone_Int_done;
  assign lizzieLet12_6QVal_Int_9QNone_Int_1_d = {lizzieLet12_6QVal_Int_9QNone_Int_d[32:1],
                                                 (lizzieLet12_6QVal_Int_9QNone_Int_d[0] && (! lizzieLet12_6QVal_Int_9QNone_Int_emitted[0]))};
  assign lizzieLet12_6QVal_Int_9QNone_Int_2_d = {lizzieLet12_6QVal_Int_9QNone_Int_d[32:1],
                                                 (lizzieLet12_6QVal_Int_9QNone_Int_d[0] && (! lizzieLet12_6QVal_Int_9QNone_Int_emitted[1]))};
  assign lizzieLet12_6QVal_Int_9QNone_Int_done = (lizzieLet12_6QVal_Int_9QNone_Int_emitted | ({lizzieLet12_6QVal_Int_9QNone_Int_2_d[0],
                                                                                               lizzieLet12_6QVal_Int_9QNone_Int_1_d[0]} & {lizzieLet12_6QVal_Int_9QNone_Int_2_r,
                                                                                                                                           lizzieLet12_6QVal_Int_9QNone_Int_1_r}));
  assign lizzieLet12_6QVal_Int_9QNone_Int_r = (& lizzieLet12_6QVal_Int_9QNone_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QVal_Int_9QNone_Int_emitted <= 2'd0;
    else
      lizzieLet12_6QVal_Int_9QNone_Int_emitted <= (lizzieLet12_6QVal_Int_9QNone_Int_r ? 2'd0 :
                                                   lizzieLet12_6QVal_Int_9QNone_Int_done);
  
  /* buf (Ty Int) : (lizzieLet12_6QVal_Int_9QNone_Int_1,Int) > (lizzieLet12_6QVal_Int_9QNone_Int_1_argbuf,Int) */
  Int_t lizzieLet12_6QVal_Int_9QNone_Int_1_bufchan_d;
  logic lizzieLet12_6QVal_Int_9QNone_Int_1_bufchan_r;
  assign lizzieLet12_6QVal_Int_9QNone_Int_1_r = ((! lizzieLet12_6QVal_Int_9QNone_Int_1_bufchan_d[0]) || lizzieLet12_6QVal_Int_9QNone_Int_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QVal_Int_9QNone_Int_1_bufchan_d <= {32'd0, 1'd0};
    else
      if (lizzieLet12_6QVal_Int_9QNone_Int_1_r)
        lizzieLet12_6QVal_Int_9QNone_Int_1_bufchan_d <= lizzieLet12_6QVal_Int_9QNone_Int_1_d;
  Int_t lizzieLet12_6QVal_Int_9QNone_Int_1_bufchan_buf;
  assign lizzieLet12_6QVal_Int_9QNone_Int_1_bufchan_r = (! lizzieLet12_6QVal_Int_9QNone_Int_1_bufchan_buf[0]);
  assign lizzieLet12_6QVal_Int_9QNone_Int_1_argbuf_d = (lizzieLet12_6QVal_Int_9QNone_Int_1_bufchan_buf[0] ? lizzieLet12_6QVal_Int_9QNone_Int_1_bufchan_buf :
                                                        lizzieLet12_6QVal_Int_9QNone_Int_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QVal_Int_9QNone_Int_1_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((lizzieLet12_6QVal_Int_9QNone_Int_1_argbuf_r && lizzieLet12_6QVal_Int_9QNone_Int_1_bufchan_buf[0]))
        lizzieLet12_6QVal_Int_9QNone_Int_1_bufchan_buf <= {32'd0, 1'd0};
      else if (((! lizzieLet12_6QVal_Int_9QNone_Int_1_argbuf_r) && (! lizzieLet12_6QVal_Int_9QNone_Int_1_bufchan_buf[0])))
        lizzieLet12_6QVal_Int_9QNone_Int_1_bufchan_buf <= lizzieLet12_6QVal_Int_9QNone_Int_1_bufchan_d;
  
  /* fork (Ty Int) : (lizzieLet12_6QVal_Int_9QVal_Int,Int) > [(lizzieLet12_6QVal_Int_9QVal_Int_1,Int),
                                                         (lizzieLet12_6QVal_Int_9QVal_Int_2,Int)] */
  logic [1:0] lizzieLet12_6QVal_Int_9QVal_Int_emitted;
  logic [1:0] lizzieLet12_6QVal_Int_9QVal_Int_done;
  assign lizzieLet12_6QVal_Int_9QVal_Int_1_d = {lizzieLet12_6QVal_Int_9QVal_Int_d[32:1],
                                                (lizzieLet12_6QVal_Int_9QVal_Int_d[0] && (! lizzieLet12_6QVal_Int_9QVal_Int_emitted[0]))};
  assign lizzieLet12_6QVal_Int_9QVal_Int_2_d = {lizzieLet12_6QVal_Int_9QVal_Int_d[32:1],
                                                (lizzieLet12_6QVal_Int_9QVal_Int_d[0] && (! lizzieLet12_6QVal_Int_9QVal_Int_emitted[1]))};
  assign lizzieLet12_6QVal_Int_9QVal_Int_done = (lizzieLet12_6QVal_Int_9QVal_Int_emitted | ({lizzieLet12_6QVal_Int_9QVal_Int_2_d[0],
                                                                                             lizzieLet12_6QVal_Int_9QVal_Int_1_d[0]} & {lizzieLet12_6QVal_Int_9QVal_Int_2_r,
                                                                                                                                        lizzieLet12_6QVal_Int_9QVal_Int_1_r}));
  assign lizzieLet12_6QVal_Int_9QVal_Int_r = (& lizzieLet12_6QVal_Int_9QVal_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QVal_Int_9QVal_Int_emitted <= 2'd0;
    else
      lizzieLet12_6QVal_Int_9QVal_Int_emitted <= (lizzieLet12_6QVal_Int_9QVal_Int_r ? 2'd0 :
                                                  lizzieLet12_6QVal_Int_9QVal_Int_done);
  
  /* buf (Ty Int) : (lizzieLet12_6QVal_Int_9QVal_Int_1,Int) > (lizzieLet12_6QVal_Int_9QVal_Int_1_argbuf,Int) */
  Int_t lizzieLet12_6QVal_Int_9QVal_Int_1_bufchan_d;
  logic lizzieLet12_6QVal_Int_9QVal_Int_1_bufchan_r;
  assign lizzieLet12_6QVal_Int_9QVal_Int_1_r = ((! lizzieLet12_6QVal_Int_9QVal_Int_1_bufchan_d[0]) || lizzieLet12_6QVal_Int_9QVal_Int_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QVal_Int_9QVal_Int_1_bufchan_d <= {32'd0, 1'd0};
    else
      if (lizzieLet12_6QVal_Int_9QVal_Int_1_r)
        lizzieLet12_6QVal_Int_9QVal_Int_1_bufchan_d <= lizzieLet12_6QVal_Int_9QVal_Int_1_d;
  Int_t lizzieLet12_6QVal_Int_9QVal_Int_1_bufchan_buf;
  assign lizzieLet12_6QVal_Int_9QVal_Int_1_bufchan_r = (! lizzieLet12_6QVal_Int_9QVal_Int_1_bufchan_buf[0]);
  assign lizzieLet12_6QVal_Int_9QVal_Int_1_argbuf_d = (lizzieLet12_6QVal_Int_9QVal_Int_1_bufchan_buf[0] ? lizzieLet12_6QVal_Int_9QVal_Int_1_bufchan_buf :
                                                       lizzieLet12_6QVal_Int_9QVal_Int_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_6QVal_Int_9QVal_Int_1_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((lizzieLet12_6QVal_Int_9QVal_Int_1_argbuf_r && lizzieLet12_6QVal_Int_9QVal_Int_1_bufchan_buf[0]))
        lizzieLet12_6QVal_Int_9QVal_Int_1_bufchan_buf <= {32'd0, 1'd0};
      else if (((! lizzieLet12_6QVal_Int_9QVal_Int_1_argbuf_r) && (! lizzieLet12_6QVal_Int_9QVal_Int_1_bufchan_buf[0])))
        lizzieLet12_6QVal_Int_9QVal_Int_1_bufchan_buf <= lizzieLet12_6QVal_Int_9QVal_Int_1_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty MyDTInt_Int_Int) : (lizzieLet12_7,QTree_Int) (op_adda8H_goMux_mux,MyDTInt_Int_Int) > [(_17,MyDTInt_Int_Int),
                                                                                                (lizzieLet12_7QVal_Int,MyDTInt_Int_Int),
                                                                                                (lizzieLet12_7QNode_Int,MyDTInt_Int_Int),
                                                                                                (_16,MyDTInt_Int_Int)] */
  logic [3:0] op_adda8H_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet12_7_d[0] && op_adda8H_goMux_mux_d[0]))
      unique case (lizzieLet12_7_d[2:1])
        2'd0: op_adda8H_goMux_mux_onehotd = 4'd1;
        2'd1: op_adda8H_goMux_mux_onehotd = 4'd2;
        2'd2: op_adda8H_goMux_mux_onehotd = 4'd4;
        2'd3: op_adda8H_goMux_mux_onehotd = 4'd8;
        default: op_adda8H_goMux_mux_onehotd = 4'd0;
      endcase
    else op_adda8H_goMux_mux_onehotd = 4'd0;
  assign _17_d = op_adda8H_goMux_mux_onehotd[0];
  assign lizzieLet12_7QVal_Int_d = op_adda8H_goMux_mux_onehotd[1];
  assign lizzieLet12_7QNode_Int_d = op_adda8H_goMux_mux_onehotd[2];
  assign _16_d = op_adda8H_goMux_mux_onehotd[3];
  assign op_adda8H_goMux_mux_r = (| (op_adda8H_goMux_mux_onehotd & {_16_r,
                                                                    lizzieLet12_7QNode_Int_r,
                                                                    lizzieLet12_7QVal_Int_r,
                                                                    _17_r}));
  assign lizzieLet12_7_r = op_adda8H_goMux_mux_r;
  
  /* demux (Ty QTree_Int,
       Ty MyDTInt_Int) : (lizzieLet12_8,QTree_Int) (op_mapa8F_goMux_mux,MyDTInt_Int) > [(lizzieLet12_8QNone_Int,MyDTInt_Int),
                                                                                        (lizzieLet12_8QVal_Int,MyDTInt_Int),
                                                                                        (lizzieLet12_8QNode_Int,MyDTInt_Int),
                                                                                        (_15,MyDTInt_Int)] */
  logic [3:0] op_mapa8F_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet12_8_d[0] && op_mapa8F_goMux_mux_d[0]))
      unique case (lizzieLet12_8_d[2:1])
        2'd0: op_mapa8F_goMux_mux_onehotd = 4'd1;
        2'd1: op_mapa8F_goMux_mux_onehotd = 4'd2;
        2'd2: op_mapa8F_goMux_mux_onehotd = 4'd4;
        2'd3: op_mapa8F_goMux_mux_onehotd = 4'd8;
        default: op_mapa8F_goMux_mux_onehotd = 4'd0;
      endcase
    else op_mapa8F_goMux_mux_onehotd = 4'd0;
  assign lizzieLet12_8QNone_Int_d = op_mapa8F_goMux_mux_onehotd[0];
  assign lizzieLet12_8QVal_Int_d = op_mapa8F_goMux_mux_onehotd[1];
  assign lizzieLet12_8QNode_Int_d = op_mapa8F_goMux_mux_onehotd[2];
  assign _15_d = op_mapa8F_goMux_mux_onehotd[3];
  assign op_mapa8F_goMux_mux_r = (| (op_mapa8F_goMux_mux_onehotd & {_15_r,
                                                                    lizzieLet12_8QNode_Int_r,
                                                                    lizzieLet12_8QVal_Int_r,
                                                                    lizzieLet12_8QNone_Int_r}));
  assign lizzieLet12_8_r = op_mapa8F_goMux_mux_r;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_CTf_f_Int_Int) : (lizzieLet12_9,QTree_Int) (sc_0_2_goMux_mux,Pointer_CTf_f_Int_Int) > [(lizzieLet12_9QNone_Int,Pointer_CTf_f_Int_Int),
                                                                                                         (lizzieLet12_9QVal_Int,Pointer_CTf_f_Int_Int),
                                                                                                         (lizzieLet12_9QNode_Int,Pointer_CTf_f_Int_Int),
                                                                                                         (lizzieLet12_9QError_Int,Pointer_CTf_f_Int_Int)] */
  logic [3:0] sc_0_2_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet12_9_d[0] && sc_0_2_goMux_mux_d[0]))
      unique case (lizzieLet12_9_d[2:1])
        2'd0: sc_0_2_goMux_mux_onehotd = 4'd1;
        2'd1: sc_0_2_goMux_mux_onehotd = 4'd2;
        2'd2: sc_0_2_goMux_mux_onehotd = 4'd4;
        2'd3: sc_0_2_goMux_mux_onehotd = 4'd8;
        default: sc_0_2_goMux_mux_onehotd = 4'd0;
      endcase
    else sc_0_2_goMux_mux_onehotd = 4'd0;
  assign lizzieLet12_9QNone_Int_d = {sc_0_2_goMux_mux_d[16:1],
                                     sc_0_2_goMux_mux_onehotd[0]};
  assign lizzieLet12_9QVal_Int_d = {sc_0_2_goMux_mux_d[16:1],
                                    sc_0_2_goMux_mux_onehotd[1]};
  assign lizzieLet12_9QNode_Int_d = {sc_0_2_goMux_mux_d[16:1],
                                     sc_0_2_goMux_mux_onehotd[2]};
  assign lizzieLet12_9QError_Int_d = {sc_0_2_goMux_mux_d[16:1],
                                      sc_0_2_goMux_mux_onehotd[3]};
  assign sc_0_2_goMux_mux_r = (| (sc_0_2_goMux_mux_onehotd & {lizzieLet12_9QError_Int_r,
                                                              lizzieLet12_9QNode_Int_r,
                                                              lizzieLet12_9QVal_Int_r,
                                                              lizzieLet12_9QNone_Int_r}));
  assign lizzieLet12_9_r = sc_0_2_goMux_mux_r;
  
  /* buf (Ty Pointer_CTf_f_Int_Int) : (lizzieLet12_9QError_Int,Pointer_CTf_f_Int_Int) > (lizzieLet12_9QError_Int_1_argbuf,Pointer_CTf_f_Int_Int) */
  Pointer_CTf_f_Int_Int_t lizzieLet12_9QError_Int_bufchan_d;
  logic lizzieLet12_9QError_Int_bufchan_r;
  assign lizzieLet12_9QError_Int_r = ((! lizzieLet12_9QError_Int_bufchan_d[0]) || lizzieLet12_9QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_9QError_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet12_9QError_Int_r)
        lizzieLet12_9QError_Int_bufchan_d <= lizzieLet12_9QError_Int_d;
  Pointer_CTf_f_Int_Int_t lizzieLet12_9QError_Int_bufchan_buf;
  assign lizzieLet12_9QError_Int_bufchan_r = (! lizzieLet12_9QError_Int_bufchan_buf[0]);
  assign lizzieLet12_9QError_Int_1_argbuf_d = (lizzieLet12_9QError_Int_bufchan_buf[0] ? lizzieLet12_9QError_Int_bufchan_buf :
                                               lizzieLet12_9QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_9QError_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet12_9QError_Int_1_argbuf_r && lizzieLet12_9QError_Int_bufchan_buf[0]))
        lizzieLet12_9QError_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet12_9QError_Int_1_argbuf_r) && (! lizzieLet12_9QError_Int_bufchan_buf[0])))
        lizzieLet12_9QError_Int_bufchan_buf <= lizzieLet12_9QError_Int_bufchan_d;
  
  /* buf (Ty Bool) : (lizzieLet1_1wild1Xr_1_Eq,Bool) > (lizzieLet2_1_argbuf,Bool) */
  Bool_t lizzieLet1_1wild1Xr_1_Eq_bufchan_d;
  logic lizzieLet1_1wild1Xr_1_Eq_bufchan_r;
  assign lizzieLet1_1wild1Xr_1_Eq_r = ((! lizzieLet1_1wild1Xr_1_Eq_bufchan_d[0]) || lizzieLet1_1wild1Xr_1_Eq_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet1_1wild1Xr_1_Eq_bufchan_d <= {1'd0, 1'd0};
    else
      if (lizzieLet1_1wild1Xr_1_Eq_r)
        lizzieLet1_1wild1Xr_1_Eq_bufchan_d <= lizzieLet1_1wild1Xr_1_Eq_d;
  Bool_t lizzieLet1_1wild1Xr_1_Eq_bufchan_buf;
  assign lizzieLet1_1wild1Xr_1_Eq_bufchan_r = (! lizzieLet1_1wild1Xr_1_Eq_bufchan_buf[0]);
  assign lizzieLet2_1_argbuf_d = (lizzieLet1_1wild1Xr_1_Eq_bufchan_buf[0] ? lizzieLet1_1wild1Xr_1_Eq_bufchan_buf :
                                  lizzieLet1_1wild1Xr_1_Eq_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet1_1wild1Xr_1_Eq_bufchan_buf <= {1'd0, 1'd0};
    else
      if ((lizzieLet2_1_argbuf_r && lizzieLet1_1wild1Xr_1_Eq_bufchan_buf[0]))
        lizzieLet1_1wild1Xr_1_Eq_bufchan_buf <= {1'd0, 1'd0};
      else if (((! lizzieLet2_1_argbuf_r) && (! lizzieLet1_1wild1Xr_1_Eq_bufchan_buf[0])))
        lizzieLet1_1wild1Xr_1_Eq_bufchan_buf <= lizzieLet1_1wild1Xr_1_Eq_bufchan_d;
  
  /* destruct (Ty CT$wnnz,
          Dcon Lcall_$wnnz0) : (lizzieLet35_1Lcall_$wnnz0,CT$wnnz) > [(wwsj0_4_destruct,Int#),
                                                                      (ww1Xju_2_destruct,Int#),
                                                                      (ww2Xjx_1_destruct,Int#),
                                                                      (sc_0_6_destruct,Pointer_CT$wnnz)] */
  logic [3:0] lizzieLet35_1Lcall_$wnnz0_emitted;
  logic [3:0] lizzieLet35_1Lcall_$wnnz0_done;
  assign wwsj0_4_destruct_d = {lizzieLet35_1Lcall_$wnnz0_d[35:4],
                               (lizzieLet35_1Lcall_$wnnz0_d[0] && (! lizzieLet35_1Lcall_$wnnz0_emitted[0]))};
  assign ww1Xju_2_destruct_d = {lizzieLet35_1Lcall_$wnnz0_d[67:36],
                                (lizzieLet35_1Lcall_$wnnz0_d[0] && (! lizzieLet35_1Lcall_$wnnz0_emitted[1]))};
  assign ww2Xjx_1_destruct_d = {lizzieLet35_1Lcall_$wnnz0_d[99:68],
                                (lizzieLet35_1Lcall_$wnnz0_d[0] && (! lizzieLet35_1Lcall_$wnnz0_emitted[2]))};
  assign sc_0_6_destruct_d = {lizzieLet35_1Lcall_$wnnz0_d[115:100],
                              (lizzieLet35_1Lcall_$wnnz0_d[0] && (! lizzieLet35_1Lcall_$wnnz0_emitted[3]))};
  assign lizzieLet35_1Lcall_$wnnz0_done = (lizzieLet35_1Lcall_$wnnz0_emitted | ({sc_0_6_destruct_d[0],
                                                                                 ww2Xjx_1_destruct_d[0],
                                                                                 ww1Xju_2_destruct_d[0],
                                                                                 wwsj0_4_destruct_d[0]} & {sc_0_6_destruct_r,
                                                                                                           ww2Xjx_1_destruct_r,
                                                                                                           ww1Xju_2_destruct_r,
                                                                                                           wwsj0_4_destruct_r}));
  assign lizzieLet35_1Lcall_$wnnz0_r = (& lizzieLet35_1Lcall_$wnnz0_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet35_1Lcall_$wnnz0_emitted <= 4'd0;
    else
      lizzieLet35_1Lcall_$wnnz0_emitted <= (lizzieLet35_1Lcall_$wnnz0_r ? 4'd0 :
                                            lizzieLet35_1Lcall_$wnnz0_done);
  
  /* destruct (Ty CT$wnnz,
          Dcon Lcall_$wnnz1) : (lizzieLet35_1Lcall_$wnnz1,CT$wnnz) > [(wwsj0_3_destruct,Int#),
                                                                      (ww1Xju_1_destruct,Int#),
                                                                      (sc_0_5_destruct,Pointer_CT$wnnz),
                                                                      (q4a87_3_destruct,Pointer_QTree_Int)] */
  logic [3:0] lizzieLet35_1Lcall_$wnnz1_emitted;
  logic [3:0] lizzieLet35_1Lcall_$wnnz1_done;
  assign wwsj0_3_destruct_d = {lizzieLet35_1Lcall_$wnnz1_d[35:4],
                               (lizzieLet35_1Lcall_$wnnz1_d[0] && (! lizzieLet35_1Lcall_$wnnz1_emitted[0]))};
  assign ww1Xju_1_destruct_d = {lizzieLet35_1Lcall_$wnnz1_d[67:36],
                                (lizzieLet35_1Lcall_$wnnz1_d[0] && (! lizzieLet35_1Lcall_$wnnz1_emitted[1]))};
  assign sc_0_5_destruct_d = {lizzieLet35_1Lcall_$wnnz1_d[83:68],
                              (lizzieLet35_1Lcall_$wnnz1_d[0] && (! lizzieLet35_1Lcall_$wnnz1_emitted[2]))};
  assign q4a87_3_destruct_d = {lizzieLet35_1Lcall_$wnnz1_d[99:84],
                               (lizzieLet35_1Lcall_$wnnz1_d[0] && (! lizzieLet35_1Lcall_$wnnz1_emitted[3]))};
  assign lizzieLet35_1Lcall_$wnnz1_done = (lizzieLet35_1Lcall_$wnnz1_emitted | ({q4a87_3_destruct_d[0],
                                                                                 sc_0_5_destruct_d[0],
                                                                                 ww1Xju_1_destruct_d[0],
                                                                                 wwsj0_3_destruct_d[0]} & {q4a87_3_destruct_r,
                                                                                                           sc_0_5_destruct_r,
                                                                                                           ww1Xju_1_destruct_r,
                                                                                                           wwsj0_3_destruct_r}));
  assign lizzieLet35_1Lcall_$wnnz1_r = (& lizzieLet35_1Lcall_$wnnz1_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet35_1Lcall_$wnnz1_emitted <= 4'd0;
    else
      lizzieLet35_1Lcall_$wnnz1_emitted <= (lizzieLet35_1Lcall_$wnnz1_r ? 4'd0 :
                                            lizzieLet35_1Lcall_$wnnz1_done);
  
  /* destruct (Ty CT$wnnz,
          Dcon Lcall_$wnnz2) : (lizzieLet35_1Lcall_$wnnz2,CT$wnnz) > [(wwsj0_2_destruct,Int#),
                                                                      (sc_0_4_destruct,Pointer_CT$wnnz),
                                                                      (q4a87_2_destruct,Pointer_QTree_Int),
                                                                      (q3a86_2_destruct,Pointer_QTree_Int)] */
  logic [3:0] lizzieLet35_1Lcall_$wnnz2_emitted;
  logic [3:0] lizzieLet35_1Lcall_$wnnz2_done;
  assign wwsj0_2_destruct_d = {lizzieLet35_1Lcall_$wnnz2_d[35:4],
                               (lizzieLet35_1Lcall_$wnnz2_d[0] && (! lizzieLet35_1Lcall_$wnnz2_emitted[0]))};
  assign sc_0_4_destruct_d = {lizzieLet35_1Lcall_$wnnz2_d[51:36],
                              (lizzieLet35_1Lcall_$wnnz2_d[0] && (! lizzieLet35_1Lcall_$wnnz2_emitted[1]))};
  assign q4a87_2_destruct_d = {lizzieLet35_1Lcall_$wnnz2_d[67:52],
                               (lizzieLet35_1Lcall_$wnnz2_d[0] && (! lizzieLet35_1Lcall_$wnnz2_emitted[2]))};
  assign q3a86_2_destruct_d = {lizzieLet35_1Lcall_$wnnz2_d[83:68],
                               (lizzieLet35_1Lcall_$wnnz2_d[0] && (! lizzieLet35_1Lcall_$wnnz2_emitted[3]))};
  assign lizzieLet35_1Lcall_$wnnz2_done = (lizzieLet35_1Lcall_$wnnz2_emitted | ({q3a86_2_destruct_d[0],
                                                                                 q4a87_2_destruct_d[0],
                                                                                 sc_0_4_destruct_d[0],
                                                                                 wwsj0_2_destruct_d[0]} & {q3a86_2_destruct_r,
                                                                                                           q4a87_2_destruct_r,
                                                                                                           sc_0_4_destruct_r,
                                                                                                           wwsj0_2_destruct_r}));
  assign lizzieLet35_1Lcall_$wnnz2_r = (& lizzieLet35_1Lcall_$wnnz2_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet35_1Lcall_$wnnz2_emitted <= 4'd0;
    else
      lizzieLet35_1Lcall_$wnnz2_emitted <= (lizzieLet35_1Lcall_$wnnz2_r ? 4'd0 :
                                            lizzieLet35_1Lcall_$wnnz2_done);
  
  /* destruct (Ty CT$wnnz,
          Dcon Lcall_$wnnz3) : (lizzieLet35_1Lcall_$wnnz3,CT$wnnz) > [(sc_0_3_destruct,Pointer_CT$wnnz),
                                                                      (q4a87_1_destruct,Pointer_QTree_Int),
                                                                      (q3a86_1_destruct,Pointer_QTree_Int),
                                                                      (q2a85_1_destruct,Pointer_QTree_Int)] */
  logic [3:0] lizzieLet35_1Lcall_$wnnz3_emitted;
  logic [3:0] lizzieLet35_1Lcall_$wnnz3_done;
  assign sc_0_3_destruct_d = {lizzieLet35_1Lcall_$wnnz3_d[19:4],
                              (lizzieLet35_1Lcall_$wnnz3_d[0] && (! lizzieLet35_1Lcall_$wnnz3_emitted[0]))};
  assign q4a87_1_destruct_d = {lizzieLet35_1Lcall_$wnnz3_d[35:20],
                               (lizzieLet35_1Lcall_$wnnz3_d[0] && (! lizzieLet35_1Lcall_$wnnz3_emitted[1]))};
  assign q3a86_1_destruct_d = {lizzieLet35_1Lcall_$wnnz3_d[51:36],
                               (lizzieLet35_1Lcall_$wnnz3_d[0] && (! lizzieLet35_1Lcall_$wnnz3_emitted[2]))};
  assign q2a85_1_destruct_d = {lizzieLet35_1Lcall_$wnnz3_d[67:52],
                               (lizzieLet35_1Lcall_$wnnz3_d[0] && (! lizzieLet35_1Lcall_$wnnz3_emitted[3]))};
  assign lizzieLet35_1Lcall_$wnnz3_done = (lizzieLet35_1Lcall_$wnnz3_emitted | ({q2a85_1_destruct_d[0],
                                                                                 q3a86_1_destruct_d[0],
                                                                                 q4a87_1_destruct_d[0],
                                                                                 sc_0_3_destruct_d[0]} & {q2a85_1_destruct_r,
                                                                                                          q3a86_1_destruct_r,
                                                                                                          q4a87_1_destruct_r,
                                                                                                          sc_0_3_destruct_r}));
  assign lizzieLet35_1Lcall_$wnnz3_r = (& lizzieLet35_1Lcall_$wnnz3_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet35_1Lcall_$wnnz3_emitted <= 4'd0;
    else
      lizzieLet35_1Lcall_$wnnz3_emitted <= (lizzieLet35_1Lcall_$wnnz3_r ? 4'd0 :
                                            lizzieLet35_1Lcall_$wnnz3_done);
  
  /* demux (Ty CT$wnnz,
       Ty CT$wnnz) : (lizzieLet35_2,CT$wnnz) (lizzieLet35_1,CT$wnnz) > [(_14,CT$wnnz),
                                                                        (lizzieLet35_1Lcall_$wnnz3,CT$wnnz),
                                                                        (lizzieLet35_1Lcall_$wnnz2,CT$wnnz),
                                                                        (lizzieLet35_1Lcall_$wnnz1,CT$wnnz),
                                                                        (lizzieLet35_1Lcall_$wnnz0,CT$wnnz)] */
  logic [4:0] lizzieLet35_1_onehotd;
  always_comb
    if ((lizzieLet35_2_d[0] && lizzieLet35_1_d[0]))
      unique case (lizzieLet35_2_d[3:1])
        3'd0: lizzieLet35_1_onehotd = 5'd1;
        3'd1: lizzieLet35_1_onehotd = 5'd2;
        3'd2: lizzieLet35_1_onehotd = 5'd4;
        3'd3: lizzieLet35_1_onehotd = 5'd8;
        3'd4: lizzieLet35_1_onehotd = 5'd16;
        default: lizzieLet35_1_onehotd = 5'd0;
      endcase
    else lizzieLet35_1_onehotd = 5'd0;
  assign _14_d = {lizzieLet35_1_d[115:1], lizzieLet35_1_onehotd[0]};
  assign lizzieLet35_1Lcall_$wnnz3_d = {lizzieLet35_1_d[115:1],
                                        lizzieLet35_1_onehotd[1]};
  assign lizzieLet35_1Lcall_$wnnz2_d = {lizzieLet35_1_d[115:1],
                                        lizzieLet35_1_onehotd[2]};
  assign lizzieLet35_1Lcall_$wnnz1_d = {lizzieLet35_1_d[115:1],
                                        lizzieLet35_1_onehotd[3]};
  assign lizzieLet35_1Lcall_$wnnz0_d = {lizzieLet35_1_d[115:1],
                                        lizzieLet35_1_onehotd[4]};
  assign lizzieLet35_1_r = (| (lizzieLet35_1_onehotd & {lizzieLet35_1Lcall_$wnnz0_r,
                                                        lizzieLet35_1Lcall_$wnnz1_r,
                                                        lizzieLet35_1Lcall_$wnnz2_r,
                                                        lizzieLet35_1Lcall_$wnnz3_r,
                                                        _14_r}));
  assign lizzieLet35_2_r = lizzieLet35_1_r;
  
  /* demux (Ty CT$wnnz,
       Ty Go) : (lizzieLet35_3,CT$wnnz) (go_15_goMux_data,Go) > [(_13,Go),
                                                                 (lizzieLet35_3Lcall_$wnnz3,Go),
                                                                 (lizzieLet35_3Lcall_$wnnz2,Go),
                                                                 (lizzieLet35_3Lcall_$wnnz1,Go),
                                                                 (lizzieLet35_3Lcall_$wnnz0,Go)] */
  logic [4:0] go_15_goMux_data_onehotd;
  always_comb
    if ((lizzieLet35_3_d[0] && go_15_goMux_data_d[0]))
      unique case (lizzieLet35_3_d[3:1])
        3'd0: go_15_goMux_data_onehotd = 5'd1;
        3'd1: go_15_goMux_data_onehotd = 5'd2;
        3'd2: go_15_goMux_data_onehotd = 5'd4;
        3'd3: go_15_goMux_data_onehotd = 5'd8;
        3'd4: go_15_goMux_data_onehotd = 5'd16;
        default: go_15_goMux_data_onehotd = 5'd0;
      endcase
    else go_15_goMux_data_onehotd = 5'd0;
  assign _13_d = go_15_goMux_data_onehotd[0];
  assign lizzieLet35_3Lcall_$wnnz3_d = go_15_goMux_data_onehotd[1];
  assign lizzieLet35_3Lcall_$wnnz2_d = go_15_goMux_data_onehotd[2];
  assign lizzieLet35_3Lcall_$wnnz1_d = go_15_goMux_data_onehotd[3];
  assign lizzieLet35_3Lcall_$wnnz0_d = go_15_goMux_data_onehotd[4];
  assign go_15_goMux_data_r = (| (go_15_goMux_data_onehotd & {lizzieLet35_3Lcall_$wnnz0_r,
                                                              lizzieLet35_3Lcall_$wnnz1_r,
                                                              lizzieLet35_3Lcall_$wnnz2_r,
                                                              lizzieLet35_3Lcall_$wnnz3_r,
                                                              _13_r}));
  assign lizzieLet35_3_r = go_15_goMux_data_r;
  
  /* buf (Ty Go) : (lizzieLet35_3Lcall_$wnnz0,Go) > (lizzieLet35_3Lcall_$wnnz0_1_argbuf,Go) */
  Go_t lizzieLet35_3Lcall_$wnnz0_bufchan_d;
  logic lizzieLet35_3Lcall_$wnnz0_bufchan_r;
  assign lizzieLet35_3Lcall_$wnnz0_r = ((! lizzieLet35_3Lcall_$wnnz0_bufchan_d[0]) || lizzieLet35_3Lcall_$wnnz0_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet35_3Lcall_$wnnz0_bufchan_d <= 1'd0;
    else
      if (lizzieLet35_3Lcall_$wnnz0_r)
        lizzieLet35_3Lcall_$wnnz0_bufchan_d <= lizzieLet35_3Lcall_$wnnz0_d;
  Go_t lizzieLet35_3Lcall_$wnnz0_bufchan_buf;
  assign lizzieLet35_3Lcall_$wnnz0_bufchan_r = (! lizzieLet35_3Lcall_$wnnz0_bufchan_buf[0]);
  assign lizzieLet35_3Lcall_$wnnz0_1_argbuf_d = (lizzieLet35_3Lcall_$wnnz0_bufchan_buf[0] ? lizzieLet35_3Lcall_$wnnz0_bufchan_buf :
                                                 lizzieLet35_3Lcall_$wnnz0_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet35_3Lcall_$wnnz0_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet35_3Lcall_$wnnz0_1_argbuf_r && lizzieLet35_3Lcall_$wnnz0_bufchan_buf[0]))
        lizzieLet35_3Lcall_$wnnz0_bufchan_buf <= 1'd0;
      else if (((! lizzieLet35_3Lcall_$wnnz0_1_argbuf_r) && (! lizzieLet35_3Lcall_$wnnz0_bufchan_buf[0])))
        lizzieLet35_3Lcall_$wnnz0_bufchan_buf <= lizzieLet35_3Lcall_$wnnz0_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet35_3Lcall_$wnnz1,Go) > (lizzieLet35_3Lcall_$wnnz1_1_argbuf,Go) */
  Go_t lizzieLet35_3Lcall_$wnnz1_bufchan_d;
  logic lizzieLet35_3Lcall_$wnnz1_bufchan_r;
  assign lizzieLet35_3Lcall_$wnnz1_r = ((! lizzieLet35_3Lcall_$wnnz1_bufchan_d[0]) || lizzieLet35_3Lcall_$wnnz1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet35_3Lcall_$wnnz1_bufchan_d <= 1'd0;
    else
      if (lizzieLet35_3Lcall_$wnnz1_r)
        lizzieLet35_3Lcall_$wnnz1_bufchan_d <= lizzieLet35_3Lcall_$wnnz1_d;
  Go_t lizzieLet35_3Lcall_$wnnz1_bufchan_buf;
  assign lizzieLet35_3Lcall_$wnnz1_bufchan_r = (! lizzieLet35_3Lcall_$wnnz1_bufchan_buf[0]);
  assign lizzieLet35_3Lcall_$wnnz1_1_argbuf_d = (lizzieLet35_3Lcall_$wnnz1_bufchan_buf[0] ? lizzieLet35_3Lcall_$wnnz1_bufchan_buf :
                                                 lizzieLet35_3Lcall_$wnnz1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet35_3Lcall_$wnnz1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet35_3Lcall_$wnnz1_1_argbuf_r && lizzieLet35_3Lcall_$wnnz1_bufchan_buf[0]))
        lizzieLet35_3Lcall_$wnnz1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet35_3Lcall_$wnnz1_1_argbuf_r) && (! lizzieLet35_3Lcall_$wnnz1_bufchan_buf[0])))
        lizzieLet35_3Lcall_$wnnz1_bufchan_buf <= lizzieLet35_3Lcall_$wnnz1_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet35_3Lcall_$wnnz2,Go) > (lizzieLet35_3Lcall_$wnnz2_1_argbuf,Go) */
  Go_t lizzieLet35_3Lcall_$wnnz2_bufchan_d;
  logic lizzieLet35_3Lcall_$wnnz2_bufchan_r;
  assign lizzieLet35_3Lcall_$wnnz2_r = ((! lizzieLet35_3Lcall_$wnnz2_bufchan_d[0]) || lizzieLet35_3Lcall_$wnnz2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet35_3Lcall_$wnnz2_bufchan_d <= 1'd0;
    else
      if (lizzieLet35_3Lcall_$wnnz2_r)
        lizzieLet35_3Lcall_$wnnz2_bufchan_d <= lizzieLet35_3Lcall_$wnnz2_d;
  Go_t lizzieLet35_3Lcall_$wnnz2_bufchan_buf;
  assign lizzieLet35_3Lcall_$wnnz2_bufchan_r = (! lizzieLet35_3Lcall_$wnnz2_bufchan_buf[0]);
  assign lizzieLet35_3Lcall_$wnnz2_1_argbuf_d = (lizzieLet35_3Lcall_$wnnz2_bufchan_buf[0] ? lizzieLet35_3Lcall_$wnnz2_bufchan_buf :
                                                 lizzieLet35_3Lcall_$wnnz2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet35_3Lcall_$wnnz2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet35_3Lcall_$wnnz2_1_argbuf_r && lizzieLet35_3Lcall_$wnnz2_bufchan_buf[0]))
        lizzieLet35_3Lcall_$wnnz2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet35_3Lcall_$wnnz2_1_argbuf_r) && (! lizzieLet35_3Lcall_$wnnz2_bufchan_buf[0])))
        lizzieLet35_3Lcall_$wnnz2_bufchan_buf <= lizzieLet35_3Lcall_$wnnz2_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet35_3Lcall_$wnnz3,Go) > (lizzieLet35_3Lcall_$wnnz3_1_argbuf,Go) */
  Go_t lizzieLet35_3Lcall_$wnnz3_bufchan_d;
  logic lizzieLet35_3Lcall_$wnnz3_bufchan_r;
  assign lizzieLet35_3Lcall_$wnnz3_r = ((! lizzieLet35_3Lcall_$wnnz3_bufchan_d[0]) || lizzieLet35_3Lcall_$wnnz3_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet35_3Lcall_$wnnz3_bufchan_d <= 1'd0;
    else
      if (lizzieLet35_3Lcall_$wnnz3_r)
        lizzieLet35_3Lcall_$wnnz3_bufchan_d <= lizzieLet35_3Lcall_$wnnz3_d;
  Go_t lizzieLet35_3Lcall_$wnnz3_bufchan_buf;
  assign lizzieLet35_3Lcall_$wnnz3_bufchan_r = (! lizzieLet35_3Lcall_$wnnz3_bufchan_buf[0]);
  assign lizzieLet35_3Lcall_$wnnz3_1_argbuf_d = (lizzieLet35_3Lcall_$wnnz3_bufchan_buf[0] ? lizzieLet35_3Lcall_$wnnz3_bufchan_buf :
                                                 lizzieLet35_3Lcall_$wnnz3_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet35_3Lcall_$wnnz3_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet35_3Lcall_$wnnz3_1_argbuf_r && lizzieLet35_3Lcall_$wnnz3_bufchan_buf[0]))
        lizzieLet35_3Lcall_$wnnz3_bufchan_buf <= 1'd0;
      else if (((! lizzieLet35_3Lcall_$wnnz3_1_argbuf_r) && (! lizzieLet35_3Lcall_$wnnz3_bufchan_buf[0])))
        lizzieLet35_3Lcall_$wnnz3_bufchan_buf <= lizzieLet35_3Lcall_$wnnz3_bufchan_d;
  
  /* demux (Ty CT$wnnz,
       Ty Int#) : (lizzieLet35_4,CT$wnnz) (srtarg_0_goMux_mux,Int#) > [(lizzieLet35_4L$wnnzsbos,Int#),
                                                                       (lizzieLet35_4Lcall_$wnnz3,Int#),
                                                                       (lizzieLet35_4Lcall_$wnnz2,Int#),
                                                                       (lizzieLet35_4Lcall_$wnnz1,Int#),
                                                                       (lizzieLet35_4Lcall_$wnnz0,Int#)] */
  logic [4:0] srtarg_0_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet35_4_d[0] && srtarg_0_goMux_mux_d[0]))
      unique case (lizzieLet35_4_d[3:1])
        3'd0: srtarg_0_goMux_mux_onehotd = 5'd1;
        3'd1: srtarg_0_goMux_mux_onehotd = 5'd2;
        3'd2: srtarg_0_goMux_mux_onehotd = 5'd4;
        3'd3: srtarg_0_goMux_mux_onehotd = 5'd8;
        3'd4: srtarg_0_goMux_mux_onehotd = 5'd16;
        default: srtarg_0_goMux_mux_onehotd = 5'd0;
      endcase
    else srtarg_0_goMux_mux_onehotd = 5'd0;
  assign lizzieLet35_4L$wnnzsbos_d = {srtarg_0_goMux_mux_d[32:1],
                                      srtarg_0_goMux_mux_onehotd[0]};
  assign lizzieLet35_4Lcall_$wnnz3_d = {srtarg_0_goMux_mux_d[32:1],
                                        srtarg_0_goMux_mux_onehotd[1]};
  assign lizzieLet35_4Lcall_$wnnz2_d = {srtarg_0_goMux_mux_d[32:1],
                                        srtarg_0_goMux_mux_onehotd[2]};
  assign lizzieLet35_4Lcall_$wnnz1_d = {srtarg_0_goMux_mux_d[32:1],
                                        srtarg_0_goMux_mux_onehotd[3]};
  assign lizzieLet35_4Lcall_$wnnz0_d = {srtarg_0_goMux_mux_d[32:1],
                                        srtarg_0_goMux_mux_onehotd[4]};
  assign srtarg_0_goMux_mux_r = (| (srtarg_0_goMux_mux_onehotd & {lizzieLet35_4Lcall_$wnnz0_r,
                                                                  lizzieLet35_4Lcall_$wnnz1_r,
                                                                  lizzieLet35_4Lcall_$wnnz2_r,
                                                                  lizzieLet35_4Lcall_$wnnz3_r,
                                                                  lizzieLet35_4L$wnnzsbos_r}));
  assign lizzieLet35_4_r = srtarg_0_goMux_mux_r;
  
  /* fork (Ty Int#) : (lizzieLet35_4L$wnnzsbos,Int#) > [(lizzieLet35_4L$wnnzsbos_1_merge_merge_fork_1,Int#),
                                                   (lizzieLet35_4L$wnnzsbos_1_merge_merge_fork_2,Int#)] */
  logic [1:0] lizzieLet35_4L$wnnzsbos_emitted;
  logic [1:0] lizzieLet35_4L$wnnzsbos_done;
  assign lizzieLet35_4L$wnnzsbos_1_merge_merge_fork_1_d = {lizzieLet35_4L$wnnzsbos_d[32:1],
                                                           (lizzieLet35_4L$wnnzsbos_d[0] && (! lizzieLet35_4L$wnnzsbos_emitted[0]))};
  assign lizzieLet35_4L$wnnzsbos_1_merge_merge_fork_2_d = {lizzieLet35_4L$wnnzsbos_d[32:1],
                                                           (lizzieLet35_4L$wnnzsbos_d[0] && (! lizzieLet35_4L$wnnzsbos_emitted[1]))};
  assign lizzieLet35_4L$wnnzsbos_done = (lizzieLet35_4L$wnnzsbos_emitted | ({lizzieLet35_4L$wnnzsbos_1_merge_merge_fork_2_d[0],
                                                                             lizzieLet35_4L$wnnzsbos_1_merge_merge_fork_1_d[0]} & {lizzieLet35_4L$wnnzsbos_1_merge_merge_fork_2_r,
                                                                                                                                   lizzieLet35_4L$wnnzsbos_1_merge_merge_fork_1_r}));
  assign lizzieLet35_4L$wnnzsbos_r = (& lizzieLet35_4L$wnnzsbos_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet35_4L$wnnzsbos_emitted <= 2'd0;
    else
      lizzieLet35_4L$wnnzsbos_emitted <= (lizzieLet35_4L$wnnzsbos_r ? 2'd0 :
                                          lizzieLet35_4L$wnnzsbos_done);
  
  /* togo (Ty Int#) : (lizzieLet35_4L$wnnzsbos_1_merge_merge_fork_1,Int#) > (call_$wnnz_goConst,Go) */
  assign call_$wnnz_goConst_d = lizzieLet35_4L$wnnzsbos_1_merge_merge_fork_1_d[0];
  assign lizzieLet35_4L$wnnzsbos_1_merge_merge_fork_1_r = call_$wnnz_goConst_r;
  
  /* buf (Ty Int#) : (lizzieLet35_4L$wnnzsbos_1_merge_merge_fork_2,Int#) > ($wnnz_resbuf,Int#) */
  \Int#_t  lizzieLet35_4L$wnnzsbos_1_merge_merge_fork_2_bufchan_d;
  logic lizzieLet35_4L$wnnzsbos_1_merge_merge_fork_2_bufchan_r;
  assign lizzieLet35_4L$wnnzsbos_1_merge_merge_fork_2_r = ((! lizzieLet35_4L$wnnzsbos_1_merge_merge_fork_2_bufchan_d[0]) || lizzieLet35_4L$wnnzsbos_1_merge_merge_fork_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet35_4L$wnnzsbos_1_merge_merge_fork_2_bufchan_d <= {32'd0,
                                                                 1'd0};
    else
      if (lizzieLet35_4L$wnnzsbos_1_merge_merge_fork_2_r)
        lizzieLet35_4L$wnnzsbos_1_merge_merge_fork_2_bufchan_d <= lizzieLet35_4L$wnnzsbos_1_merge_merge_fork_2_d;
  \Int#_t  lizzieLet35_4L$wnnzsbos_1_merge_merge_fork_2_bufchan_buf;
  assign lizzieLet35_4L$wnnzsbos_1_merge_merge_fork_2_bufchan_r = (! lizzieLet35_4L$wnnzsbos_1_merge_merge_fork_2_bufchan_buf[0]);
  assign \$wnnz_resbuf_d  = (lizzieLet35_4L$wnnzsbos_1_merge_merge_fork_2_bufchan_buf[0] ? lizzieLet35_4L$wnnzsbos_1_merge_merge_fork_2_bufchan_buf :
                             lizzieLet35_4L$wnnzsbos_1_merge_merge_fork_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet35_4L$wnnzsbos_1_merge_merge_fork_2_bufchan_buf <= {32'd0,
                                                                   1'd0};
    else
      if ((\$wnnz_resbuf_r  && lizzieLet35_4L$wnnzsbos_1_merge_merge_fork_2_bufchan_buf[0]))
        lizzieLet35_4L$wnnzsbos_1_merge_merge_fork_2_bufchan_buf <= {32'd0,
                                                                     1'd0};
      else if (((! \$wnnz_resbuf_r ) && (! lizzieLet35_4L$wnnzsbos_1_merge_merge_fork_2_bufchan_buf[0])))
        lizzieLet35_4L$wnnzsbos_1_merge_merge_fork_2_bufchan_buf <= lizzieLet35_4L$wnnzsbos_1_merge_merge_fork_2_bufchan_d;
  
  /* dcon (Ty CT$wnnz,
      Dcon Lcall_$wnnz2) : [(lizzieLet35_4Lcall_$wnnz3,Int#),
                            (sc_0_3_destruct,Pointer_CT$wnnz),
                            (q4a87_1_destruct,Pointer_QTree_Int),
                            (q3a86_1_destruct,Pointer_QTree_Int)] > (lizzieLet35_4Lcall_$wnnz3_1sc_0_3_1q4a87_1_1q3a86_1_1Lcall_$wnnz2,CT$wnnz) */
  assign lizzieLet35_4Lcall_$wnnz3_1sc_0_3_1q4a87_1_1q3a86_1_1Lcall_$wnnz2_d = Lcall_$wnnz2_dc((& {lizzieLet35_4Lcall_$wnnz3_d[0],
                                                                                                   sc_0_3_destruct_d[0],
                                                                                                   q4a87_1_destruct_d[0],
                                                                                                   q3a86_1_destruct_d[0]}), lizzieLet35_4Lcall_$wnnz3_d, sc_0_3_destruct_d, q4a87_1_destruct_d, q3a86_1_destruct_d);
  assign {lizzieLet35_4Lcall_$wnnz3_r,
          sc_0_3_destruct_r,
          q4a87_1_destruct_r,
          q3a86_1_destruct_r} = {4 {(lizzieLet35_4Lcall_$wnnz3_1sc_0_3_1q4a87_1_1q3a86_1_1Lcall_$wnnz2_r && lizzieLet35_4Lcall_$wnnz3_1sc_0_3_1q4a87_1_1q3a86_1_1Lcall_$wnnz2_d[0])}};
  
  /* buf (Ty CT$wnnz) : (lizzieLet35_4Lcall_$wnnz3_1sc_0_3_1q4a87_1_1q3a86_1_1Lcall_$wnnz2,CT$wnnz) > (lizzieLet36_1_argbuf,CT$wnnz) */
  CT$wnnz_t lizzieLet35_4Lcall_$wnnz3_1sc_0_3_1q4a87_1_1q3a86_1_1Lcall_$wnnz2_bufchan_d;
  logic lizzieLet35_4Lcall_$wnnz3_1sc_0_3_1q4a87_1_1q3a86_1_1Lcall_$wnnz2_bufchan_r;
  assign lizzieLet35_4Lcall_$wnnz3_1sc_0_3_1q4a87_1_1q3a86_1_1Lcall_$wnnz2_r = ((! lizzieLet35_4Lcall_$wnnz3_1sc_0_3_1q4a87_1_1q3a86_1_1Lcall_$wnnz2_bufchan_d[0]) || lizzieLet35_4Lcall_$wnnz3_1sc_0_3_1q4a87_1_1q3a86_1_1Lcall_$wnnz2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet35_4Lcall_$wnnz3_1sc_0_3_1q4a87_1_1q3a86_1_1Lcall_$wnnz2_bufchan_d <= {115'd0,
                                                                                      1'd0};
    else
      if (lizzieLet35_4Lcall_$wnnz3_1sc_0_3_1q4a87_1_1q3a86_1_1Lcall_$wnnz2_r)
        lizzieLet35_4Lcall_$wnnz3_1sc_0_3_1q4a87_1_1q3a86_1_1Lcall_$wnnz2_bufchan_d <= lizzieLet35_4Lcall_$wnnz3_1sc_0_3_1q4a87_1_1q3a86_1_1Lcall_$wnnz2_d;
  CT$wnnz_t lizzieLet35_4Lcall_$wnnz3_1sc_0_3_1q4a87_1_1q3a86_1_1Lcall_$wnnz2_bufchan_buf;
  assign lizzieLet35_4Lcall_$wnnz3_1sc_0_3_1q4a87_1_1q3a86_1_1Lcall_$wnnz2_bufchan_r = (! lizzieLet35_4Lcall_$wnnz3_1sc_0_3_1q4a87_1_1q3a86_1_1Lcall_$wnnz2_bufchan_buf[0]);
  assign lizzieLet36_1_argbuf_d = (lizzieLet35_4Lcall_$wnnz3_1sc_0_3_1q4a87_1_1q3a86_1_1Lcall_$wnnz2_bufchan_buf[0] ? lizzieLet35_4Lcall_$wnnz3_1sc_0_3_1q4a87_1_1q3a86_1_1Lcall_$wnnz2_bufchan_buf :
                                   lizzieLet35_4Lcall_$wnnz3_1sc_0_3_1q4a87_1_1q3a86_1_1Lcall_$wnnz2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet35_4Lcall_$wnnz3_1sc_0_3_1q4a87_1_1q3a86_1_1Lcall_$wnnz2_bufchan_buf <= {115'd0,
                                                                                        1'd0};
    else
      if ((lizzieLet36_1_argbuf_r && lizzieLet35_4Lcall_$wnnz3_1sc_0_3_1q4a87_1_1q3a86_1_1Lcall_$wnnz2_bufchan_buf[0]))
        lizzieLet35_4Lcall_$wnnz3_1sc_0_3_1q4a87_1_1q3a86_1_1Lcall_$wnnz2_bufchan_buf <= {115'd0,
                                                                                          1'd0};
      else if (((! lizzieLet36_1_argbuf_r) && (! lizzieLet35_4Lcall_$wnnz3_1sc_0_3_1q4a87_1_1q3a86_1_1Lcall_$wnnz2_bufchan_buf[0])))
        lizzieLet35_4Lcall_$wnnz3_1sc_0_3_1q4a87_1_1q3a86_1_1Lcall_$wnnz2_bufchan_buf <= lizzieLet35_4Lcall_$wnnz3_1sc_0_3_1q4a87_1_1q3a86_1_1Lcall_$wnnz2_bufchan_d;
  
  /* destruct (Ty CTf''''''''_f''''''''_Int_Int,
          Dcon Lcall_f''''''''_f''''''''_Int_Int0) : (lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int0,CTf''''''''_f''''''''_Int_Int) > [(es_5_2_destruct,Pointer_QTree_Int),
                                                                                                                                        (es_6_4_destruct,Pointer_QTree_Int),
                                                                                                                                        (es_7_4_destruct,Pointer_QTree_Int),
                                                                                                                                        (sc_0_10_destruct,Pointer_CTf''''''''_f''''''''_Int_Int)] */
  logic [3:0] \lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int0_emitted ;
  logic [3:0] \lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int0_done ;
  assign es_5_2_destruct_d = {\lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int0_d [19:4],
                              (\lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int0_d [0] && (! \lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int0_emitted [0]))};
  assign es_6_4_destruct_d = {\lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int0_d [35:20],
                              (\lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int0_d [0] && (! \lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int0_emitted [1]))};
  assign es_7_4_destruct_d = {\lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int0_d [51:36],
                              (\lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int0_d [0] && (! \lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int0_emitted [2]))};
  assign sc_0_10_destruct_d = {\lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int0_d [67:52],
                               (\lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int0_d [0] && (! \lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int0_emitted [3]))};
  assign \lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int0_done  = (\lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int0_emitted  | ({sc_0_10_destruct_d[0],
                                                                                                                                 es_7_4_destruct_d[0],
                                                                                                                                 es_6_4_destruct_d[0],
                                                                                                                                 es_5_2_destruct_d[0]} & {sc_0_10_destruct_r,
                                                                                                                                                          es_7_4_destruct_r,
                                                                                                                                                          es_6_4_destruct_r,
                                                                                                                                                          es_5_2_destruct_r}));
  assign \lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int0_r  = (& \lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int0_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int0_emitted  <= 4'd0;
    else
      \lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int0_emitted  <= (\lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int0_r  ? 4'd0 :
                                                                    \lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int0_done );
  
  /* destruct (Ty CTf''''''''_f''''''''_Int_Int,
          Dcon Lcall_f''''''''_f''''''''_Int_Int1) : (lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int1,CTf''''''''_f''''''''_Int_Int) > [(es_6_3_destruct,Pointer_QTree_Int),
                                                                                                                                        (es_7_3_destruct,Pointer_QTree_Int),
                                                                                                                                        (sc_0_9_destruct,Pointer_CTf''''''''_f''''''''_Int_Int),
                                                                                                                                        (tla8y_3_destruct,Pointer_QTree_Int),
                                                                                                                                        (is_z_mapa8v_4_destruct,MyDTInt_Bool),
                                                                                                                                        (op_mapa8w_4_destruct,MyDTInt_Int)] */
  logic [5:0] \lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int1_emitted ;
  logic [5:0] \lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int1_done ;
  assign es_6_3_destruct_d = {\lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int1_d [19:4],
                              (\lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int1_d [0] && (! \lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int1_emitted [0]))};
  assign es_7_3_destruct_d = {\lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int1_d [35:20],
                              (\lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int1_d [0] && (! \lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int1_emitted [1]))};
  assign sc_0_9_destruct_d = {\lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int1_d [51:36],
                              (\lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int1_d [0] && (! \lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int1_emitted [2]))};
  assign tla8y_3_destruct_d = {\lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int1_d [67:52],
                               (\lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int1_d [0] && (! \lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int1_emitted [3]))};
  assign is_z_mapa8v_4_destruct_d = (\lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int1_d [0] && (! \lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int1_emitted [4]));
  assign op_mapa8w_4_destruct_d = (\lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int1_d [0] && (! \lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int1_emitted [5]));
  assign \lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int1_done  = (\lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int1_emitted  | ({op_mapa8w_4_destruct_d[0],
                                                                                                                                 is_z_mapa8v_4_destruct_d[0],
                                                                                                                                 tla8y_3_destruct_d[0],
                                                                                                                                 sc_0_9_destruct_d[0],
                                                                                                                                 es_7_3_destruct_d[0],
                                                                                                                                 es_6_3_destruct_d[0]} & {op_mapa8w_4_destruct_r,
                                                                                                                                                          is_z_mapa8v_4_destruct_r,
                                                                                                                                                          tla8y_3_destruct_r,
                                                                                                                                                          sc_0_9_destruct_r,
                                                                                                                                                          es_7_3_destruct_r,
                                                                                                                                                          es_6_3_destruct_r}));
  assign \lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int1_r  = (& \lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int1_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int1_emitted  <= 6'd0;
    else
      \lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int1_emitted  <= (\lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int1_r  ? 6'd0 :
                                                                    \lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int1_done );
  
  /* destruct (Ty CTf''''''''_f''''''''_Int_Int,
          Dcon Lcall_f''''''''_f''''''''_Int_Int2) : (lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int2,CTf''''''''_f''''''''_Int_Int) > [(es_7_2_destruct,Pointer_QTree_Int),
                                                                                                                                        (sc_0_8_destruct,Pointer_CTf''''''''_f''''''''_Int_Int),
                                                                                                                                        (tla8y_2_destruct,Pointer_QTree_Int),
                                                                                                                                        (is_z_mapa8v_3_destruct,MyDTInt_Bool),
                                                                                                                                        (op_mapa8w_3_destruct,MyDTInt_Int),
                                                                                                                                        (tra8z_2_destruct,Pointer_QTree_Int)] */
  logic [5:0] \lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int2_emitted ;
  logic [5:0] \lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int2_done ;
  assign es_7_2_destruct_d = {\lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int2_d [19:4],
                              (\lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int2_d [0] && (! \lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int2_emitted [0]))};
  assign sc_0_8_destruct_d = {\lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int2_d [35:20],
                              (\lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int2_d [0] && (! \lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int2_emitted [1]))};
  assign tla8y_2_destruct_d = {\lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int2_d [51:36],
                               (\lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int2_d [0] && (! \lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int2_emitted [2]))};
  assign is_z_mapa8v_3_destruct_d = (\lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int2_d [0] && (! \lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int2_emitted [3]));
  assign op_mapa8w_3_destruct_d = (\lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int2_d [0] && (! \lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int2_emitted [4]));
  assign tra8z_2_destruct_d = {\lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int2_d [67:52],
                               (\lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int2_d [0] && (! \lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int2_emitted [5]))};
  assign \lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int2_done  = (\lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int2_emitted  | ({tra8z_2_destruct_d[0],
                                                                                                                                 op_mapa8w_3_destruct_d[0],
                                                                                                                                 is_z_mapa8v_3_destruct_d[0],
                                                                                                                                 tla8y_2_destruct_d[0],
                                                                                                                                 sc_0_8_destruct_d[0],
                                                                                                                                 es_7_2_destruct_d[0]} & {tra8z_2_destruct_r,
                                                                                                                                                          op_mapa8w_3_destruct_r,
                                                                                                                                                          is_z_mapa8v_3_destruct_r,
                                                                                                                                                          tla8y_2_destruct_r,
                                                                                                                                                          sc_0_8_destruct_r,
                                                                                                                                                          es_7_2_destruct_r}));
  assign \lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int2_r  = (& \lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int2_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int2_emitted  <= 6'd0;
    else
      \lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int2_emitted  <= (\lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int2_r  ? 6'd0 :
                                                                    \lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int2_done );
  
  /* destruct (Ty CTf''''''''_f''''''''_Int_Int,
          Dcon Lcall_f''''''''_f''''''''_Int_Int3) : (lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int3,CTf''''''''_f''''''''_Int_Int) > [(sc_0_7_destruct,Pointer_CTf''''''''_f''''''''_Int_Int),
                                                                                                                                        (tla8y_1_destruct,Pointer_QTree_Int),
                                                                                                                                        (is_z_mapa8v_2_destruct,MyDTInt_Bool),
                                                                                                                                        (op_mapa8w_2_destruct,MyDTInt_Int),
                                                                                                                                        (tra8z_1_destruct,Pointer_QTree_Int),
                                                                                                                                        (bla8A_1_destruct,Pointer_QTree_Int)] */
  logic [5:0] \lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int3_emitted ;
  logic [5:0] \lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int3_done ;
  assign sc_0_7_destruct_d = {\lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int3_d [19:4],
                              (\lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int3_d [0] && (! \lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int3_emitted [0]))};
  assign tla8y_1_destruct_d = {\lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int3_d [35:20],
                               (\lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int3_d [0] && (! \lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int3_emitted [1]))};
  assign is_z_mapa8v_2_destruct_d = (\lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int3_d [0] && (! \lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int3_emitted [2]));
  assign op_mapa8w_2_destruct_d = (\lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int3_d [0] && (! \lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int3_emitted [3]));
  assign tra8z_1_destruct_d = {\lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int3_d [51:36],
                               (\lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int3_d [0] && (! \lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int3_emitted [4]))};
  assign bla8A_1_destruct_d = {\lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int3_d [67:52],
                               (\lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int3_d [0] && (! \lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int3_emitted [5]))};
  assign \lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int3_done  = (\lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int3_emitted  | ({bla8A_1_destruct_d[0],
                                                                                                                                 tra8z_1_destruct_d[0],
                                                                                                                                 op_mapa8w_2_destruct_d[0],
                                                                                                                                 is_z_mapa8v_2_destruct_d[0],
                                                                                                                                 tla8y_1_destruct_d[0],
                                                                                                                                 sc_0_7_destruct_d[0]} & {bla8A_1_destruct_r,
                                                                                                                                                          tra8z_1_destruct_r,
                                                                                                                                                          op_mapa8w_2_destruct_r,
                                                                                                                                                          is_z_mapa8v_2_destruct_r,
                                                                                                                                                          tla8y_1_destruct_r,
                                                                                                                                                          sc_0_7_destruct_r}));
  assign \lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int3_r  = (& \lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int3_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int3_emitted  <= 6'd0;
    else
      \lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int3_emitted  <= (\lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int3_r  ? 6'd0 :
                                                                    \lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int3_done );
  
  /* demux (Ty CTf''''''''_f''''''''_Int_Int,
       Ty CTf''''''''_f''''''''_Int_Int) : (lizzieLet39_2,CTf''''''''_f''''''''_Int_Int) (lizzieLet39_1,CTf''''''''_f''''''''_Int_Int) > [(_12,CTf''''''''_f''''''''_Int_Int),
                                                                                                                                          (lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int3,CTf''''''''_f''''''''_Int_Int),
                                                                                                                                          (lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int2,CTf''''''''_f''''''''_Int_Int),
                                                                                                                                          (lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int1,CTf''''''''_f''''''''_Int_Int),
                                                                                                                                          (lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int0,CTf''''''''_f''''''''_Int_Int)] */
  logic [4:0] lizzieLet39_1_onehotd;
  always_comb
    if ((lizzieLet39_2_d[0] && lizzieLet39_1_d[0]))
      unique case (lizzieLet39_2_d[3:1])
        3'd0: lizzieLet39_1_onehotd = 5'd1;
        3'd1: lizzieLet39_1_onehotd = 5'd2;
        3'd2: lizzieLet39_1_onehotd = 5'd4;
        3'd3: lizzieLet39_1_onehotd = 5'd8;
        3'd4: lizzieLet39_1_onehotd = 5'd16;
        default: lizzieLet39_1_onehotd = 5'd0;
      endcase
    else lizzieLet39_1_onehotd = 5'd0;
  assign _12_d = {lizzieLet39_1_d[67:1], lizzieLet39_1_onehotd[0]};
  assign \lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int3_d  = {lizzieLet39_1_d[67:1],
                                                                lizzieLet39_1_onehotd[1]};
  assign \lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int2_d  = {lizzieLet39_1_d[67:1],
                                                                lizzieLet39_1_onehotd[2]};
  assign \lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int1_d  = {lizzieLet39_1_d[67:1],
                                                                lizzieLet39_1_onehotd[3]};
  assign \lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int0_d  = {lizzieLet39_1_d[67:1],
                                                                lizzieLet39_1_onehotd[4]};
  assign lizzieLet39_1_r = (| (lizzieLet39_1_onehotd & {\lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int0_r ,
                                                        \lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int1_r ,
                                                        \lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int2_r ,
                                                        \lizzieLet39_1Lcall_f''''''''_f''''''''_Int_Int3_r ,
                                                        _12_r}));
  assign lizzieLet39_2_r = lizzieLet39_1_r;
  
  /* demux (Ty CTf''''''''_f''''''''_Int_Int,
       Ty Go) : (lizzieLet39_3,CTf''''''''_f''''''''_Int_Int) (go_16_goMux_data,Go) > [(_11,Go),
                                                                                       (lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int3,Go),
                                                                                       (lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int2,Go),
                                                                                       (lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int1,Go),
                                                                                       (lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int0,Go)] */
  logic [4:0] go_16_goMux_data_onehotd;
  always_comb
    if ((lizzieLet39_3_d[0] && go_16_goMux_data_d[0]))
      unique case (lizzieLet39_3_d[3:1])
        3'd0: go_16_goMux_data_onehotd = 5'd1;
        3'd1: go_16_goMux_data_onehotd = 5'd2;
        3'd2: go_16_goMux_data_onehotd = 5'd4;
        3'd3: go_16_goMux_data_onehotd = 5'd8;
        3'd4: go_16_goMux_data_onehotd = 5'd16;
        default: go_16_goMux_data_onehotd = 5'd0;
      endcase
    else go_16_goMux_data_onehotd = 5'd0;
  assign _11_d = go_16_goMux_data_onehotd[0];
  assign \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int3_d  = go_16_goMux_data_onehotd[1];
  assign \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int2_d  = go_16_goMux_data_onehotd[2];
  assign \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int1_d  = go_16_goMux_data_onehotd[3];
  assign \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int0_d  = go_16_goMux_data_onehotd[4];
  assign go_16_goMux_data_r = (| (go_16_goMux_data_onehotd & {\lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int0_r ,
                                                              \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int1_r ,
                                                              \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int2_r ,
                                                              \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int3_r ,
                                                              _11_r}));
  assign lizzieLet39_3_r = go_16_goMux_data_r;
  
  /* buf (Ty Go) : (lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int0,Go) > (lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int0_1_argbuf,Go) */
  Go_t \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int0_bufchan_d ;
  logic \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int0_bufchan_r ;
  assign \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int0_r  = ((! \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int0_bufchan_d [0]) || \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int0_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int0_bufchan_d  <= 1'd0;
    else
      if (\lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int0_r )
        \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int0_bufchan_d  <= \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int0_d ;
  Go_t \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int0_bufchan_buf ;
  assign \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int0_bufchan_r  = (! \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int0_bufchan_buf [0]);
  assign \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int0_1_argbuf_d  = (\lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int0_bufchan_buf [0] ? \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int0_bufchan_buf  :
                                                                         \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int0_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int0_bufchan_buf  <= 1'd0;
    else
      if ((\lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int0_1_argbuf_r  && \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int0_bufchan_buf [0]))
        \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int0_bufchan_buf  <= 1'd0;
      else if (((! \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int0_1_argbuf_r ) && (! \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int0_bufchan_buf [0])))
        \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int0_bufchan_buf  <= \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int0_bufchan_d ;
  
  /* buf (Ty Go) : (lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int1,Go) > (lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int1_1_argbuf,Go) */
  Go_t \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int1_bufchan_d ;
  logic \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int1_bufchan_r ;
  assign \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int1_r  = ((! \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int1_bufchan_d [0]) || \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int1_bufchan_d  <= 1'd0;
    else
      if (\lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int1_r )
        \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int1_bufchan_d  <= \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int1_d ;
  Go_t \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int1_bufchan_buf ;
  assign \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int1_bufchan_r  = (! \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int1_bufchan_buf [0]);
  assign \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int1_1_argbuf_d  = (\lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int1_bufchan_buf [0] ? \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int1_bufchan_buf  :
                                                                         \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int1_bufchan_buf  <= 1'd0;
    else
      if ((\lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int1_1_argbuf_r  && \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int1_bufchan_buf [0]))
        \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int1_bufchan_buf  <= 1'd0;
      else if (((! \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int1_1_argbuf_r ) && (! \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int1_bufchan_buf [0])))
        \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int1_bufchan_buf  <= \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int1_bufchan_d ;
  
  /* buf (Ty Go) : (lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int2,Go) > (lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int2_1_argbuf,Go) */
  Go_t \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int2_bufchan_d ;
  logic \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int2_bufchan_r ;
  assign \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int2_r  = ((! \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int2_bufchan_d [0]) || \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int2_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int2_bufchan_d  <= 1'd0;
    else
      if (\lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int2_r )
        \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int2_bufchan_d  <= \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int2_d ;
  Go_t \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int2_bufchan_buf ;
  assign \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int2_bufchan_r  = (! \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int2_bufchan_buf [0]);
  assign \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int2_1_argbuf_d  = (\lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int2_bufchan_buf [0] ? \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int2_bufchan_buf  :
                                                                         \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int2_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int2_bufchan_buf  <= 1'd0;
    else
      if ((\lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int2_1_argbuf_r  && \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int2_bufchan_buf [0]))
        \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int2_bufchan_buf  <= 1'd0;
      else if (((! \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int2_1_argbuf_r ) && (! \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int2_bufchan_buf [0])))
        \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int2_bufchan_buf  <= \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int2_bufchan_d ;
  
  /* buf (Ty Go) : (lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int3,Go) > (lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int3_1_argbuf,Go) */
  Go_t \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int3_bufchan_d ;
  logic \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int3_bufchan_r ;
  assign \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int3_r  = ((! \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int3_bufchan_d [0]) || \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int3_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int3_bufchan_d  <= 1'd0;
    else
      if (\lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int3_r )
        \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int3_bufchan_d  <= \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int3_d ;
  Go_t \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int3_bufchan_buf ;
  assign \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int3_bufchan_r  = (! \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int3_bufchan_buf [0]);
  assign \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int3_1_argbuf_d  = (\lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int3_bufchan_buf [0] ? \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int3_bufchan_buf  :
                                                                         \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int3_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int3_bufchan_buf  <= 1'd0;
    else
      if ((\lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int3_1_argbuf_r  && \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int3_bufchan_buf [0]))
        \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int3_bufchan_buf  <= 1'd0;
      else if (((! \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int3_1_argbuf_r ) && (! \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int3_bufchan_buf [0])))
        \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int3_bufchan_buf  <= \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int3_bufchan_d ;
  
  /* demux (Ty CTf''''''''_f''''''''_Int_Int,
       Ty Pointer_QTree_Int) : (lizzieLet39_4,CTf''''''''_f''''''''_Int_Int) (srtarg_0_1_goMux_mux,Pointer_QTree_Int) > [(lizzieLet39_4Lf''''''''_f''''''''_Int_Intsbos,Pointer_QTree_Int),
                                                                                                                         (lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int3,Pointer_QTree_Int),
                                                                                                                         (lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int2,Pointer_QTree_Int),
                                                                                                                         (lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int1,Pointer_QTree_Int),
                                                                                                                         (lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int0,Pointer_QTree_Int)] */
  logic [4:0] srtarg_0_1_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet39_4_d[0] && srtarg_0_1_goMux_mux_d[0]))
      unique case (lizzieLet39_4_d[3:1])
        3'd0: srtarg_0_1_goMux_mux_onehotd = 5'd1;
        3'd1: srtarg_0_1_goMux_mux_onehotd = 5'd2;
        3'd2: srtarg_0_1_goMux_mux_onehotd = 5'd4;
        3'd3: srtarg_0_1_goMux_mux_onehotd = 5'd8;
        3'd4: srtarg_0_1_goMux_mux_onehotd = 5'd16;
        default: srtarg_0_1_goMux_mux_onehotd = 5'd0;
      endcase
    else srtarg_0_1_goMux_mux_onehotd = 5'd0;
  assign \lizzieLet39_4Lf''''''''_f''''''''_Int_Intsbos_d  = {srtarg_0_1_goMux_mux_d[16:1],
                                                              srtarg_0_1_goMux_mux_onehotd[0]};
  assign \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int3_d  = {srtarg_0_1_goMux_mux_d[16:1],
                                                                srtarg_0_1_goMux_mux_onehotd[1]};
  assign \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int2_d  = {srtarg_0_1_goMux_mux_d[16:1],
                                                                srtarg_0_1_goMux_mux_onehotd[2]};
  assign \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int1_d  = {srtarg_0_1_goMux_mux_d[16:1],
                                                                srtarg_0_1_goMux_mux_onehotd[3]};
  assign \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int0_d  = {srtarg_0_1_goMux_mux_d[16:1],
                                                                srtarg_0_1_goMux_mux_onehotd[4]};
  assign srtarg_0_1_goMux_mux_r = (| (srtarg_0_1_goMux_mux_onehotd & {\lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int0_r ,
                                                                      \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int1_r ,
                                                                      \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int2_r ,
                                                                      \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int3_r ,
                                                                      \lizzieLet39_4Lf''''''''_f''''''''_Int_Intsbos_r }));
  assign lizzieLet39_4_r = srtarg_0_1_goMux_mux_r;
  
  /* dcon (Ty QTree_Int,
      Dcon QNode_Int) : [(lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int0,Pointer_QTree_Int),
                         (es_5_2_destruct,Pointer_QTree_Int),
                         (es_6_4_destruct,Pointer_QTree_Int),
                         (es_7_4_destruct,Pointer_QTree_Int)] > (lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int0_1es_5_2_1es_6_4_1es_7_4_1QNode_Int,QTree_Int) */
  assign \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int0_1es_5_2_1es_6_4_1es_7_4_1QNode_Int_d  = QNode_Int_dc((& {\lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int0_d [0],
                                                                                                                   es_5_2_destruct_d[0],
                                                                                                                   es_6_4_destruct_d[0],
                                                                                                                   es_7_4_destruct_d[0]}), \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int0_d , es_5_2_destruct_d, es_6_4_destruct_d, es_7_4_destruct_d);
  assign {\lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int0_r ,
          es_5_2_destruct_r,
          es_6_4_destruct_r,
          es_7_4_destruct_r} = {4 {(\lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int0_1es_5_2_1es_6_4_1es_7_4_1QNode_Int_r  && \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int0_1es_5_2_1es_6_4_1es_7_4_1QNode_Int_d [0])}};
  
  /* buf (Ty QTree_Int) : (lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int0_1es_5_2_1es_6_4_1es_7_4_1QNode_Int,QTree_Int) > (lizzieLet43_1_argbuf,QTree_Int) */
  QTree_Int_t \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int0_1es_5_2_1es_6_4_1es_7_4_1QNode_Int_bufchan_d ;
  logic \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int0_1es_5_2_1es_6_4_1es_7_4_1QNode_Int_bufchan_r ;
  assign \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int0_1es_5_2_1es_6_4_1es_7_4_1QNode_Int_r  = ((! \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int0_1es_5_2_1es_6_4_1es_7_4_1QNode_Int_bufchan_d [0]) || \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int0_1es_5_2_1es_6_4_1es_7_4_1QNode_Int_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int0_1es_5_2_1es_6_4_1es_7_4_1QNode_Int_bufchan_d  <= {66'd0,
                                                                                                         1'd0};
    else
      if (\lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int0_1es_5_2_1es_6_4_1es_7_4_1QNode_Int_r )
        \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int0_1es_5_2_1es_6_4_1es_7_4_1QNode_Int_bufchan_d  <= \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int0_1es_5_2_1es_6_4_1es_7_4_1QNode_Int_d ;
  QTree_Int_t \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int0_1es_5_2_1es_6_4_1es_7_4_1QNode_Int_bufchan_buf ;
  assign \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int0_1es_5_2_1es_6_4_1es_7_4_1QNode_Int_bufchan_r  = (! \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int0_1es_5_2_1es_6_4_1es_7_4_1QNode_Int_bufchan_buf [0]);
  assign lizzieLet43_1_argbuf_d = (\lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int0_1es_5_2_1es_6_4_1es_7_4_1QNode_Int_bufchan_buf [0] ? \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int0_1es_5_2_1es_6_4_1es_7_4_1QNode_Int_bufchan_buf  :
                                   \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int0_1es_5_2_1es_6_4_1es_7_4_1QNode_Int_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int0_1es_5_2_1es_6_4_1es_7_4_1QNode_Int_bufchan_buf  <= {66'd0,
                                                                                                           1'd0};
    else
      if ((lizzieLet43_1_argbuf_r && \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int0_1es_5_2_1es_6_4_1es_7_4_1QNode_Int_bufchan_buf [0]))
        \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int0_1es_5_2_1es_6_4_1es_7_4_1QNode_Int_bufchan_buf  <= {66'd0,
                                                                                                             1'd0};
      else if (((! lizzieLet43_1_argbuf_r) && (! \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int0_1es_5_2_1es_6_4_1es_7_4_1QNode_Int_bufchan_buf [0])))
        \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int0_1es_5_2_1es_6_4_1es_7_4_1QNode_Int_bufchan_buf  <= \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int0_1es_5_2_1es_6_4_1es_7_4_1QNode_Int_bufchan_d ;
  
  /* dcon (Ty CTf''''''''_f''''''''_Int_Int,
      Dcon Lcall_f''''''''_f''''''''_Int_Int0) : [(lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int1,Pointer_QTree_Int),
                                                  (es_6_3_destruct,Pointer_QTree_Int),
                                                  (es_7_3_destruct,Pointer_QTree_Int),
                                                  (sc_0_9_destruct,Pointer_CTf''''''''_f''''''''_Int_Int)] > (lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int1_1es_6_3_1es_7_3_1sc_0_9_1Lcall_f''''''''_f''''''''_Int_Int0,CTf''''''''_f''''''''_Int_Int) */
  assign \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int1_1es_6_3_1es_7_3_1sc_0_9_1Lcall_f''''''''_f''''''''_Int_Int0_d  = \Lcall_f''''''''_f''''''''_Int_Int0_dc ((& {\lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int1_d [0],
                                                                                                                                                                       es_6_3_destruct_d[0],
                                                                                                                                                                       es_7_3_destruct_d[0],
                                                                                                                                                                       sc_0_9_destruct_d[0]}), \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int1_d , es_6_3_destruct_d, es_7_3_destruct_d, sc_0_9_destruct_d);
  assign {\lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int1_r ,
          es_6_3_destruct_r,
          es_7_3_destruct_r,
          sc_0_9_destruct_r} = {4 {(\lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int1_1es_6_3_1es_7_3_1sc_0_9_1Lcall_f''''''''_f''''''''_Int_Int0_r  && \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int1_1es_6_3_1es_7_3_1sc_0_9_1Lcall_f''''''''_f''''''''_Int_Int0_d [0])}};
  
  /* buf (Ty CTf''''''''_f''''''''_Int_Int) : (lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int1_1es_6_3_1es_7_3_1sc_0_9_1Lcall_f''''''''_f''''''''_Int_Int0,CTf''''''''_f''''''''_Int_Int) > (lizzieLet42_1_argbuf,CTf''''''''_f''''''''_Int_Int) */
  \CTf''''''''_f''''''''_Int_Int_t  \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int1_1es_6_3_1es_7_3_1sc_0_9_1Lcall_f''''''''_f''''''''_Int_Int0_bufchan_d ;
  logic \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int1_1es_6_3_1es_7_3_1sc_0_9_1Lcall_f''''''''_f''''''''_Int_Int0_bufchan_r ;
  assign \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int1_1es_6_3_1es_7_3_1sc_0_9_1Lcall_f''''''''_f''''''''_Int_Int0_r  = ((! \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int1_1es_6_3_1es_7_3_1sc_0_9_1Lcall_f''''''''_f''''''''_Int_Int0_bufchan_d [0]) || \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int1_1es_6_3_1es_7_3_1sc_0_9_1Lcall_f''''''''_f''''''''_Int_Int0_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int1_1es_6_3_1es_7_3_1sc_0_9_1Lcall_f''''''''_f''''''''_Int_Int0_bufchan_d  <= {67'd0,
                                                                                                                                  1'd0};
    else
      if (\lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int1_1es_6_3_1es_7_3_1sc_0_9_1Lcall_f''''''''_f''''''''_Int_Int0_r )
        \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int1_1es_6_3_1es_7_3_1sc_0_9_1Lcall_f''''''''_f''''''''_Int_Int0_bufchan_d  <= \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int1_1es_6_3_1es_7_3_1sc_0_9_1Lcall_f''''''''_f''''''''_Int_Int0_d ;
  \CTf''''''''_f''''''''_Int_Int_t  \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int1_1es_6_3_1es_7_3_1sc_0_9_1Lcall_f''''''''_f''''''''_Int_Int0_bufchan_buf ;
  assign \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int1_1es_6_3_1es_7_3_1sc_0_9_1Lcall_f''''''''_f''''''''_Int_Int0_bufchan_r  = (! \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int1_1es_6_3_1es_7_3_1sc_0_9_1Lcall_f''''''''_f''''''''_Int_Int0_bufchan_buf [0]);
  assign lizzieLet42_1_argbuf_d = (\lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int1_1es_6_3_1es_7_3_1sc_0_9_1Lcall_f''''''''_f''''''''_Int_Int0_bufchan_buf [0] ? \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int1_1es_6_3_1es_7_3_1sc_0_9_1Lcall_f''''''''_f''''''''_Int_Int0_bufchan_buf  :
                                   \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int1_1es_6_3_1es_7_3_1sc_0_9_1Lcall_f''''''''_f''''''''_Int_Int0_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int1_1es_6_3_1es_7_3_1sc_0_9_1Lcall_f''''''''_f''''''''_Int_Int0_bufchan_buf  <= {67'd0,
                                                                                                                                    1'd0};
    else
      if ((lizzieLet42_1_argbuf_r && \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int1_1es_6_3_1es_7_3_1sc_0_9_1Lcall_f''''''''_f''''''''_Int_Int0_bufchan_buf [0]))
        \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int1_1es_6_3_1es_7_3_1sc_0_9_1Lcall_f''''''''_f''''''''_Int_Int0_bufchan_buf  <= {67'd0,
                                                                                                                                      1'd0};
      else if (((! lizzieLet42_1_argbuf_r) && (! \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int1_1es_6_3_1es_7_3_1sc_0_9_1Lcall_f''''''''_f''''''''_Int_Int0_bufchan_buf [0])))
        \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int1_1es_6_3_1es_7_3_1sc_0_9_1Lcall_f''''''''_f''''''''_Int_Int0_bufchan_buf  <= \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int1_1es_6_3_1es_7_3_1sc_0_9_1Lcall_f''''''''_f''''''''_Int_Int0_bufchan_d ;
  
  /* dcon (Ty CTf''''''''_f''''''''_Int_Int,
      Dcon Lcall_f''''''''_f''''''''_Int_Int1) : [(lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int2,Pointer_QTree_Int),
                                                  (es_7_2_destruct,Pointer_QTree_Int),
                                                  (sc_0_8_destruct,Pointer_CTf''''''''_f''''''''_Int_Int),
                                                  (tla8y_2_destruct,Pointer_QTree_Int),
                                                  (is_z_mapa8v_3_1,MyDTInt_Bool),
                                                  (op_mapa8w_3_1,MyDTInt_Int)] > (lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int2_1es_7_2_1sc_0_8_1tla8y_2_1is_z_mapa8v_3_1op_mapa8w_3_1Lcall_f''''''''_f''''''''_Int_Int1,CTf''''''''_f''''''''_Int_Int) */
  assign \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int2_1es_7_2_1sc_0_8_1tla8y_2_1is_z_mapa8v_3_1op_mapa8w_3_1Lcall_f''''''''_f''''''''_Int_Int1_d  = \Lcall_f''''''''_f''''''''_Int_Int1_dc ((& {\lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int2_d [0],
                                                                                                                                                                                                    es_7_2_destruct_d[0],
                                                                                                                                                                                                    sc_0_8_destruct_d[0],
                                                                                                                                                                                                    tla8y_2_destruct_d[0],
                                                                                                                                                                                                    is_z_mapa8v_3_1_d[0],
                                                                                                                                                                                                    op_mapa8w_3_1_d[0]}), \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int2_d , es_7_2_destruct_d, sc_0_8_destruct_d, tla8y_2_destruct_d, is_z_mapa8v_3_1_d, op_mapa8w_3_1_d);
  assign {\lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int2_r ,
          es_7_2_destruct_r,
          sc_0_8_destruct_r,
          tla8y_2_destruct_r,
          is_z_mapa8v_3_1_r,
          op_mapa8w_3_1_r} = {6 {(\lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int2_1es_7_2_1sc_0_8_1tla8y_2_1is_z_mapa8v_3_1op_mapa8w_3_1Lcall_f''''''''_f''''''''_Int_Int1_r  && \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int2_1es_7_2_1sc_0_8_1tla8y_2_1is_z_mapa8v_3_1op_mapa8w_3_1Lcall_f''''''''_f''''''''_Int_Int1_d [0])}};
  
  /* buf (Ty CTf''''''''_f''''''''_Int_Int) : (lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int2_1es_7_2_1sc_0_8_1tla8y_2_1is_z_mapa8v_3_1op_mapa8w_3_1Lcall_f''''''''_f''''''''_Int_Int1,CTf''''''''_f''''''''_Int_Int) > (lizzieLet41_1_argbuf,CTf''''''''_f''''''''_Int_Int) */
  \CTf''''''''_f''''''''_Int_Int_t  \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int2_1es_7_2_1sc_0_8_1tla8y_2_1is_z_mapa8v_3_1op_mapa8w_3_1Lcall_f''''''''_f''''''''_Int_Int1_bufchan_d ;
  logic \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int2_1es_7_2_1sc_0_8_1tla8y_2_1is_z_mapa8v_3_1op_mapa8w_3_1Lcall_f''''''''_f''''''''_Int_Int1_bufchan_r ;
  assign \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int2_1es_7_2_1sc_0_8_1tla8y_2_1is_z_mapa8v_3_1op_mapa8w_3_1Lcall_f''''''''_f''''''''_Int_Int1_r  = ((! \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int2_1es_7_2_1sc_0_8_1tla8y_2_1is_z_mapa8v_3_1op_mapa8w_3_1Lcall_f''''''''_f''''''''_Int_Int1_bufchan_d [0]) || \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int2_1es_7_2_1sc_0_8_1tla8y_2_1is_z_mapa8v_3_1op_mapa8w_3_1Lcall_f''''''''_f''''''''_Int_Int1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int2_1es_7_2_1sc_0_8_1tla8y_2_1is_z_mapa8v_3_1op_mapa8w_3_1Lcall_f''''''''_f''''''''_Int_Int1_bufchan_d  <= {67'd0,
                                                                                                                                                               1'd0};
    else
      if (\lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int2_1es_7_2_1sc_0_8_1tla8y_2_1is_z_mapa8v_3_1op_mapa8w_3_1Lcall_f''''''''_f''''''''_Int_Int1_r )
        \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int2_1es_7_2_1sc_0_8_1tla8y_2_1is_z_mapa8v_3_1op_mapa8w_3_1Lcall_f''''''''_f''''''''_Int_Int1_bufchan_d  <= \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int2_1es_7_2_1sc_0_8_1tla8y_2_1is_z_mapa8v_3_1op_mapa8w_3_1Lcall_f''''''''_f''''''''_Int_Int1_d ;
  \CTf''''''''_f''''''''_Int_Int_t  \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int2_1es_7_2_1sc_0_8_1tla8y_2_1is_z_mapa8v_3_1op_mapa8w_3_1Lcall_f''''''''_f''''''''_Int_Int1_bufchan_buf ;
  assign \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int2_1es_7_2_1sc_0_8_1tla8y_2_1is_z_mapa8v_3_1op_mapa8w_3_1Lcall_f''''''''_f''''''''_Int_Int1_bufchan_r  = (! \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int2_1es_7_2_1sc_0_8_1tla8y_2_1is_z_mapa8v_3_1op_mapa8w_3_1Lcall_f''''''''_f''''''''_Int_Int1_bufchan_buf [0]);
  assign lizzieLet41_1_argbuf_d = (\lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int2_1es_7_2_1sc_0_8_1tla8y_2_1is_z_mapa8v_3_1op_mapa8w_3_1Lcall_f''''''''_f''''''''_Int_Int1_bufchan_buf [0] ? \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int2_1es_7_2_1sc_0_8_1tla8y_2_1is_z_mapa8v_3_1op_mapa8w_3_1Lcall_f''''''''_f''''''''_Int_Int1_bufchan_buf  :
                                   \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int2_1es_7_2_1sc_0_8_1tla8y_2_1is_z_mapa8v_3_1op_mapa8w_3_1Lcall_f''''''''_f''''''''_Int_Int1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int2_1es_7_2_1sc_0_8_1tla8y_2_1is_z_mapa8v_3_1op_mapa8w_3_1Lcall_f''''''''_f''''''''_Int_Int1_bufchan_buf  <= {67'd0,
                                                                                                                                                                 1'd0};
    else
      if ((lizzieLet41_1_argbuf_r && \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int2_1es_7_2_1sc_0_8_1tla8y_2_1is_z_mapa8v_3_1op_mapa8w_3_1Lcall_f''''''''_f''''''''_Int_Int1_bufchan_buf [0]))
        \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int2_1es_7_2_1sc_0_8_1tla8y_2_1is_z_mapa8v_3_1op_mapa8w_3_1Lcall_f''''''''_f''''''''_Int_Int1_bufchan_buf  <= {67'd0,
                                                                                                                                                                   1'd0};
      else if (((! lizzieLet41_1_argbuf_r) && (! \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int2_1es_7_2_1sc_0_8_1tla8y_2_1is_z_mapa8v_3_1op_mapa8w_3_1Lcall_f''''''''_f''''''''_Int_Int1_bufchan_buf [0])))
        \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int2_1es_7_2_1sc_0_8_1tla8y_2_1is_z_mapa8v_3_1op_mapa8w_3_1Lcall_f''''''''_f''''''''_Int_Int1_bufchan_buf  <= \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int2_1es_7_2_1sc_0_8_1tla8y_2_1is_z_mapa8v_3_1op_mapa8w_3_1Lcall_f''''''''_f''''''''_Int_Int1_bufchan_d ;
  
  /* dcon (Ty CTf''''''''_f''''''''_Int_Int,
      Dcon Lcall_f''''''''_f''''''''_Int_Int2) : [(lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int3,Pointer_QTree_Int),
                                                  (sc_0_7_destruct,Pointer_CTf''''''''_f''''''''_Int_Int),
                                                  (tla8y_1_destruct,Pointer_QTree_Int),
                                                  (is_z_mapa8v_2_1,MyDTInt_Bool),
                                                  (op_mapa8w_2_1,MyDTInt_Int),
                                                  (tra8z_1_destruct,Pointer_QTree_Int)] > (lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int3_1sc_0_7_1tla8y_1_1is_z_mapa8v_2_1op_mapa8w_2_1tra8z_1_1Lcall_f''''''''_f''''''''_Int_Int2,CTf''''''''_f''''''''_Int_Int) */
  assign \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int3_1sc_0_7_1tla8y_1_1is_z_mapa8v_2_1op_mapa8w_2_1tra8z_1_1Lcall_f''''''''_f''''''''_Int_Int2_d  = \Lcall_f''''''''_f''''''''_Int_Int2_dc ((& {\lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int3_d [0],
                                                                                                                                                                                                     sc_0_7_destruct_d[0],
                                                                                                                                                                                                     tla8y_1_destruct_d[0],
                                                                                                                                                                                                     is_z_mapa8v_2_1_d[0],
                                                                                                                                                                                                     op_mapa8w_2_1_d[0],
                                                                                                                                                                                                     tra8z_1_destruct_d[0]}), \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int3_d , sc_0_7_destruct_d, tla8y_1_destruct_d, is_z_mapa8v_2_1_d, op_mapa8w_2_1_d, tra8z_1_destruct_d);
  assign {\lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int3_r ,
          sc_0_7_destruct_r,
          tla8y_1_destruct_r,
          is_z_mapa8v_2_1_r,
          op_mapa8w_2_1_r,
          tra8z_1_destruct_r} = {6 {(\lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int3_1sc_0_7_1tla8y_1_1is_z_mapa8v_2_1op_mapa8w_2_1tra8z_1_1Lcall_f''''''''_f''''''''_Int_Int2_r  && \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int3_1sc_0_7_1tla8y_1_1is_z_mapa8v_2_1op_mapa8w_2_1tra8z_1_1Lcall_f''''''''_f''''''''_Int_Int2_d [0])}};
  
  /* buf (Ty CTf''''''''_f''''''''_Int_Int) : (lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int3_1sc_0_7_1tla8y_1_1is_z_mapa8v_2_1op_mapa8w_2_1tra8z_1_1Lcall_f''''''''_f''''''''_Int_Int2,CTf''''''''_f''''''''_Int_Int) > (lizzieLet40_1_argbuf,CTf''''''''_f''''''''_Int_Int) */
  \CTf''''''''_f''''''''_Int_Int_t  \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int3_1sc_0_7_1tla8y_1_1is_z_mapa8v_2_1op_mapa8w_2_1tra8z_1_1Lcall_f''''''''_f''''''''_Int_Int2_bufchan_d ;
  logic \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int3_1sc_0_7_1tla8y_1_1is_z_mapa8v_2_1op_mapa8w_2_1tra8z_1_1Lcall_f''''''''_f''''''''_Int_Int2_bufchan_r ;
  assign \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int3_1sc_0_7_1tla8y_1_1is_z_mapa8v_2_1op_mapa8w_2_1tra8z_1_1Lcall_f''''''''_f''''''''_Int_Int2_r  = ((! \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int3_1sc_0_7_1tla8y_1_1is_z_mapa8v_2_1op_mapa8w_2_1tra8z_1_1Lcall_f''''''''_f''''''''_Int_Int2_bufchan_d [0]) || \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int3_1sc_0_7_1tla8y_1_1is_z_mapa8v_2_1op_mapa8w_2_1tra8z_1_1Lcall_f''''''''_f''''''''_Int_Int2_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int3_1sc_0_7_1tla8y_1_1is_z_mapa8v_2_1op_mapa8w_2_1tra8z_1_1Lcall_f''''''''_f''''''''_Int_Int2_bufchan_d  <= {67'd0,
                                                                                                                                                                1'd0};
    else
      if (\lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int3_1sc_0_7_1tla8y_1_1is_z_mapa8v_2_1op_mapa8w_2_1tra8z_1_1Lcall_f''''''''_f''''''''_Int_Int2_r )
        \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int3_1sc_0_7_1tla8y_1_1is_z_mapa8v_2_1op_mapa8w_2_1tra8z_1_1Lcall_f''''''''_f''''''''_Int_Int2_bufchan_d  <= \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int3_1sc_0_7_1tla8y_1_1is_z_mapa8v_2_1op_mapa8w_2_1tra8z_1_1Lcall_f''''''''_f''''''''_Int_Int2_d ;
  \CTf''''''''_f''''''''_Int_Int_t  \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int3_1sc_0_7_1tla8y_1_1is_z_mapa8v_2_1op_mapa8w_2_1tra8z_1_1Lcall_f''''''''_f''''''''_Int_Int2_bufchan_buf ;
  assign \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int3_1sc_0_7_1tla8y_1_1is_z_mapa8v_2_1op_mapa8w_2_1tra8z_1_1Lcall_f''''''''_f''''''''_Int_Int2_bufchan_r  = (! \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int3_1sc_0_7_1tla8y_1_1is_z_mapa8v_2_1op_mapa8w_2_1tra8z_1_1Lcall_f''''''''_f''''''''_Int_Int2_bufchan_buf [0]);
  assign lizzieLet40_1_argbuf_d = (\lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int3_1sc_0_7_1tla8y_1_1is_z_mapa8v_2_1op_mapa8w_2_1tra8z_1_1Lcall_f''''''''_f''''''''_Int_Int2_bufchan_buf [0] ? \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int3_1sc_0_7_1tla8y_1_1is_z_mapa8v_2_1op_mapa8w_2_1tra8z_1_1Lcall_f''''''''_f''''''''_Int_Int2_bufchan_buf  :
                                   \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int3_1sc_0_7_1tla8y_1_1is_z_mapa8v_2_1op_mapa8w_2_1tra8z_1_1Lcall_f''''''''_f''''''''_Int_Int2_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int3_1sc_0_7_1tla8y_1_1is_z_mapa8v_2_1op_mapa8w_2_1tra8z_1_1Lcall_f''''''''_f''''''''_Int_Int2_bufchan_buf  <= {67'd0,
                                                                                                                                                                  1'd0};
    else
      if ((lizzieLet40_1_argbuf_r && \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int3_1sc_0_7_1tla8y_1_1is_z_mapa8v_2_1op_mapa8w_2_1tra8z_1_1Lcall_f''''''''_f''''''''_Int_Int2_bufchan_buf [0]))
        \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int3_1sc_0_7_1tla8y_1_1is_z_mapa8v_2_1op_mapa8w_2_1tra8z_1_1Lcall_f''''''''_f''''''''_Int_Int2_bufchan_buf  <= {67'd0,
                                                                                                                                                                    1'd0};
      else if (((! lizzieLet40_1_argbuf_r) && (! \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int3_1sc_0_7_1tla8y_1_1is_z_mapa8v_2_1op_mapa8w_2_1tra8z_1_1Lcall_f''''''''_f''''''''_Int_Int2_bufchan_buf [0])))
        \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int3_1sc_0_7_1tla8y_1_1is_z_mapa8v_2_1op_mapa8w_2_1tra8z_1_1Lcall_f''''''''_f''''''''_Int_Int2_bufchan_buf  <= \lizzieLet39_4Lcall_f''''''''_f''''''''_Int_Int3_1sc_0_7_1tla8y_1_1is_z_mapa8v_2_1op_mapa8w_2_1tra8z_1_1Lcall_f''''''''_f''''''''_Int_Int2_bufchan_d ;
  
  /* fork (Ty Pointer_QTree_Int) : (lizzieLet39_4Lf''''''''_f''''''''_Int_Intsbos,Pointer_QTree_Int) > [(lizzieLet39_4Lf''''''''_f''''''''_Int_Intsbos_1_merge_merge_fork_1,Pointer_QTree_Int),
                                                                                                   (lizzieLet39_4Lf''''''''_f''''''''_Int_Intsbos_1_merge_merge_fork_2,Pointer_QTree_Int)] */
  logic [1:0] \lizzieLet39_4Lf''''''''_f''''''''_Int_Intsbos_emitted ;
  logic [1:0] \lizzieLet39_4Lf''''''''_f''''''''_Int_Intsbos_done ;
  assign \lizzieLet39_4Lf''''''''_f''''''''_Int_Intsbos_1_merge_merge_fork_1_d  = {\lizzieLet39_4Lf''''''''_f''''''''_Int_Intsbos_d [16:1],
                                                                                   (\lizzieLet39_4Lf''''''''_f''''''''_Int_Intsbos_d [0] && (! \lizzieLet39_4Lf''''''''_f''''''''_Int_Intsbos_emitted [0]))};
  assign \lizzieLet39_4Lf''''''''_f''''''''_Int_Intsbos_1_merge_merge_fork_2_d  = {\lizzieLet39_4Lf''''''''_f''''''''_Int_Intsbos_d [16:1],
                                                                                   (\lizzieLet39_4Lf''''''''_f''''''''_Int_Intsbos_d [0] && (! \lizzieLet39_4Lf''''''''_f''''''''_Int_Intsbos_emitted [1]))};
  assign \lizzieLet39_4Lf''''''''_f''''''''_Int_Intsbos_done  = (\lizzieLet39_4Lf''''''''_f''''''''_Int_Intsbos_emitted  | ({\lizzieLet39_4Lf''''''''_f''''''''_Int_Intsbos_1_merge_merge_fork_2_d [0],
                                                                                                                             \lizzieLet39_4Lf''''''''_f''''''''_Int_Intsbos_1_merge_merge_fork_1_d [0]} & {\lizzieLet39_4Lf''''''''_f''''''''_Int_Intsbos_1_merge_merge_fork_2_r ,
                                                                                                                                                                                                           \lizzieLet39_4Lf''''''''_f''''''''_Int_Intsbos_1_merge_merge_fork_1_r }));
  assign \lizzieLet39_4Lf''''''''_f''''''''_Int_Intsbos_r  = (& \lizzieLet39_4Lf''''''''_f''''''''_Int_Intsbos_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet39_4Lf''''''''_f''''''''_Int_Intsbos_emitted  <= 2'd0;
    else
      \lizzieLet39_4Lf''''''''_f''''''''_Int_Intsbos_emitted  <= (\lizzieLet39_4Lf''''''''_f''''''''_Int_Intsbos_r  ? 2'd0 :
                                                                  \lizzieLet39_4Lf''''''''_f''''''''_Int_Intsbos_done );
  
  /* togo (Ty Pointer_QTree_Int) : (lizzieLet39_4Lf''''''''_f''''''''_Int_Intsbos_1_merge_merge_fork_1,Pointer_QTree_Int) > (call_f''''''''_f''''''''_Int_Int_goConst,Go) */
  assign \call_f''''''''_f''''''''_Int_Int_goConst_d  = \lizzieLet39_4Lf''''''''_f''''''''_Int_Intsbos_1_merge_merge_fork_1_d [0];
  assign \lizzieLet39_4Lf''''''''_f''''''''_Int_Intsbos_1_merge_merge_fork_1_r  = \call_f''''''''_f''''''''_Int_Int_goConst_r ;
  
  /* demux (Ty MyBool,
       Ty Go) : (lizzieLet3_1,MyBool) (arg0_1Dcon_is_z_1_3I#_3,Go) > [(lizzieLet3_1MyFalse,Go),
                                                                      (lizzieLet3_1MyTrue,Go)] */
  logic [1:0] \arg0_1Dcon_is_z_1_3I#_3_onehotd ;
  always_comb
    if ((lizzieLet3_1_d[0] && \arg0_1Dcon_is_z_1_3I#_3_d [0]))
      unique case (lizzieLet3_1_d[1:1])
        1'd0: \arg0_1Dcon_is_z_1_3I#_3_onehotd  = 2'd1;
        1'd1: \arg0_1Dcon_is_z_1_3I#_3_onehotd  = 2'd2;
        default: \arg0_1Dcon_is_z_1_3I#_3_onehotd  = 2'd0;
      endcase
    else \arg0_1Dcon_is_z_1_3I#_3_onehotd  = 2'd0;
  assign lizzieLet3_1MyFalse_d = \arg0_1Dcon_is_z_1_3I#_3_onehotd [0];
  assign lizzieLet3_1MyTrue_d = \arg0_1Dcon_is_z_1_3I#_3_onehotd [1];
  assign \arg0_1Dcon_is_z_1_3I#_3_r  = (| (\arg0_1Dcon_is_z_1_3I#_3_onehotd  & {lizzieLet3_1MyTrue_r,
                                                                                lizzieLet3_1MyFalse_r}));
  assign lizzieLet3_1_r = \arg0_1Dcon_is_z_1_3I#_3_r ;
  
  /* dcon (Ty MyBool,
      Dcon MyFalse) : [(lizzieLet3_1MyFalse,Go)] > (lizzieLet3_1MyFalse_1MyFalse,MyBool) */
  assign lizzieLet3_1MyFalse_1MyFalse_d = MyFalse_dc((& {lizzieLet3_1MyFalse_d[0]}), lizzieLet3_1MyFalse_d);
  assign {lizzieLet3_1MyFalse_r} = {1 {(lizzieLet3_1MyFalse_1MyFalse_r && lizzieLet3_1MyFalse_1MyFalse_d[0])}};
  
  /* dcon (Ty MyBool,
      Dcon MyTrue) : [(lizzieLet3_1MyTrue,Go)] > (lizzieLet3_1MyTrue_1MyTrue,MyBool) */
  assign lizzieLet3_1MyTrue_1MyTrue_d = MyTrue_dc((& {lizzieLet3_1MyTrue_d[0]}), lizzieLet3_1MyTrue_d);
  assign {lizzieLet3_1MyTrue_r} = {1 {(lizzieLet3_1MyTrue_1MyTrue_r && lizzieLet3_1MyTrue_1MyTrue_d[0])}};
  
  /* mux (Ty MyBool,
     Ty MyBool) : (lizzieLet3_2,MyBool) [(lizzieLet3_1MyFalse_1MyFalse,MyBool),
                                         (lizzieLet3_1MyTrue_1MyTrue,MyBool)] > (lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux,MyBool) */
  logic [1:0] lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux;
  logic [1:0] lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_onehot;
  always_comb
    unique case (lizzieLet3_2_d[1:1])
      1'd0:
        {lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_onehot,
         lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux} = {2'd1,
                                                                            lizzieLet3_1MyFalse_1MyFalse_d};
      1'd1:
        {lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_onehot,
         lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux} = {2'd2,
                                                                            lizzieLet3_1MyTrue_1MyTrue_d};
      default:
        {lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_onehot,
         lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux} = {2'd0,
                                                                            {1'd0, 1'd0}};
    endcase
  assign lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_d = {lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux[1:1],
                                                                         (lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux[0] && lizzieLet3_2_d[0])};
  assign lizzieLet3_2_r = (lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_d[0] && lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_r);
  assign {lizzieLet3_1MyTrue_1MyTrue_r,
          lizzieLet3_1MyFalse_1MyFalse_r} = (lizzieLet3_2_r ? lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_onehot :
                                             2'd0);
  
  /* destruct (Ty CTf_f_Int_Int,
          Dcon Lcall_f_f_Int_Int0) : (lizzieLet44_1Lcall_f_f_Int_Int0,CTf_f_Int_Int) > [(es_28_destruct,Pointer_QTree_Int),
                                                                                        (es_29_1_destruct,Pointer_QTree_Int),
                                                                                        (es_30_2_destruct,Pointer_QTree_Int),
                                                                                        (sc_0_14_destruct,Pointer_CTf_f_Int_Int)] */
  logic [3:0] lizzieLet44_1Lcall_f_f_Int_Int0_emitted;
  logic [3:0] lizzieLet44_1Lcall_f_f_Int_Int0_done;
  assign es_28_destruct_d = {lizzieLet44_1Lcall_f_f_Int_Int0_d[19:4],
                             (lizzieLet44_1Lcall_f_f_Int_Int0_d[0] && (! lizzieLet44_1Lcall_f_f_Int_Int0_emitted[0]))};
  assign es_29_1_destruct_d = {lizzieLet44_1Lcall_f_f_Int_Int0_d[35:20],
                               (lizzieLet44_1Lcall_f_f_Int_Int0_d[0] && (! lizzieLet44_1Lcall_f_f_Int_Int0_emitted[1]))};
  assign es_30_2_destruct_d = {lizzieLet44_1Lcall_f_f_Int_Int0_d[51:36],
                               (lizzieLet44_1Lcall_f_f_Int_Int0_d[0] && (! lizzieLet44_1Lcall_f_f_Int_Int0_emitted[2]))};
  assign sc_0_14_destruct_d = {lizzieLet44_1Lcall_f_f_Int_Int0_d[67:52],
                               (lizzieLet44_1Lcall_f_f_Int_Int0_d[0] && (! lizzieLet44_1Lcall_f_f_Int_Int0_emitted[3]))};
  assign lizzieLet44_1Lcall_f_f_Int_Int0_done = (lizzieLet44_1Lcall_f_f_Int_Int0_emitted | ({sc_0_14_destruct_d[0],
                                                                                             es_30_2_destruct_d[0],
                                                                                             es_29_1_destruct_d[0],
                                                                                             es_28_destruct_d[0]} & {sc_0_14_destruct_r,
                                                                                                                     es_30_2_destruct_r,
                                                                                                                     es_29_1_destruct_r,
                                                                                                                     es_28_destruct_r}));
  assign lizzieLet44_1Lcall_f_f_Int_Int0_r = (& lizzieLet44_1Lcall_f_f_Int_Int0_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet44_1Lcall_f_f_Int_Int0_emitted <= 4'd0;
    else
      lizzieLet44_1Lcall_f_f_Int_Int0_emitted <= (lizzieLet44_1Lcall_f_f_Int_Int0_r ? 4'd0 :
                                                  lizzieLet44_1Lcall_f_f_Int_Int0_done);
  
  /* destruct (Ty CTf_f_Int_Int,
          Dcon Lcall_f_f_Int_Int1) : (lizzieLet44_1Lcall_f_f_Int_Int1,CTf_f_Int_Int) > [(es_29_destruct,Pointer_QTree_Int),
                                                                                        (es_30_1_destruct,Pointer_QTree_Int),
                                                                                        (sc_0_13_destruct,Pointer_CTf_f_Int_Int),
                                                                                        (q1a8T_3_destruct,Pointer_QTree_Int),
                                                                                        (t1a8Y_3_destruct,Pointer_QTree_Int),
                                                                                        (is_z_mapa8E_4_destruct,MyDTInt_Bool),
                                                                                        (op_mapa8F_4_destruct,MyDTInt_Int),
                                                                                        (is_z_adda8G_4_destruct,MyDTInt_Bool),
                                                                                        (op_adda8H_4_destruct,MyDTInt_Int_Int)] */
  logic [8:0] lizzieLet44_1Lcall_f_f_Int_Int1_emitted;
  logic [8:0] lizzieLet44_1Lcall_f_f_Int_Int1_done;
  assign es_29_destruct_d = {lizzieLet44_1Lcall_f_f_Int_Int1_d[19:4],
                             (lizzieLet44_1Lcall_f_f_Int_Int1_d[0] && (! lizzieLet44_1Lcall_f_f_Int_Int1_emitted[0]))};
  assign es_30_1_destruct_d = {lizzieLet44_1Lcall_f_f_Int_Int1_d[35:20],
                               (lizzieLet44_1Lcall_f_f_Int_Int1_d[0] && (! lizzieLet44_1Lcall_f_f_Int_Int1_emitted[1]))};
  assign sc_0_13_destruct_d = {lizzieLet44_1Lcall_f_f_Int_Int1_d[51:36],
                               (lizzieLet44_1Lcall_f_f_Int_Int1_d[0] && (! lizzieLet44_1Lcall_f_f_Int_Int1_emitted[2]))};
  assign q1a8T_3_destruct_d = {lizzieLet44_1Lcall_f_f_Int_Int1_d[67:52],
                               (lizzieLet44_1Lcall_f_f_Int_Int1_d[0] && (! lizzieLet44_1Lcall_f_f_Int_Int1_emitted[3]))};
  assign t1a8Y_3_destruct_d = {lizzieLet44_1Lcall_f_f_Int_Int1_d[83:68],
                               (lizzieLet44_1Lcall_f_f_Int_Int1_d[0] && (! lizzieLet44_1Lcall_f_f_Int_Int1_emitted[4]))};
  assign is_z_mapa8E_4_destruct_d = (lizzieLet44_1Lcall_f_f_Int_Int1_d[0] && (! lizzieLet44_1Lcall_f_f_Int_Int1_emitted[5]));
  assign op_mapa8F_4_destruct_d = (lizzieLet44_1Lcall_f_f_Int_Int1_d[0] && (! lizzieLet44_1Lcall_f_f_Int_Int1_emitted[6]));
  assign is_z_adda8G_4_destruct_d = (lizzieLet44_1Lcall_f_f_Int_Int1_d[0] && (! lizzieLet44_1Lcall_f_f_Int_Int1_emitted[7]));
  assign op_adda8H_4_destruct_d = (lizzieLet44_1Lcall_f_f_Int_Int1_d[0] && (! lizzieLet44_1Lcall_f_f_Int_Int1_emitted[8]));
  assign lizzieLet44_1Lcall_f_f_Int_Int1_done = (lizzieLet44_1Lcall_f_f_Int_Int1_emitted | ({op_adda8H_4_destruct_d[0],
                                                                                             is_z_adda8G_4_destruct_d[0],
                                                                                             op_mapa8F_4_destruct_d[0],
                                                                                             is_z_mapa8E_4_destruct_d[0],
                                                                                             t1a8Y_3_destruct_d[0],
                                                                                             q1a8T_3_destruct_d[0],
                                                                                             sc_0_13_destruct_d[0],
                                                                                             es_30_1_destruct_d[0],
                                                                                             es_29_destruct_d[0]} & {op_adda8H_4_destruct_r,
                                                                                                                     is_z_adda8G_4_destruct_r,
                                                                                                                     op_mapa8F_4_destruct_r,
                                                                                                                     is_z_mapa8E_4_destruct_r,
                                                                                                                     t1a8Y_3_destruct_r,
                                                                                                                     q1a8T_3_destruct_r,
                                                                                                                     sc_0_13_destruct_r,
                                                                                                                     es_30_1_destruct_r,
                                                                                                                     es_29_destruct_r}));
  assign lizzieLet44_1Lcall_f_f_Int_Int1_r = (& lizzieLet44_1Lcall_f_f_Int_Int1_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet44_1Lcall_f_f_Int_Int1_emitted <= 9'd0;
    else
      lizzieLet44_1Lcall_f_f_Int_Int1_emitted <= (lizzieLet44_1Lcall_f_f_Int_Int1_r ? 9'd0 :
                                                  lizzieLet44_1Lcall_f_f_Int_Int1_done);
  
  /* destruct (Ty CTf_f_Int_Int,
          Dcon Lcall_f_f_Int_Int2) : (lizzieLet44_1Lcall_f_f_Int_Int2,CTf_f_Int_Int) > [(es_30_destruct,Pointer_QTree_Int),
                                                                                        (sc_0_12_destruct,Pointer_CTf_f_Int_Int),
                                                                                        (q1a8T_2_destruct,Pointer_QTree_Int),
                                                                                        (t1a8Y_2_destruct,Pointer_QTree_Int),
                                                                                        (is_z_mapa8E_3_destruct,MyDTInt_Bool),
                                                                                        (op_mapa8F_3_destruct,MyDTInt_Int),
                                                                                        (is_z_adda8G_3_destruct,MyDTInt_Bool),
                                                                                        (op_adda8H_3_destruct,MyDTInt_Int_Int),
                                                                                        (q2a8U_2_destruct,Pointer_QTree_Int),
                                                                                        (t2a8Z_2_destruct,Pointer_QTree_Int)] */
  logic [9:0] lizzieLet44_1Lcall_f_f_Int_Int2_emitted;
  logic [9:0] lizzieLet44_1Lcall_f_f_Int_Int2_done;
  assign es_30_destruct_d = {lizzieLet44_1Lcall_f_f_Int_Int2_d[19:4],
                             (lizzieLet44_1Lcall_f_f_Int_Int2_d[0] && (! lizzieLet44_1Lcall_f_f_Int_Int2_emitted[0]))};
  assign sc_0_12_destruct_d = {lizzieLet44_1Lcall_f_f_Int_Int2_d[35:20],
                               (lizzieLet44_1Lcall_f_f_Int_Int2_d[0] && (! lizzieLet44_1Lcall_f_f_Int_Int2_emitted[1]))};
  assign q1a8T_2_destruct_d = {lizzieLet44_1Lcall_f_f_Int_Int2_d[51:36],
                               (lizzieLet44_1Lcall_f_f_Int_Int2_d[0] && (! lizzieLet44_1Lcall_f_f_Int_Int2_emitted[2]))};
  assign t1a8Y_2_destruct_d = {lizzieLet44_1Lcall_f_f_Int_Int2_d[67:52],
                               (lizzieLet44_1Lcall_f_f_Int_Int2_d[0] && (! lizzieLet44_1Lcall_f_f_Int_Int2_emitted[3]))};
  assign is_z_mapa8E_3_destruct_d = (lizzieLet44_1Lcall_f_f_Int_Int2_d[0] && (! lizzieLet44_1Lcall_f_f_Int_Int2_emitted[4]));
  assign op_mapa8F_3_destruct_d = (lizzieLet44_1Lcall_f_f_Int_Int2_d[0] && (! lizzieLet44_1Lcall_f_f_Int_Int2_emitted[5]));
  assign is_z_adda8G_3_destruct_d = (lizzieLet44_1Lcall_f_f_Int_Int2_d[0] && (! lizzieLet44_1Lcall_f_f_Int_Int2_emitted[6]));
  assign op_adda8H_3_destruct_d = (lizzieLet44_1Lcall_f_f_Int_Int2_d[0] && (! lizzieLet44_1Lcall_f_f_Int_Int2_emitted[7]));
  assign q2a8U_2_destruct_d = {lizzieLet44_1Lcall_f_f_Int_Int2_d[83:68],
                               (lizzieLet44_1Lcall_f_f_Int_Int2_d[0] && (! lizzieLet44_1Lcall_f_f_Int_Int2_emitted[8]))};
  assign t2a8Z_2_destruct_d = {lizzieLet44_1Lcall_f_f_Int_Int2_d[99:84],
                               (lizzieLet44_1Lcall_f_f_Int_Int2_d[0] && (! lizzieLet44_1Lcall_f_f_Int_Int2_emitted[9]))};
  assign lizzieLet44_1Lcall_f_f_Int_Int2_done = (lizzieLet44_1Lcall_f_f_Int_Int2_emitted | ({t2a8Z_2_destruct_d[0],
                                                                                             q2a8U_2_destruct_d[0],
                                                                                             op_adda8H_3_destruct_d[0],
                                                                                             is_z_adda8G_3_destruct_d[0],
                                                                                             op_mapa8F_3_destruct_d[0],
                                                                                             is_z_mapa8E_3_destruct_d[0],
                                                                                             t1a8Y_2_destruct_d[0],
                                                                                             q1a8T_2_destruct_d[0],
                                                                                             sc_0_12_destruct_d[0],
                                                                                             es_30_destruct_d[0]} & {t2a8Z_2_destruct_r,
                                                                                                                     q2a8U_2_destruct_r,
                                                                                                                     op_adda8H_3_destruct_r,
                                                                                                                     is_z_adda8G_3_destruct_r,
                                                                                                                     op_mapa8F_3_destruct_r,
                                                                                                                     is_z_mapa8E_3_destruct_r,
                                                                                                                     t1a8Y_2_destruct_r,
                                                                                                                     q1a8T_2_destruct_r,
                                                                                                                     sc_0_12_destruct_r,
                                                                                                                     es_30_destruct_r}));
  assign lizzieLet44_1Lcall_f_f_Int_Int2_r = (& lizzieLet44_1Lcall_f_f_Int_Int2_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet44_1Lcall_f_f_Int_Int2_emitted <= 10'd0;
    else
      lizzieLet44_1Lcall_f_f_Int_Int2_emitted <= (lizzieLet44_1Lcall_f_f_Int_Int2_r ? 10'd0 :
                                                  lizzieLet44_1Lcall_f_f_Int_Int2_done);
  
  /* destruct (Ty CTf_f_Int_Int,
          Dcon Lcall_f_f_Int_Int3) : (lizzieLet44_1Lcall_f_f_Int_Int3,CTf_f_Int_Int) > [(sc_0_11_destruct,Pointer_CTf_f_Int_Int),
                                                                                        (q1a8T_1_destruct,Pointer_QTree_Int),
                                                                                        (t1a8Y_1_destruct,Pointer_QTree_Int),
                                                                                        (is_z_mapa8E_2_destruct,MyDTInt_Bool),
                                                                                        (op_mapa8F_2_destruct,MyDTInt_Int),
                                                                                        (is_z_adda8G_2_destruct,MyDTInt_Bool),
                                                                                        (op_adda8H_2_destruct,MyDTInt_Int_Int),
                                                                                        (q2a8U_1_destruct,Pointer_QTree_Int),
                                                                                        (t2a8Z_1_destruct,Pointer_QTree_Int),
                                                                                        (q3a8V_1_destruct,Pointer_QTree_Int),
                                                                                        (t3a90_1_destruct,Pointer_QTree_Int)] */
  logic [10:0] lizzieLet44_1Lcall_f_f_Int_Int3_emitted;
  logic [10:0] lizzieLet44_1Lcall_f_f_Int_Int3_done;
  assign sc_0_11_destruct_d = {lizzieLet44_1Lcall_f_f_Int_Int3_d[19:4],
                               (lizzieLet44_1Lcall_f_f_Int_Int3_d[0] && (! lizzieLet44_1Lcall_f_f_Int_Int3_emitted[0]))};
  assign q1a8T_1_destruct_d = {lizzieLet44_1Lcall_f_f_Int_Int3_d[35:20],
                               (lizzieLet44_1Lcall_f_f_Int_Int3_d[0] && (! lizzieLet44_1Lcall_f_f_Int_Int3_emitted[1]))};
  assign t1a8Y_1_destruct_d = {lizzieLet44_1Lcall_f_f_Int_Int3_d[51:36],
                               (lizzieLet44_1Lcall_f_f_Int_Int3_d[0] && (! lizzieLet44_1Lcall_f_f_Int_Int3_emitted[2]))};
  assign is_z_mapa8E_2_destruct_d = (lizzieLet44_1Lcall_f_f_Int_Int3_d[0] && (! lizzieLet44_1Lcall_f_f_Int_Int3_emitted[3]));
  assign op_mapa8F_2_destruct_d = (lizzieLet44_1Lcall_f_f_Int_Int3_d[0] && (! lizzieLet44_1Lcall_f_f_Int_Int3_emitted[4]));
  assign is_z_adda8G_2_destruct_d = (lizzieLet44_1Lcall_f_f_Int_Int3_d[0] && (! lizzieLet44_1Lcall_f_f_Int_Int3_emitted[5]));
  assign op_adda8H_2_destruct_d = (lizzieLet44_1Lcall_f_f_Int_Int3_d[0] && (! lizzieLet44_1Lcall_f_f_Int_Int3_emitted[6]));
  assign q2a8U_1_destruct_d = {lizzieLet44_1Lcall_f_f_Int_Int3_d[67:52],
                               (lizzieLet44_1Lcall_f_f_Int_Int3_d[0] && (! lizzieLet44_1Lcall_f_f_Int_Int3_emitted[7]))};
  assign t2a8Z_1_destruct_d = {lizzieLet44_1Lcall_f_f_Int_Int3_d[83:68],
                               (lizzieLet44_1Lcall_f_f_Int_Int3_d[0] && (! lizzieLet44_1Lcall_f_f_Int_Int3_emitted[8]))};
  assign q3a8V_1_destruct_d = {lizzieLet44_1Lcall_f_f_Int_Int3_d[99:84],
                               (lizzieLet44_1Lcall_f_f_Int_Int3_d[0] && (! lizzieLet44_1Lcall_f_f_Int_Int3_emitted[9]))};
  assign t3a90_1_destruct_d = {lizzieLet44_1Lcall_f_f_Int_Int3_d[115:100],
                               (lizzieLet44_1Lcall_f_f_Int_Int3_d[0] && (! lizzieLet44_1Lcall_f_f_Int_Int3_emitted[10]))};
  assign lizzieLet44_1Lcall_f_f_Int_Int3_done = (lizzieLet44_1Lcall_f_f_Int_Int3_emitted | ({t3a90_1_destruct_d[0],
                                                                                             q3a8V_1_destruct_d[0],
                                                                                             t2a8Z_1_destruct_d[0],
                                                                                             q2a8U_1_destruct_d[0],
                                                                                             op_adda8H_2_destruct_d[0],
                                                                                             is_z_adda8G_2_destruct_d[0],
                                                                                             op_mapa8F_2_destruct_d[0],
                                                                                             is_z_mapa8E_2_destruct_d[0],
                                                                                             t1a8Y_1_destruct_d[0],
                                                                                             q1a8T_1_destruct_d[0],
                                                                                             sc_0_11_destruct_d[0]} & {t3a90_1_destruct_r,
                                                                                                                       q3a8V_1_destruct_r,
                                                                                                                       t2a8Z_1_destruct_r,
                                                                                                                       q2a8U_1_destruct_r,
                                                                                                                       op_adda8H_2_destruct_r,
                                                                                                                       is_z_adda8G_2_destruct_r,
                                                                                                                       op_mapa8F_2_destruct_r,
                                                                                                                       is_z_mapa8E_2_destruct_r,
                                                                                                                       t1a8Y_1_destruct_r,
                                                                                                                       q1a8T_1_destruct_r,
                                                                                                                       sc_0_11_destruct_r}));
  assign lizzieLet44_1Lcall_f_f_Int_Int3_r = (& lizzieLet44_1Lcall_f_f_Int_Int3_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet44_1Lcall_f_f_Int_Int3_emitted <= 11'd0;
    else
      lizzieLet44_1Lcall_f_f_Int_Int3_emitted <= (lizzieLet44_1Lcall_f_f_Int_Int3_r ? 11'd0 :
                                                  lizzieLet44_1Lcall_f_f_Int_Int3_done);
  
  /* demux (Ty CTf_f_Int_Int,
       Ty CTf_f_Int_Int) : (lizzieLet44_2,CTf_f_Int_Int) (lizzieLet44_1,CTf_f_Int_Int) > [(_10,CTf_f_Int_Int),
                                                                                          (lizzieLet44_1Lcall_f_f_Int_Int3,CTf_f_Int_Int),
                                                                                          (lizzieLet44_1Lcall_f_f_Int_Int2,CTf_f_Int_Int),
                                                                                          (lizzieLet44_1Lcall_f_f_Int_Int1,CTf_f_Int_Int),
                                                                                          (lizzieLet44_1Lcall_f_f_Int_Int0,CTf_f_Int_Int)] */
  logic [4:0] lizzieLet44_1_onehotd;
  always_comb
    if ((lizzieLet44_2_d[0] && lizzieLet44_1_d[0]))
      unique case (lizzieLet44_2_d[3:1])
        3'd0: lizzieLet44_1_onehotd = 5'd1;
        3'd1: lizzieLet44_1_onehotd = 5'd2;
        3'd2: lizzieLet44_1_onehotd = 5'd4;
        3'd3: lizzieLet44_1_onehotd = 5'd8;
        3'd4: lizzieLet44_1_onehotd = 5'd16;
        default: lizzieLet44_1_onehotd = 5'd0;
      endcase
    else lizzieLet44_1_onehotd = 5'd0;
  assign _10_d = {lizzieLet44_1_d[115:1], lizzieLet44_1_onehotd[0]};
  assign lizzieLet44_1Lcall_f_f_Int_Int3_d = {lizzieLet44_1_d[115:1],
                                              lizzieLet44_1_onehotd[1]};
  assign lizzieLet44_1Lcall_f_f_Int_Int2_d = {lizzieLet44_1_d[115:1],
                                              lizzieLet44_1_onehotd[2]};
  assign lizzieLet44_1Lcall_f_f_Int_Int1_d = {lizzieLet44_1_d[115:1],
                                              lizzieLet44_1_onehotd[3]};
  assign lizzieLet44_1Lcall_f_f_Int_Int0_d = {lizzieLet44_1_d[115:1],
                                              lizzieLet44_1_onehotd[4]};
  assign lizzieLet44_1_r = (| (lizzieLet44_1_onehotd & {lizzieLet44_1Lcall_f_f_Int_Int0_r,
                                                        lizzieLet44_1Lcall_f_f_Int_Int1_r,
                                                        lizzieLet44_1Lcall_f_f_Int_Int2_r,
                                                        lizzieLet44_1Lcall_f_f_Int_Int3_r,
                                                        _10_r}));
  assign lizzieLet44_2_r = lizzieLet44_1_r;
  
  /* demux (Ty CTf_f_Int_Int,
       Ty Go) : (lizzieLet44_3,CTf_f_Int_Int) (go_17_goMux_data,Go) > [(_9,Go),
                                                                       (lizzieLet44_3Lcall_f_f_Int_Int3,Go),
                                                                       (lizzieLet44_3Lcall_f_f_Int_Int2,Go),
                                                                       (lizzieLet44_3Lcall_f_f_Int_Int1,Go),
                                                                       (lizzieLet44_3Lcall_f_f_Int_Int0,Go)] */
  logic [4:0] go_17_goMux_data_onehotd;
  always_comb
    if ((lizzieLet44_3_d[0] && go_17_goMux_data_d[0]))
      unique case (lizzieLet44_3_d[3:1])
        3'd0: go_17_goMux_data_onehotd = 5'd1;
        3'd1: go_17_goMux_data_onehotd = 5'd2;
        3'd2: go_17_goMux_data_onehotd = 5'd4;
        3'd3: go_17_goMux_data_onehotd = 5'd8;
        3'd4: go_17_goMux_data_onehotd = 5'd16;
        default: go_17_goMux_data_onehotd = 5'd0;
      endcase
    else go_17_goMux_data_onehotd = 5'd0;
  assign _9_d = go_17_goMux_data_onehotd[0];
  assign lizzieLet44_3Lcall_f_f_Int_Int3_d = go_17_goMux_data_onehotd[1];
  assign lizzieLet44_3Lcall_f_f_Int_Int2_d = go_17_goMux_data_onehotd[2];
  assign lizzieLet44_3Lcall_f_f_Int_Int1_d = go_17_goMux_data_onehotd[3];
  assign lizzieLet44_3Lcall_f_f_Int_Int0_d = go_17_goMux_data_onehotd[4];
  assign go_17_goMux_data_r = (| (go_17_goMux_data_onehotd & {lizzieLet44_3Lcall_f_f_Int_Int0_r,
                                                              lizzieLet44_3Lcall_f_f_Int_Int1_r,
                                                              lizzieLet44_3Lcall_f_f_Int_Int2_r,
                                                              lizzieLet44_3Lcall_f_f_Int_Int3_r,
                                                              _9_r}));
  assign lizzieLet44_3_r = go_17_goMux_data_r;
  
  /* buf (Ty Go) : (lizzieLet44_3Lcall_f_f_Int_Int0,Go) > (lizzieLet44_3Lcall_f_f_Int_Int0_1_argbuf,Go) */
  Go_t lizzieLet44_3Lcall_f_f_Int_Int0_bufchan_d;
  logic lizzieLet44_3Lcall_f_f_Int_Int0_bufchan_r;
  assign lizzieLet44_3Lcall_f_f_Int_Int0_r = ((! lizzieLet44_3Lcall_f_f_Int_Int0_bufchan_d[0]) || lizzieLet44_3Lcall_f_f_Int_Int0_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet44_3Lcall_f_f_Int_Int0_bufchan_d <= 1'd0;
    else
      if (lizzieLet44_3Lcall_f_f_Int_Int0_r)
        lizzieLet44_3Lcall_f_f_Int_Int0_bufchan_d <= lizzieLet44_3Lcall_f_f_Int_Int0_d;
  Go_t lizzieLet44_3Lcall_f_f_Int_Int0_bufchan_buf;
  assign lizzieLet44_3Lcall_f_f_Int_Int0_bufchan_r = (! lizzieLet44_3Lcall_f_f_Int_Int0_bufchan_buf[0]);
  assign lizzieLet44_3Lcall_f_f_Int_Int0_1_argbuf_d = (lizzieLet44_3Lcall_f_f_Int_Int0_bufchan_buf[0] ? lizzieLet44_3Lcall_f_f_Int_Int0_bufchan_buf :
                                                       lizzieLet44_3Lcall_f_f_Int_Int0_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet44_3Lcall_f_f_Int_Int0_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet44_3Lcall_f_f_Int_Int0_1_argbuf_r && lizzieLet44_3Lcall_f_f_Int_Int0_bufchan_buf[0]))
        lizzieLet44_3Lcall_f_f_Int_Int0_bufchan_buf <= 1'd0;
      else if (((! lizzieLet44_3Lcall_f_f_Int_Int0_1_argbuf_r) && (! lizzieLet44_3Lcall_f_f_Int_Int0_bufchan_buf[0])))
        lizzieLet44_3Lcall_f_f_Int_Int0_bufchan_buf <= lizzieLet44_3Lcall_f_f_Int_Int0_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet44_3Lcall_f_f_Int_Int1,Go) > (lizzieLet44_3Lcall_f_f_Int_Int1_1_argbuf,Go) */
  Go_t lizzieLet44_3Lcall_f_f_Int_Int1_bufchan_d;
  logic lizzieLet44_3Lcall_f_f_Int_Int1_bufchan_r;
  assign lizzieLet44_3Lcall_f_f_Int_Int1_r = ((! lizzieLet44_3Lcall_f_f_Int_Int1_bufchan_d[0]) || lizzieLet44_3Lcall_f_f_Int_Int1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet44_3Lcall_f_f_Int_Int1_bufchan_d <= 1'd0;
    else
      if (lizzieLet44_3Lcall_f_f_Int_Int1_r)
        lizzieLet44_3Lcall_f_f_Int_Int1_bufchan_d <= lizzieLet44_3Lcall_f_f_Int_Int1_d;
  Go_t lizzieLet44_3Lcall_f_f_Int_Int1_bufchan_buf;
  assign lizzieLet44_3Lcall_f_f_Int_Int1_bufchan_r = (! lizzieLet44_3Lcall_f_f_Int_Int1_bufchan_buf[0]);
  assign lizzieLet44_3Lcall_f_f_Int_Int1_1_argbuf_d = (lizzieLet44_3Lcall_f_f_Int_Int1_bufchan_buf[0] ? lizzieLet44_3Lcall_f_f_Int_Int1_bufchan_buf :
                                                       lizzieLet44_3Lcall_f_f_Int_Int1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet44_3Lcall_f_f_Int_Int1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet44_3Lcall_f_f_Int_Int1_1_argbuf_r && lizzieLet44_3Lcall_f_f_Int_Int1_bufchan_buf[0]))
        lizzieLet44_3Lcall_f_f_Int_Int1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet44_3Lcall_f_f_Int_Int1_1_argbuf_r) && (! lizzieLet44_3Lcall_f_f_Int_Int1_bufchan_buf[0])))
        lizzieLet44_3Lcall_f_f_Int_Int1_bufchan_buf <= lizzieLet44_3Lcall_f_f_Int_Int1_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet44_3Lcall_f_f_Int_Int2,Go) > (lizzieLet44_3Lcall_f_f_Int_Int2_1_argbuf,Go) */
  Go_t lizzieLet44_3Lcall_f_f_Int_Int2_bufchan_d;
  logic lizzieLet44_3Lcall_f_f_Int_Int2_bufchan_r;
  assign lizzieLet44_3Lcall_f_f_Int_Int2_r = ((! lizzieLet44_3Lcall_f_f_Int_Int2_bufchan_d[0]) || lizzieLet44_3Lcall_f_f_Int_Int2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet44_3Lcall_f_f_Int_Int2_bufchan_d <= 1'd0;
    else
      if (lizzieLet44_3Lcall_f_f_Int_Int2_r)
        lizzieLet44_3Lcall_f_f_Int_Int2_bufchan_d <= lizzieLet44_3Lcall_f_f_Int_Int2_d;
  Go_t lizzieLet44_3Lcall_f_f_Int_Int2_bufchan_buf;
  assign lizzieLet44_3Lcall_f_f_Int_Int2_bufchan_r = (! lizzieLet44_3Lcall_f_f_Int_Int2_bufchan_buf[0]);
  assign lizzieLet44_3Lcall_f_f_Int_Int2_1_argbuf_d = (lizzieLet44_3Lcall_f_f_Int_Int2_bufchan_buf[0] ? lizzieLet44_3Lcall_f_f_Int_Int2_bufchan_buf :
                                                       lizzieLet44_3Lcall_f_f_Int_Int2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet44_3Lcall_f_f_Int_Int2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet44_3Lcall_f_f_Int_Int2_1_argbuf_r && lizzieLet44_3Lcall_f_f_Int_Int2_bufchan_buf[0]))
        lizzieLet44_3Lcall_f_f_Int_Int2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet44_3Lcall_f_f_Int_Int2_1_argbuf_r) && (! lizzieLet44_3Lcall_f_f_Int_Int2_bufchan_buf[0])))
        lizzieLet44_3Lcall_f_f_Int_Int2_bufchan_buf <= lizzieLet44_3Lcall_f_f_Int_Int2_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet44_3Lcall_f_f_Int_Int3,Go) > (lizzieLet44_3Lcall_f_f_Int_Int3_1_argbuf,Go) */
  Go_t lizzieLet44_3Lcall_f_f_Int_Int3_bufchan_d;
  logic lizzieLet44_3Lcall_f_f_Int_Int3_bufchan_r;
  assign lizzieLet44_3Lcall_f_f_Int_Int3_r = ((! lizzieLet44_3Lcall_f_f_Int_Int3_bufchan_d[0]) || lizzieLet44_3Lcall_f_f_Int_Int3_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet44_3Lcall_f_f_Int_Int3_bufchan_d <= 1'd0;
    else
      if (lizzieLet44_3Lcall_f_f_Int_Int3_r)
        lizzieLet44_3Lcall_f_f_Int_Int3_bufchan_d <= lizzieLet44_3Lcall_f_f_Int_Int3_d;
  Go_t lizzieLet44_3Lcall_f_f_Int_Int3_bufchan_buf;
  assign lizzieLet44_3Lcall_f_f_Int_Int3_bufchan_r = (! lizzieLet44_3Lcall_f_f_Int_Int3_bufchan_buf[0]);
  assign lizzieLet44_3Lcall_f_f_Int_Int3_1_argbuf_d = (lizzieLet44_3Lcall_f_f_Int_Int3_bufchan_buf[0] ? lizzieLet44_3Lcall_f_f_Int_Int3_bufchan_buf :
                                                       lizzieLet44_3Lcall_f_f_Int_Int3_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet44_3Lcall_f_f_Int_Int3_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet44_3Lcall_f_f_Int_Int3_1_argbuf_r && lizzieLet44_3Lcall_f_f_Int_Int3_bufchan_buf[0]))
        lizzieLet44_3Lcall_f_f_Int_Int3_bufchan_buf <= 1'd0;
      else if (((! lizzieLet44_3Lcall_f_f_Int_Int3_1_argbuf_r) && (! lizzieLet44_3Lcall_f_f_Int_Int3_bufchan_buf[0])))
        lizzieLet44_3Lcall_f_f_Int_Int3_bufchan_buf <= lizzieLet44_3Lcall_f_f_Int_Int3_bufchan_d;
  
  /* demux (Ty CTf_f_Int_Int,
       Ty Pointer_QTree_Int) : (lizzieLet44_4,CTf_f_Int_Int) (srtarg_0_2_goMux_mux,Pointer_QTree_Int) > [(lizzieLet44_4Lf_f_Int_Intsbos,Pointer_QTree_Int),
                                                                                                         (lizzieLet44_4Lcall_f_f_Int_Int3,Pointer_QTree_Int),
                                                                                                         (lizzieLet44_4Lcall_f_f_Int_Int2,Pointer_QTree_Int),
                                                                                                         (lizzieLet44_4Lcall_f_f_Int_Int1,Pointer_QTree_Int),
                                                                                                         (lizzieLet44_4Lcall_f_f_Int_Int0,Pointer_QTree_Int)] */
  logic [4:0] srtarg_0_2_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet44_4_d[0] && srtarg_0_2_goMux_mux_d[0]))
      unique case (lizzieLet44_4_d[3:1])
        3'd0: srtarg_0_2_goMux_mux_onehotd = 5'd1;
        3'd1: srtarg_0_2_goMux_mux_onehotd = 5'd2;
        3'd2: srtarg_0_2_goMux_mux_onehotd = 5'd4;
        3'd3: srtarg_0_2_goMux_mux_onehotd = 5'd8;
        3'd4: srtarg_0_2_goMux_mux_onehotd = 5'd16;
        default: srtarg_0_2_goMux_mux_onehotd = 5'd0;
      endcase
    else srtarg_0_2_goMux_mux_onehotd = 5'd0;
  assign lizzieLet44_4Lf_f_Int_Intsbos_d = {srtarg_0_2_goMux_mux_d[16:1],
                                            srtarg_0_2_goMux_mux_onehotd[0]};
  assign lizzieLet44_4Lcall_f_f_Int_Int3_d = {srtarg_0_2_goMux_mux_d[16:1],
                                              srtarg_0_2_goMux_mux_onehotd[1]};
  assign lizzieLet44_4Lcall_f_f_Int_Int2_d = {srtarg_0_2_goMux_mux_d[16:1],
                                              srtarg_0_2_goMux_mux_onehotd[2]};
  assign lizzieLet44_4Lcall_f_f_Int_Int1_d = {srtarg_0_2_goMux_mux_d[16:1],
                                              srtarg_0_2_goMux_mux_onehotd[3]};
  assign lizzieLet44_4Lcall_f_f_Int_Int0_d = {srtarg_0_2_goMux_mux_d[16:1],
                                              srtarg_0_2_goMux_mux_onehotd[4]};
  assign srtarg_0_2_goMux_mux_r = (| (srtarg_0_2_goMux_mux_onehotd & {lizzieLet44_4Lcall_f_f_Int_Int0_r,
                                                                      lizzieLet44_4Lcall_f_f_Int_Int1_r,
                                                                      lizzieLet44_4Lcall_f_f_Int_Int2_r,
                                                                      lizzieLet44_4Lcall_f_f_Int_Int3_r,
                                                                      lizzieLet44_4Lf_f_Int_Intsbos_r}));
  assign lizzieLet44_4_r = srtarg_0_2_goMux_mux_r;
  
  /* dcon (Ty QTree_Int,
      Dcon QNode_Int) : [(lizzieLet44_4Lcall_f_f_Int_Int0,Pointer_QTree_Int),
                         (es_28_destruct,Pointer_QTree_Int),
                         (es_29_1_destruct,Pointer_QTree_Int),
                         (es_30_2_destruct,Pointer_QTree_Int)] > (lizzieLet44_4Lcall_f_f_Int_Int0_1es_28_1es_29_1_1es_30_2_1QNode_Int,QTree_Int) */
  assign lizzieLet44_4Lcall_f_f_Int_Int0_1es_28_1es_29_1_1es_30_2_1QNode_Int_d = QNode_Int_dc((& {lizzieLet44_4Lcall_f_f_Int_Int0_d[0],
                                                                                                  es_28_destruct_d[0],
                                                                                                  es_29_1_destruct_d[0],
                                                                                                  es_30_2_destruct_d[0]}), lizzieLet44_4Lcall_f_f_Int_Int0_d, es_28_destruct_d, es_29_1_destruct_d, es_30_2_destruct_d);
  assign {lizzieLet44_4Lcall_f_f_Int_Int0_r,
          es_28_destruct_r,
          es_29_1_destruct_r,
          es_30_2_destruct_r} = {4 {(lizzieLet44_4Lcall_f_f_Int_Int0_1es_28_1es_29_1_1es_30_2_1QNode_Int_r && lizzieLet44_4Lcall_f_f_Int_Int0_1es_28_1es_29_1_1es_30_2_1QNode_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (lizzieLet44_4Lcall_f_f_Int_Int0_1es_28_1es_29_1_1es_30_2_1QNode_Int,QTree_Int) > (lizzieLet48_1_argbuf,QTree_Int) */
  QTree_Int_t lizzieLet44_4Lcall_f_f_Int_Int0_1es_28_1es_29_1_1es_30_2_1QNode_Int_bufchan_d;
  logic lizzieLet44_4Lcall_f_f_Int_Int0_1es_28_1es_29_1_1es_30_2_1QNode_Int_bufchan_r;
  assign lizzieLet44_4Lcall_f_f_Int_Int0_1es_28_1es_29_1_1es_30_2_1QNode_Int_r = ((! lizzieLet44_4Lcall_f_f_Int_Int0_1es_28_1es_29_1_1es_30_2_1QNode_Int_bufchan_d[0]) || lizzieLet44_4Lcall_f_f_Int_Int0_1es_28_1es_29_1_1es_30_2_1QNode_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet44_4Lcall_f_f_Int_Int0_1es_28_1es_29_1_1es_30_2_1QNode_Int_bufchan_d <= {66'd0,
                                                                                        1'd0};
    else
      if (lizzieLet44_4Lcall_f_f_Int_Int0_1es_28_1es_29_1_1es_30_2_1QNode_Int_r)
        lizzieLet44_4Lcall_f_f_Int_Int0_1es_28_1es_29_1_1es_30_2_1QNode_Int_bufchan_d <= lizzieLet44_4Lcall_f_f_Int_Int0_1es_28_1es_29_1_1es_30_2_1QNode_Int_d;
  QTree_Int_t lizzieLet44_4Lcall_f_f_Int_Int0_1es_28_1es_29_1_1es_30_2_1QNode_Int_bufchan_buf;
  assign lizzieLet44_4Lcall_f_f_Int_Int0_1es_28_1es_29_1_1es_30_2_1QNode_Int_bufchan_r = (! lizzieLet44_4Lcall_f_f_Int_Int0_1es_28_1es_29_1_1es_30_2_1QNode_Int_bufchan_buf[0]);
  assign lizzieLet48_1_argbuf_d = (lizzieLet44_4Lcall_f_f_Int_Int0_1es_28_1es_29_1_1es_30_2_1QNode_Int_bufchan_buf[0] ? lizzieLet44_4Lcall_f_f_Int_Int0_1es_28_1es_29_1_1es_30_2_1QNode_Int_bufchan_buf :
                                   lizzieLet44_4Lcall_f_f_Int_Int0_1es_28_1es_29_1_1es_30_2_1QNode_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet44_4Lcall_f_f_Int_Int0_1es_28_1es_29_1_1es_30_2_1QNode_Int_bufchan_buf <= {66'd0,
                                                                                          1'd0};
    else
      if ((lizzieLet48_1_argbuf_r && lizzieLet44_4Lcall_f_f_Int_Int0_1es_28_1es_29_1_1es_30_2_1QNode_Int_bufchan_buf[0]))
        lizzieLet44_4Lcall_f_f_Int_Int0_1es_28_1es_29_1_1es_30_2_1QNode_Int_bufchan_buf <= {66'd0,
                                                                                            1'd0};
      else if (((! lizzieLet48_1_argbuf_r) && (! lizzieLet44_4Lcall_f_f_Int_Int0_1es_28_1es_29_1_1es_30_2_1QNode_Int_bufchan_buf[0])))
        lizzieLet44_4Lcall_f_f_Int_Int0_1es_28_1es_29_1_1es_30_2_1QNode_Int_bufchan_buf <= lizzieLet44_4Lcall_f_f_Int_Int0_1es_28_1es_29_1_1es_30_2_1QNode_Int_bufchan_d;
  
  /* dcon (Ty CTf_f_Int_Int,
      Dcon Lcall_f_f_Int_Int0) : [(lizzieLet44_4Lcall_f_f_Int_Int1,Pointer_QTree_Int),
                                  (es_29_destruct,Pointer_QTree_Int),
                                  (es_30_1_destruct,Pointer_QTree_Int),
                                  (sc_0_13_destruct,Pointer_CTf_f_Int_Int)] > (lizzieLet44_4Lcall_f_f_Int_Int1_1es_29_1es_30_1_1sc_0_13_1Lcall_f_f_Int_Int0,CTf_f_Int_Int) */
  assign lizzieLet44_4Lcall_f_f_Int_Int1_1es_29_1es_30_1_1sc_0_13_1Lcall_f_f_Int_Int0_d = Lcall_f_f_Int_Int0_dc((& {lizzieLet44_4Lcall_f_f_Int_Int1_d[0],
                                                                                                                    es_29_destruct_d[0],
                                                                                                                    es_30_1_destruct_d[0],
                                                                                                                    sc_0_13_destruct_d[0]}), lizzieLet44_4Lcall_f_f_Int_Int1_d, es_29_destruct_d, es_30_1_destruct_d, sc_0_13_destruct_d);
  assign {lizzieLet44_4Lcall_f_f_Int_Int1_r,
          es_29_destruct_r,
          es_30_1_destruct_r,
          sc_0_13_destruct_r} = {4 {(lizzieLet44_4Lcall_f_f_Int_Int1_1es_29_1es_30_1_1sc_0_13_1Lcall_f_f_Int_Int0_r && lizzieLet44_4Lcall_f_f_Int_Int1_1es_29_1es_30_1_1sc_0_13_1Lcall_f_f_Int_Int0_d[0])}};
  
  /* buf (Ty CTf_f_Int_Int) : (lizzieLet44_4Lcall_f_f_Int_Int1_1es_29_1es_30_1_1sc_0_13_1Lcall_f_f_Int_Int0,CTf_f_Int_Int) > (lizzieLet47_1_argbuf,CTf_f_Int_Int) */
  CTf_f_Int_Int_t lizzieLet44_4Lcall_f_f_Int_Int1_1es_29_1es_30_1_1sc_0_13_1Lcall_f_f_Int_Int0_bufchan_d;
  logic lizzieLet44_4Lcall_f_f_Int_Int1_1es_29_1es_30_1_1sc_0_13_1Lcall_f_f_Int_Int0_bufchan_r;
  assign lizzieLet44_4Lcall_f_f_Int_Int1_1es_29_1es_30_1_1sc_0_13_1Lcall_f_f_Int_Int0_r = ((! lizzieLet44_4Lcall_f_f_Int_Int1_1es_29_1es_30_1_1sc_0_13_1Lcall_f_f_Int_Int0_bufchan_d[0]) || lizzieLet44_4Lcall_f_f_Int_Int1_1es_29_1es_30_1_1sc_0_13_1Lcall_f_f_Int_Int0_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet44_4Lcall_f_f_Int_Int1_1es_29_1es_30_1_1sc_0_13_1Lcall_f_f_Int_Int0_bufchan_d <= {115'd0,
                                                                                                 1'd0};
    else
      if (lizzieLet44_4Lcall_f_f_Int_Int1_1es_29_1es_30_1_1sc_0_13_1Lcall_f_f_Int_Int0_r)
        lizzieLet44_4Lcall_f_f_Int_Int1_1es_29_1es_30_1_1sc_0_13_1Lcall_f_f_Int_Int0_bufchan_d <= lizzieLet44_4Lcall_f_f_Int_Int1_1es_29_1es_30_1_1sc_0_13_1Lcall_f_f_Int_Int0_d;
  CTf_f_Int_Int_t lizzieLet44_4Lcall_f_f_Int_Int1_1es_29_1es_30_1_1sc_0_13_1Lcall_f_f_Int_Int0_bufchan_buf;
  assign lizzieLet44_4Lcall_f_f_Int_Int1_1es_29_1es_30_1_1sc_0_13_1Lcall_f_f_Int_Int0_bufchan_r = (! lizzieLet44_4Lcall_f_f_Int_Int1_1es_29_1es_30_1_1sc_0_13_1Lcall_f_f_Int_Int0_bufchan_buf[0]);
  assign lizzieLet47_1_argbuf_d = (lizzieLet44_4Lcall_f_f_Int_Int1_1es_29_1es_30_1_1sc_0_13_1Lcall_f_f_Int_Int0_bufchan_buf[0] ? lizzieLet44_4Lcall_f_f_Int_Int1_1es_29_1es_30_1_1sc_0_13_1Lcall_f_f_Int_Int0_bufchan_buf :
                                   lizzieLet44_4Lcall_f_f_Int_Int1_1es_29_1es_30_1_1sc_0_13_1Lcall_f_f_Int_Int0_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet44_4Lcall_f_f_Int_Int1_1es_29_1es_30_1_1sc_0_13_1Lcall_f_f_Int_Int0_bufchan_buf <= {115'd0,
                                                                                                   1'd0};
    else
      if ((lizzieLet47_1_argbuf_r && lizzieLet44_4Lcall_f_f_Int_Int1_1es_29_1es_30_1_1sc_0_13_1Lcall_f_f_Int_Int0_bufchan_buf[0]))
        lizzieLet44_4Lcall_f_f_Int_Int1_1es_29_1es_30_1_1sc_0_13_1Lcall_f_f_Int_Int0_bufchan_buf <= {115'd0,
                                                                                                     1'd0};
      else if (((! lizzieLet47_1_argbuf_r) && (! lizzieLet44_4Lcall_f_f_Int_Int1_1es_29_1es_30_1_1sc_0_13_1Lcall_f_f_Int_Int0_bufchan_buf[0])))
        lizzieLet44_4Lcall_f_f_Int_Int1_1es_29_1es_30_1_1sc_0_13_1Lcall_f_f_Int_Int0_bufchan_buf <= lizzieLet44_4Lcall_f_f_Int_Int1_1es_29_1es_30_1_1sc_0_13_1Lcall_f_f_Int_Int0_bufchan_d;
  
  /* dcon (Ty CTf_f_Int_Int,
      Dcon Lcall_f_f_Int_Int1) : [(lizzieLet44_4Lcall_f_f_Int_Int2,Pointer_QTree_Int),
                                  (es_30_destruct,Pointer_QTree_Int),
                                  (sc_0_12_destruct,Pointer_CTf_f_Int_Int),
                                  (q1a8T_2_destruct,Pointer_QTree_Int),
                                  (t1a8Y_2_destruct,Pointer_QTree_Int),
                                  (is_z_mapa8E_3_1,MyDTInt_Bool),
                                  (op_mapa8F_3_1,MyDTInt_Int),
                                  (is_z_adda8G_3_1,MyDTInt_Bool),
                                  (op_adda8H_3_1,MyDTInt_Int_Int)] > (lizzieLet44_4Lcall_f_f_Int_Int2_1es_30_1sc_0_12_1q1a8T_2_1t1a8Y_2_1is_z_mapa8E_3_1op_mapa8F_3_1is_z_adda8G_3_1op_adda8H_3_1Lcall_f_f_Int_Int1,CTf_f_Int_Int) */
  assign lizzieLet44_4Lcall_f_f_Int_Int2_1es_30_1sc_0_12_1q1a8T_2_1t1a8Y_2_1is_z_mapa8E_3_1op_mapa8F_3_1is_z_adda8G_3_1op_adda8H_3_1Lcall_f_f_Int_Int1_d = Lcall_f_f_Int_Int1_dc((& {lizzieLet44_4Lcall_f_f_Int_Int2_d[0],
                                                                                                                                                                                     es_30_destruct_d[0],
                                                                                                                                                                                     sc_0_12_destruct_d[0],
                                                                                                                                                                                     q1a8T_2_destruct_d[0],
                                                                                                                                                                                     t1a8Y_2_destruct_d[0],
                                                                                                                                                                                     is_z_mapa8E_3_1_d[0],
                                                                                                                                                                                     op_mapa8F_3_1_d[0],
                                                                                                                                                                                     is_z_adda8G_3_1_d[0],
                                                                                                                                                                                     op_adda8H_3_1_d[0]}), lizzieLet44_4Lcall_f_f_Int_Int2_d, es_30_destruct_d, sc_0_12_destruct_d, q1a8T_2_destruct_d, t1a8Y_2_destruct_d, is_z_mapa8E_3_1_d, op_mapa8F_3_1_d, is_z_adda8G_3_1_d, op_adda8H_3_1_d);
  assign {lizzieLet44_4Lcall_f_f_Int_Int2_r,
          es_30_destruct_r,
          sc_0_12_destruct_r,
          q1a8T_2_destruct_r,
          t1a8Y_2_destruct_r,
          is_z_mapa8E_3_1_r,
          op_mapa8F_3_1_r,
          is_z_adda8G_3_1_r,
          op_adda8H_3_1_r} = {9 {(lizzieLet44_4Lcall_f_f_Int_Int2_1es_30_1sc_0_12_1q1a8T_2_1t1a8Y_2_1is_z_mapa8E_3_1op_mapa8F_3_1is_z_adda8G_3_1op_adda8H_3_1Lcall_f_f_Int_Int1_r && lizzieLet44_4Lcall_f_f_Int_Int2_1es_30_1sc_0_12_1q1a8T_2_1t1a8Y_2_1is_z_mapa8E_3_1op_mapa8F_3_1is_z_adda8G_3_1op_adda8H_3_1Lcall_f_f_Int_Int1_d[0])}};
  
  /* buf (Ty CTf_f_Int_Int) : (lizzieLet44_4Lcall_f_f_Int_Int2_1es_30_1sc_0_12_1q1a8T_2_1t1a8Y_2_1is_z_mapa8E_3_1op_mapa8F_3_1is_z_adda8G_3_1op_adda8H_3_1Lcall_f_f_Int_Int1,CTf_f_Int_Int) > (lizzieLet46_1_argbuf,CTf_f_Int_Int) */
  CTf_f_Int_Int_t lizzieLet44_4Lcall_f_f_Int_Int2_1es_30_1sc_0_12_1q1a8T_2_1t1a8Y_2_1is_z_mapa8E_3_1op_mapa8F_3_1is_z_adda8G_3_1op_adda8H_3_1Lcall_f_f_Int_Int1_bufchan_d;
  logic lizzieLet44_4Lcall_f_f_Int_Int2_1es_30_1sc_0_12_1q1a8T_2_1t1a8Y_2_1is_z_mapa8E_3_1op_mapa8F_3_1is_z_adda8G_3_1op_adda8H_3_1Lcall_f_f_Int_Int1_bufchan_r;
  assign lizzieLet44_4Lcall_f_f_Int_Int2_1es_30_1sc_0_12_1q1a8T_2_1t1a8Y_2_1is_z_mapa8E_3_1op_mapa8F_3_1is_z_adda8G_3_1op_adda8H_3_1Lcall_f_f_Int_Int1_r = ((! lizzieLet44_4Lcall_f_f_Int_Int2_1es_30_1sc_0_12_1q1a8T_2_1t1a8Y_2_1is_z_mapa8E_3_1op_mapa8F_3_1is_z_adda8G_3_1op_adda8H_3_1Lcall_f_f_Int_Int1_bufchan_d[0]) || lizzieLet44_4Lcall_f_f_Int_Int2_1es_30_1sc_0_12_1q1a8T_2_1t1a8Y_2_1is_z_mapa8E_3_1op_mapa8F_3_1is_z_adda8G_3_1op_adda8H_3_1Lcall_f_f_Int_Int1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet44_4Lcall_f_f_Int_Int2_1es_30_1sc_0_12_1q1a8T_2_1t1a8Y_2_1is_z_mapa8E_3_1op_mapa8F_3_1is_z_adda8G_3_1op_adda8H_3_1Lcall_f_f_Int_Int1_bufchan_d <= {115'd0,
                                                                                                                                                                  1'd0};
    else
      if (lizzieLet44_4Lcall_f_f_Int_Int2_1es_30_1sc_0_12_1q1a8T_2_1t1a8Y_2_1is_z_mapa8E_3_1op_mapa8F_3_1is_z_adda8G_3_1op_adda8H_3_1Lcall_f_f_Int_Int1_r)
        lizzieLet44_4Lcall_f_f_Int_Int2_1es_30_1sc_0_12_1q1a8T_2_1t1a8Y_2_1is_z_mapa8E_3_1op_mapa8F_3_1is_z_adda8G_3_1op_adda8H_3_1Lcall_f_f_Int_Int1_bufchan_d <= lizzieLet44_4Lcall_f_f_Int_Int2_1es_30_1sc_0_12_1q1a8T_2_1t1a8Y_2_1is_z_mapa8E_3_1op_mapa8F_3_1is_z_adda8G_3_1op_adda8H_3_1Lcall_f_f_Int_Int1_d;
  CTf_f_Int_Int_t lizzieLet44_4Lcall_f_f_Int_Int2_1es_30_1sc_0_12_1q1a8T_2_1t1a8Y_2_1is_z_mapa8E_3_1op_mapa8F_3_1is_z_adda8G_3_1op_adda8H_3_1Lcall_f_f_Int_Int1_bufchan_buf;
  assign lizzieLet44_4Lcall_f_f_Int_Int2_1es_30_1sc_0_12_1q1a8T_2_1t1a8Y_2_1is_z_mapa8E_3_1op_mapa8F_3_1is_z_adda8G_3_1op_adda8H_3_1Lcall_f_f_Int_Int1_bufchan_r = (! lizzieLet44_4Lcall_f_f_Int_Int2_1es_30_1sc_0_12_1q1a8T_2_1t1a8Y_2_1is_z_mapa8E_3_1op_mapa8F_3_1is_z_adda8G_3_1op_adda8H_3_1Lcall_f_f_Int_Int1_bufchan_buf[0]);
  assign lizzieLet46_1_argbuf_d = (lizzieLet44_4Lcall_f_f_Int_Int2_1es_30_1sc_0_12_1q1a8T_2_1t1a8Y_2_1is_z_mapa8E_3_1op_mapa8F_3_1is_z_adda8G_3_1op_adda8H_3_1Lcall_f_f_Int_Int1_bufchan_buf[0] ? lizzieLet44_4Lcall_f_f_Int_Int2_1es_30_1sc_0_12_1q1a8T_2_1t1a8Y_2_1is_z_mapa8E_3_1op_mapa8F_3_1is_z_adda8G_3_1op_adda8H_3_1Lcall_f_f_Int_Int1_bufchan_buf :
                                   lizzieLet44_4Lcall_f_f_Int_Int2_1es_30_1sc_0_12_1q1a8T_2_1t1a8Y_2_1is_z_mapa8E_3_1op_mapa8F_3_1is_z_adda8G_3_1op_adda8H_3_1Lcall_f_f_Int_Int1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet44_4Lcall_f_f_Int_Int2_1es_30_1sc_0_12_1q1a8T_2_1t1a8Y_2_1is_z_mapa8E_3_1op_mapa8F_3_1is_z_adda8G_3_1op_adda8H_3_1Lcall_f_f_Int_Int1_bufchan_buf <= {115'd0,
                                                                                                                                                                    1'd0};
    else
      if ((lizzieLet46_1_argbuf_r && lizzieLet44_4Lcall_f_f_Int_Int2_1es_30_1sc_0_12_1q1a8T_2_1t1a8Y_2_1is_z_mapa8E_3_1op_mapa8F_3_1is_z_adda8G_3_1op_adda8H_3_1Lcall_f_f_Int_Int1_bufchan_buf[0]))
        lizzieLet44_4Lcall_f_f_Int_Int2_1es_30_1sc_0_12_1q1a8T_2_1t1a8Y_2_1is_z_mapa8E_3_1op_mapa8F_3_1is_z_adda8G_3_1op_adda8H_3_1Lcall_f_f_Int_Int1_bufchan_buf <= {115'd0,
                                                                                                                                                                      1'd0};
      else if (((! lizzieLet46_1_argbuf_r) && (! lizzieLet44_4Lcall_f_f_Int_Int2_1es_30_1sc_0_12_1q1a8T_2_1t1a8Y_2_1is_z_mapa8E_3_1op_mapa8F_3_1is_z_adda8G_3_1op_adda8H_3_1Lcall_f_f_Int_Int1_bufchan_buf[0])))
        lizzieLet44_4Lcall_f_f_Int_Int2_1es_30_1sc_0_12_1q1a8T_2_1t1a8Y_2_1is_z_mapa8E_3_1op_mapa8F_3_1is_z_adda8G_3_1op_adda8H_3_1Lcall_f_f_Int_Int1_bufchan_buf <= lizzieLet44_4Lcall_f_f_Int_Int2_1es_30_1sc_0_12_1q1a8T_2_1t1a8Y_2_1is_z_mapa8E_3_1op_mapa8F_3_1is_z_adda8G_3_1op_adda8H_3_1Lcall_f_f_Int_Int1_bufchan_d;
  
  /* dcon (Ty CTf_f_Int_Int,
      Dcon Lcall_f_f_Int_Int2) : [(lizzieLet44_4Lcall_f_f_Int_Int3,Pointer_QTree_Int),
                                  (sc_0_11_destruct,Pointer_CTf_f_Int_Int),
                                  (q1a8T_1_destruct,Pointer_QTree_Int),
                                  (t1a8Y_1_destruct,Pointer_QTree_Int),
                                  (is_z_mapa8E_2_1,MyDTInt_Bool),
                                  (op_mapa8F_2_1,MyDTInt_Int),
                                  (is_z_adda8G_2_1,MyDTInt_Bool),
                                  (op_adda8H_2_1,MyDTInt_Int_Int),
                                  (q2a8U_1_destruct,Pointer_QTree_Int),
                                  (t2a8Z_1_destruct,Pointer_QTree_Int)] > (lizzieLet44_4Lcall_f_f_Int_Int3_1sc_0_11_1q1a8T_1_1t1a8Y_1_1is_z_mapa8E_2_1op_mapa8F_2_1is_z_adda8G_2_1op_adda8H_2_1q2a8U_1_1t2a8Z_1_1Lcall_f_f_Int_Int2,CTf_f_Int_Int) */
  assign lizzieLet44_4Lcall_f_f_Int_Int3_1sc_0_11_1q1a8T_1_1t1a8Y_1_1is_z_mapa8E_2_1op_mapa8F_2_1is_z_adda8G_2_1op_adda8H_2_1q2a8U_1_1t2a8Z_1_1Lcall_f_f_Int_Int2_d = Lcall_f_f_Int_Int2_dc((& {lizzieLet44_4Lcall_f_f_Int_Int3_d[0],
                                                                                                                                                                                                sc_0_11_destruct_d[0],
                                                                                                                                                                                                q1a8T_1_destruct_d[0],
                                                                                                                                                                                                t1a8Y_1_destruct_d[0],
                                                                                                                                                                                                is_z_mapa8E_2_1_d[0],
                                                                                                                                                                                                op_mapa8F_2_1_d[0],
                                                                                                                                                                                                is_z_adda8G_2_1_d[0],
                                                                                                                                                                                                op_adda8H_2_1_d[0],
                                                                                                                                                                                                q2a8U_1_destruct_d[0],
                                                                                                                                                                                                t2a8Z_1_destruct_d[0]}), lizzieLet44_4Lcall_f_f_Int_Int3_d, sc_0_11_destruct_d, q1a8T_1_destruct_d, t1a8Y_1_destruct_d, is_z_mapa8E_2_1_d, op_mapa8F_2_1_d, is_z_adda8G_2_1_d, op_adda8H_2_1_d, q2a8U_1_destruct_d, t2a8Z_1_destruct_d);
  assign {lizzieLet44_4Lcall_f_f_Int_Int3_r,
          sc_0_11_destruct_r,
          q1a8T_1_destruct_r,
          t1a8Y_1_destruct_r,
          is_z_mapa8E_2_1_r,
          op_mapa8F_2_1_r,
          is_z_adda8G_2_1_r,
          op_adda8H_2_1_r,
          q2a8U_1_destruct_r,
          t2a8Z_1_destruct_r} = {10 {(lizzieLet44_4Lcall_f_f_Int_Int3_1sc_0_11_1q1a8T_1_1t1a8Y_1_1is_z_mapa8E_2_1op_mapa8F_2_1is_z_adda8G_2_1op_adda8H_2_1q2a8U_1_1t2a8Z_1_1Lcall_f_f_Int_Int2_r && lizzieLet44_4Lcall_f_f_Int_Int3_1sc_0_11_1q1a8T_1_1t1a8Y_1_1is_z_mapa8E_2_1op_mapa8F_2_1is_z_adda8G_2_1op_adda8H_2_1q2a8U_1_1t2a8Z_1_1Lcall_f_f_Int_Int2_d[0])}};
  
  /* buf (Ty CTf_f_Int_Int) : (lizzieLet44_4Lcall_f_f_Int_Int3_1sc_0_11_1q1a8T_1_1t1a8Y_1_1is_z_mapa8E_2_1op_mapa8F_2_1is_z_adda8G_2_1op_adda8H_2_1q2a8U_1_1t2a8Z_1_1Lcall_f_f_Int_Int2,CTf_f_Int_Int) > (lizzieLet45_1_argbuf,CTf_f_Int_Int) */
  CTf_f_Int_Int_t lizzieLet44_4Lcall_f_f_Int_Int3_1sc_0_11_1q1a8T_1_1t1a8Y_1_1is_z_mapa8E_2_1op_mapa8F_2_1is_z_adda8G_2_1op_adda8H_2_1q2a8U_1_1t2a8Z_1_1Lcall_f_f_Int_Int2_bufchan_d;
  logic lizzieLet44_4Lcall_f_f_Int_Int3_1sc_0_11_1q1a8T_1_1t1a8Y_1_1is_z_mapa8E_2_1op_mapa8F_2_1is_z_adda8G_2_1op_adda8H_2_1q2a8U_1_1t2a8Z_1_1Lcall_f_f_Int_Int2_bufchan_r;
  assign lizzieLet44_4Lcall_f_f_Int_Int3_1sc_0_11_1q1a8T_1_1t1a8Y_1_1is_z_mapa8E_2_1op_mapa8F_2_1is_z_adda8G_2_1op_adda8H_2_1q2a8U_1_1t2a8Z_1_1Lcall_f_f_Int_Int2_r = ((! lizzieLet44_4Lcall_f_f_Int_Int3_1sc_0_11_1q1a8T_1_1t1a8Y_1_1is_z_mapa8E_2_1op_mapa8F_2_1is_z_adda8G_2_1op_adda8H_2_1q2a8U_1_1t2a8Z_1_1Lcall_f_f_Int_Int2_bufchan_d[0]) || lizzieLet44_4Lcall_f_f_Int_Int3_1sc_0_11_1q1a8T_1_1t1a8Y_1_1is_z_mapa8E_2_1op_mapa8F_2_1is_z_adda8G_2_1op_adda8H_2_1q2a8U_1_1t2a8Z_1_1Lcall_f_f_Int_Int2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet44_4Lcall_f_f_Int_Int3_1sc_0_11_1q1a8T_1_1t1a8Y_1_1is_z_mapa8E_2_1op_mapa8F_2_1is_z_adda8G_2_1op_adda8H_2_1q2a8U_1_1t2a8Z_1_1Lcall_f_f_Int_Int2_bufchan_d <= {115'd0,
                                                                                                                                                                             1'd0};
    else
      if (lizzieLet44_4Lcall_f_f_Int_Int3_1sc_0_11_1q1a8T_1_1t1a8Y_1_1is_z_mapa8E_2_1op_mapa8F_2_1is_z_adda8G_2_1op_adda8H_2_1q2a8U_1_1t2a8Z_1_1Lcall_f_f_Int_Int2_r)
        lizzieLet44_4Lcall_f_f_Int_Int3_1sc_0_11_1q1a8T_1_1t1a8Y_1_1is_z_mapa8E_2_1op_mapa8F_2_1is_z_adda8G_2_1op_adda8H_2_1q2a8U_1_1t2a8Z_1_1Lcall_f_f_Int_Int2_bufchan_d <= lizzieLet44_4Lcall_f_f_Int_Int3_1sc_0_11_1q1a8T_1_1t1a8Y_1_1is_z_mapa8E_2_1op_mapa8F_2_1is_z_adda8G_2_1op_adda8H_2_1q2a8U_1_1t2a8Z_1_1Lcall_f_f_Int_Int2_d;
  CTf_f_Int_Int_t lizzieLet44_4Lcall_f_f_Int_Int3_1sc_0_11_1q1a8T_1_1t1a8Y_1_1is_z_mapa8E_2_1op_mapa8F_2_1is_z_adda8G_2_1op_adda8H_2_1q2a8U_1_1t2a8Z_1_1Lcall_f_f_Int_Int2_bufchan_buf;
  assign lizzieLet44_4Lcall_f_f_Int_Int3_1sc_0_11_1q1a8T_1_1t1a8Y_1_1is_z_mapa8E_2_1op_mapa8F_2_1is_z_adda8G_2_1op_adda8H_2_1q2a8U_1_1t2a8Z_1_1Lcall_f_f_Int_Int2_bufchan_r = (! lizzieLet44_4Lcall_f_f_Int_Int3_1sc_0_11_1q1a8T_1_1t1a8Y_1_1is_z_mapa8E_2_1op_mapa8F_2_1is_z_adda8G_2_1op_adda8H_2_1q2a8U_1_1t2a8Z_1_1Lcall_f_f_Int_Int2_bufchan_buf[0]);
  assign lizzieLet45_1_argbuf_d = (lizzieLet44_4Lcall_f_f_Int_Int3_1sc_0_11_1q1a8T_1_1t1a8Y_1_1is_z_mapa8E_2_1op_mapa8F_2_1is_z_adda8G_2_1op_adda8H_2_1q2a8U_1_1t2a8Z_1_1Lcall_f_f_Int_Int2_bufchan_buf[0] ? lizzieLet44_4Lcall_f_f_Int_Int3_1sc_0_11_1q1a8T_1_1t1a8Y_1_1is_z_mapa8E_2_1op_mapa8F_2_1is_z_adda8G_2_1op_adda8H_2_1q2a8U_1_1t2a8Z_1_1Lcall_f_f_Int_Int2_bufchan_buf :
                                   lizzieLet44_4Lcall_f_f_Int_Int3_1sc_0_11_1q1a8T_1_1t1a8Y_1_1is_z_mapa8E_2_1op_mapa8F_2_1is_z_adda8G_2_1op_adda8H_2_1q2a8U_1_1t2a8Z_1_1Lcall_f_f_Int_Int2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet44_4Lcall_f_f_Int_Int3_1sc_0_11_1q1a8T_1_1t1a8Y_1_1is_z_mapa8E_2_1op_mapa8F_2_1is_z_adda8G_2_1op_adda8H_2_1q2a8U_1_1t2a8Z_1_1Lcall_f_f_Int_Int2_bufchan_buf <= {115'd0,
                                                                                                                                                                               1'd0};
    else
      if ((lizzieLet45_1_argbuf_r && lizzieLet44_4Lcall_f_f_Int_Int3_1sc_0_11_1q1a8T_1_1t1a8Y_1_1is_z_mapa8E_2_1op_mapa8F_2_1is_z_adda8G_2_1op_adda8H_2_1q2a8U_1_1t2a8Z_1_1Lcall_f_f_Int_Int2_bufchan_buf[0]))
        lizzieLet44_4Lcall_f_f_Int_Int3_1sc_0_11_1q1a8T_1_1t1a8Y_1_1is_z_mapa8E_2_1op_mapa8F_2_1is_z_adda8G_2_1op_adda8H_2_1q2a8U_1_1t2a8Z_1_1Lcall_f_f_Int_Int2_bufchan_buf <= {115'd0,
                                                                                                                                                                                 1'd0};
      else if (((! lizzieLet45_1_argbuf_r) && (! lizzieLet44_4Lcall_f_f_Int_Int3_1sc_0_11_1q1a8T_1_1t1a8Y_1_1is_z_mapa8E_2_1op_mapa8F_2_1is_z_adda8G_2_1op_adda8H_2_1q2a8U_1_1t2a8Z_1_1Lcall_f_f_Int_Int2_bufchan_buf[0])))
        lizzieLet44_4Lcall_f_f_Int_Int3_1sc_0_11_1q1a8T_1_1t1a8Y_1_1is_z_mapa8E_2_1op_mapa8F_2_1is_z_adda8G_2_1op_adda8H_2_1q2a8U_1_1t2a8Z_1_1Lcall_f_f_Int_Int2_bufchan_buf <= lizzieLet44_4Lcall_f_f_Int_Int3_1sc_0_11_1q1a8T_1_1t1a8Y_1_1is_z_mapa8E_2_1op_mapa8F_2_1is_z_adda8G_2_1op_adda8H_2_1q2a8U_1_1t2a8Z_1_1Lcall_f_f_Int_Int2_bufchan_d;
  
  /* fork (Ty Pointer_QTree_Int) : (lizzieLet44_4Lf_f_Int_Intsbos,Pointer_QTree_Int) > [(lizzieLet44_4Lf_f_Int_Intsbos_1_merge_merge_merge_fork_1,Pointer_QTree_Int),
                                                                                   (lizzieLet44_4Lf_f_Int_Intsbos_1_merge_merge_merge_fork_2,Pointer_QTree_Int)] */
  logic [1:0] lizzieLet44_4Lf_f_Int_Intsbos_emitted;
  logic [1:0] lizzieLet44_4Lf_f_Int_Intsbos_done;
  assign lizzieLet44_4Lf_f_Int_Intsbos_1_merge_merge_merge_fork_1_d = {lizzieLet44_4Lf_f_Int_Intsbos_d[16:1],
                                                                       (lizzieLet44_4Lf_f_Int_Intsbos_d[0] && (! lizzieLet44_4Lf_f_Int_Intsbos_emitted[0]))};
  assign lizzieLet44_4Lf_f_Int_Intsbos_1_merge_merge_merge_fork_2_d = {lizzieLet44_4Lf_f_Int_Intsbos_d[16:1],
                                                                       (lizzieLet44_4Lf_f_Int_Intsbos_d[0] && (! lizzieLet44_4Lf_f_Int_Intsbos_emitted[1]))};
  assign lizzieLet44_4Lf_f_Int_Intsbos_done = (lizzieLet44_4Lf_f_Int_Intsbos_emitted | ({lizzieLet44_4Lf_f_Int_Intsbos_1_merge_merge_merge_fork_2_d[0],
                                                                                         lizzieLet44_4Lf_f_Int_Intsbos_1_merge_merge_merge_fork_1_d[0]} & {lizzieLet44_4Lf_f_Int_Intsbos_1_merge_merge_merge_fork_2_r,
                                                                                                                                                           lizzieLet44_4Lf_f_Int_Intsbos_1_merge_merge_merge_fork_1_r}));
  assign lizzieLet44_4Lf_f_Int_Intsbos_r = (& lizzieLet44_4Lf_f_Int_Intsbos_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet44_4Lf_f_Int_Intsbos_emitted <= 2'd0;
    else
      lizzieLet44_4Lf_f_Int_Intsbos_emitted <= (lizzieLet44_4Lf_f_Int_Intsbos_r ? 2'd0 :
                                                lizzieLet44_4Lf_f_Int_Intsbos_done);
  
  /* togo (Ty Pointer_QTree_Int) : (lizzieLet44_4Lf_f_Int_Intsbos_1_merge_merge_merge_fork_1,Pointer_QTree_Int) > (call_f_f_Int_Int_goConst,Go) */
  assign call_f_f_Int_Int_goConst_d = lizzieLet44_4Lf_f_Int_Intsbos_1_merge_merge_merge_fork_1_d[0];
  assign lizzieLet44_4Lf_f_Int_Intsbos_1_merge_merge_merge_fork_1_r = call_f_f_Int_Int_goConst_r;
  
  /* buf (Ty Pointer_QTree_Int) : (lizzieLet44_4Lf_f_Int_Intsbos_1_merge_merge_merge_fork_2,Pointer_QTree_Int) > (f_f_Int_Int_resbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t lizzieLet44_4Lf_f_Int_Intsbos_1_merge_merge_merge_fork_2_bufchan_d;
  logic lizzieLet44_4Lf_f_Int_Intsbos_1_merge_merge_merge_fork_2_bufchan_r;
  assign lizzieLet44_4Lf_f_Int_Intsbos_1_merge_merge_merge_fork_2_r = ((! lizzieLet44_4Lf_f_Int_Intsbos_1_merge_merge_merge_fork_2_bufchan_d[0]) || lizzieLet44_4Lf_f_Int_Intsbos_1_merge_merge_merge_fork_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet44_4Lf_f_Int_Intsbos_1_merge_merge_merge_fork_2_bufchan_d <= {16'd0,
                                                                             1'd0};
    else
      if (lizzieLet44_4Lf_f_Int_Intsbos_1_merge_merge_merge_fork_2_r)
        lizzieLet44_4Lf_f_Int_Intsbos_1_merge_merge_merge_fork_2_bufchan_d <= lizzieLet44_4Lf_f_Int_Intsbos_1_merge_merge_merge_fork_2_d;
  Pointer_QTree_Int_t lizzieLet44_4Lf_f_Int_Intsbos_1_merge_merge_merge_fork_2_bufchan_buf;
  assign lizzieLet44_4Lf_f_Int_Intsbos_1_merge_merge_merge_fork_2_bufchan_r = (! lizzieLet44_4Lf_f_Int_Intsbos_1_merge_merge_merge_fork_2_bufchan_buf[0]);
  assign f_f_Int_Int_resbuf_d = (lizzieLet44_4Lf_f_Int_Intsbos_1_merge_merge_merge_fork_2_bufchan_buf[0] ? lizzieLet44_4Lf_f_Int_Intsbos_1_merge_merge_merge_fork_2_bufchan_buf :
                                 lizzieLet44_4Lf_f_Int_Intsbos_1_merge_merge_merge_fork_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet44_4Lf_f_Int_Intsbos_1_merge_merge_merge_fork_2_bufchan_buf <= {16'd0,
                                                                               1'd0};
    else
      if ((f_f_Int_Int_resbuf_r && lizzieLet44_4Lf_f_Int_Intsbos_1_merge_merge_merge_fork_2_bufchan_buf[0]))
        lizzieLet44_4Lf_f_Int_Intsbos_1_merge_merge_merge_fork_2_bufchan_buf <= {16'd0,
                                                                                 1'd0};
      else if (((! f_f_Int_Int_resbuf_r) && (! lizzieLet44_4Lf_f_Int_Intsbos_1_merge_merge_merge_fork_2_bufchan_buf[0])))
        lizzieLet44_4Lf_f_Int_Intsbos_1_merge_merge_merge_fork_2_bufchan_buf <= lizzieLet44_4Lf_f_Int_Intsbos_1_merge_merge_merge_fork_2_bufchan_d;
  
  /* destruct (Ty QTree_Int,
          Dcon QNode_Int) : (lizzieLet4_1QNode_Int,QTree_Int) > [(q1a84_destruct,Pointer_QTree_Int),
                                                                 (q2a85_destruct,Pointer_QTree_Int),
                                                                 (q3a86_destruct,Pointer_QTree_Int),
                                                                 (q4a87_destruct,Pointer_QTree_Int)] */
  logic [3:0] lizzieLet4_1QNode_Int_emitted;
  logic [3:0] lizzieLet4_1QNode_Int_done;
  assign q1a84_destruct_d = {lizzieLet4_1QNode_Int_d[18:3],
                             (lizzieLet4_1QNode_Int_d[0] && (! lizzieLet4_1QNode_Int_emitted[0]))};
  assign q2a85_destruct_d = {lizzieLet4_1QNode_Int_d[34:19],
                             (lizzieLet4_1QNode_Int_d[0] && (! lizzieLet4_1QNode_Int_emitted[1]))};
  assign q3a86_destruct_d = {lizzieLet4_1QNode_Int_d[50:35],
                             (lizzieLet4_1QNode_Int_d[0] && (! lizzieLet4_1QNode_Int_emitted[2]))};
  assign q4a87_destruct_d = {lizzieLet4_1QNode_Int_d[66:51],
                             (lizzieLet4_1QNode_Int_d[0] && (! lizzieLet4_1QNode_Int_emitted[3]))};
  assign lizzieLet4_1QNode_Int_done = (lizzieLet4_1QNode_Int_emitted | ({q4a87_destruct_d[0],
                                                                         q3a86_destruct_d[0],
                                                                         q2a85_destruct_d[0],
                                                                         q1a84_destruct_d[0]} & {q4a87_destruct_r,
                                                                                                 q3a86_destruct_r,
                                                                                                 q2a85_destruct_r,
                                                                                                 q1a84_destruct_r}));
  assign lizzieLet4_1QNode_Int_r = (& lizzieLet4_1QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_1QNode_Int_emitted <= 4'd0;
    else
      lizzieLet4_1QNode_Int_emitted <= (lizzieLet4_1QNode_Int_r ? 4'd0 :
                                        lizzieLet4_1QNode_Int_done);
  
  /* demux (Ty QTree_Int,
       Ty QTree_Int) : (lizzieLet4_2,QTree_Int) (lizzieLet4_1,QTree_Int) > [(_8,QTree_Int),
                                                                            (_7,QTree_Int),
                                                                            (lizzieLet4_1QNode_Int,QTree_Int),
                                                                            (_6,QTree_Int)] */
  logic [3:0] lizzieLet4_1_onehotd;
  always_comb
    if ((lizzieLet4_2_d[0] && lizzieLet4_1_d[0]))
      unique case (lizzieLet4_2_d[2:1])
        2'd0: lizzieLet4_1_onehotd = 4'd1;
        2'd1: lizzieLet4_1_onehotd = 4'd2;
        2'd2: lizzieLet4_1_onehotd = 4'd4;
        2'd3: lizzieLet4_1_onehotd = 4'd8;
        default: lizzieLet4_1_onehotd = 4'd0;
      endcase
    else lizzieLet4_1_onehotd = 4'd0;
  assign _8_d = {lizzieLet4_1_d[66:1], lizzieLet4_1_onehotd[0]};
  assign _7_d = {lizzieLet4_1_d[66:1], lizzieLet4_1_onehotd[1]};
  assign lizzieLet4_1QNode_Int_d = {lizzieLet4_1_d[66:1],
                                    lizzieLet4_1_onehotd[2]};
  assign _6_d = {lizzieLet4_1_d[66:1], lizzieLet4_1_onehotd[3]};
  assign lizzieLet4_1_r = (| (lizzieLet4_1_onehotd & {_6_r,
                                                      lizzieLet4_1QNode_Int_r,
                                                      _7_r,
                                                      _8_r}));
  assign lizzieLet4_2_r = lizzieLet4_1_r;
  
  /* demux (Ty QTree_Int,
       Ty Go) : (lizzieLet4_3,QTree_Int) (go_10_goMux_data,Go) > [(lizzieLet4_3QNone_Int,Go),
                                                                  (lizzieLet4_3QVal_Int,Go),
                                                                  (lizzieLet4_3QNode_Int,Go),
                                                                  (lizzieLet4_3QError_Int,Go)] */
  logic [3:0] go_10_goMux_data_onehotd;
  always_comb
    if ((lizzieLet4_3_d[0] && go_10_goMux_data_d[0]))
      unique case (lizzieLet4_3_d[2:1])
        2'd0: go_10_goMux_data_onehotd = 4'd1;
        2'd1: go_10_goMux_data_onehotd = 4'd2;
        2'd2: go_10_goMux_data_onehotd = 4'd4;
        2'd3: go_10_goMux_data_onehotd = 4'd8;
        default: go_10_goMux_data_onehotd = 4'd0;
      endcase
    else go_10_goMux_data_onehotd = 4'd0;
  assign lizzieLet4_3QNone_Int_d = go_10_goMux_data_onehotd[0];
  assign lizzieLet4_3QVal_Int_d = go_10_goMux_data_onehotd[1];
  assign lizzieLet4_3QNode_Int_d = go_10_goMux_data_onehotd[2];
  assign lizzieLet4_3QError_Int_d = go_10_goMux_data_onehotd[3];
  assign go_10_goMux_data_r = (| (go_10_goMux_data_onehotd & {lizzieLet4_3QError_Int_r,
                                                              lizzieLet4_3QNode_Int_r,
                                                              lizzieLet4_3QVal_Int_r,
                                                              lizzieLet4_3QNone_Int_r}));
  assign lizzieLet4_3_r = go_10_goMux_data_r;
  
  /* fork (Ty Go) : (lizzieLet4_3QError_Int,Go) > [(lizzieLet4_3QError_Int_1,Go),
                                              (lizzieLet4_3QError_Int_2,Go)] */
  logic [1:0] lizzieLet4_3QError_Int_emitted;
  logic [1:0] lizzieLet4_3QError_Int_done;
  assign lizzieLet4_3QError_Int_1_d = (lizzieLet4_3QError_Int_d[0] && (! lizzieLet4_3QError_Int_emitted[0]));
  assign lizzieLet4_3QError_Int_2_d = (lizzieLet4_3QError_Int_d[0] && (! lizzieLet4_3QError_Int_emitted[1]));
  assign lizzieLet4_3QError_Int_done = (lizzieLet4_3QError_Int_emitted | ({lizzieLet4_3QError_Int_2_d[0],
                                                                           lizzieLet4_3QError_Int_1_d[0]} & {lizzieLet4_3QError_Int_2_r,
                                                                                                             lizzieLet4_3QError_Int_1_r}));
  assign lizzieLet4_3QError_Int_r = (& lizzieLet4_3QError_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3QError_Int_emitted <= 2'd0;
    else
      lizzieLet4_3QError_Int_emitted <= (lizzieLet4_3QError_Int_r ? 2'd0 :
                                         lizzieLet4_3QError_Int_done);
  
  /* buf (Ty Go) : (lizzieLet4_3QError_Int_1,Go) > (lizzieLet4_3QError_Int_1_argbuf,Go) */
  Go_t lizzieLet4_3QError_Int_1_bufchan_d;
  logic lizzieLet4_3QError_Int_1_bufchan_r;
  assign lizzieLet4_3QError_Int_1_r = ((! lizzieLet4_3QError_Int_1_bufchan_d[0]) || lizzieLet4_3QError_Int_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3QError_Int_1_bufchan_d <= 1'd0;
    else
      if (lizzieLet4_3QError_Int_1_r)
        lizzieLet4_3QError_Int_1_bufchan_d <= lizzieLet4_3QError_Int_1_d;
  Go_t lizzieLet4_3QError_Int_1_bufchan_buf;
  assign lizzieLet4_3QError_Int_1_bufchan_r = (! lizzieLet4_3QError_Int_1_bufchan_buf[0]);
  assign lizzieLet4_3QError_Int_1_argbuf_d = (lizzieLet4_3QError_Int_1_bufchan_buf[0] ? lizzieLet4_3QError_Int_1_bufchan_buf :
                                              lizzieLet4_3QError_Int_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3QError_Int_1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet4_3QError_Int_1_argbuf_r && lizzieLet4_3QError_Int_1_bufchan_buf[0]))
        lizzieLet4_3QError_Int_1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet4_3QError_Int_1_argbuf_r) && (! lizzieLet4_3QError_Int_1_bufchan_buf[0])))
        lizzieLet4_3QError_Int_1_bufchan_buf <= lizzieLet4_3QError_Int_1_bufchan_d;
  
  /* const (Ty Int#,
       Lit 0) : (lizzieLet4_3QError_Int_1_argbuf,Go) > (lizzieLet4_3QError_Int_1_argbuf_0,Int#) */
  assign lizzieLet4_3QError_Int_1_argbuf_0_d = {32'd0,
                                                lizzieLet4_3QError_Int_1_argbuf_d[0]};
  assign lizzieLet4_3QError_Int_1_argbuf_r = lizzieLet4_3QError_Int_1_argbuf_0_r;
  
  /* buf (Ty Int#) : (lizzieLet4_3QError_Int_1_argbuf_0,Int#) > (lizzieLet23_1_1_argbuf,Int#) */
  \Int#_t  lizzieLet4_3QError_Int_1_argbuf_0_bufchan_d;
  logic lizzieLet4_3QError_Int_1_argbuf_0_bufchan_r;
  assign lizzieLet4_3QError_Int_1_argbuf_0_r = ((! lizzieLet4_3QError_Int_1_argbuf_0_bufchan_d[0]) || lizzieLet4_3QError_Int_1_argbuf_0_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_3QError_Int_1_argbuf_0_bufchan_d <= {32'd0, 1'd0};
    else
      if (lizzieLet4_3QError_Int_1_argbuf_0_r)
        lizzieLet4_3QError_Int_1_argbuf_0_bufchan_d <= lizzieLet4_3QError_Int_1_argbuf_0_d;
  \Int#_t  lizzieLet4_3QError_Int_1_argbuf_0_bufchan_buf;
  assign lizzieLet4_3QError_Int_1_argbuf_0_bufchan_r = (! lizzieLet4_3QError_Int_1_argbuf_0_bufchan_buf[0]);
  assign lizzieLet23_1_1_argbuf_d = (lizzieLet4_3QError_Int_1_argbuf_0_bufchan_buf[0] ? lizzieLet4_3QError_Int_1_argbuf_0_bufchan_buf :
                                     lizzieLet4_3QError_Int_1_argbuf_0_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_3QError_Int_1_argbuf_0_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((lizzieLet23_1_1_argbuf_r && lizzieLet4_3QError_Int_1_argbuf_0_bufchan_buf[0]))
        lizzieLet4_3QError_Int_1_argbuf_0_bufchan_buf <= {32'd0, 1'd0};
      else if (((! lizzieLet23_1_1_argbuf_r) && (! lizzieLet4_3QError_Int_1_argbuf_0_bufchan_buf[0])))
        lizzieLet4_3QError_Int_1_argbuf_0_bufchan_buf <= lizzieLet4_3QError_Int_1_argbuf_0_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet4_3QError_Int_2,Go) > (lizzieLet4_3QError_Int_2_argbuf,Go) */
  Go_t lizzieLet4_3QError_Int_2_bufchan_d;
  logic lizzieLet4_3QError_Int_2_bufchan_r;
  assign lizzieLet4_3QError_Int_2_r = ((! lizzieLet4_3QError_Int_2_bufchan_d[0]) || lizzieLet4_3QError_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3QError_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet4_3QError_Int_2_r)
        lizzieLet4_3QError_Int_2_bufchan_d <= lizzieLet4_3QError_Int_2_d;
  Go_t lizzieLet4_3QError_Int_2_bufchan_buf;
  assign lizzieLet4_3QError_Int_2_bufchan_r = (! lizzieLet4_3QError_Int_2_bufchan_buf[0]);
  assign lizzieLet4_3QError_Int_2_argbuf_d = (lizzieLet4_3QError_Int_2_bufchan_buf[0] ? lizzieLet4_3QError_Int_2_bufchan_buf :
                                              lizzieLet4_3QError_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3QError_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet4_3QError_Int_2_argbuf_r && lizzieLet4_3QError_Int_2_bufchan_buf[0]))
        lizzieLet4_3QError_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet4_3QError_Int_2_argbuf_r) && (! lizzieLet4_3QError_Int_2_bufchan_buf[0])))
        lizzieLet4_3QError_Int_2_bufchan_buf <= lizzieLet4_3QError_Int_2_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet4_3QNode_Int,Go) > (lizzieLet4_3QNode_Int_1_argbuf,Go) */
  Go_t lizzieLet4_3QNode_Int_bufchan_d;
  logic lizzieLet4_3QNode_Int_bufchan_r;
  assign lizzieLet4_3QNode_Int_r = ((! lizzieLet4_3QNode_Int_bufchan_d[0]) || lizzieLet4_3QNode_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3QNode_Int_bufchan_d <= 1'd0;
    else
      if (lizzieLet4_3QNode_Int_r)
        lizzieLet4_3QNode_Int_bufchan_d <= lizzieLet4_3QNode_Int_d;
  Go_t lizzieLet4_3QNode_Int_bufchan_buf;
  assign lizzieLet4_3QNode_Int_bufchan_r = (! lizzieLet4_3QNode_Int_bufchan_buf[0]);
  assign lizzieLet4_3QNode_Int_1_argbuf_d = (lizzieLet4_3QNode_Int_bufchan_buf[0] ? lizzieLet4_3QNode_Int_bufchan_buf :
                                             lizzieLet4_3QNode_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3QNode_Int_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet4_3QNode_Int_1_argbuf_r && lizzieLet4_3QNode_Int_bufchan_buf[0]))
        lizzieLet4_3QNode_Int_bufchan_buf <= 1'd0;
      else if (((! lizzieLet4_3QNode_Int_1_argbuf_r) && (! lizzieLet4_3QNode_Int_bufchan_buf[0])))
        lizzieLet4_3QNode_Int_bufchan_buf <= lizzieLet4_3QNode_Int_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet4_3QNone_Int,Go) > [(lizzieLet4_3QNone_Int_1,Go),
                                             (lizzieLet4_3QNone_Int_2,Go)] */
  logic [1:0] lizzieLet4_3QNone_Int_emitted;
  logic [1:0] lizzieLet4_3QNone_Int_done;
  assign lizzieLet4_3QNone_Int_1_d = (lizzieLet4_3QNone_Int_d[0] && (! lizzieLet4_3QNone_Int_emitted[0]));
  assign lizzieLet4_3QNone_Int_2_d = (lizzieLet4_3QNone_Int_d[0] && (! lizzieLet4_3QNone_Int_emitted[1]));
  assign lizzieLet4_3QNone_Int_done = (lizzieLet4_3QNone_Int_emitted | ({lizzieLet4_3QNone_Int_2_d[0],
                                                                         lizzieLet4_3QNone_Int_1_d[0]} & {lizzieLet4_3QNone_Int_2_r,
                                                                                                          lizzieLet4_3QNone_Int_1_r}));
  assign lizzieLet4_3QNone_Int_r = (& lizzieLet4_3QNone_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3QNone_Int_emitted <= 2'd0;
    else
      lizzieLet4_3QNone_Int_emitted <= (lizzieLet4_3QNone_Int_r ? 2'd0 :
                                        lizzieLet4_3QNone_Int_done);
  
  /* buf (Ty Go) : (lizzieLet4_3QNone_Int_1,Go) > (lizzieLet4_3QNone_Int_1_argbuf,Go) */
  Go_t lizzieLet4_3QNone_Int_1_bufchan_d;
  logic lizzieLet4_3QNone_Int_1_bufchan_r;
  assign lizzieLet4_3QNone_Int_1_r = ((! lizzieLet4_3QNone_Int_1_bufchan_d[0]) || lizzieLet4_3QNone_Int_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3QNone_Int_1_bufchan_d <= 1'd0;
    else
      if (lizzieLet4_3QNone_Int_1_r)
        lizzieLet4_3QNone_Int_1_bufchan_d <= lizzieLet4_3QNone_Int_1_d;
  Go_t lizzieLet4_3QNone_Int_1_bufchan_buf;
  assign lizzieLet4_3QNone_Int_1_bufchan_r = (! lizzieLet4_3QNone_Int_1_bufchan_buf[0]);
  assign lizzieLet4_3QNone_Int_1_argbuf_d = (lizzieLet4_3QNone_Int_1_bufchan_buf[0] ? lizzieLet4_3QNone_Int_1_bufchan_buf :
                                             lizzieLet4_3QNone_Int_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3QNone_Int_1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet4_3QNone_Int_1_argbuf_r && lizzieLet4_3QNone_Int_1_bufchan_buf[0]))
        lizzieLet4_3QNone_Int_1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet4_3QNone_Int_1_argbuf_r) && (! lizzieLet4_3QNone_Int_1_bufchan_buf[0])))
        lizzieLet4_3QNone_Int_1_bufchan_buf <= lizzieLet4_3QNone_Int_1_bufchan_d;
  
  /* const (Ty Int#,
       Lit 0) : (lizzieLet4_3QNone_Int_1_argbuf,Go) > (lizzieLet4_3QNone_Int_1_argbuf_0,Int#) */
  assign lizzieLet4_3QNone_Int_1_argbuf_0_d = {32'd0,
                                               lizzieLet4_3QNone_Int_1_argbuf_d[0]};
  assign lizzieLet4_3QNone_Int_1_argbuf_r = lizzieLet4_3QNone_Int_1_argbuf_0_r;
  
  /* buf (Ty Int#) : (lizzieLet4_3QNone_Int_1_argbuf_0,Int#) > (lizzieLet23_1_argbuf,Int#) */
  \Int#_t  lizzieLet4_3QNone_Int_1_argbuf_0_bufchan_d;
  logic lizzieLet4_3QNone_Int_1_argbuf_0_bufchan_r;
  assign lizzieLet4_3QNone_Int_1_argbuf_0_r = ((! lizzieLet4_3QNone_Int_1_argbuf_0_bufchan_d[0]) || lizzieLet4_3QNone_Int_1_argbuf_0_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_3QNone_Int_1_argbuf_0_bufchan_d <= {32'd0, 1'd0};
    else
      if (lizzieLet4_3QNone_Int_1_argbuf_0_r)
        lizzieLet4_3QNone_Int_1_argbuf_0_bufchan_d <= lizzieLet4_3QNone_Int_1_argbuf_0_d;
  \Int#_t  lizzieLet4_3QNone_Int_1_argbuf_0_bufchan_buf;
  assign lizzieLet4_3QNone_Int_1_argbuf_0_bufchan_r = (! lizzieLet4_3QNone_Int_1_argbuf_0_bufchan_buf[0]);
  assign lizzieLet23_1_argbuf_d = (lizzieLet4_3QNone_Int_1_argbuf_0_bufchan_buf[0] ? lizzieLet4_3QNone_Int_1_argbuf_0_bufchan_buf :
                                   lizzieLet4_3QNone_Int_1_argbuf_0_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_3QNone_Int_1_argbuf_0_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((lizzieLet23_1_argbuf_r && lizzieLet4_3QNone_Int_1_argbuf_0_bufchan_buf[0]))
        lizzieLet4_3QNone_Int_1_argbuf_0_bufchan_buf <= {32'd0, 1'd0};
      else if (((! lizzieLet23_1_argbuf_r) && (! lizzieLet4_3QNone_Int_1_argbuf_0_bufchan_buf[0])))
        lizzieLet4_3QNone_Int_1_argbuf_0_bufchan_buf <= lizzieLet4_3QNone_Int_1_argbuf_0_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet4_3QNone_Int_2,Go) > (lizzieLet4_3QNone_Int_2_argbuf,Go) */
  Go_t lizzieLet4_3QNone_Int_2_bufchan_d;
  logic lizzieLet4_3QNone_Int_2_bufchan_r;
  assign lizzieLet4_3QNone_Int_2_r = ((! lizzieLet4_3QNone_Int_2_bufchan_d[0]) || lizzieLet4_3QNone_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3QNone_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet4_3QNone_Int_2_r)
        lizzieLet4_3QNone_Int_2_bufchan_d <= lizzieLet4_3QNone_Int_2_d;
  Go_t lizzieLet4_3QNone_Int_2_bufchan_buf;
  assign lizzieLet4_3QNone_Int_2_bufchan_r = (! lizzieLet4_3QNone_Int_2_bufchan_buf[0]);
  assign lizzieLet4_3QNone_Int_2_argbuf_d = (lizzieLet4_3QNone_Int_2_bufchan_buf[0] ? lizzieLet4_3QNone_Int_2_bufchan_buf :
                                             lizzieLet4_3QNone_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3QNone_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet4_3QNone_Int_2_argbuf_r && lizzieLet4_3QNone_Int_2_bufchan_buf[0]))
        lizzieLet4_3QNone_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet4_3QNone_Int_2_argbuf_r) && (! lizzieLet4_3QNone_Int_2_bufchan_buf[0])))
        lizzieLet4_3QNone_Int_2_bufchan_buf <= lizzieLet4_3QNone_Int_2_bufchan_d;
  
  /* mergectrl (Ty C4,Ty Go) : [(lizzieLet4_3QNone_Int_2_argbuf,Go),
                           (lizzieLet35_3Lcall_$wnnz0_1_argbuf,Go),
                           (lizzieLet4_3QVal_Int_2_argbuf,Go),
                           (lizzieLet4_3QError_Int_2_argbuf,Go)] > (go_15_goMux_choice,C4) (go_15_goMux_data,Go) */
  logic [3:0] lizzieLet4_3QNone_Int_2_argbuf_select_d;
  assign lizzieLet4_3QNone_Int_2_argbuf_select_d = ((| lizzieLet4_3QNone_Int_2_argbuf_select_q) ? lizzieLet4_3QNone_Int_2_argbuf_select_q :
                                                    (lizzieLet4_3QNone_Int_2_argbuf_d[0] ? 4'd1 :
                                                     (lizzieLet35_3Lcall_$wnnz0_1_argbuf_d[0] ? 4'd2 :
                                                      (lizzieLet4_3QVal_Int_2_argbuf_d[0] ? 4'd4 :
                                                       (lizzieLet4_3QError_Int_2_argbuf_d[0] ? 4'd8 :
                                                        4'd0)))));
  logic [3:0] lizzieLet4_3QNone_Int_2_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_3QNone_Int_2_argbuf_select_q <= 4'd0;
    else
      lizzieLet4_3QNone_Int_2_argbuf_select_q <= (lizzieLet4_3QNone_Int_2_argbuf_done ? 4'd0 :
                                                  lizzieLet4_3QNone_Int_2_argbuf_select_d);
  logic [1:0] lizzieLet4_3QNone_Int_2_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3QNone_Int_2_argbuf_emit_q <= 2'd0;
    else
      lizzieLet4_3QNone_Int_2_argbuf_emit_q <= (lizzieLet4_3QNone_Int_2_argbuf_done ? 2'd0 :
                                                lizzieLet4_3QNone_Int_2_argbuf_emit_d);
  logic [1:0] lizzieLet4_3QNone_Int_2_argbuf_emit_d;
  assign lizzieLet4_3QNone_Int_2_argbuf_emit_d = (lizzieLet4_3QNone_Int_2_argbuf_emit_q | ({go_15_goMux_choice_d[0],
                                                                                            go_15_goMux_data_d[0]} & {go_15_goMux_choice_r,
                                                                                                                      go_15_goMux_data_r}));
  logic lizzieLet4_3QNone_Int_2_argbuf_done;
  assign lizzieLet4_3QNone_Int_2_argbuf_done = (& lizzieLet4_3QNone_Int_2_argbuf_emit_d);
  assign {lizzieLet4_3QError_Int_2_argbuf_r,
          lizzieLet4_3QVal_Int_2_argbuf_r,
          lizzieLet35_3Lcall_$wnnz0_1_argbuf_r,
          lizzieLet4_3QNone_Int_2_argbuf_r} = (lizzieLet4_3QNone_Int_2_argbuf_done ? lizzieLet4_3QNone_Int_2_argbuf_select_d :
                                               4'd0);
  assign go_15_goMux_data_d = ((lizzieLet4_3QNone_Int_2_argbuf_select_d[0] && (! lizzieLet4_3QNone_Int_2_argbuf_emit_q[0])) ? lizzieLet4_3QNone_Int_2_argbuf_d :
                               ((lizzieLet4_3QNone_Int_2_argbuf_select_d[1] && (! lizzieLet4_3QNone_Int_2_argbuf_emit_q[0])) ? lizzieLet35_3Lcall_$wnnz0_1_argbuf_d :
                                ((lizzieLet4_3QNone_Int_2_argbuf_select_d[2] && (! lizzieLet4_3QNone_Int_2_argbuf_emit_q[0])) ? lizzieLet4_3QVal_Int_2_argbuf_d :
                                 ((lizzieLet4_3QNone_Int_2_argbuf_select_d[3] && (! lizzieLet4_3QNone_Int_2_argbuf_emit_q[0])) ? lizzieLet4_3QError_Int_2_argbuf_d :
                                  1'd0))));
  assign go_15_goMux_choice_d = ((lizzieLet4_3QNone_Int_2_argbuf_select_d[0] && (! lizzieLet4_3QNone_Int_2_argbuf_emit_q[1])) ? C1_4_dc(1'd1) :
                                 ((lizzieLet4_3QNone_Int_2_argbuf_select_d[1] && (! lizzieLet4_3QNone_Int_2_argbuf_emit_q[1])) ? C2_4_dc(1'd1) :
                                  ((lizzieLet4_3QNone_Int_2_argbuf_select_d[2] && (! lizzieLet4_3QNone_Int_2_argbuf_emit_q[1])) ? C3_4_dc(1'd1) :
                                   ((lizzieLet4_3QNone_Int_2_argbuf_select_d[3] && (! lizzieLet4_3QNone_Int_2_argbuf_emit_q[1])) ? C4_4_dc(1'd1) :
                                    {2'd0, 1'd0}))));
  
  /* fork (Ty Go) : (lizzieLet4_3QVal_Int,Go) > [(lizzieLet4_3QVal_Int_1,Go),
                                            (lizzieLet4_3QVal_Int_2,Go)] */
  logic [1:0] lizzieLet4_3QVal_Int_emitted;
  logic [1:0] lizzieLet4_3QVal_Int_done;
  assign lizzieLet4_3QVal_Int_1_d = (lizzieLet4_3QVal_Int_d[0] && (! lizzieLet4_3QVal_Int_emitted[0]));
  assign lizzieLet4_3QVal_Int_2_d = (lizzieLet4_3QVal_Int_d[0] && (! lizzieLet4_3QVal_Int_emitted[1]));
  assign lizzieLet4_3QVal_Int_done = (lizzieLet4_3QVal_Int_emitted | ({lizzieLet4_3QVal_Int_2_d[0],
                                                                       lizzieLet4_3QVal_Int_1_d[0]} & {lizzieLet4_3QVal_Int_2_r,
                                                                                                       lizzieLet4_3QVal_Int_1_r}));
  assign lizzieLet4_3QVal_Int_r = (& lizzieLet4_3QVal_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3QVal_Int_emitted <= 2'd0;
    else
      lizzieLet4_3QVal_Int_emitted <= (lizzieLet4_3QVal_Int_r ? 2'd0 :
                                       lizzieLet4_3QVal_Int_done);
  
  /* buf (Ty Go) : (lizzieLet4_3QVal_Int_1,Go) > (lizzieLet4_3QVal_Int_1_argbuf,Go) */
  Go_t lizzieLet4_3QVal_Int_1_bufchan_d;
  logic lizzieLet4_3QVal_Int_1_bufchan_r;
  assign lizzieLet4_3QVal_Int_1_r = ((! lizzieLet4_3QVal_Int_1_bufchan_d[0]) || lizzieLet4_3QVal_Int_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3QVal_Int_1_bufchan_d <= 1'd0;
    else
      if (lizzieLet4_3QVal_Int_1_r)
        lizzieLet4_3QVal_Int_1_bufchan_d <= lizzieLet4_3QVal_Int_1_d;
  Go_t lizzieLet4_3QVal_Int_1_bufchan_buf;
  assign lizzieLet4_3QVal_Int_1_bufchan_r = (! lizzieLet4_3QVal_Int_1_bufchan_buf[0]);
  assign lizzieLet4_3QVal_Int_1_argbuf_d = (lizzieLet4_3QVal_Int_1_bufchan_buf[0] ? lizzieLet4_3QVal_Int_1_bufchan_buf :
                                            lizzieLet4_3QVal_Int_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3QVal_Int_1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet4_3QVal_Int_1_argbuf_r && lizzieLet4_3QVal_Int_1_bufchan_buf[0]))
        lizzieLet4_3QVal_Int_1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet4_3QVal_Int_1_argbuf_r) && (! lizzieLet4_3QVal_Int_1_bufchan_buf[0])))
        lizzieLet4_3QVal_Int_1_bufchan_buf <= lizzieLet4_3QVal_Int_1_bufchan_d;
  
  /* const (Ty Int#,
       Lit 1) : (lizzieLet4_3QVal_Int_1_argbuf,Go) > (lizzieLet4_3QVal_Int_1_argbuf_1,Int#) */
  assign lizzieLet4_3QVal_Int_1_argbuf_1_d = {32'd1,
                                              lizzieLet4_3QVal_Int_1_argbuf_d[0]};
  assign lizzieLet4_3QVal_Int_1_argbuf_r = lizzieLet4_3QVal_Int_1_argbuf_1_r;
  
  /* buf (Ty Int#) : (lizzieLet4_3QVal_Int_1_argbuf_1,Int#) > (lizzieLet24_1_argbuf,Int#) */
  \Int#_t  lizzieLet4_3QVal_Int_1_argbuf_1_bufchan_d;
  logic lizzieLet4_3QVal_Int_1_argbuf_1_bufchan_r;
  assign lizzieLet4_3QVal_Int_1_argbuf_1_r = ((! lizzieLet4_3QVal_Int_1_argbuf_1_bufchan_d[0]) || lizzieLet4_3QVal_Int_1_argbuf_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_3QVal_Int_1_argbuf_1_bufchan_d <= {32'd0, 1'd0};
    else
      if (lizzieLet4_3QVal_Int_1_argbuf_1_r)
        lizzieLet4_3QVal_Int_1_argbuf_1_bufchan_d <= lizzieLet4_3QVal_Int_1_argbuf_1_d;
  \Int#_t  lizzieLet4_3QVal_Int_1_argbuf_1_bufchan_buf;
  assign lizzieLet4_3QVal_Int_1_argbuf_1_bufchan_r = (! lizzieLet4_3QVal_Int_1_argbuf_1_bufchan_buf[0]);
  assign lizzieLet24_1_argbuf_d = (lizzieLet4_3QVal_Int_1_argbuf_1_bufchan_buf[0] ? lizzieLet4_3QVal_Int_1_argbuf_1_bufchan_buf :
                                   lizzieLet4_3QVal_Int_1_argbuf_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_3QVal_Int_1_argbuf_1_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((lizzieLet24_1_argbuf_r && lizzieLet4_3QVal_Int_1_argbuf_1_bufchan_buf[0]))
        lizzieLet4_3QVal_Int_1_argbuf_1_bufchan_buf <= {32'd0, 1'd0};
      else if (((! lizzieLet24_1_argbuf_r) && (! lizzieLet4_3QVal_Int_1_argbuf_1_bufchan_buf[0])))
        lizzieLet4_3QVal_Int_1_argbuf_1_bufchan_buf <= lizzieLet4_3QVal_Int_1_argbuf_1_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet4_3QVal_Int_2,Go) > (lizzieLet4_3QVal_Int_2_argbuf,Go) */
  Go_t lizzieLet4_3QVal_Int_2_bufchan_d;
  logic lizzieLet4_3QVal_Int_2_bufchan_r;
  assign lizzieLet4_3QVal_Int_2_r = ((! lizzieLet4_3QVal_Int_2_bufchan_d[0]) || lizzieLet4_3QVal_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3QVal_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet4_3QVal_Int_2_r)
        lizzieLet4_3QVal_Int_2_bufchan_d <= lizzieLet4_3QVal_Int_2_d;
  Go_t lizzieLet4_3QVal_Int_2_bufchan_buf;
  assign lizzieLet4_3QVal_Int_2_bufchan_r = (! lizzieLet4_3QVal_Int_2_bufchan_buf[0]);
  assign lizzieLet4_3QVal_Int_2_argbuf_d = (lizzieLet4_3QVal_Int_2_bufchan_buf[0] ? lizzieLet4_3QVal_Int_2_bufchan_buf :
                                            lizzieLet4_3QVal_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3QVal_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet4_3QVal_Int_2_argbuf_r && lizzieLet4_3QVal_Int_2_bufchan_buf[0]))
        lizzieLet4_3QVal_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet4_3QVal_Int_2_argbuf_r) && (! lizzieLet4_3QVal_Int_2_bufchan_buf[0])))
        lizzieLet4_3QVal_Int_2_bufchan_buf <= lizzieLet4_3QVal_Int_2_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_CT$wnnz) : (lizzieLet4_4,QTree_Int) (sc_0_goMux_mux,Pointer_CT$wnnz) > [(lizzieLet4_4QNone_Int,Pointer_CT$wnnz),
                                                                                          (lizzieLet4_4QVal_Int,Pointer_CT$wnnz),
                                                                                          (lizzieLet4_4QNode_Int,Pointer_CT$wnnz),
                                                                                          (lizzieLet4_4QError_Int,Pointer_CT$wnnz)] */
  logic [3:0] sc_0_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet4_4_d[0] && sc_0_goMux_mux_d[0]))
      unique case (lizzieLet4_4_d[2:1])
        2'd0: sc_0_goMux_mux_onehotd = 4'd1;
        2'd1: sc_0_goMux_mux_onehotd = 4'd2;
        2'd2: sc_0_goMux_mux_onehotd = 4'd4;
        2'd3: sc_0_goMux_mux_onehotd = 4'd8;
        default: sc_0_goMux_mux_onehotd = 4'd0;
      endcase
    else sc_0_goMux_mux_onehotd = 4'd0;
  assign lizzieLet4_4QNone_Int_d = {sc_0_goMux_mux_d[16:1],
                                    sc_0_goMux_mux_onehotd[0]};
  assign lizzieLet4_4QVal_Int_d = {sc_0_goMux_mux_d[16:1],
                                   sc_0_goMux_mux_onehotd[1]};
  assign lizzieLet4_4QNode_Int_d = {sc_0_goMux_mux_d[16:1],
                                    sc_0_goMux_mux_onehotd[2]};
  assign lizzieLet4_4QError_Int_d = {sc_0_goMux_mux_d[16:1],
                                     sc_0_goMux_mux_onehotd[3]};
  assign sc_0_goMux_mux_r = (| (sc_0_goMux_mux_onehotd & {lizzieLet4_4QError_Int_r,
                                                          lizzieLet4_4QNode_Int_r,
                                                          lizzieLet4_4QVal_Int_r,
                                                          lizzieLet4_4QNone_Int_r}));
  assign lizzieLet4_4_r = sc_0_goMux_mux_r;
  
  /* buf (Ty Pointer_CT$wnnz) : (lizzieLet4_4QError_Int,Pointer_CT$wnnz) > (lizzieLet4_4QError_Int_1_argbuf,Pointer_CT$wnnz) */
  Pointer_CT$wnnz_t lizzieLet4_4QError_Int_bufchan_d;
  logic lizzieLet4_4QError_Int_bufchan_r;
  assign lizzieLet4_4QError_Int_r = ((! lizzieLet4_4QError_Int_bufchan_d[0]) || lizzieLet4_4QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_4QError_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet4_4QError_Int_r)
        lizzieLet4_4QError_Int_bufchan_d <= lizzieLet4_4QError_Int_d;
  Pointer_CT$wnnz_t lizzieLet4_4QError_Int_bufchan_buf;
  assign lizzieLet4_4QError_Int_bufchan_r = (! lizzieLet4_4QError_Int_bufchan_buf[0]);
  assign lizzieLet4_4QError_Int_1_argbuf_d = (lizzieLet4_4QError_Int_bufchan_buf[0] ? lizzieLet4_4QError_Int_bufchan_buf :
                                              lizzieLet4_4QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_4QError_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet4_4QError_Int_1_argbuf_r && lizzieLet4_4QError_Int_bufchan_buf[0]))
        lizzieLet4_4QError_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet4_4QError_Int_1_argbuf_r) && (! lizzieLet4_4QError_Int_bufchan_buf[0])))
        lizzieLet4_4QError_Int_bufchan_buf <= lizzieLet4_4QError_Int_bufchan_d;
  
  /* dcon (Ty CT$wnnz,
      Dcon Lcall_$wnnz3) : [(lizzieLet4_4QNode_Int,Pointer_CT$wnnz),
                            (q4a87_destruct,Pointer_QTree_Int),
                            (q3a86_destruct,Pointer_QTree_Int),
                            (q2a85_destruct,Pointer_QTree_Int)] > (lizzieLet4_4QNode_Int_1q4a87_1q3a86_1q2a85_1Lcall_$wnnz3,CT$wnnz) */
  assign lizzieLet4_4QNode_Int_1q4a87_1q3a86_1q2a85_1Lcall_$wnnz3_d = Lcall_$wnnz3_dc((& {lizzieLet4_4QNode_Int_d[0],
                                                                                          q4a87_destruct_d[0],
                                                                                          q3a86_destruct_d[0],
                                                                                          q2a85_destruct_d[0]}), lizzieLet4_4QNode_Int_d, q4a87_destruct_d, q3a86_destruct_d, q2a85_destruct_d);
  assign {lizzieLet4_4QNode_Int_r,
          q4a87_destruct_r,
          q3a86_destruct_r,
          q2a85_destruct_r} = {4 {(lizzieLet4_4QNode_Int_1q4a87_1q3a86_1q2a85_1Lcall_$wnnz3_r && lizzieLet4_4QNode_Int_1q4a87_1q3a86_1q2a85_1Lcall_$wnnz3_d[0])}};
  
  /* buf (Ty CT$wnnz) : (lizzieLet4_4QNode_Int_1q4a87_1q3a86_1q2a85_1Lcall_$wnnz3,CT$wnnz) > (lizzieLet5_1_argbuf,CT$wnnz) */
  CT$wnnz_t lizzieLet4_4QNode_Int_1q4a87_1q3a86_1q2a85_1Lcall_$wnnz3_bufchan_d;
  logic lizzieLet4_4QNode_Int_1q4a87_1q3a86_1q2a85_1Lcall_$wnnz3_bufchan_r;
  assign lizzieLet4_4QNode_Int_1q4a87_1q3a86_1q2a85_1Lcall_$wnnz3_r = ((! lizzieLet4_4QNode_Int_1q4a87_1q3a86_1q2a85_1Lcall_$wnnz3_bufchan_d[0]) || lizzieLet4_4QNode_Int_1q4a87_1q3a86_1q2a85_1Lcall_$wnnz3_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_4QNode_Int_1q4a87_1q3a86_1q2a85_1Lcall_$wnnz3_bufchan_d <= {115'd0,
                                                                             1'd0};
    else
      if (lizzieLet4_4QNode_Int_1q4a87_1q3a86_1q2a85_1Lcall_$wnnz3_r)
        lizzieLet4_4QNode_Int_1q4a87_1q3a86_1q2a85_1Lcall_$wnnz3_bufchan_d <= lizzieLet4_4QNode_Int_1q4a87_1q3a86_1q2a85_1Lcall_$wnnz3_d;
  CT$wnnz_t lizzieLet4_4QNode_Int_1q4a87_1q3a86_1q2a85_1Lcall_$wnnz3_bufchan_buf;
  assign lizzieLet4_4QNode_Int_1q4a87_1q3a86_1q2a85_1Lcall_$wnnz3_bufchan_r = (! lizzieLet4_4QNode_Int_1q4a87_1q3a86_1q2a85_1Lcall_$wnnz3_bufchan_buf[0]);
  assign lizzieLet5_1_argbuf_d = (lizzieLet4_4QNode_Int_1q4a87_1q3a86_1q2a85_1Lcall_$wnnz3_bufchan_buf[0] ? lizzieLet4_4QNode_Int_1q4a87_1q3a86_1q2a85_1Lcall_$wnnz3_bufchan_buf :
                                  lizzieLet4_4QNode_Int_1q4a87_1q3a86_1q2a85_1Lcall_$wnnz3_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_4QNode_Int_1q4a87_1q3a86_1q2a85_1Lcall_$wnnz3_bufchan_buf <= {115'd0,
                                                                               1'd0};
    else
      if ((lizzieLet5_1_argbuf_r && lizzieLet4_4QNode_Int_1q4a87_1q3a86_1q2a85_1Lcall_$wnnz3_bufchan_buf[0]))
        lizzieLet4_4QNode_Int_1q4a87_1q3a86_1q2a85_1Lcall_$wnnz3_bufchan_buf <= {115'd0,
                                                                                 1'd0};
      else if (((! lizzieLet5_1_argbuf_r) && (! lizzieLet4_4QNode_Int_1q4a87_1q3a86_1q2a85_1Lcall_$wnnz3_bufchan_buf[0])))
        lizzieLet4_4QNode_Int_1q4a87_1q3a86_1q2a85_1Lcall_$wnnz3_bufchan_buf <= lizzieLet4_4QNode_Int_1q4a87_1q3a86_1q2a85_1Lcall_$wnnz3_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz) : (lizzieLet4_4QNone_Int,Pointer_CT$wnnz) > (lizzieLet4_4QNone_Int_1_argbuf,Pointer_CT$wnnz) */
  Pointer_CT$wnnz_t lizzieLet4_4QNone_Int_bufchan_d;
  logic lizzieLet4_4QNone_Int_bufchan_r;
  assign lizzieLet4_4QNone_Int_r = ((! lizzieLet4_4QNone_Int_bufchan_d[0]) || lizzieLet4_4QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_4QNone_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet4_4QNone_Int_r)
        lizzieLet4_4QNone_Int_bufchan_d <= lizzieLet4_4QNone_Int_d;
  Pointer_CT$wnnz_t lizzieLet4_4QNone_Int_bufchan_buf;
  assign lizzieLet4_4QNone_Int_bufchan_r = (! lizzieLet4_4QNone_Int_bufchan_buf[0]);
  assign lizzieLet4_4QNone_Int_1_argbuf_d = (lizzieLet4_4QNone_Int_bufchan_buf[0] ? lizzieLet4_4QNone_Int_bufchan_buf :
                                             lizzieLet4_4QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_4QNone_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet4_4QNone_Int_1_argbuf_r && lizzieLet4_4QNone_Int_bufchan_buf[0]))
        lizzieLet4_4QNone_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet4_4QNone_Int_1_argbuf_r) && (! lizzieLet4_4QNone_Int_bufchan_buf[0])))
        lizzieLet4_4QNone_Int_bufchan_buf <= lizzieLet4_4QNone_Int_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz) : (lizzieLet4_4QVal_Int,Pointer_CT$wnnz) > (lizzieLet4_4QVal_Int_1_argbuf,Pointer_CT$wnnz) */
  Pointer_CT$wnnz_t lizzieLet4_4QVal_Int_bufchan_d;
  logic lizzieLet4_4QVal_Int_bufchan_r;
  assign lizzieLet4_4QVal_Int_r = ((! lizzieLet4_4QVal_Int_bufchan_d[0]) || lizzieLet4_4QVal_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_4QVal_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet4_4QVal_Int_r)
        lizzieLet4_4QVal_Int_bufchan_d <= lizzieLet4_4QVal_Int_d;
  Pointer_CT$wnnz_t lizzieLet4_4QVal_Int_bufchan_buf;
  assign lizzieLet4_4QVal_Int_bufchan_r = (! lizzieLet4_4QVal_Int_bufchan_buf[0]);
  assign lizzieLet4_4QVal_Int_1_argbuf_d = (lizzieLet4_4QVal_Int_bufchan_buf[0] ? lizzieLet4_4QVal_Int_bufchan_buf :
                                            lizzieLet4_4QVal_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_4QVal_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet4_4QVal_Int_1_argbuf_r && lizzieLet4_4QVal_Int_bufchan_buf[0]))
        lizzieLet4_4QVal_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet4_4QVal_Int_1_argbuf_r) && (! lizzieLet4_4QVal_Int_bufchan_buf[0])))
        lizzieLet4_4QVal_Int_bufchan_buf <= lizzieLet4_4QVal_Int_bufchan_d;
  
  /* destruct (Ty QTree_Int,
          Dcon QNode_Int) : (lizzieLet6_1QNode_Int,QTree_Int) > [(tla8y_destruct,Pointer_QTree_Int),
                                                                 (tra8z_destruct,Pointer_QTree_Int),
                                                                 (bla8A_destruct,Pointer_QTree_Int),
                                                                 (bra8B_destruct,Pointer_QTree_Int)] */
  logic [3:0] lizzieLet6_1QNode_Int_emitted;
  logic [3:0] lizzieLet6_1QNode_Int_done;
  assign tla8y_destruct_d = {lizzieLet6_1QNode_Int_d[18:3],
                             (lizzieLet6_1QNode_Int_d[0] && (! lizzieLet6_1QNode_Int_emitted[0]))};
  assign tra8z_destruct_d = {lizzieLet6_1QNode_Int_d[34:19],
                             (lizzieLet6_1QNode_Int_d[0] && (! lizzieLet6_1QNode_Int_emitted[1]))};
  assign bla8A_destruct_d = {lizzieLet6_1QNode_Int_d[50:35],
                             (lizzieLet6_1QNode_Int_d[0] && (! lizzieLet6_1QNode_Int_emitted[2]))};
  assign bra8B_destruct_d = {lizzieLet6_1QNode_Int_d[66:51],
                             (lizzieLet6_1QNode_Int_d[0] && (! lizzieLet6_1QNode_Int_emitted[3]))};
  assign lizzieLet6_1QNode_Int_done = (lizzieLet6_1QNode_Int_emitted | ({bra8B_destruct_d[0],
                                                                         bla8A_destruct_d[0],
                                                                         tra8z_destruct_d[0],
                                                                         tla8y_destruct_d[0]} & {bra8B_destruct_r,
                                                                                                 bla8A_destruct_r,
                                                                                                 tra8z_destruct_r,
                                                                                                 tla8y_destruct_r}));
  assign lizzieLet6_1QNode_Int_r = (& lizzieLet6_1QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_1QNode_Int_emitted <= 4'd0;
    else
      lizzieLet6_1QNode_Int_emitted <= (lizzieLet6_1QNode_Int_r ? 4'd0 :
                                        lizzieLet6_1QNode_Int_done);
  
  /* destruct (Ty QTree_Int,
          Dcon QVal_Int) : (lizzieLet6_1QVal_Int,QTree_Int) > [(va8x_destruct,Int)] */
  assign va8x_destruct_d = {lizzieLet6_1QVal_Int_d[34:3],
                            lizzieLet6_1QVal_Int_d[0]};
  assign lizzieLet6_1QVal_Int_r = va8x_destruct_r;
  
  /* demux (Ty QTree_Int,
       Ty QTree_Int) : (lizzieLet6_2,QTree_Int) (lizzieLet6_1,QTree_Int) > [(_5,QTree_Int),
                                                                            (lizzieLet6_1QVal_Int,QTree_Int),
                                                                            (lizzieLet6_1QNode_Int,QTree_Int),
                                                                            (_4,QTree_Int)] */
  logic [3:0] lizzieLet6_1_onehotd;
  always_comb
    if ((lizzieLet6_2_d[0] && lizzieLet6_1_d[0]))
      unique case (lizzieLet6_2_d[2:1])
        2'd0: lizzieLet6_1_onehotd = 4'd1;
        2'd1: lizzieLet6_1_onehotd = 4'd2;
        2'd2: lizzieLet6_1_onehotd = 4'd4;
        2'd3: lizzieLet6_1_onehotd = 4'd8;
        default: lizzieLet6_1_onehotd = 4'd0;
      endcase
    else lizzieLet6_1_onehotd = 4'd0;
  assign _5_d = {lizzieLet6_1_d[66:1], lizzieLet6_1_onehotd[0]};
  assign lizzieLet6_1QVal_Int_d = {lizzieLet6_1_d[66:1],
                                   lizzieLet6_1_onehotd[1]};
  assign lizzieLet6_1QNode_Int_d = {lizzieLet6_1_d[66:1],
                                    lizzieLet6_1_onehotd[2]};
  assign _4_d = {lizzieLet6_1_d[66:1], lizzieLet6_1_onehotd[3]};
  assign lizzieLet6_1_r = (| (lizzieLet6_1_onehotd & {_4_r,
                                                      lizzieLet6_1QNode_Int_r,
                                                      lizzieLet6_1QVal_Int_r,
                                                      _5_r}));
  assign lizzieLet6_2_r = lizzieLet6_1_r;
  
  /* demux (Ty QTree_Int,
       Ty Go) : (lizzieLet6_3,QTree_Int) (go_11_goMux_data,Go) > [(lizzieLet6_3QNone_Int,Go),
                                                                  (lizzieLet6_3QVal_Int,Go),
                                                                  (lizzieLet6_3QNode_Int,Go),
                                                                  (lizzieLet6_3QError_Int,Go)] */
  logic [3:0] go_11_goMux_data_onehotd;
  always_comb
    if ((lizzieLet6_3_d[0] && go_11_goMux_data_d[0]))
      unique case (lizzieLet6_3_d[2:1])
        2'd0: go_11_goMux_data_onehotd = 4'd1;
        2'd1: go_11_goMux_data_onehotd = 4'd2;
        2'd2: go_11_goMux_data_onehotd = 4'd4;
        2'd3: go_11_goMux_data_onehotd = 4'd8;
        default: go_11_goMux_data_onehotd = 4'd0;
      endcase
    else go_11_goMux_data_onehotd = 4'd0;
  assign lizzieLet6_3QNone_Int_d = go_11_goMux_data_onehotd[0];
  assign lizzieLet6_3QVal_Int_d = go_11_goMux_data_onehotd[1];
  assign lizzieLet6_3QNode_Int_d = go_11_goMux_data_onehotd[2];
  assign lizzieLet6_3QError_Int_d = go_11_goMux_data_onehotd[3];
  assign go_11_goMux_data_r = (| (go_11_goMux_data_onehotd & {lizzieLet6_3QError_Int_r,
                                                              lizzieLet6_3QNode_Int_r,
                                                              lizzieLet6_3QVal_Int_r,
                                                              lizzieLet6_3QNone_Int_r}));
  assign lizzieLet6_3_r = go_11_goMux_data_r;
  
  /* fork (Ty Go) : (lizzieLet6_3QError_Int,Go) > [(lizzieLet6_3QError_Int_1,Go),
                                              (lizzieLet6_3QError_Int_2,Go)] */
  logic [1:0] lizzieLet6_3QError_Int_emitted;
  logic [1:0] lizzieLet6_3QError_Int_done;
  assign lizzieLet6_3QError_Int_1_d = (lizzieLet6_3QError_Int_d[0] && (! lizzieLet6_3QError_Int_emitted[0]));
  assign lizzieLet6_3QError_Int_2_d = (lizzieLet6_3QError_Int_d[0] && (! lizzieLet6_3QError_Int_emitted[1]));
  assign lizzieLet6_3QError_Int_done = (lizzieLet6_3QError_Int_emitted | ({lizzieLet6_3QError_Int_2_d[0],
                                                                           lizzieLet6_3QError_Int_1_d[0]} & {lizzieLet6_3QError_Int_2_r,
                                                                                                             lizzieLet6_3QError_Int_1_r}));
  assign lizzieLet6_3QError_Int_r = (& lizzieLet6_3QError_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_3QError_Int_emitted <= 2'd0;
    else
      lizzieLet6_3QError_Int_emitted <= (lizzieLet6_3QError_Int_r ? 2'd0 :
                                         lizzieLet6_3QError_Int_done);
  
  /* dcon (Ty QTree_Int,
      Dcon QError_Int) : [(lizzieLet6_3QError_Int_1,Go)] > (lizzieLet6_3QError_Int_1QError_Int,QTree_Int) */
  assign lizzieLet6_3QError_Int_1QError_Int_d = QError_Int_dc((& {lizzieLet6_3QError_Int_1_d[0]}), lizzieLet6_3QError_Int_1_d);
  assign {lizzieLet6_3QError_Int_1_r} = {1 {(lizzieLet6_3QError_Int_1QError_Int_r && lizzieLet6_3QError_Int_1QError_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (lizzieLet6_3QError_Int_1QError_Int,QTree_Int) > (lizzieLet11_1_argbuf,QTree_Int) */
  QTree_Int_t lizzieLet6_3QError_Int_1QError_Int_bufchan_d;
  logic lizzieLet6_3QError_Int_1QError_Int_bufchan_r;
  assign lizzieLet6_3QError_Int_1QError_Int_r = ((! lizzieLet6_3QError_Int_1QError_Int_bufchan_d[0]) || lizzieLet6_3QError_Int_1QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_3QError_Int_1QError_Int_bufchan_d <= {66'd0, 1'd0};
    else
      if (lizzieLet6_3QError_Int_1QError_Int_r)
        lizzieLet6_3QError_Int_1QError_Int_bufchan_d <= lizzieLet6_3QError_Int_1QError_Int_d;
  QTree_Int_t lizzieLet6_3QError_Int_1QError_Int_bufchan_buf;
  assign lizzieLet6_3QError_Int_1QError_Int_bufchan_r = (! lizzieLet6_3QError_Int_1QError_Int_bufchan_buf[0]);
  assign lizzieLet11_1_argbuf_d = (lizzieLet6_3QError_Int_1QError_Int_bufchan_buf[0] ? lizzieLet6_3QError_Int_1QError_Int_bufchan_buf :
                                   lizzieLet6_3QError_Int_1QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_3QError_Int_1QError_Int_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((lizzieLet11_1_argbuf_r && lizzieLet6_3QError_Int_1QError_Int_bufchan_buf[0]))
        lizzieLet6_3QError_Int_1QError_Int_bufchan_buf <= {66'd0, 1'd0};
      else if (((! lizzieLet11_1_argbuf_r) && (! lizzieLet6_3QError_Int_1QError_Int_bufchan_buf[0])))
        lizzieLet6_3QError_Int_1QError_Int_bufchan_buf <= lizzieLet6_3QError_Int_1QError_Int_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet6_3QError_Int_2,Go) > (lizzieLet6_3QError_Int_2_argbuf,Go) */
  Go_t lizzieLet6_3QError_Int_2_bufchan_d;
  logic lizzieLet6_3QError_Int_2_bufchan_r;
  assign lizzieLet6_3QError_Int_2_r = ((! lizzieLet6_3QError_Int_2_bufchan_d[0]) || lizzieLet6_3QError_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_3QError_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet6_3QError_Int_2_r)
        lizzieLet6_3QError_Int_2_bufchan_d <= lizzieLet6_3QError_Int_2_d;
  Go_t lizzieLet6_3QError_Int_2_bufchan_buf;
  assign lizzieLet6_3QError_Int_2_bufchan_r = (! lizzieLet6_3QError_Int_2_bufchan_buf[0]);
  assign lizzieLet6_3QError_Int_2_argbuf_d = (lizzieLet6_3QError_Int_2_bufchan_buf[0] ? lizzieLet6_3QError_Int_2_bufchan_buf :
                                              lizzieLet6_3QError_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_3QError_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet6_3QError_Int_2_argbuf_r && lizzieLet6_3QError_Int_2_bufchan_buf[0]))
        lizzieLet6_3QError_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet6_3QError_Int_2_argbuf_r) && (! lizzieLet6_3QError_Int_2_bufchan_buf[0])))
        lizzieLet6_3QError_Int_2_bufchan_buf <= lizzieLet6_3QError_Int_2_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet6_3QNode_Int,Go) > (lizzieLet6_3QNode_Int_1_argbuf,Go) */
  Go_t lizzieLet6_3QNode_Int_bufchan_d;
  logic lizzieLet6_3QNode_Int_bufchan_r;
  assign lizzieLet6_3QNode_Int_r = ((! lizzieLet6_3QNode_Int_bufchan_d[0]) || lizzieLet6_3QNode_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_3QNode_Int_bufchan_d <= 1'd0;
    else
      if (lizzieLet6_3QNode_Int_r)
        lizzieLet6_3QNode_Int_bufchan_d <= lizzieLet6_3QNode_Int_d;
  Go_t lizzieLet6_3QNode_Int_bufchan_buf;
  assign lizzieLet6_3QNode_Int_bufchan_r = (! lizzieLet6_3QNode_Int_bufchan_buf[0]);
  assign lizzieLet6_3QNode_Int_1_argbuf_d = (lizzieLet6_3QNode_Int_bufchan_buf[0] ? lizzieLet6_3QNode_Int_bufchan_buf :
                                             lizzieLet6_3QNode_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_3QNode_Int_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet6_3QNode_Int_1_argbuf_r && lizzieLet6_3QNode_Int_bufchan_buf[0]))
        lizzieLet6_3QNode_Int_bufchan_buf <= 1'd0;
      else if (((! lizzieLet6_3QNode_Int_1_argbuf_r) && (! lizzieLet6_3QNode_Int_bufchan_buf[0])))
        lizzieLet6_3QNode_Int_bufchan_buf <= lizzieLet6_3QNode_Int_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet6_3QNone_Int,Go) > [(lizzieLet6_3QNone_Int_1,Go),
                                             (lizzieLet6_3QNone_Int_2,Go)] */
  logic [1:0] lizzieLet6_3QNone_Int_emitted;
  logic [1:0] lizzieLet6_3QNone_Int_done;
  assign lizzieLet6_3QNone_Int_1_d = (lizzieLet6_3QNone_Int_d[0] && (! lizzieLet6_3QNone_Int_emitted[0]));
  assign lizzieLet6_3QNone_Int_2_d = (lizzieLet6_3QNone_Int_d[0] && (! lizzieLet6_3QNone_Int_emitted[1]));
  assign lizzieLet6_3QNone_Int_done = (lizzieLet6_3QNone_Int_emitted | ({lizzieLet6_3QNone_Int_2_d[0],
                                                                         lizzieLet6_3QNone_Int_1_d[0]} & {lizzieLet6_3QNone_Int_2_r,
                                                                                                          lizzieLet6_3QNone_Int_1_r}));
  assign lizzieLet6_3QNone_Int_r = (& lizzieLet6_3QNone_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_3QNone_Int_emitted <= 2'd0;
    else
      lizzieLet6_3QNone_Int_emitted <= (lizzieLet6_3QNone_Int_r ? 2'd0 :
                                        lizzieLet6_3QNone_Int_done);
  
  /* dcon (Ty QTree_Int,
      Dcon QNone_Int) : [(lizzieLet6_3QNone_Int_1,Go)] > (lizzieLet6_3QNone_Int_1QNone_Int,QTree_Int) */
  assign lizzieLet6_3QNone_Int_1QNone_Int_d = QNone_Int_dc((& {lizzieLet6_3QNone_Int_1_d[0]}), lizzieLet6_3QNone_Int_1_d);
  assign {lizzieLet6_3QNone_Int_1_r} = {1 {(lizzieLet6_3QNone_Int_1QNone_Int_r && lizzieLet6_3QNone_Int_1QNone_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (lizzieLet6_3QNone_Int_1QNone_Int,QTree_Int) > (lizzieLet7_1_argbuf,QTree_Int) */
  QTree_Int_t lizzieLet6_3QNone_Int_1QNone_Int_bufchan_d;
  logic lizzieLet6_3QNone_Int_1QNone_Int_bufchan_r;
  assign lizzieLet6_3QNone_Int_1QNone_Int_r = ((! lizzieLet6_3QNone_Int_1QNone_Int_bufchan_d[0]) || lizzieLet6_3QNone_Int_1QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_3QNone_Int_1QNone_Int_bufchan_d <= {66'd0, 1'd0};
    else
      if (lizzieLet6_3QNone_Int_1QNone_Int_r)
        lizzieLet6_3QNone_Int_1QNone_Int_bufchan_d <= lizzieLet6_3QNone_Int_1QNone_Int_d;
  QTree_Int_t lizzieLet6_3QNone_Int_1QNone_Int_bufchan_buf;
  assign lizzieLet6_3QNone_Int_1QNone_Int_bufchan_r = (! lizzieLet6_3QNone_Int_1QNone_Int_bufchan_buf[0]);
  assign lizzieLet7_1_argbuf_d = (lizzieLet6_3QNone_Int_1QNone_Int_bufchan_buf[0] ? lizzieLet6_3QNone_Int_1QNone_Int_bufchan_buf :
                                  lizzieLet6_3QNone_Int_1QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_3QNone_Int_1QNone_Int_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((lizzieLet7_1_argbuf_r && lizzieLet6_3QNone_Int_1QNone_Int_bufchan_buf[0]))
        lizzieLet6_3QNone_Int_1QNone_Int_bufchan_buf <= {66'd0, 1'd0};
      else if (((! lizzieLet7_1_argbuf_r) && (! lizzieLet6_3QNone_Int_1QNone_Int_bufchan_buf[0])))
        lizzieLet6_3QNone_Int_1QNone_Int_bufchan_buf <= lizzieLet6_3QNone_Int_1QNone_Int_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet6_3QNone_Int_2,Go) > (lizzieLet6_3QNone_Int_2_argbuf,Go) */
  Go_t lizzieLet6_3QNone_Int_2_bufchan_d;
  logic lizzieLet6_3QNone_Int_2_bufchan_r;
  assign lizzieLet6_3QNone_Int_2_r = ((! lizzieLet6_3QNone_Int_2_bufchan_d[0]) || lizzieLet6_3QNone_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_3QNone_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet6_3QNone_Int_2_r)
        lizzieLet6_3QNone_Int_2_bufchan_d <= lizzieLet6_3QNone_Int_2_d;
  Go_t lizzieLet6_3QNone_Int_2_bufchan_buf;
  assign lizzieLet6_3QNone_Int_2_bufchan_r = (! lizzieLet6_3QNone_Int_2_bufchan_buf[0]);
  assign lizzieLet6_3QNone_Int_2_argbuf_d = (lizzieLet6_3QNone_Int_2_bufchan_buf[0] ? lizzieLet6_3QNone_Int_2_bufchan_buf :
                                             lizzieLet6_3QNone_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_3QNone_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet6_3QNone_Int_2_argbuf_r && lizzieLet6_3QNone_Int_2_bufchan_buf[0]))
        lizzieLet6_3QNone_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet6_3QNone_Int_2_argbuf_r) && (! lizzieLet6_3QNone_Int_2_bufchan_buf[0])))
        lizzieLet6_3QNone_Int_2_bufchan_buf <= lizzieLet6_3QNone_Int_2_bufchan_d;
  
  /* mergectrl (Ty C5,Ty Go) : [(lizzieLet6_3QNone_Int_2_argbuf,Go),
                           (lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int0_1_argbuf,Go),
                           (es_2_1MyFalse_2_argbuf,Go),
                           (es_2_1MyTrue_2_argbuf,Go),
                           (lizzieLet6_3QError_Int_2_argbuf,Go)] > (go_16_goMux_choice,C5) (go_16_goMux_data,Go) */
  logic [4:0] lizzieLet6_3QNone_Int_2_argbuf_select_d;
  assign lizzieLet6_3QNone_Int_2_argbuf_select_d = ((| lizzieLet6_3QNone_Int_2_argbuf_select_q) ? lizzieLet6_3QNone_Int_2_argbuf_select_q :
                                                    (lizzieLet6_3QNone_Int_2_argbuf_d[0] ? 5'd1 :
                                                     (\lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int0_1_argbuf_d [0] ? 5'd2 :
                                                      (es_2_1MyFalse_2_argbuf_d[0] ? 5'd4 :
                                                       (es_2_1MyTrue_2_argbuf_d[0] ? 5'd8 :
                                                        (lizzieLet6_3QError_Int_2_argbuf_d[0] ? 5'd16 :
                                                         5'd0))))));
  logic [4:0] lizzieLet6_3QNone_Int_2_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_3QNone_Int_2_argbuf_select_q <= 5'd0;
    else
      lizzieLet6_3QNone_Int_2_argbuf_select_q <= (lizzieLet6_3QNone_Int_2_argbuf_done ? 5'd0 :
                                                  lizzieLet6_3QNone_Int_2_argbuf_select_d);
  logic [1:0] lizzieLet6_3QNone_Int_2_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_3QNone_Int_2_argbuf_emit_q <= 2'd0;
    else
      lizzieLet6_3QNone_Int_2_argbuf_emit_q <= (lizzieLet6_3QNone_Int_2_argbuf_done ? 2'd0 :
                                                lizzieLet6_3QNone_Int_2_argbuf_emit_d);
  logic [1:0] lizzieLet6_3QNone_Int_2_argbuf_emit_d;
  assign lizzieLet6_3QNone_Int_2_argbuf_emit_d = (lizzieLet6_3QNone_Int_2_argbuf_emit_q | ({go_16_goMux_choice_d[0],
                                                                                            go_16_goMux_data_d[0]} & {go_16_goMux_choice_r,
                                                                                                                      go_16_goMux_data_r}));
  logic lizzieLet6_3QNone_Int_2_argbuf_done;
  assign lizzieLet6_3QNone_Int_2_argbuf_done = (& lizzieLet6_3QNone_Int_2_argbuf_emit_d);
  assign {lizzieLet6_3QError_Int_2_argbuf_r,
          es_2_1MyTrue_2_argbuf_r,
          es_2_1MyFalse_2_argbuf_r,
          \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int0_1_argbuf_r ,
          lizzieLet6_3QNone_Int_2_argbuf_r} = (lizzieLet6_3QNone_Int_2_argbuf_done ? lizzieLet6_3QNone_Int_2_argbuf_select_d :
                                               5'd0);
  assign go_16_goMux_data_d = ((lizzieLet6_3QNone_Int_2_argbuf_select_d[0] && (! lizzieLet6_3QNone_Int_2_argbuf_emit_q[0])) ? lizzieLet6_3QNone_Int_2_argbuf_d :
                               ((lizzieLet6_3QNone_Int_2_argbuf_select_d[1] && (! lizzieLet6_3QNone_Int_2_argbuf_emit_q[0])) ? \lizzieLet39_3Lcall_f''''''''_f''''''''_Int_Int0_1_argbuf_d  :
                                ((lizzieLet6_3QNone_Int_2_argbuf_select_d[2] && (! lizzieLet6_3QNone_Int_2_argbuf_emit_q[0])) ? es_2_1MyFalse_2_argbuf_d :
                                 ((lizzieLet6_3QNone_Int_2_argbuf_select_d[3] && (! lizzieLet6_3QNone_Int_2_argbuf_emit_q[0])) ? es_2_1MyTrue_2_argbuf_d :
                                  ((lizzieLet6_3QNone_Int_2_argbuf_select_d[4] && (! lizzieLet6_3QNone_Int_2_argbuf_emit_q[0])) ? lizzieLet6_3QError_Int_2_argbuf_d :
                                   1'd0)))));
  assign go_16_goMux_choice_d = ((lizzieLet6_3QNone_Int_2_argbuf_select_d[0] && (! lizzieLet6_3QNone_Int_2_argbuf_emit_q[1])) ? C1_5_dc(1'd1) :
                                 ((lizzieLet6_3QNone_Int_2_argbuf_select_d[1] && (! lizzieLet6_3QNone_Int_2_argbuf_emit_q[1])) ? C2_5_dc(1'd1) :
                                  ((lizzieLet6_3QNone_Int_2_argbuf_select_d[2] && (! lizzieLet6_3QNone_Int_2_argbuf_emit_q[1])) ? C3_5_dc(1'd1) :
                                   ((lizzieLet6_3QNone_Int_2_argbuf_select_d[3] && (! lizzieLet6_3QNone_Int_2_argbuf_emit_q[1])) ? C4_5_dc(1'd1) :
                                    ((lizzieLet6_3QNone_Int_2_argbuf_select_d[4] && (! lizzieLet6_3QNone_Int_2_argbuf_emit_q[1])) ? C5_5_dc(1'd1) :
                                     {3'd0, 1'd0})))));
  
  /* fork (Ty Go) : (lizzieLet6_3QVal_Int,Go) > [(lizzieLet6_3QVal_Int_1,Go),
                                            (lizzieLet6_3QVal_Int_2,Go),
                                            (lizzieLet6_3QVal_Int_3,Go)] */
  logic [2:0] lizzieLet6_3QVal_Int_emitted;
  logic [2:0] lizzieLet6_3QVal_Int_done;
  assign lizzieLet6_3QVal_Int_1_d = (lizzieLet6_3QVal_Int_d[0] && (! lizzieLet6_3QVal_Int_emitted[0]));
  assign lizzieLet6_3QVal_Int_2_d = (lizzieLet6_3QVal_Int_d[0] && (! lizzieLet6_3QVal_Int_emitted[1]));
  assign lizzieLet6_3QVal_Int_3_d = (lizzieLet6_3QVal_Int_d[0] && (! lizzieLet6_3QVal_Int_emitted[2]));
  assign lizzieLet6_3QVal_Int_done = (lizzieLet6_3QVal_Int_emitted | ({lizzieLet6_3QVal_Int_3_d[0],
                                                                       lizzieLet6_3QVal_Int_2_d[0],
                                                                       lizzieLet6_3QVal_Int_1_d[0]} & {lizzieLet6_3QVal_Int_3_r,
                                                                                                       lizzieLet6_3QVal_Int_2_r,
                                                                                                       lizzieLet6_3QVal_Int_1_r}));
  assign lizzieLet6_3QVal_Int_r = (& lizzieLet6_3QVal_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_3QVal_Int_emitted <= 3'd0;
    else
      lizzieLet6_3QVal_Int_emitted <= (lizzieLet6_3QVal_Int_r ? 3'd0 :
                                       lizzieLet6_3QVal_Int_done);
  
  /* buf (Ty Go) : (lizzieLet6_3QVal_Int_1,Go) > (lizzieLet6_3QVal_Int_1_argbuf,Go) */
  Go_t lizzieLet6_3QVal_Int_1_bufchan_d;
  logic lizzieLet6_3QVal_Int_1_bufchan_r;
  assign lizzieLet6_3QVal_Int_1_r = ((! lizzieLet6_3QVal_Int_1_bufchan_d[0]) || lizzieLet6_3QVal_Int_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_3QVal_Int_1_bufchan_d <= 1'd0;
    else
      if (lizzieLet6_3QVal_Int_1_r)
        lizzieLet6_3QVal_Int_1_bufchan_d <= lizzieLet6_3QVal_Int_1_d;
  Go_t lizzieLet6_3QVal_Int_1_bufchan_buf;
  assign lizzieLet6_3QVal_Int_1_bufchan_r = (! lizzieLet6_3QVal_Int_1_bufchan_buf[0]);
  assign lizzieLet6_3QVal_Int_1_argbuf_d = (lizzieLet6_3QVal_Int_1_bufchan_buf[0] ? lizzieLet6_3QVal_Int_1_bufchan_buf :
                                            lizzieLet6_3QVal_Int_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_3QVal_Int_1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet6_3QVal_Int_1_argbuf_r && lizzieLet6_3QVal_Int_1_bufchan_buf[0]))
        lizzieLet6_3QVal_Int_1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet6_3QVal_Int_1_argbuf_r) && (! lizzieLet6_3QVal_Int_1_bufchan_buf[0])))
        lizzieLet6_3QVal_Int_1_bufchan_buf <= lizzieLet6_3QVal_Int_1_bufchan_d;
  
  /* dcon (Ty TupGo___MyDTInt_Int___Int,
      Dcon TupGo___MyDTInt_Int___Int) : [(lizzieLet6_3QVal_Int_1_argbuf,Go),
                                         (lizzieLet6_5QVal_Int_1_argbuf,MyDTInt_Int),
                                         (va8x_1_argbuf,Int)] > (applyfnInt_Int_5TupGo___MyDTInt_Int___Int3,TupGo___MyDTInt_Int___Int) */
  assign applyfnInt_Int_5TupGo___MyDTInt_Int___Int3_d = TupGo___MyDTInt_Int___Int_dc((& {lizzieLet6_3QVal_Int_1_argbuf_d[0],
                                                                                         lizzieLet6_5QVal_Int_1_argbuf_d[0],
                                                                                         va8x_1_argbuf_d[0]}), lizzieLet6_3QVal_Int_1_argbuf_d, lizzieLet6_5QVal_Int_1_argbuf_d, va8x_1_argbuf_d);
  assign {lizzieLet6_3QVal_Int_1_argbuf_r,
          lizzieLet6_5QVal_Int_1_argbuf_r,
          va8x_1_argbuf_r} = {3 {(applyfnInt_Int_5TupGo___MyDTInt_Int___Int3_r && applyfnInt_Int_5TupGo___MyDTInt_Int___Int3_d[0])}};
  
  /* buf (Ty Go) : (lizzieLet6_3QVal_Int_2,Go) > (lizzieLet6_3QVal_Int_2_argbuf,Go) */
  Go_t lizzieLet6_3QVal_Int_2_bufchan_d;
  logic lizzieLet6_3QVal_Int_2_bufchan_r;
  assign lizzieLet6_3QVal_Int_2_r = ((! lizzieLet6_3QVal_Int_2_bufchan_d[0]) || lizzieLet6_3QVal_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_3QVal_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet6_3QVal_Int_2_r)
        lizzieLet6_3QVal_Int_2_bufchan_d <= lizzieLet6_3QVal_Int_2_d;
  Go_t lizzieLet6_3QVal_Int_2_bufchan_buf;
  assign lizzieLet6_3QVal_Int_2_bufchan_r = (! lizzieLet6_3QVal_Int_2_bufchan_buf[0]);
  assign lizzieLet6_3QVal_Int_2_argbuf_d = (lizzieLet6_3QVal_Int_2_bufchan_buf[0] ? lizzieLet6_3QVal_Int_2_bufchan_buf :
                                            lizzieLet6_3QVal_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_3QVal_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet6_3QVal_Int_2_argbuf_r && lizzieLet6_3QVal_Int_2_bufchan_buf[0]))
        lizzieLet6_3QVal_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet6_3QVal_Int_2_argbuf_r) && (! lizzieLet6_3QVal_Int_2_bufchan_buf[0])))
        lizzieLet6_3QVal_Int_2_bufchan_buf <= lizzieLet6_3QVal_Int_2_bufchan_d;
  
  /* dcon (Ty TupGo___MyDTInt_Bool___Int,
      Dcon TupGo___MyDTInt_Bool___Int) : [(lizzieLet6_3QVal_Int_2_argbuf,Go),
                                          (lizzieLet6_4QVal_Int_1_argbuf,MyDTInt_Bool),
                                          (es_1_1_argbuf,Int)] > (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int2,TupGo___MyDTInt_Bool___Int) */
  assign applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int2_d = TupGo___MyDTInt_Bool___Int_dc((& {lizzieLet6_3QVal_Int_2_argbuf_d[0],
                                                                                            lizzieLet6_4QVal_Int_1_argbuf_d[0],
                                                                                            es_1_1_argbuf_d[0]}), lizzieLet6_3QVal_Int_2_argbuf_d, lizzieLet6_4QVal_Int_1_argbuf_d, es_1_1_argbuf_d);
  assign {lizzieLet6_3QVal_Int_2_argbuf_r,
          lizzieLet6_4QVal_Int_1_argbuf_r,
          es_1_1_argbuf_r} = {3 {(applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int2_r && applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int2_d[0])}};
  
  /* demux (Ty QTree_Int,
       Ty MyDTInt_Bool) : (lizzieLet6_4,QTree_Int) (is_z_mapa8v_goMux_mux,MyDTInt_Bool) > [(_3,MyDTInt_Bool),
                                                                                           (lizzieLet6_4QVal_Int,MyDTInt_Bool),
                                                                                           (lizzieLet6_4QNode_Int,MyDTInt_Bool),
                                                                                           (_2,MyDTInt_Bool)] */
  logic [3:0] is_z_mapa8v_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet6_4_d[0] && is_z_mapa8v_goMux_mux_d[0]))
      unique case (lizzieLet6_4_d[2:1])
        2'd0: is_z_mapa8v_goMux_mux_onehotd = 4'd1;
        2'd1: is_z_mapa8v_goMux_mux_onehotd = 4'd2;
        2'd2: is_z_mapa8v_goMux_mux_onehotd = 4'd4;
        2'd3: is_z_mapa8v_goMux_mux_onehotd = 4'd8;
        default: is_z_mapa8v_goMux_mux_onehotd = 4'd0;
      endcase
    else is_z_mapa8v_goMux_mux_onehotd = 4'd0;
  assign _3_d = is_z_mapa8v_goMux_mux_onehotd[0];
  assign lizzieLet6_4QVal_Int_d = is_z_mapa8v_goMux_mux_onehotd[1];
  assign lizzieLet6_4QNode_Int_d = is_z_mapa8v_goMux_mux_onehotd[2];
  assign _2_d = is_z_mapa8v_goMux_mux_onehotd[3];
  assign is_z_mapa8v_goMux_mux_r = (| (is_z_mapa8v_goMux_mux_onehotd & {_2_r,
                                                                        lizzieLet6_4QNode_Int_r,
                                                                        lizzieLet6_4QVal_Int_r,
                                                                        _3_r}));
  assign lizzieLet6_4_r = is_z_mapa8v_goMux_mux_r;
  
  /* fork (Ty MyDTInt_Bool) : (lizzieLet6_4QNode_Int,MyDTInt_Bool) > [(lizzieLet6_4QNode_Int_1,MyDTInt_Bool),
                                                                 (lizzieLet6_4QNode_Int_2,MyDTInt_Bool)] */
  logic [1:0] lizzieLet6_4QNode_Int_emitted;
  logic [1:0] lizzieLet6_4QNode_Int_done;
  assign lizzieLet6_4QNode_Int_1_d = (lizzieLet6_4QNode_Int_d[0] && (! lizzieLet6_4QNode_Int_emitted[0]));
  assign lizzieLet6_4QNode_Int_2_d = (lizzieLet6_4QNode_Int_d[0] && (! lizzieLet6_4QNode_Int_emitted[1]));
  assign lizzieLet6_4QNode_Int_done = (lizzieLet6_4QNode_Int_emitted | ({lizzieLet6_4QNode_Int_2_d[0],
                                                                         lizzieLet6_4QNode_Int_1_d[0]} & {lizzieLet6_4QNode_Int_2_r,
                                                                                                          lizzieLet6_4QNode_Int_1_r}));
  assign lizzieLet6_4QNode_Int_r = (& lizzieLet6_4QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_4QNode_Int_emitted <= 2'd0;
    else
      lizzieLet6_4QNode_Int_emitted <= (lizzieLet6_4QNode_Int_r ? 2'd0 :
                                        lizzieLet6_4QNode_Int_done);
  
  /* buf (Ty MyDTInt_Bool) : (lizzieLet6_4QNode_Int_2,MyDTInt_Bool) > (lizzieLet6_4QNode_Int_2_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t lizzieLet6_4QNode_Int_2_bufchan_d;
  logic lizzieLet6_4QNode_Int_2_bufchan_r;
  assign lizzieLet6_4QNode_Int_2_r = ((! lizzieLet6_4QNode_Int_2_bufchan_d[0]) || lizzieLet6_4QNode_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_4QNode_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet6_4QNode_Int_2_r)
        lizzieLet6_4QNode_Int_2_bufchan_d <= lizzieLet6_4QNode_Int_2_d;
  MyDTInt_Bool_t lizzieLet6_4QNode_Int_2_bufchan_buf;
  assign lizzieLet6_4QNode_Int_2_bufchan_r = (! lizzieLet6_4QNode_Int_2_bufchan_buf[0]);
  assign lizzieLet6_4QNode_Int_2_argbuf_d = (lizzieLet6_4QNode_Int_2_bufchan_buf[0] ? lizzieLet6_4QNode_Int_2_bufchan_buf :
                                             lizzieLet6_4QNode_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_4QNode_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet6_4QNode_Int_2_argbuf_r && lizzieLet6_4QNode_Int_2_bufchan_buf[0]))
        lizzieLet6_4QNode_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet6_4QNode_Int_2_argbuf_r) && (! lizzieLet6_4QNode_Int_2_bufchan_buf[0])))
        lizzieLet6_4QNode_Int_2_bufchan_buf <= lizzieLet6_4QNode_Int_2_bufchan_d;
  
  /* buf (Ty MyDTInt_Bool) : (lizzieLet6_4QVal_Int,MyDTInt_Bool) > (lizzieLet6_4QVal_Int_1_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t lizzieLet6_4QVal_Int_bufchan_d;
  logic lizzieLet6_4QVal_Int_bufchan_r;
  assign lizzieLet6_4QVal_Int_r = ((! lizzieLet6_4QVal_Int_bufchan_d[0]) || lizzieLet6_4QVal_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_4QVal_Int_bufchan_d <= 1'd0;
    else
      if (lizzieLet6_4QVal_Int_r)
        lizzieLet6_4QVal_Int_bufchan_d <= lizzieLet6_4QVal_Int_d;
  MyDTInt_Bool_t lizzieLet6_4QVal_Int_bufchan_buf;
  assign lizzieLet6_4QVal_Int_bufchan_r = (! lizzieLet6_4QVal_Int_bufchan_buf[0]);
  assign lizzieLet6_4QVal_Int_1_argbuf_d = (lizzieLet6_4QVal_Int_bufchan_buf[0] ? lizzieLet6_4QVal_Int_bufchan_buf :
                                            lizzieLet6_4QVal_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_4QVal_Int_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet6_4QVal_Int_1_argbuf_r && lizzieLet6_4QVal_Int_bufchan_buf[0]))
        lizzieLet6_4QVal_Int_bufchan_buf <= 1'd0;
      else if (((! lizzieLet6_4QVal_Int_1_argbuf_r) && (! lizzieLet6_4QVal_Int_bufchan_buf[0])))
        lizzieLet6_4QVal_Int_bufchan_buf <= lizzieLet6_4QVal_Int_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty MyDTInt_Int) : (lizzieLet6_5,QTree_Int) (op_mapa8w_goMux_mux,MyDTInt_Int) > [(_1,MyDTInt_Int),
                                                                                       (lizzieLet6_5QVal_Int,MyDTInt_Int),
                                                                                       (lizzieLet6_5QNode_Int,MyDTInt_Int),
                                                                                       (_0,MyDTInt_Int)] */
  logic [3:0] op_mapa8w_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet6_5_d[0] && op_mapa8w_goMux_mux_d[0]))
      unique case (lizzieLet6_5_d[2:1])
        2'd0: op_mapa8w_goMux_mux_onehotd = 4'd1;
        2'd1: op_mapa8w_goMux_mux_onehotd = 4'd2;
        2'd2: op_mapa8w_goMux_mux_onehotd = 4'd4;
        2'd3: op_mapa8w_goMux_mux_onehotd = 4'd8;
        default: op_mapa8w_goMux_mux_onehotd = 4'd0;
      endcase
    else op_mapa8w_goMux_mux_onehotd = 4'd0;
  assign _1_d = op_mapa8w_goMux_mux_onehotd[0];
  assign lizzieLet6_5QVal_Int_d = op_mapa8w_goMux_mux_onehotd[1];
  assign lizzieLet6_5QNode_Int_d = op_mapa8w_goMux_mux_onehotd[2];
  assign _0_d = op_mapa8w_goMux_mux_onehotd[3];
  assign op_mapa8w_goMux_mux_r = (| (op_mapa8w_goMux_mux_onehotd & {_0_r,
                                                                    lizzieLet6_5QNode_Int_r,
                                                                    lizzieLet6_5QVal_Int_r,
                                                                    _1_r}));
  assign lizzieLet6_5_r = op_mapa8w_goMux_mux_r;
  
  /* fork (Ty MyDTInt_Int) : (lizzieLet6_5QNode_Int,MyDTInt_Int) > [(lizzieLet6_5QNode_Int_1,MyDTInt_Int),
                                                               (lizzieLet6_5QNode_Int_2,MyDTInt_Int)] */
  logic [1:0] lizzieLet6_5QNode_Int_emitted;
  logic [1:0] lizzieLet6_5QNode_Int_done;
  assign lizzieLet6_5QNode_Int_1_d = (lizzieLet6_5QNode_Int_d[0] && (! lizzieLet6_5QNode_Int_emitted[0]));
  assign lizzieLet6_5QNode_Int_2_d = (lizzieLet6_5QNode_Int_d[0] && (! lizzieLet6_5QNode_Int_emitted[1]));
  assign lizzieLet6_5QNode_Int_done = (lizzieLet6_5QNode_Int_emitted | ({lizzieLet6_5QNode_Int_2_d[0],
                                                                         lizzieLet6_5QNode_Int_1_d[0]} & {lizzieLet6_5QNode_Int_2_r,
                                                                                                          lizzieLet6_5QNode_Int_1_r}));
  assign lizzieLet6_5QNode_Int_r = (& lizzieLet6_5QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_5QNode_Int_emitted <= 2'd0;
    else
      lizzieLet6_5QNode_Int_emitted <= (lizzieLet6_5QNode_Int_r ? 2'd0 :
                                        lizzieLet6_5QNode_Int_done);
  
  /* buf (Ty MyDTInt_Int) : (lizzieLet6_5QNode_Int_2,MyDTInt_Int) > (lizzieLet6_5QNode_Int_2_argbuf,MyDTInt_Int) */
  MyDTInt_Int_t lizzieLet6_5QNode_Int_2_bufchan_d;
  logic lizzieLet6_5QNode_Int_2_bufchan_r;
  assign lizzieLet6_5QNode_Int_2_r = ((! lizzieLet6_5QNode_Int_2_bufchan_d[0]) || lizzieLet6_5QNode_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_5QNode_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet6_5QNode_Int_2_r)
        lizzieLet6_5QNode_Int_2_bufchan_d <= lizzieLet6_5QNode_Int_2_d;
  MyDTInt_Int_t lizzieLet6_5QNode_Int_2_bufchan_buf;
  assign lizzieLet6_5QNode_Int_2_bufchan_r = (! lizzieLet6_5QNode_Int_2_bufchan_buf[0]);
  assign lizzieLet6_5QNode_Int_2_argbuf_d = (lizzieLet6_5QNode_Int_2_bufchan_buf[0] ? lizzieLet6_5QNode_Int_2_bufchan_buf :
                                             lizzieLet6_5QNode_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_5QNode_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet6_5QNode_Int_2_argbuf_r && lizzieLet6_5QNode_Int_2_bufchan_buf[0]))
        lizzieLet6_5QNode_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet6_5QNode_Int_2_argbuf_r) && (! lizzieLet6_5QNode_Int_2_bufchan_buf[0])))
        lizzieLet6_5QNode_Int_2_bufchan_buf <= lizzieLet6_5QNode_Int_2_bufchan_d;
  
  /* fork (Ty MyDTInt_Int) : (lizzieLet6_5QVal_Int,MyDTInt_Int) > [(lizzieLet6_5QVal_Int_1,MyDTInt_Int),
                                                              (lizzieLet6_5QVal_Int_2,MyDTInt_Int)] */
  logic [1:0] lizzieLet6_5QVal_Int_emitted;
  logic [1:0] lizzieLet6_5QVal_Int_done;
  assign lizzieLet6_5QVal_Int_1_d = (lizzieLet6_5QVal_Int_d[0] && (! lizzieLet6_5QVal_Int_emitted[0]));
  assign lizzieLet6_5QVal_Int_2_d = (lizzieLet6_5QVal_Int_d[0] && (! lizzieLet6_5QVal_Int_emitted[1]));
  assign lizzieLet6_5QVal_Int_done = (lizzieLet6_5QVal_Int_emitted | ({lizzieLet6_5QVal_Int_2_d[0],
                                                                       lizzieLet6_5QVal_Int_1_d[0]} & {lizzieLet6_5QVal_Int_2_r,
                                                                                                       lizzieLet6_5QVal_Int_1_r}));
  assign lizzieLet6_5QVal_Int_r = (& lizzieLet6_5QVal_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_5QVal_Int_emitted <= 2'd0;
    else
      lizzieLet6_5QVal_Int_emitted <= (lizzieLet6_5QVal_Int_r ? 2'd0 :
                                       lizzieLet6_5QVal_Int_done);
  
  /* buf (Ty MyDTInt_Int) : (lizzieLet6_5QVal_Int_1,MyDTInt_Int) > (lizzieLet6_5QVal_Int_1_argbuf,MyDTInt_Int) */
  MyDTInt_Int_t lizzieLet6_5QVal_Int_1_bufchan_d;
  logic lizzieLet6_5QVal_Int_1_bufchan_r;
  assign lizzieLet6_5QVal_Int_1_r = ((! lizzieLet6_5QVal_Int_1_bufchan_d[0]) || lizzieLet6_5QVal_Int_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_5QVal_Int_1_bufchan_d <= 1'd0;
    else
      if (lizzieLet6_5QVal_Int_1_r)
        lizzieLet6_5QVal_Int_1_bufchan_d <= lizzieLet6_5QVal_Int_1_d;
  MyDTInt_Int_t lizzieLet6_5QVal_Int_1_bufchan_buf;
  assign lizzieLet6_5QVal_Int_1_bufchan_r = (! lizzieLet6_5QVal_Int_1_bufchan_buf[0]);
  assign lizzieLet6_5QVal_Int_1_argbuf_d = (lizzieLet6_5QVal_Int_1_bufchan_buf[0] ? lizzieLet6_5QVal_Int_1_bufchan_buf :
                                            lizzieLet6_5QVal_Int_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_5QVal_Int_1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet6_5QVal_Int_1_argbuf_r && lizzieLet6_5QVal_Int_1_bufchan_buf[0]))
        lizzieLet6_5QVal_Int_1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet6_5QVal_Int_1_argbuf_r) && (! lizzieLet6_5QVal_Int_1_bufchan_buf[0])))
        lizzieLet6_5QVal_Int_1_bufchan_buf <= lizzieLet6_5QVal_Int_1_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_CTf''''''''_f''''''''_Int_Int) : (lizzieLet6_6,QTree_Int) (sc_0_1_goMux_mux,Pointer_CTf''''''''_f''''''''_Int_Int) > [(lizzieLet6_6QNone_Int,Pointer_CTf''''''''_f''''''''_Int_Int),
                                                                                                                                        (lizzieLet6_6QVal_Int,Pointer_CTf''''''''_f''''''''_Int_Int),
                                                                                                                                        (lizzieLet6_6QNode_Int,Pointer_CTf''''''''_f''''''''_Int_Int),
                                                                                                                                        (lizzieLet6_6QError_Int,Pointer_CTf''''''''_f''''''''_Int_Int)] */
  logic [3:0] sc_0_1_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet6_6_d[0] && sc_0_1_goMux_mux_d[0]))
      unique case (lizzieLet6_6_d[2:1])
        2'd0: sc_0_1_goMux_mux_onehotd = 4'd1;
        2'd1: sc_0_1_goMux_mux_onehotd = 4'd2;
        2'd2: sc_0_1_goMux_mux_onehotd = 4'd4;
        2'd3: sc_0_1_goMux_mux_onehotd = 4'd8;
        default: sc_0_1_goMux_mux_onehotd = 4'd0;
      endcase
    else sc_0_1_goMux_mux_onehotd = 4'd0;
  assign lizzieLet6_6QNone_Int_d = {sc_0_1_goMux_mux_d[16:1],
                                    sc_0_1_goMux_mux_onehotd[0]};
  assign lizzieLet6_6QVal_Int_d = {sc_0_1_goMux_mux_d[16:1],
                                   sc_0_1_goMux_mux_onehotd[1]};
  assign lizzieLet6_6QNode_Int_d = {sc_0_1_goMux_mux_d[16:1],
                                    sc_0_1_goMux_mux_onehotd[2]};
  assign lizzieLet6_6QError_Int_d = {sc_0_1_goMux_mux_d[16:1],
                                     sc_0_1_goMux_mux_onehotd[3]};
  assign sc_0_1_goMux_mux_r = (| (sc_0_1_goMux_mux_onehotd & {lizzieLet6_6QError_Int_r,
                                                              lizzieLet6_6QNode_Int_r,
                                                              lizzieLet6_6QVal_Int_r,
                                                              lizzieLet6_6QNone_Int_r}));
  assign lizzieLet6_6_r = sc_0_1_goMux_mux_r;
  
  /* buf (Ty Pointer_CTf''''''''_f''''''''_Int_Int) : (lizzieLet6_6QError_Int,Pointer_CTf''''''''_f''''''''_Int_Int) > (lizzieLet6_6QError_Int_1_argbuf,Pointer_CTf''''''''_f''''''''_Int_Int) */
  \Pointer_CTf''''''''_f''''''''_Int_Int_t  lizzieLet6_6QError_Int_bufchan_d;
  logic lizzieLet6_6QError_Int_bufchan_r;
  assign lizzieLet6_6QError_Int_r = ((! lizzieLet6_6QError_Int_bufchan_d[0]) || lizzieLet6_6QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_6QError_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet6_6QError_Int_r)
        lizzieLet6_6QError_Int_bufchan_d <= lizzieLet6_6QError_Int_d;
  \Pointer_CTf''''''''_f''''''''_Int_Int_t  lizzieLet6_6QError_Int_bufchan_buf;
  assign lizzieLet6_6QError_Int_bufchan_r = (! lizzieLet6_6QError_Int_bufchan_buf[0]);
  assign lizzieLet6_6QError_Int_1_argbuf_d = (lizzieLet6_6QError_Int_bufchan_buf[0] ? lizzieLet6_6QError_Int_bufchan_buf :
                                              lizzieLet6_6QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_6QError_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet6_6QError_Int_1_argbuf_r && lizzieLet6_6QError_Int_bufchan_buf[0]))
        lizzieLet6_6QError_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet6_6QError_Int_1_argbuf_r) && (! lizzieLet6_6QError_Int_bufchan_buf[0])))
        lizzieLet6_6QError_Int_bufchan_buf <= lizzieLet6_6QError_Int_bufchan_d;
  
  /* dcon (Ty CTf''''''''_f''''''''_Int_Int,
      Dcon Lcall_f''''''''_f''''''''_Int_Int3) : [(lizzieLet6_6QNode_Int,Pointer_CTf''''''''_f''''''''_Int_Int),
                                                  (tla8y_destruct,Pointer_QTree_Int),
                                                  (lizzieLet6_4QNode_Int_1,MyDTInt_Bool),
                                                  (lizzieLet6_5QNode_Int_1,MyDTInt_Int),
                                                  (tra8z_destruct,Pointer_QTree_Int),
                                                  (bla8A_destruct,Pointer_QTree_Int)] > (lizzieLet6_6QNode_Int_1tla8y_1lizzieLet6_4QNode_Int_1lizzieLet6_5QNode_Int_1tra8z_1bla8A_1Lcall_f''''''''_f''''''''_Int_Int3,CTf''''''''_f''''''''_Int_Int) */
  assign \lizzieLet6_6QNode_Int_1tla8y_1lizzieLet6_4QNode_Int_1lizzieLet6_5QNode_Int_1tra8z_1bla8A_1Lcall_f''''''''_f''''''''_Int_Int3_d  = \Lcall_f''''''''_f''''''''_Int_Int3_dc ((& {lizzieLet6_6QNode_Int_d[0],
                                                                                                                                                                                        tla8y_destruct_d[0],
                                                                                                                                                                                        lizzieLet6_4QNode_Int_1_d[0],
                                                                                                                                                                                        lizzieLet6_5QNode_Int_1_d[0],
                                                                                                                                                                                        tra8z_destruct_d[0],
                                                                                                                                                                                        bla8A_destruct_d[0]}), lizzieLet6_6QNode_Int_d, tla8y_destruct_d, lizzieLet6_4QNode_Int_1_d, lizzieLet6_5QNode_Int_1_d, tra8z_destruct_d, bla8A_destruct_d);
  assign {lizzieLet6_6QNode_Int_r,
          tla8y_destruct_r,
          lizzieLet6_4QNode_Int_1_r,
          lizzieLet6_5QNode_Int_1_r,
          tra8z_destruct_r,
          bla8A_destruct_r} = {6 {(\lizzieLet6_6QNode_Int_1tla8y_1lizzieLet6_4QNode_Int_1lizzieLet6_5QNode_Int_1tra8z_1bla8A_1Lcall_f''''''''_f''''''''_Int_Int3_r  && \lizzieLet6_6QNode_Int_1tla8y_1lizzieLet6_4QNode_Int_1lizzieLet6_5QNode_Int_1tra8z_1bla8A_1Lcall_f''''''''_f''''''''_Int_Int3_d [0])}};
  
  /* buf (Ty CTf''''''''_f''''''''_Int_Int) : (lizzieLet6_6QNode_Int_1tla8y_1lizzieLet6_4QNode_Int_1lizzieLet6_5QNode_Int_1tra8z_1bla8A_1Lcall_f''''''''_f''''''''_Int_Int3,CTf''''''''_f''''''''_Int_Int) > (lizzieLet10_1_argbuf,CTf''''''''_f''''''''_Int_Int) */
  \CTf''''''''_f''''''''_Int_Int_t  \lizzieLet6_6QNode_Int_1tla8y_1lizzieLet6_4QNode_Int_1lizzieLet6_5QNode_Int_1tra8z_1bla8A_1Lcall_f''''''''_f''''''''_Int_Int3_bufchan_d ;
  logic \lizzieLet6_6QNode_Int_1tla8y_1lizzieLet6_4QNode_Int_1lizzieLet6_5QNode_Int_1tra8z_1bla8A_1Lcall_f''''''''_f''''''''_Int_Int3_bufchan_r ;
  assign \lizzieLet6_6QNode_Int_1tla8y_1lizzieLet6_4QNode_Int_1lizzieLet6_5QNode_Int_1tra8z_1bla8A_1Lcall_f''''''''_f''''''''_Int_Int3_r  = ((! \lizzieLet6_6QNode_Int_1tla8y_1lizzieLet6_4QNode_Int_1lizzieLet6_5QNode_Int_1tra8z_1bla8A_1Lcall_f''''''''_f''''''''_Int_Int3_bufchan_d [0]) || \lizzieLet6_6QNode_Int_1tla8y_1lizzieLet6_4QNode_Int_1lizzieLet6_5QNode_Int_1tra8z_1bla8A_1Lcall_f''''''''_f''''''''_Int_Int3_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet6_6QNode_Int_1tla8y_1lizzieLet6_4QNode_Int_1lizzieLet6_5QNode_Int_1tra8z_1bla8A_1Lcall_f''''''''_f''''''''_Int_Int3_bufchan_d  <= {67'd0,
                                                                                                                                                   1'd0};
    else
      if (\lizzieLet6_6QNode_Int_1tla8y_1lizzieLet6_4QNode_Int_1lizzieLet6_5QNode_Int_1tra8z_1bla8A_1Lcall_f''''''''_f''''''''_Int_Int3_r )
        \lizzieLet6_6QNode_Int_1tla8y_1lizzieLet6_4QNode_Int_1lizzieLet6_5QNode_Int_1tra8z_1bla8A_1Lcall_f''''''''_f''''''''_Int_Int3_bufchan_d  <= \lizzieLet6_6QNode_Int_1tla8y_1lizzieLet6_4QNode_Int_1lizzieLet6_5QNode_Int_1tra8z_1bla8A_1Lcall_f''''''''_f''''''''_Int_Int3_d ;
  \CTf''''''''_f''''''''_Int_Int_t  \lizzieLet6_6QNode_Int_1tla8y_1lizzieLet6_4QNode_Int_1lizzieLet6_5QNode_Int_1tra8z_1bla8A_1Lcall_f''''''''_f''''''''_Int_Int3_bufchan_buf ;
  assign \lizzieLet6_6QNode_Int_1tla8y_1lizzieLet6_4QNode_Int_1lizzieLet6_5QNode_Int_1tra8z_1bla8A_1Lcall_f''''''''_f''''''''_Int_Int3_bufchan_r  = (! \lizzieLet6_6QNode_Int_1tla8y_1lizzieLet6_4QNode_Int_1lizzieLet6_5QNode_Int_1tra8z_1bla8A_1Lcall_f''''''''_f''''''''_Int_Int3_bufchan_buf [0]);
  assign lizzieLet10_1_argbuf_d = (\lizzieLet6_6QNode_Int_1tla8y_1lizzieLet6_4QNode_Int_1lizzieLet6_5QNode_Int_1tra8z_1bla8A_1Lcall_f''''''''_f''''''''_Int_Int3_bufchan_buf [0] ? \lizzieLet6_6QNode_Int_1tla8y_1lizzieLet6_4QNode_Int_1lizzieLet6_5QNode_Int_1tra8z_1bla8A_1Lcall_f''''''''_f''''''''_Int_Int3_bufchan_buf  :
                                   \lizzieLet6_6QNode_Int_1tla8y_1lizzieLet6_4QNode_Int_1lizzieLet6_5QNode_Int_1tra8z_1bla8A_1Lcall_f''''''''_f''''''''_Int_Int3_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet6_6QNode_Int_1tla8y_1lizzieLet6_4QNode_Int_1lizzieLet6_5QNode_Int_1tra8z_1bla8A_1Lcall_f''''''''_f''''''''_Int_Int3_bufchan_buf  <= {67'd0,
                                                                                                                                                     1'd0};
    else
      if ((lizzieLet10_1_argbuf_r && \lizzieLet6_6QNode_Int_1tla8y_1lizzieLet6_4QNode_Int_1lizzieLet6_5QNode_Int_1tra8z_1bla8A_1Lcall_f''''''''_f''''''''_Int_Int3_bufchan_buf [0]))
        \lizzieLet6_6QNode_Int_1tla8y_1lizzieLet6_4QNode_Int_1lizzieLet6_5QNode_Int_1tra8z_1bla8A_1Lcall_f''''''''_f''''''''_Int_Int3_bufchan_buf  <= {67'd0,
                                                                                                                                                       1'd0};
      else if (((! lizzieLet10_1_argbuf_r) && (! \lizzieLet6_6QNode_Int_1tla8y_1lizzieLet6_4QNode_Int_1lizzieLet6_5QNode_Int_1tra8z_1bla8A_1Lcall_f''''''''_f''''''''_Int_Int3_bufchan_buf [0])))
        \lizzieLet6_6QNode_Int_1tla8y_1lizzieLet6_4QNode_Int_1lizzieLet6_5QNode_Int_1tra8z_1bla8A_1Lcall_f''''''''_f''''''''_Int_Int3_bufchan_buf  <= \lizzieLet6_6QNode_Int_1tla8y_1lizzieLet6_4QNode_Int_1lizzieLet6_5QNode_Int_1tra8z_1bla8A_1Lcall_f''''''''_f''''''''_Int_Int3_bufchan_d ;
  
  /* buf (Ty Pointer_CTf''''''''_f''''''''_Int_Int) : (lizzieLet6_6QNone_Int,Pointer_CTf''''''''_f''''''''_Int_Int) > (lizzieLet6_6QNone_Int_1_argbuf,Pointer_CTf''''''''_f''''''''_Int_Int) */
  \Pointer_CTf''''''''_f''''''''_Int_Int_t  lizzieLet6_6QNone_Int_bufchan_d;
  logic lizzieLet6_6QNone_Int_bufchan_r;
  assign lizzieLet6_6QNone_Int_r = ((! lizzieLet6_6QNone_Int_bufchan_d[0]) || lizzieLet6_6QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_6QNone_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet6_6QNone_Int_r)
        lizzieLet6_6QNone_Int_bufchan_d <= lizzieLet6_6QNone_Int_d;
  \Pointer_CTf''''''''_f''''''''_Int_Int_t  lizzieLet6_6QNone_Int_bufchan_buf;
  assign lizzieLet6_6QNone_Int_bufchan_r = (! lizzieLet6_6QNone_Int_bufchan_buf[0]);
  assign lizzieLet6_6QNone_Int_1_argbuf_d = (lizzieLet6_6QNone_Int_bufchan_buf[0] ? lizzieLet6_6QNone_Int_bufchan_buf :
                                             lizzieLet6_6QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_6QNone_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet6_6QNone_Int_1_argbuf_r && lizzieLet6_6QNone_Int_bufchan_buf[0]))
        lizzieLet6_6QNone_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet6_6QNone_Int_1_argbuf_r) && (! lizzieLet6_6QNone_Int_bufchan_buf[0])))
        lizzieLet6_6QNone_Int_bufchan_buf <= lizzieLet6_6QNone_Int_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (m1a8C_goMux_mux,Pointer_QTree_Int) > (m1a8C_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t m1a8C_goMux_mux_bufchan_d;
  logic m1a8C_goMux_mux_bufchan_r;
  assign m1a8C_goMux_mux_r = ((! m1a8C_goMux_mux_bufchan_d[0]) || m1a8C_goMux_mux_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m1a8C_goMux_mux_bufchan_d <= {16'd0, 1'd0};
    else
      if (m1a8C_goMux_mux_r)
        m1a8C_goMux_mux_bufchan_d <= m1a8C_goMux_mux_d;
  Pointer_QTree_Int_t m1a8C_goMux_mux_bufchan_buf;
  assign m1a8C_goMux_mux_bufchan_r = (! m1a8C_goMux_mux_bufchan_buf[0]);
  assign m1a8C_1_argbuf_d = (m1a8C_goMux_mux_bufchan_buf[0] ? m1a8C_goMux_mux_bufchan_buf :
                             m1a8C_goMux_mux_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m1a8C_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((m1a8C_1_argbuf_r && m1a8C_goMux_mux_bufchan_buf[0]))
        m1a8C_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
      else if (((! m1a8C_1_argbuf_r) && (! m1a8C_goMux_mux_bufchan_buf[0])))
        m1a8C_goMux_mux_bufchan_buf <= m1a8C_goMux_mux_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (m2a8D_goMux_mux,Pointer_QTree_Int) > (m2a8D_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t m2a8D_goMux_mux_bufchan_d;
  logic m2a8D_goMux_mux_bufchan_r;
  assign m2a8D_goMux_mux_r = ((! m2a8D_goMux_mux_bufchan_d[0]) || m2a8D_goMux_mux_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m2a8D_goMux_mux_bufchan_d <= {16'd0, 1'd0};
    else
      if (m2a8D_goMux_mux_r)
        m2a8D_goMux_mux_bufchan_d <= m2a8D_goMux_mux_d;
  Pointer_QTree_Int_t m2a8D_goMux_mux_bufchan_buf;
  assign m2a8D_goMux_mux_bufchan_r = (! m2a8D_goMux_mux_bufchan_buf[0]);
  assign m2a8D_1_argbuf_d = (m2a8D_goMux_mux_bufchan_buf[0] ? m2a8D_goMux_mux_bufchan_buf :
                             m2a8D_goMux_mux_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m2a8D_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((m2a8D_1_argbuf_r && m2a8D_goMux_mux_bufchan_buf[0]))
        m2a8D_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
      else if (((! m2a8D_1_argbuf_r) && (! m2a8D_goMux_mux_bufchan_buf[0])))
        m2a8D_goMux_mux_bufchan_buf <= m2a8D_goMux_mux_bufchan_d;
  
  /* buf (Ty MyDTInt_Int_Int) : (op_adda8H_2_2,MyDTInt_Int_Int) > (op_adda8H_2_2_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t op_adda8H_2_2_bufchan_d;
  logic op_adda8H_2_2_bufchan_r;
  assign op_adda8H_2_2_r = ((! op_adda8H_2_2_bufchan_d[0]) || op_adda8H_2_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) op_adda8H_2_2_bufchan_d <= 1'd0;
    else
      if (op_adda8H_2_2_r) op_adda8H_2_2_bufchan_d <= op_adda8H_2_2_d;
  MyDTInt_Int_Int_t op_adda8H_2_2_bufchan_buf;
  assign op_adda8H_2_2_bufchan_r = (! op_adda8H_2_2_bufchan_buf[0]);
  assign op_adda8H_2_2_argbuf_d = (op_adda8H_2_2_bufchan_buf[0] ? op_adda8H_2_2_bufchan_buf :
                                   op_adda8H_2_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) op_adda8H_2_2_bufchan_buf <= 1'd0;
    else
      if ((op_adda8H_2_2_argbuf_r && op_adda8H_2_2_bufchan_buf[0]))
        op_adda8H_2_2_bufchan_buf <= 1'd0;
      else if (((! op_adda8H_2_2_argbuf_r) && (! op_adda8H_2_2_bufchan_buf[0])))
        op_adda8H_2_2_bufchan_buf <= op_adda8H_2_2_bufchan_d;
  
  /* fork (Ty MyDTInt_Int_Int) : (op_adda8H_2_destruct,MyDTInt_Int_Int) > [(op_adda8H_2_1,MyDTInt_Int_Int),
                                                                      (op_adda8H_2_2,MyDTInt_Int_Int)] */
  logic [1:0] op_adda8H_2_destruct_emitted;
  logic [1:0] op_adda8H_2_destruct_done;
  assign op_adda8H_2_1_d = (op_adda8H_2_destruct_d[0] && (! op_adda8H_2_destruct_emitted[0]));
  assign op_adda8H_2_2_d = (op_adda8H_2_destruct_d[0] && (! op_adda8H_2_destruct_emitted[1]));
  assign op_adda8H_2_destruct_done = (op_adda8H_2_destruct_emitted | ({op_adda8H_2_2_d[0],
                                                                       op_adda8H_2_1_d[0]} & {op_adda8H_2_2_r,
                                                                                              op_adda8H_2_1_r}));
  assign op_adda8H_2_destruct_r = (& op_adda8H_2_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) op_adda8H_2_destruct_emitted <= 2'd0;
    else
      op_adda8H_2_destruct_emitted <= (op_adda8H_2_destruct_r ? 2'd0 :
                                       op_adda8H_2_destruct_done);
  
  /* buf (Ty MyDTInt_Int_Int) : (op_adda8H_3_2,MyDTInt_Int_Int) > (op_adda8H_3_2_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t op_adda8H_3_2_bufchan_d;
  logic op_adda8H_3_2_bufchan_r;
  assign op_adda8H_3_2_r = ((! op_adda8H_3_2_bufchan_d[0]) || op_adda8H_3_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) op_adda8H_3_2_bufchan_d <= 1'd0;
    else
      if (op_adda8H_3_2_r) op_adda8H_3_2_bufchan_d <= op_adda8H_3_2_d;
  MyDTInt_Int_Int_t op_adda8H_3_2_bufchan_buf;
  assign op_adda8H_3_2_bufchan_r = (! op_adda8H_3_2_bufchan_buf[0]);
  assign op_adda8H_3_2_argbuf_d = (op_adda8H_3_2_bufchan_buf[0] ? op_adda8H_3_2_bufchan_buf :
                                   op_adda8H_3_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) op_adda8H_3_2_bufchan_buf <= 1'd0;
    else
      if ((op_adda8H_3_2_argbuf_r && op_adda8H_3_2_bufchan_buf[0]))
        op_adda8H_3_2_bufchan_buf <= 1'd0;
      else if (((! op_adda8H_3_2_argbuf_r) && (! op_adda8H_3_2_bufchan_buf[0])))
        op_adda8H_3_2_bufchan_buf <= op_adda8H_3_2_bufchan_d;
  
  /* fork (Ty MyDTInt_Int_Int) : (op_adda8H_3_destruct,MyDTInt_Int_Int) > [(op_adda8H_3_1,MyDTInt_Int_Int),
                                                                      (op_adda8H_3_2,MyDTInt_Int_Int)] */
  logic [1:0] op_adda8H_3_destruct_emitted;
  logic [1:0] op_adda8H_3_destruct_done;
  assign op_adda8H_3_1_d = (op_adda8H_3_destruct_d[0] && (! op_adda8H_3_destruct_emitted[0]));
  assign op_adda8H_3_2_d = (op_adda8H_3_destruct_d[0] && (! op_adda8H_3_destruct_emitted[1]));
  assign op_adda8H_3_destruct_done = (op_adda8H_3_destruct_emitted | ({op_adda8H_3_2_d[0],
                                                                       op_adda8H_3_1_d[0]} & {op_adda8H_3_2_r,
                                                                                              op_adda8H_3_1_r}));
  assign op_adda8H_3_destruct_r = (& op_adda8H_3_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) op_adda8H_3_destruct_emitted <= 2'd0;
    else
      op_adda8H_3_destruct_emitted <= (op_adda8H_3_destruct_r ? 2'd0 :
                                       op_adda8H_3_destruct_done);
  
  /* buf (Ty MyDTInt_Int_Int) : (op_adda8H_4_destruct,MyDTInt_Int_Int) > (op_adda8H_4_1_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t op_adda8H_4_destruct_bufchan_d;
  logic op_adda8H_4_destruct_bufchan_r;
  assign op_adda8H_4_destruct_r = ((! op_adda8H_4_destruct_bufchan_d[0]) || op_adda8H_4_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) op_adda8H_4_destruct_bufchan_d <= 1'd0;
    else
      if (op_adda8H_4_destruct_r)
        op_adda8H_4_destruct_bufchan_d <= op_adda8H_4_destruct_d;
  MyDTInt_Int_Int_t op_adda8H_4_destruct_bufchan_buf;
  assign op_adda8H_4_destruct_bufchan_r = (! op_adda8H_4_destruct_bufchan_buf[0]);
  assign op_adda8H_4_1_argbuf_d = (op_adda8H_4_destruct_bufchan_buf[0] ? op_adda8H_4_destruct_bufchan_buf :
                                   op_adda8H_4_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) op_adda8H_4_destruct_bufchan_buf <= 1'd0;
    else
      if ((op_adda8H_4_1_argbuf_r && op_adda8H_4_destruct_bufchan_buf[0]))
        op_adda8H_4_destruct_bufchan_buf <= 1'd0;
      else if (((! op_adda8H_4_1_argbuf_r) && (! op_adda8H_4_destruct_bufchan_buf[0])))
        op_adda8H_4_destruct_bufchan_buf <= op_adda8H_4_destruct_bufchan_d;
  
  /* buf (Ty MyDTInt_Int) : (op_mapa8F_2_2,MyDTInt_Int) > (op_mapa8F_2_2_argbuf,MyDTInt_Int) */
  MyDTInt_Int_t op_mapa8F_2_2_bufchan_d;
  logic op_mapa8F_2_2_bufchan_r;
  assign op_mapa8F_2_2_r = ((! op_mapa8F_2_2_bufchan_d[0]) || op_mapa8F_2_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) op_mapa8F_2_2_bufchan_d <= 1'd0;
    else
      if (op_mapa8F_2_2_r) op_mapa8F_2_2_bufchan_d <= op_mapa8F_2_2_d;
  MyDTInt_Int_t op_mapa8F_2_2_bufchan_buf;
  assign op_mapa8F_2_2_bufchan_r = (! op_mapa8F_2_2_bufchan_buf[0]);
  assign op_mapa8F_2_2_argbuf_d = (op_mapa8F_2_2_bufchan_buf[0] ? op_mapa8F_2_2_bufchan_buf :
                                   op_mapa8F_2_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) op_mapa8F_2_2_bufchan_buf <= 1'd0;
    else
      if ((op_mapa8F_2_2_argbuf_r && op_mapa8F_2_2_bufchan_buf[0]))
        op_mapa8F_2_2_bufchan_buf <= 1'd0;
      else if (((! op_mapa8F_2_2_argbuf_r) && (! op_mapa8F_2_2_bufchan_buf[0])))
        op_mapa8F_2_2_bufchan_buf <= op_mapa8F_2_2_bufchan_d;
  
  /* fork (Ty MyDTInt_Int) : (op_mapa8F_2_destruct,MyDTInt_Int) > [(op_mapa8F_2_1,MyDTInt_Int),
                                                              (op_mapa8F_2_2,MyDTInt_Int)] */
  logic [1:0] op_mapa8F_2_destruct_emitted;
  logic [1:0] op_mapa8F_2_destruct_done;
  assign op_mapa8F_2_1_d = (op_mapa8F_2_destruct_d[0] && (! op_mapa8F_2_destruct_emitted[0]));
  assign op_mapa8F_2_2_d = (op_mapa8F_2_destruct_d[0] && (! op_mapa8F_2_destruct_emitted[1]));
  assign op_mapa8F_2_destruct_done = (op_mapa8F_2_destruct_emitted | ({op_mapa8F_2_2_d[0],
                                                                       op_mapa8F_2_1_d[0]} & {op_mapa8F_2_2_r,
                                                                                              op_mapa8F_2_1_r}));
  assign op_mapa8F_2_destruct_r = (& op_mapa8F_2_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) op_mapa8F_2_destruct_emitted <= 2'd0;
    else
      op_mapa8F_2_destruct_emitted <= (op_mapa8F_2_destruct_r ? 2'd0 :
                                       op_mapa8F_2_destruct_done);
  
  /* buf (Ty MyDTInt_Int) : (op_mapa8F_3_2,MyDTInt_Int) > (op_mapa8F_3_2_argbuf,MyDTInt_Int) */
  MyDTInt_Int_t op_mapa8F_3_2_bufchan_d;
  logic op_mapa8F_3_2_bufchan_r;
  assign op_mapa8F_3_2_r = ((! op_mapa8F_3_2_bufchan_d[0]) || op_mapa8F_3_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) op_mapa8F_3_2_bufchan_d <= 1'd0;
    else
      if (op_mapa8F_3_2_r) op_mapa8F_3_2_bufchan_d <= op_mapa8F_3_2_d;
  MyDTInt_Int_t op_mapa8F_3_2_bufchan_buf;
  assign op_mapa8F_3_2_bufchan_r = (! op_mapa8F_3_2_bufchan_buf[0]);
  assign op_mapa8F_3_2_argbuf_d = (op_mapa8F_3_2_bufchan_buf[0] ? op_mapa8F_3_2_bufchan_buf :
                                   op_mapa8F_3_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) op_mapa8F_3_2_bufchan_buf <= 1'd0;
    else
      if ((op_mapa8F_3_2_argbuf_r && op_mapa8F_3_2_bufchan_buf[0]))
        op_mapa8F_3_2_bufchan_buf <= 1'd0;
      else if (((! op_mapa8F_3_2_argbuf_r) && (! op_mapa8F_3_2_bufchan_buf[0])))
        op_mapa8F_3_2_bufchan_buf <= op_mapa8F_3_2_bufchan_d;
  
  /* fork (Ty MyDTInt_Int) : (op_mapa8F_3_destruct,MyDTInt_Int) > [(op_mapa8F_3_1,MyDTInt_Int),
                                                              (op_mapa8F_3_2,MyDTInt_Int)] */
  logic [1:0] op_mapa8F_3_destruct_emitted;
  logic [1:0] op_mapa8F_3_destruct_done;
  assign op_mapa8F_3_1_d = (op_mapa8F_3_destruct_d[0] && (! op_mapa8F_3_destruct_emitted[0]));
  assign op_mapa8F_3_2_d = (op_mapa8F_3_destruct_d[0] && (! op_mapa8F_3_destruct_emitted[1]));
  assign op_mapa8F_3_destruct_done = (op_mapa8F_3_destruct_emitted | ({op_mapa8F_3_2_d[0],
                                                                       op_mapa8F_3_1_d[0]} & {op_mapa8F_3_2_r,
                                                                                              op_mapa8F_3_1_r}));
  assign op_mapa8F_3_destruct_r = (& op_mapa8F_3_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) op_mapa8F_3_destruct_emitted <= 2'd0;
    else
      op_mapa8F_3_destruct_emitted <= (op_mapa8F_3_destruct_r ? 2'd0 :
                                       op_mapa8F_3_destruct_done);
  
  /* buf (Ty MyDTInt_Int) : (op_mapa8F_4_destruct,MyDTInt_Int) > (op_mapa8F_4_1_argbuf,MyDTInt_Int) */
  MyDTInt_Int_t op_mapa8F_4_destruct_bufchan_d;
  logic op_mapa8F_4_destruct_bufchan_r;
  assign op_mapa8F_4_destruct_r = ((! op_mapa8F_4_destruct_bufchan_d[0]) || op_mapa8F_4_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) op_mapa8F_4_destruct_bufchan_d <= 1'd0;
    else
      if (op_mapa8F_4_destruct_r)
        op_mapa8F_4_destruct_bufchan_d <= op_mapa8F_4_destruct_d;
  MyDTInt_Int_t op_mapa8F_4_destruct_bufchan_buf;
  assign op_mapa8F_4_destruct_bufchan_r = (! op_mapa8F_4_destruct_bufchan_buf[0]);
  assign op_mapa8F_4_1_argbuf_d = (op_mapa8F_4_destruct_bufchan_buf[0] ? op_mapa8F_4_destruct_bufchan_buf :
                                   op_mapa8F_4_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) op_mapa8F_4_destruct_bufchan_buf <= 1'd0;
    else
      if ((op_mapa8F_4_1_argbuf_r && op_mapa8F_4_destruct_bufchan_buf[0]))
        op_mapa8F_4_destruct_bufchan_buf <= 1'd0;
      else if (((! op_mapa8F_4_1_argbuf_r) && (! op_mapa8F_4_destruct_bufchan_buf[0])))
        op_mapa8F_4_destruct_bufchan_buf <= op_mapa8F_4_destruct_bufchan_d;
  
  /* buf (Ty MyDTInt_Int) : (op_mapa8w_2_2,MyDTInt_Int) > (op_mapa8w_2_2_argbuf,MyDTInt_Int) */
  MyDTInt_Int_t op_mapa8w_2_2_bufchan_d;
  logic op_mapa8w_2_2_bufchan_r;
  assign op_mapa8w_2_2_r = ((! op_mapa8w_2_2_bufchan_d[0]) || op_mapa8w_2_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) op_mapa8w_2_2_bufchan_d <= 1'd0;
    else
      if (op_mapa8w_2_2_r) op_mapa8w_2_2_bufchan_d <= op_mapa8w_2_2_d;
  MyDTInt_Int_t op_mapa8w_2_2_bufchan_buf;
  assign op_mapa8w_2_2_bufchan_r = (! op_mapa8w_2_2_bufchan_buf[0]);
  assign op_mapa8w_2_2_argbuf_d = (op_mapa8w_2_2_bufchan_buf[0] ? op_mapa8w_2_2_bufchan_buf :
                                   op_mapa8w_2_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) op_mapa8w_2_2_bufchan_buf <= 1'd0;
    else
      if ((op_mapa8w_2_2_argbuf_r && op_mapa8w_2_2_bufchan_buf[0]))
        op_mapa8w_2_2_bufchan_buf <= 1'd0;
      else if (((! op_mapa8w_2_2_argbuf_r) && (! op_mapa8w_2_2_bufchan_buf[0])))
        op_mapa8w_2_2_bufchan_buf <= op_mapa8w_2_2_bufchan_d;
  
  /* fork (Ty MyDTInt_Int) : (op_mapa8w_2_destruct,MyDTInt_Int) > [(op_mapa8w_2_1,MyDTInt_Int),
                                                              (op_mapa8w_2_2,MyDTInt_Int)] */
  logic [1:0] op_mapa8w_2_destruct_emitted;
  logic [1:0] op_mapa8w_2_destruct_done;
  assign op_mapa8w_2_1_d = (op_mapa8w_2_destruct_d[0] && (! op_mapa8w_2_destruct_emitted[0]));
  assign op_mapa8w_2_2_d = (op_mapa8w_2_destruct_d[0] && (! op_mapa8w_2_destruct_emitted[1]));
  assign op_mapa8w_2_destruct_done = (op_mapa8w_2_destruct_emitted | ({op_mapa8w_2_2_d[0],
                                                                       op_mapa8w_2_1_d[0]} & {op_mapa8w_2_2_r,
                                                                                              op_mapa8w_2_1_r}));
  assign op_mapa8w_2_destruct_r = (& op_mapa8w_2_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) op_mapa8w_2_destruct_emitted <= 2'd0;
    else
      op_mapa8w_2_destruct_emitted <= (op_mapa8w_2_destruct_r ? 2'd0 :
                                       op_mapa8w_2_destruct_done);
  
  /* buf (Ty MyDTInt_Int) : (op_mapa8w_3_2,MyDTInt_Int) > (op_mapa8w_3_2_argbuf,MyDTInt_Int) */
  MyDTInt_Int_t op_mapa8w_3_2_bufchan_d;
  logic op_mapa8w_3_2_bufchan_r;
  assign op_mapa8w_3_2_r = ((! op_mapa8w_3_2_bufchan_d[0]) || op_mapa8w_3_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) op_mapa8w_3_2_bufchan_d <= 1'd0;
    else
      if (op_mapa8w_3_2_r) op_mapa8w_3_2_bufchan_d <= op_mapa8w_3_2_d;
  MyDTInt_Int_t op_mapa8w_3_2_bufchan_buf;
  assign op_mapa8w_3_2_bufchan_r = (! op_mapa8w_3_2_bufchan_buf[0]);
  assign op_mapa8w_3_2_argbuf_d = (op_mapa8w_3_2_bufchan_buf[0] ? op_mapa8w_3_2_bufchan_buf :
                                   op_mapa8w_3_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) op_mapa8w_3_2_bufchan_buf <= 1'd0;
    else
      if ((op_mapa8w_3_2_argbuf_r && op_mapa8w_3_2_bufchan_buf[0]))
        op_mapa8w_3_2_bufchan_buf <= 1'd0;
      else if (((! op_mapa8w_3_2_argbuf_r) && (! op_mapa8w_3_2_bufchan_buf[0])))
        op_mapa8w_3_2_bufchan_buf <= op_mapa8w_3_2_bufchan_d;
  
  /* fork (Ty MyDTInt_Int) : (op_mapa8w_3_destruct,MyDTInt_Int) > [(op_mapa8w_3_1,MyDTInt_Int),
                                                              (op_mapa8w_3_2,MyDTInt_Int)] */
  logic [1:0] op_mapa8w_3_destruct_emitted;
  logic [1:0] op_mapa8w_3_destruct_done;
  assign op_mapa8w_3_1_d = (op_mapa8w_3_destruct_d[0] && (! op_mapa8w_3_destruct_emitted[0]));
  assign op_mapa8w_3_2_d = (op_mapa8w_3_destruct_d[0] && (! op_mapa8w_3_destruct_emitted[1]));
  assign op_mapa8w_3_destruct_done = (op_mapa8w_3_destruct_emitted | ({op_mapa8w_3_2_d[0],
                                                                       op_mapa8w_3_1_d[0]} & {op_mapa8w_3_2_r,
                                                                                              op_mapa8w_3_1_r}));
  assign op_mapa8w_3_destruct_r = (& op_mapa8w_3_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) op_mapa8w_3_destruct_emitted <= 2'd0;
    else
      op_mapa8w_3_destruct_emitted <= (op_mapa8w_3_destruct_r ? 2'd0 :
                                       op_mapa8w_3_destruct_done);
  
  /* buf (Ty MyDTInt_Int) : (op_mapa8w_4_destruct,MyDTInt_Int) > (op_mapa8w_4_1_argbuf,MyDTInt_Int) */
  MyDTInt_Int_t op_mapa8w_4_destruct_bufchan_d;
  logic op_mapa8w_4_destruct_bufchan_r;
  assign op_mapa8w_4_destruct_r = ((! op_mapa8w_4_destruct_bufchan_d[0]) || op_mapa8w_4_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) op_mapa8w_4_destruct_bufchan_d <= 1'd0;
    else
      if (op_mapa8w_4_destruct_r)
        op_mapa8w_4_destruct_bufchan_d <= op_mapa8w_4_destruct_d;
  MyDTInt_Int_t op_mapa8w_4_destruct_bufchan_buf;
  assign op_mapa8w_4_destruct_bufchan_r = (! op_mapa8w_4_destruct_bufchan_buf[0]);
  assign op_mapa8w_4_1_argbuf_d = (op_mapa8w_4_destruct_bufchan_buf[0] ? op_mapa8w_4_destruct_bufchan_buf :
                                   op_mapa8w_4_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) op_mapa8w_4_destruct_bufchan_buf <= 1'd0;
    else
      if ((op_mapa8w_4_1_argbuf_r && op_mapa8w_4_destruct_bufchan_buf[0]))
        op_mapa8w_4_destruct_bufchan_buf <= 1'd0;
      else if (((! op_mapa8w_4_1_argbuf_r) && (! op_mapa8w_4_destruct_bufchan_buf[0])))
        op_mapa8w_4_destruct_bufchan_buf <= op_mapa8w_4_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (q1a84_destruct,Pointer_QTree_Int) > (q1a84_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t q1a84_destruct_bufchan_d;
  logic q1a84_destruct_bufchan_r;
  assign q1a84_destruct_r = ((! q1a84_destruct_bufchan_d[0]) || q1a84_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q1a84_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q1a84_destruct_r) q1a84_destruct_bufchan_d <= q1a84_destruct_d;
  Pointer_QTree_Int_t q1a84_destruct_bufchan_buf;
  assign q1a84_destruct_bufchan_r = (! q1a84_destruct_bufchan_buf[0]);
  assign q1a84_1_argbuf_d = (q1a84_destruct_bufchan_buf[0] ? q1a84_destruct_bufchan_buf :
                             q1a84_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q1a84_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q1a84_1_argbuf_r && q1a84_destruct_bufchan_buf[0]))
        q1a84_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q1a84_1_argbuf_r) && (! q1a84_destruct_bufchan_buf[0])))
        q1a84_destruct_bufchan_buf <= q1a84_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (q1a8T_3_destruct,Pointer_QTree_Int) > (q1a8T_3_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t q1a8T_3_destruct_bufchan_d;
  logic q1a8T_3_destruct_bufchan_r;
  assign q1a8T_3_destruct_r = ((! q1a8T_3_destruct_bufchan_d[0]) || q1a8T_3_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q1a8T_3_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q1a8T_3_destruct_r)
        q1a8T_3_destruct_bufchan_d <= q1a8T_3_destruct_d;
  Pointer_QTree_Int_t q1a8T_3_destruct_bufchan_buf;
  assign q1a8T_3_destruct_bufchan_r = (! q1a8T_3_destruct_bufchan_buf[0]);
  assign q1a8T_3_1_argbuf_d = (q1a8T_3_destruct_bufchan_buf[0] ? q1a8T_3_destruct_bufchan_buf :
                               q1a8T_3_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q1a8T_3_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q1a8T_3_1_argbuf_r && q1a8T_3_destruct_bufchan_buf[0]))
        q1a8T_3_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q1a8T_3_1_argbuf_r) && (! q1a8T_3_destruct_bufchan_buf[0])))
        q1a8T_3_destruct_bufchan_buf <= q1a8T_3_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (q2a85_1_destruct,Pointer_QTree_Int) > (q2a85_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t q2a85_1_destruct_bufchan_d;
  logic q2a85_1_destruct_bufchan_r;
  assign q2a85_1_destruct_r = ((! q2a85_1_destruct_bufchan_d[0]) || q2a85_1_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q2a85_1_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q2a85_1_destruct_r)
        q2a85_1_destruct_bufchan_d <= q2a85_1_destruct_d;
  Pointer_QTree_Int_t q2a85_1_destruct_bufchan_buf;
  assign q2a85_1_destruct_bufchan_r = (! q2a85_1_destruct_bufchan_buf[0]);
  assign q2a85_1_1_argbuf_d = (q2a85_1_destruct_bufchan_buf[0] ? q2a85_1_destruct_bufchan_buf :
                               q2a85_1_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q2a85_1_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q2a85_1_1_argbuf_r && q2a85_1_destruct_bufchan_buf[0]))
        q2a85_1_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q2a85_1_1_argbuf_r) && (! q2a85_1_destruct_bufchan_buf[0])))
        q2a85_1_destruct_bufchan_buf <= q2a85_1_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (q2a8U_2_destruct,Pointer_QTree_Int) > (q2a8U_2_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t q2a8U_2_destruct_bufchan_d;
  logic q2a8U_2_destruct_bufchan_r;
  assign q2a8U_2_destruct_r = ((! q2a8U_2_destruct_bufchan_d[0]) || q2a8U_2_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q2a8U_2_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q2a8U_2_destruct_r)
        q2a8U_2_destruct_bufchan_d <= q2a8U_2_destruct_d;
  Pointer_QTree_Int_t q2a8U_2_destruct_bufchan_buf;
  assign q2a8U_2_destruct_bufchan_r = (! q2a8U_2_destruct_bufchan_buf[0]);
  assign q2a8U_2_1_argbuf_d = (q2a8U_2_destruct_bufchan_buf[0] ? q2a8U_2_destruct_bufchan_buf :
                               q2a8U_2_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q2a8U_2_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q2a8U_2_1_argbuf_r && q2a8U_2_destruct_bufchan_buf[0]))
        q2a8U_2_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q2a8U_2_1_argbuf_r) && (! q2a8U_2_destruct_bufchan_buf[0])))
        q2a8U_2_destruct_bufchan_buf <= q2a8U_2_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (q3a86_2_destruct,Pointer_QTree_Int) > (q3a86_2_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t q3a86_2_destruct_bufchan_d;
  logic q3a86_2_destruct_bufchan_r;
  assign q3a86_2_destruct_r = ((! q3a86_2_destruct_bufchan_d[0]) || q3a86_2_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q3a86_2_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q3a86_2_destruct_r)
        q3a86_2_destruct_bufchan_d <= q3a86_2_destruct_d;
  Pointer_QTree_Int_t q3a86_2_destruct_bufchan_buf;
  assign q3a86_2_destruct_bufchan_r = (! q3a86_2_destruct_bufchan_buf[0]);
  assign q3a86_2_1_argbuf_d = (q3a86_2_destruct_bufchan_buf[0] ? q3a86_2_destruct_bufchan_buf :
                               q3a86_2_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q3a86_2_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q3a86_2_1_argbuf_r && q3a86_2_destruct_bufchan_buf[0]))
        q3a86_2_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q3a86_2_1_argbuf_r) && (! q3a86_2_destruct_bufchan_buf[0])))
        q3a86_2_destruct_bufchan_buf <= q3a86_2_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (q3a8V_1_destruct,Pointer_QTree_Int) > (q3a8V_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t q3a8V_1_destruct_bufchan_d;
  logic q3a8V_1_destruct_bufchan_r;
  assign q3a8V_1_destruct_r = ((! q3a8V_1_destruct_bufchan_d[0]) || q3a8V_1_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q3a8V_1_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q3a8V_1_destruct_r)
        q3a8V_1_destruct_bufchan_d <= q3a8V_1_destruct_d;
  Pointer_QTree_Int_t q3a8V_1_destruct_bufchan_buf;
  assign q3a8V_1_destruct_bufchan_r = (! q3a8V_1_destruct_bufchan_buf[0]);
  assign q3a8V_1_1_argbuf_d = (q3a8V_1_destruct_bufchan_buf[0] ? q3a8V_1_destruct_bufchan_buf :
                               q3a8V_1_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q3a8V_1_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q3a8V_1_1_argbuf_r && q3a8V_1_destruct_bufchan_buf[0]))
        q3a8V_1_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q3a8V_1_1_argbuf_r) && (! q3a8V_1_destruct_bufchan_buf[0])))
        q3a8V_1_destruct_bufchan_buf <= q3a8V_1_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (q4a87_3_destruct,Pointer_QTree_Int) > (q4a87_3_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t q4a87_3_destruct_bufchan_d;
  logic q4a87_3_destruct_bufchan_r;
  assign q4a87_3_destruct_r = ((! q4a87_3_destruct_bufchan_d[0]) || q4a87_3_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q4a87_3_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q4a87_3_destruct_r)
        q4a87_3_destruct_bufchan_d <= q4a87_3_destruct_d;
  Pointer_QTree_Int_t q4a87_3_destruct_bufchan_buf;
  assign q4a87_3_destruct_bufchan_r = (! q4a87_3_destruct_bufchan_buf[0]);
  assign q4a87_3_1_argbuf_d = (q4a87_3_destruct_bufchan_buf[0] ? q4a87_3_destruct_bufchan_buf :
                               q4a87_3_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q4a87_3_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q4a87_3_1_argbuf_r && q4a87_3_destruct_bufchan_buf[0]))
        q4a87_3_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q4a87_3_1_argbuf_r) && (! q4a87_3_destruct_bufchan_buf[0])))
        q4a87_3_destruct_bufchan_buf <= q4a87_3_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (q4a8u_goMux_mux,Pointer_QTree_Int) > (q4a8u_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t q4a8u_goMux_mux_bufchan_d;
  logic q4a8u_goMux_mux_bufchan_r;
  assign q4a8u_goMux_mux_r = ((! q4a8u_goMux_mux_bufchan_d[0]) || q4a8u_goMux_mux_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q4a8u_goMux_mux_bufchan_d <= {16'd0, 1'd0};
    else
      if (q4a8u_goMux_mux_r)
        q4a8u_goMux_mux_bufchan_d <= q4a8u_goMux_mux_d;
  Pointer_QTree_Int_t q4a8u_goMux_mux_bufchan_buf;
  assign q4a8u_goMux_mux_bufchan_r = (! q4a8u_goMux_mux_bufchan_buf[0]);
  assign q4a8u_1_argbuf_d = (q4a8u_goMux_mux_bufchan_buf[0] ? q4a8u_goMux_mux_bufchan_buf :
                             q4a8u_goMux_mux_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q4a8u_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q4a8u_1_argbuf_r && q4a8u_goMux_mux_bufchan_buf[0]))
        q4a8u_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q4a8u_1_argbuf_r) && (! q4a8u_goMux_mux_bufchan_buf[0])))
        q4a8u_goMux_mux_bufchan_buf <= q4a8u_goMux_mux_bufchan_d;
  
  /* buf (Ty CT$wnnz) : (readPointer_CT$wnnzscfarg_0_1_argbuf,CT$wnnz) > (readPointer_CT$wnnzscfarg_0_1_argbuf_rwb,CT$wnnz) */
  CT$wnnz_t readPointer_CT$wnnzscfarg_0_1_argbuf_bufchan_d;
  logic readPointer_CT$wnnzscfarg_0_1_argbuf_bufchan_r;
  assign readPointer_CT$wnnzscfarg_0_1_argbuf_r = ((! readPointer_CT$wnnzscfarg_0_1_argbuf_bufchan_d[0]) || readPointer_CT$wnnzscfarg_0_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_CT$wnnzscfarg_0_1_argbuf_bufchan_d <= {115'd0, 1'd0};
    else
      if (readPointer_CT$wnnzscfarg_0_1_argbuf_r)
        readPointer_CT$wnnzscfarg_0_1_argbuf_bufchan_d <= readPointer_CT$wnnzscfarg_0_1_argbuf_d;
  CT$wnnz_t readPointer_CT$wnnzscfarg_0_1_argbuf_bufchan_buf;
  assign readPointer_CT$wnnzscfarg_0_1_argbuf_bufchan_r = (! readPointer_CT$wnnzscfarg_0_1_argbuf_bufchan_buf[0]);
  assign readPointer_CT$wnnzscfarg_0_1_argbuf_rwb_d = (readPointer_CT$wnnzscfarg_0_1_argbuf_bufchan_buf[0] ? readPointer_CT$wnnzscfarg_0_1_argbuf_bufchan_buf :
                                                       readPointer_CT$wnnzscfarg_0_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_CT$wnnzscfarg_0_1_argbuf_bufchan_buf <= {115'd0, 1'd0};
    else
      if ((readPointer_CT$wnnzscfarg_0_1_argbuf_rwb_r && readPointer_CT$wnnzscfarg_0_1_argbuf_bufchan_buf[0]))
        readPointer_CT$wnnzscfarg_0_1_argbuf_bufchan_buf <= {115'd0, 1'd0};
      else if (((! readPointer_CT$wnnzscfarg_0_1_argbuf_rwb_r) && (! readPointer_CT$wnnzscfarg_0_1_argbuf_bufchan_buf[0])))
        readPointer_CT$wnnzscfarg_0_1_argbuf_bufchan_buf <= readPointer_CT$wnnzscfarg_0_1_argbuf_bufchan_d;
  
  /* fork (Ty CT$wnnz) : (readPointer_CT$wnnzscfarg_0_1_argbuf_rwb,CT$wnnz) > [(lizzieLet35_1,CT$wnnz),
                                                                          (lizzieLet35_2,CT$wnnz),
                                                                          (lizzieLet35_3,CT$wnnz),
                                                                          (lizzieLet35_4,CT$wnnz)] */
  logic [3:0] readPointer_CT$wnnzscfarg_0_1_argbuf_rwb_emitted;
  logic [3:0] readPointer_CT$wnnzscfarg_0_1_argbuf_rwb_done;
  assign lizzieLet35_1_d = {readPointer_CT$wnnzscfarg_0_1_argbuf_rwb_d[115:1],
                            (readPointer_CT$wnnzscfarg_0_1_argbuf_rwb_d[0] && (! readPointer_CT$wnnzscfarg_0_1_argbuf_rwb_emitted[0]))};
  assign lizzieLet35_2_d = {readPointer_CT$wnnzscfarg_0_1_argbuf_rwb_d[115:1],
                            (readPointer_CT$wnnzscfarg_0_1_argbuf_rwb_d[0] && (! readPointer_CT$wnnzscfarg_0_1_argbuf_rwb_emitted[1]))};
  assign lizzieLet35_3_d = {readPointer_CT$wnnzscfarg_0_1_argbuf_rwb_d[115:1],
                            (readPointer_CT$wnnzscfarg_0_1_argbuf_rwb_d[0] && (! readPointer_CT$wnnzscfarg_0_1_argbuf_rwb_emitted[2]))};
  assign lizzieLet35_4_d = {readPointer_CT$wnnzscfarg_0_1_argbuf_rwb_d[115:1],
                            (readPointer_CT$wnnzscfarg_0_1_argbuf_rwb_d[0] && (! readPointer_CT$wnnzscfarg_0_1_argbuf_rwb_emitted[3]))};
  assign readPointer_CT$wnnzscfarg_0_1_argbuf_rwb_done = (readPointer_CT$wnnzscfarg_0_1_argbuf_rwb_emitted | ({lizzieLet35_4_d[0],
                                                                                                               lizzieLet35_3_d[0],
                                                                                                               lizzieLet35_2_d[0],
                                                                                                               lizzieLet35_1_d[0]} & {lizzieLet35_4_r,
                                                                                                                                      lizzieLet35_3_r,
                                                                                                                                      lizzieLet35_2_r,
                                                                                                                                      lizzieLet35_1_r}));
  assign readPointer_CT$wnnzscfarg_0_1_argbuf_rwb_r = (& readPointer_CT$wnnzscfarg_0_1_argbuf_rwb_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_CT$wnnzscfarg_0_1_argbuf_rwb_emitted <= 4'd0;
    else
      readPointer_CT$wnnzscfarg_0_1_argbuf_rwb_emitted <= (readPointer_CT$wnnzscfarg_0_1_argbuf_rwb_r ? 4'd0 :
                                                           readPointer_CT$wnnzscfarg_0_1_argbuf_rwb_done);
  
  /* buf (Ty CTf''''''''_f''''''''_Int_Int) : (readPointer_CTf''''''''_f''''''''_Int_Intscfarg_0_1_1_argbuf,CTf''''''''_f''''''''_Int_Int) > (readPointer_CTf''''''''_f''''''''_Int_Intscfarg_0_1_1_argbuf_rwb,CTf''''''''_f''''''''_Int_Int) */
  \CTf''''''''_f''''''''_Int_Int_t  \readPointer_CTf''''''''_f''''''''_Int_Intscfarg_0_1_1_argbuf_bufchan_d ;
  logic \readPointer_CTf''''''''_f''''''''_Int_Intscfarg_0_1_1_argbuf_bufchan_r ;
  assign \readPointer_CTf''''''''_f''''''''_Int_Intscfarg_0_1_1_argbuf_r  = ((! \readPointer_CTf''''''''_f''''''''_Int_Intscfarg_0_1_1_argbuf_bufchan_d [0]) || \readPointer_CTf''''''''_f''''''''_Int_Intscfarg_0_1_1_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \readPointer_CTf''''''''_f''''''''_Int_Intscfarg_0_1_1_argbuf_bufchan_d  <= {67'd0,
                                                                                   1'd0};
    else
      if (\readPointer_CTf''''''''_f''''''''_Int_Intscfarg_0_1_1_argbuf_r )
        \readPointer_CTf''''''''_f''''''''_Int_Intscfarg_0_1_1_argbuf_bufchan_d  <= \readPointer_CTf''''''''_f''''''''_Int_Intscfarg_0_1_1_argbuf_d ;
  \CTf''''''''_f''''''''_Int_Int_t  \readPointer_CTf''''''''_f''''''''_Int_Intscfarg_0_1_1_argbuf_bufchan_buf ;
  assign \readPointer_CTf''''''''_f''''''''_Int_Intscfarg_0_1_1_argbuf_bufchan_r  = (! \readPointer_CTf''''''''_f''''''''_Int_Intscfarg_0_1_1_argbuf_bufchan_buf [0]);
  assign \readPointer_CTf''''''''_f''''''''_Int_Intscfarg_0_1_1_argbuf_rwb_d  = (\readPointer_CTf''''''''_f''''''''_Int_Intscfarg_0_1_1_argbuf_bufchan_buf [0] ? \readPointer_CTf''''''''_f''''''''_Int_Intscfarg_0_1_1_argbuf_bufchan_buf  :
                                                                                 \readPointer_CTf''''''''_f''''''''_Int_Intscfarg_0_1_1_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \readPointer_CTf''''''''_f''''''''_Int_Intscfarg_0_1_1_argbuf_bufchan_buf  <= {67'd0,
                                                                                     1'd0};
    else
      if ((\readPointer_CTf''''''''_f''''''''_Int_Intscfarg_0_1_1_argbuf_rwb_r  && \readPointer_CTf''''''''_f''''''''_Int_Intscfarg_0_1_1_argbuf_bufchan_buf [0]))
        \readPointer_CTf''''''''_f''''''''_Int_Intscfarg_0_1_1_argbuf_bufchan_buf  <= {67'd0,
                                                                                       1'd0};
      else if (((! \readPointer_CTf''''''''_f''''''''_Int_Intscfarg_0_1_1_argbuf_rwb_r ) && (! \readPointer_CTf''''''''_f''''''''_Int_Intscfarg_0_1_1_argbuf_bufchan_buf [0])))
        \readPointer_CTf''''''''_f''''''''_Int_Intscfarg_0_1_1_argbuf_bufchan_buf  <= \readPointer_CTf''''''''_f''''''''_Int_Intscfarg_0_1_1_argbuf_bufchan_d ;
  
  /* fork (Ty CTf''''''''_f''''''''_Int_Int) : (readPointer_CTf''''''''_f''''''''_Int_Intscfarg_0_1_1_argbuf_rwb,CTf''''''''_f''''''''_Int_Int) > [(lizzieLet39_1,CTf''''''''_f''''''''_Int_Int),
                                                                                                                                              (lizzieLet39_2,CTf''''''''_f''''''''_Int_Int),
                                                                                                                                              (lizzieLet39_3,CTf''''''''_f''''''''_Int_Int),
                                                                                                                                              (lizzieLet39_4,CTf''''''''_f''''''''_Int_Int)] */
  logic [3:0] \readPointer_CTf''''''''_f''''''''_Int_Intscfarg_0_1_1_argbuf_rwb_emitted ;
  logic [3:0] \readPointer_CTf''''''''_f''''''''_Int_Intscfarg_0_1_1_argbuf_rwb_done ;
  assign lizzieLet39_1_d = {\readPointer_CTf''''''''_f''''''''_Int_Intscfarg_0_1_1_argbuf_rwb_d [67:1],
                            (\readPointer_CTf''''''''_f''''''''_Int_Intscfarg_0_1_1_argbuf_rwb_d [0] && (! \readPointer_CTf''''''''_f''''''''_Int_Intscfarg_0_1_1_argbuf_rwb_emitted [0]))};
  assign lizzieLet39_2_d = {\readPointer_CTf''''''''_f''''''''_Int_Intscfarg_0_1_1_argbuf_rwb_d [67:1],
                            (\readPointer_CTf''''''''_f''''''''_Int_Intscfarg_0_1_1_argbuf_rwb_d [0] && (! \readPointer_CTf''''''''_f''''''''_Int_Intscfarg_0_1_1_argbuf_rwb_emitted [1]))};
  assign lizzieLet39_3_d = {\readPointer_CTf''''''''_f''''''''_Int_Intscfarg_0_1_1_argbuf_rwb_d [67:1],
                            (\readPointer_CTf''''''''_f''''''''_Int_Intscfarg_0_1_1_argbuf_rwb_d [0] && (! \readPointer_CTf''''''''_f''''''''_Int_Intscfarg_0_1_1_argbuf_rwb_emitted [2]))};
  assign lizzieLet39_4_d = {\readPointer_CTf''''''''_f''''''''_Int_Intscfarg_0_1_1_argbuf_rwb_d [67:1],
                            (\readPointer_CTf''''''''_f''''''''_Int_Intscfarg_0_1_1_argbuf_rwb_d [0] && (! \readPointer_CTf''''''''_f''''''''_Int_Intscfarg_0_1_1_argbuf_rwb_emitted [3]))};
  assign \readPointer_CTf''''''''_f''''''''_Int_Intscfarg_0_1_1_argbuf_rwb_done  = (\readPointer_CTf''''''''_f''''''''_Int_Intscfarg_0_1_1_argbuf_rwb_emitted  | ({lizzieLet39_4_d[0],
                                                                                                                                                                   lizzieLet39_3_d[0],
                                                                                                                                                                   lizzieLet39_2_d[0],
                                                                                                                                                                   lizzieLet39_1_d[0]} & {lizzieLet39_4_r,
                                                                                                                                                                                          lizzieLet39_3_r,
                                                                                                                                                                                          lizzieLet39_2_r,
                                                                                                                                                                                          lizzieLet39_1_r}));
  assign \readPointer_CTf''''''''_f''''''''_Int_Intscfarg_0_1_1_argbuf_rwb_r  = (& \readPointer_CTf''''''''_f''''''''_Int_Intscfarg_0_1_1_argbuf_rwb_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \readPointer_CTf''''''''_f''''''''_Int_Intscfarg_0_1_1_argbuf_rwb_emitted  <= 4'd0;
    else
      \readPointer_CTf''''''''_f''''''''_Int_Intscfarg_0_1_1_argbuf_rwb_emitted  <= (\readPointer_CTf''''''''_f''''''''_Int_Intscfarg_0_1_1_argbuf_rwb_r  ? 4'd0 :
                                                                                     \readPointer_CTf''''''''_f''''''''_Int_Intscfarg_0_1_1_argbuf_rwb_done );
  
  /* buf (Ty CTf_f_Int_Int) : (readPointer_CTf_f_Int_Intscfarg_0_2_1_argbuf,CTf_f_Int_Int) > (readPointer_CTf_f_Int_Intscfarg_0_2_1_argbuf_rwb,CTf_f_Int_Int) */
  CTf_f_Int_Int_t readPointer_CTf_f_Int_Intscfarg_0_2_1_argbuf_bufchan_d;
  logic readPointer_CTf_f_Int_Intscfarg_0_2_1_argbuf_bufchan_r;
  assign readPointer_CTf_f_Int_Intscfarg_0_2_1_argbuf_r = ((! readPointer_CTf_f_Int_Intscfarg_0_2_1_argbuf_bufchan_d[0]) || readPointer_CTf_f_Int_Intscfarg_0_2_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_CTf_f_Int_Intscfarg_0_2_1_argbuf_bufchan_d <= {115'd0,
                                                                 1'd0};
    else
      if (readPointer_CTf_f_Int_Intscfarg_0_2_1_argbuf_r)
        readPointer_CTf_f_Int_Intscfarg_0_2_1_argbuf_bufchan_d <= readPointer_CTf_f_Int_Intscfarg_0_2_1_argbuf_d;
  CTf_f_Int_Int_t readPointer_CTf_f_Int_Intscfarg_0_2_1_argbuf_bufchan_buf;
  assign readPointer_CTf_f_Int_Intscfarg_0_2_1_argbuf_bufchan_r = (! readPointer_CTf_f_Int_Intscfarg_0_2_1_argbuf_bufchan_buf[0]);
  assign readPointer_CTf_f_Int_Intscfarg_0_2_1_argbuf_rwb_d = (readPointer_CTf_f_Int_Intscfarg_0_2_1_argbuf_bufchan_buf[0] ? readPointer_CTf_f_Int_Intscfarg_0_2_1_argbuf_bufchan_buf :
                                                               readPointer_CTf_f_Int_Intscfarg_0_2_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_CTf_f_Int_Intscfarg_0_2_1_argbuf_bufchan_buf <= {115'd0,
                                                                   1'd0};
    else
      if ((readPointer_CTf_f_Int_Intscfarg_0_2_1_argbuf_rwb_r && readPointer_CTf_f_Int_Intscfarg_0_2_1_argbuf_bufchan_buf[0]))
        readPointer_CTf_f_Int_Intscfarg_0_2_1_argbuf_bufchan_buf <= {115'd0,
                                                                     1'd0};
      else if (((! readPointer_CTf_f_Int_Intscfarg_0_2_1_argbuf_rwb_r) && (! readPointer_CTf_f_Int_Intscfarg_0_2_1_argbuf_bufchan_buf[0])))
        readPointer_CTf_f_Int_Intscfarg_0_2_1_argbuf_bufchan_buf <= readPointer_CTf_f_Int_Intscfarg_0_2_1_argbuf_bufchan_d;
  
  /* fork (Ty CTf_f_Int_Int) : (readPointer_CTf_f_Int_Intscfarg_0_2_1_argbuf_rwb,CTf_f_Int_Int) > [(lizzieLet44_1,CTf_f_Int_Int),
                                                                                              (lizzieLet44_2,CTf_f_Int_Int),
                                                                                              (lizzieLet44_3,CTf_f_Int_Int),
                                                                                              (lizzieLet44_4,CTf_f_Int_Int)] */
  logic [3:0] readPointer_CTf_f_Int_Intscfarg_0_2_1_argbuf_rwb_emitted;
  logic [3:0] readPointer_CTf_f_Int_Intscfarg_0_2_1_argbuf_rwb_done;
  assign lizzieLet44_1_d = {readPointer_CTf_f_Int_Intscfarg_0_2_1_argbuf_rwb_d[115:1],
                            (readPointer_CTf_f_Int_Intscfarg_0_2_1_argbuf_rwb_d[0] && (! readPointer_CTf_f_Int_Intscfarg_0_2_1_argbuf_rwb_emitted[0]))};
  assign lizzieLet44_2_d = {readPointer_CTf_f_Int_Intscfarg_0_2_1_argbuf_rwb_d[115:1],
                            (readPointer_CTf_f_Int_Intscfarg_0_2_1_argbuf_rwb_d[0] && (! readPointer_CTf_f_Int_Intscfarg_0_2_1_argbuf_rwb_emitted[1]))};
  assign lizzieLet44_3_d = {readPointer_CTf_f_Int_Intscfarg_0_2_1_argbuf_rwb_d[115:1],
                            (readPointer_CTf_f_Int_Intscfarg_0_2_1_argbuf_rwb_d[0] && (! readPointer_CTf_f_Int_Intscfarg_0_2_1_argbuf_rwb_emitted[2]))};
  assign lizzieLet44_4_d = {readPointer_CTf_f_Int_Intscfarg_0_2_1_argbuf_rwb_d[115:1],
                            (readPointer_CTf_f_Int_Intscfarg_0_2_1_argbuf_rwb_d[0] && (! readPointer_CTf_f_Int_Intscfarg_0_2_1_argbuf_rwb_emitted[3]))};
  assign readPointer_CTf_f_Int_Intscfarg_0_2_1_argbuf_rwb_done = (readPointer_CTf_f_Int_Intscfarg_0_2_1_argbuf_rwb_emitted | ({lizzieLet44_4_d[0],
                                                                                                                               lizzieLet44_3_d[0],
                                                                                                                               lizzieLet44_2_d[0],
                                                                                                                               lizzieLet44_1_d[0]} & {lizzieLet44_4_r,
                                                                                                                                                      lizzieLet44_3_r,
                                                                                                                                                      lizzieLet44_2_r,
                                                                                                                                                      lizzieLet44_1_r}));
  assign readPointer_CTf_f_Int_Intscfarg_0_2_1_argbuf_rwb_r = (& readPointer_CTf_f_Int_Intscfarg_0_2_1_argbuf_rwb_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_CTf_f_Int_Intscfarg_0_2_1_argbuf_rwb_emitted <= 4'd0;
    else
      readPointer_CTf_f_Int_Intscfarg_0_2_1_argbuf_rwb_emitted <= (readPointer_CTf_f_Int_Intscfarg_0_2_1_argbuf_rwb_r ? 4'd0 :
                                                                   readPointer_CTf_f_Int_Intscfarg_0_2_1_argbuf_rwb_done);
  
  /* buf (Ty QTree_Int) : (readPointer_QTree_Intm1a8C_1_argbuf,QTree_Int) > (readPointer_QTree_Intm1a8C_1_argbuf_rwb,QTree_Int) */
  QTree_Int_t readPointer_QTree_Intm1a8C_1_argbuf_bufchan_d;
  logic readPointer_QTree_Intm1a8C_1_argbuf_bufchan_r;
  assign readPointer_QTree_Intm1a8C_1_argbuf_r = ((! readPointer_QTree_Intm1a8C_1_argbuf_bufchan_d[0]) || readPointer_QTree_Intm1a8C_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Intm1a8C_1_argbuf_bufchan_d <= {66'd0, 1'd0};
    else
      if (readPointer_QTree_Intm1a8C_1_argbuf_r)
        readPointer_QTree_Intm1a8C_1_argbuf_bufchan_d <= readPointer_QTree_Intm1a8C_1_argbuf_d;
  QTree_Int_t readPointer_QTree_Intm1a8C_1_argbuf_bufchan_buf;
  assign readPointer_QTree_Intm1a8C_1_argbuf_bufchan_r = (! readPointer_QTree_Intm1a8C_1_argbuf_bufchan_buf[0]);
  assign readPointer_QTree_Intm1a8C_1_argbuf_rwb_d = (readPointer_QTree_Intm1a8C_1_argbuf_bufchan_buf[0] ? readPointer_QTree_Intm1a8C_1_argbuf_bufchan_buf :
                                                      readPointer_QTree_Intm1a8C_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Intm1a8C_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((readPointer_QTree_Intm1a8C_1_argbuf_rwb_r && readPointer_QTree_Intm1a8C_1_argbuf_bufchan_buf[0]))
        readPointer_QTree_Intm1a8C_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
      else if (((! readPointer_QTree_Intm1a8C_1_argbuf_rwb_r) && (! readPointer_QTree_Intm1a8C_1_argbuf_bufchan_buf[0])))
        readPointer_QTree_Intm1a8C_1_argbuf_bufchan_buf <= readPointer_QTree_Intm1a8C_1_argbuf_bufchan_d;
  
  /* fork (Ty QTree_Int) : (readPointer_QTree_Intm1a8C_1_argbuf_rwb,QTree_Int) > [(lizzieLet12_1,QTree_Int),
                                                                             (lizzieLet12_2,QTree_Int),
                                                                             (lizzieLet12_3,QTree_Int),
                                                                             (lizzieLet12_4,QTree_Int),
                                                                             (lizzieLet12_5,QTree_Int),
                                                                             (lizzieLet12_6,QTree_Int),
                                                                             (lizzieLet12_7,QTree_Int),
                                                                             (lizzieLet12_8,QTree_Int),
                                                                             (lizzieLet12_9,QTree_Int)] */
  logic [8:0] readPointer_QTree_Intm1a8C_1_argbuf_rwb_emitted;
  logic [8:0] readPointer_QTree_Intm1a8C_1_argbuf_rwb_done;
  assign lizzieLet12_1_d = {readPointer_QTree_Intm1a8C_1_argbuf_rwb_d[66:1],
                            (readPointer_QTree_Intm1a8C_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intm1a8C_1_argbuf_rwb_emitted[0]))};
  assign lizzieLet12_2_d = {readPointer_QTree_Intm1a8C_1_argbuf_rwb_d[66:1],
                            (readPointer_QTree_Intm1a8C_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intm1a8C_1_argbuf_rwb_emitted[1]))};
  assign lizzieLet12_3_d = {readPointer_QTree_Intm1a8C_1_argbuf_rwb_d[66:1],
                            (readPointer_QTree_Intm1a8C_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intm1a8C_1_argbuf_rwb_emitted[2]))};
  assign lizzieLet12_4_d = {readPointer_QTree_Intm1a8C_1_argbuf_rwb_d[66:1],
                            (readPointer_QTree_Intm1a8C_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intm1a8C_1_argbuf_rwb_emitted[3]))};
  assign lizzieLet12_5_d = {readPointer_QTree_Intm1a8C_1_argbuf_rwb_d[66:1],
                            (readPointer_QTree_Intm1a8C_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intm1a8C_1_argbuf_rwb_emitted[4]))};
  assign lizzieLet12_6_d = {readPointer_QTree_Intm1a8C_1_argbuf_rwb_d[66:1],
                            (readPointer_QTree_Intm1a8C_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intm1a8C_1_argbuf_rwb_emitted[5]))};
  assign lizzieLet12_7_d = {readPointer_QTree_Intm1a8C_1_argbuf_rwb_d[66:1],
                            (readPointer_QTree_Intm1a8C_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intm1a8C_1_argbuf_rwb_emitted[6]))};
  assign lizzieLet12_8_d = {readPointer_QTree_Intm1a8C_1_argbuf_rwb_d[66:1],
                            (readPointer_QTree_Intm1a8C_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intm1a8C_1_argbuf_rwb_emitted[7]))};
  assign lizzieLet12_9_d = {readPointer_QTree_Intm1a8C_1_argbuf_rwb_d[66:1],
                            (readPointer_QTree_Intm1a8C_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intm1a8C_1_argbuf_rwb_emitted[8]))};
  assign readPointer_QTree_Intm1a8C_1_argbuf_rwb_done = (readPointer_QTree_Intm1a8C_1_argbuf_rwb_emitted | ({lizzieLet12_9_d[0],
                                                                                                             lizzieLet12_8_d[0],
                                                                                                             lizzieLet12_7_d[0],
                                                                                                             lizzieLet12_6_d[0],
                                                                                                             lizzieLet12_5_d[0],
                                                                                                             lizzieLet12_4_d[0],
                                                                                                             lizzieLet12_3_d[0],
                                                                                                             lizzieLet12_2_d[0],
                                                                                                             lizzieLet12_1_d[0]} & {lizzieLet12_9_r,
                                                                                                                                    lizzieLet12_8_r,
                                                                                                                                    lizzieLet12_7_r,
                                                                                                                                    lizzieLet12_6_r,
                                                                                                                                    lizzieLet12_5_r,
                                                                                                                                    lizzieLet12_4_r,
                                                                                                                                    lizzieLet12_3_r,
                                                                                                                                    lizzieLet12_2_r,
                                                                                                                                    lizzieLet12_1_r}));
  assign readPointer_QTree_Intm1a8C_1_argbuf_rwb_r = (& readPointer_QTree_Intm1a8C_1_argbuf_rwb_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Intm1a8C_1_argbuf_rwb_emitted <= 9'd0;
    else
      readPointer_QTree_Intm1a8C_1_argbuf_rwb_emitted <= (readPointer_QTree_Intm1a8C_1_argbuf_rwb_r ? 9'd0 :
                                                          readPointer_QTree_Intm1a8C_1_argbuf_rwb_done);
  
  /* buf (Ty QTree_Int) : (readPointer_QTree_Intm2a8D_1_argbuf,QTree_Int) > (readPointer_QTree_Intm2a8D_1_argbuf_rwb,QTree_Int) */
  QTree_Int_t readPointer_QTree_Intm2a8D_1_argbuf_bufchan_d;
  logic readPointer_QTree_Intm2a8D_1_argbuf_bufchan_r;
  assign readPointer_QTree_Intm2a8D_1_argbuf_r = ((! readPointer_QTree_Intm2a8D_1_argbuf_bufchan_d[0]) || readPointer_QTree_Intm2a8D_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Intm2a8D_1_argbuf_bufchan_d <= {66'd0, 1'd0};
    else
      if (readPointer_QTree_Intm2a8D_1_argbuf_r)
        readPointer_QTree_Intm2a8D_1_argbuf_bufchan_d <= readPointer_QTree_Intm2a8D_1_argbuf_d;
  QTree_Int_t readPointer_QTree_Intm2a8D_1_argbuf_bufchan_buf;
  assign readPointer_QTree_Intm2a8D_1_argbuf_bufchan_r = (! readPointer_QTree_Intm2a8D_1_argbuf_bufchan_buf[0]);
  assign readPointer_QTree_Intm2a8D_1_argbuf_rwb_d = (readPointer_QTree_Intm2a8D_1_argbuf_bufchan_buf[0] ? readPointer_QTree_Intm2a8D_1_argbuf_bufchan_buf :
                                                      readPointer_QTree_Intm2a8D_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Intm2a8D_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((readPointer_QTree_Intm2a8D_1_argbuf_rwb_r && readPointer_QTree_Intm2a8D_1_argbuf_bufchan_buf[0]))
        readPointer_QTree_Intm2a8D_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
      else if (((! readPointer_QTree_Intm2a8D_1_argbuf_rwb_r) && (! readPointer_QTree_Intm2a8D_1_argbuf_bufchan_buf[0])))
        readPointer_QTree_Intm2a8D_1_argbuf_bufchan_buf <= readPointer_QTree_Intm2a8D_1_argbuf_bufchan_d;
  
  /* buf (Ty QTree_Int) : (readPointer_QTree_Intq4a8u_1_argbuf,QTree_Int) > (readPointer_QTree_Intq4a8u_1_argbuf_rwb,QTree_Int) */
  QTree_Int_t readPointer_QTree_Intq4a8u_1_argbuf_bufchan_d;
  logic readPointer_QTree_Intq4a8u_1_argbuf_bufchan_r;
  assign readPointer_QTree_Intq4a8u_1_argbuf_r = ((! readPointer_QTree_Intq4a8u_1_argbuf_bufchan_d[0]) || readPointer_QTree_Intq4a8u_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Intq4a8u_1_argbuf_bufchan_d <= {66'd0, 1'd0};
    else
      if (readPointer_QTree_Intq4a8u_1_argbuf_r)
        readPointer_QTree_Intq4a8u_1_argbuf_bufchan_d <= readPointer_QTree_Intq4a8u_1_argbuf_d;
  QTree_Int_t readPointer_QTree_Intq4a8u_1_argbuf_bufchan_buf;
  assign readPointer_QTree_Intq4a8u_1_argbuf_bufchan_r = (! readPointer_QTree_Intq4a8u_1_argbuf_bufchan_buf[0]);
  assign readPointer_QTree_Intq4a8u_1_argbuf_rwb_d = (readPointer_QTree_Intq4a8u_1_argbuf_bufchan_buf[0] ? readPointer_QTree_Intq4a8u_1_argbuf_bufchan_buf :
                                                      readPointer_QTree_Intq4a8u_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Intq4a8u_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((readPointer_QTree_Intq4a8u_1_argbuf_rwb_r && readPointer_QTree_Intq4a8u_1_argbuf_bufchan_buf[0]))
        readPointer_QTree_Intq4a8u_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
      else if (((! readPointer_QTree_Intq4a8u_1_argbuf_rwb_r) && (! readPointer_QTree_Intq4a8u_1_argbuf_bufchan_buf[0])))
        readPointer_QTree_Intq4a8u_1_argbuf_bufchan_buf <= readPointer_QTree_Intq4a8u_1_argbuf_bufchan_d;
  
  /* fork (Ty QTree_Int) : (readPointer_QTree_Intq4a8u_1_argbuf_rwb,QTree_Int) > [(lizzieLet6_1,QTree_Int),
                                                                             (lizzieLet6_2,QTree_Int),
                                                                             (lizzieLet6_3,QTree_Int),
                                                                             (lizzieLet6_4,QTree_Int),
                                                                             (lizzieLet6_5,QTree_Int),
                                                                             (lizzieLet6_6,QTree_Int)] */
  logic [5:0] readPointer_QTree_Intq4a8u_1_argbuf_rwb_emitted;
  logic [5:0] readPointer_QTree_Intq4a8u_1_argbuf_rwb_done;
  assign lizzieLet6_1_d = {readPointer_QTree_Intq4a8u_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_Intq4a8u_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intq4a8u_1_argbuf_rwb_emitted[0]))};
  assign lizzieLet6_2_d = {readPointer_QTree_Intq4a8u_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_Intq4a8u_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intq4a8u_1_argbuf_rwb_emitted[1]))};
  assign lizzieLet6_3_d = {readPointer_QTree_Intq4a8u_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_Intq4a8u_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intq4a8u_1_argbuf_rwb_emitted[2]))};
  assign lizzieLet6_4_d = {readPointer_QTree_Intq4a8u_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_Intq4a8u_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intq4a8u_1_argbuf_rwb_emitted[3]))};
  assign lizzieLet6_5_d = {readPointer_QTree_Intq4a8u_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_Intq4a8u_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intq4a8u_1_argbuf_rwb_emitted[4]))};
  assign lizzieLet6_6_d = {readPointer_QTree_Intq4a8u_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_Intq4a8u_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intq4a8u_1_argbuf_rwb_emitted[5]))};
  assign readPointer_QTree_Intq4a8u_1_argbuf_rwb_done = (readPointer_QTree_Intq4a8u_1_argbuf_rwb_emitted | ({lizzieLet6_6_d[0],
                                                                                                             lizzieLet6_5_d[0],
                                                                                                             lizzieLet6_4_d[0],
                                                                                                             lizzieLet6_3_d[0],
                                                                                                             lizzieLet6_2_d[0],
                                                                                                             lizzieLet6_1_d[0]} & {lizzieLet6_6_r,
                                                                                                                                   lizzieLet6_5_r,
                                                                                                                                   lizzieLet6_4_r,
                                                                                                                                   lizzieLet6_3_r,
                                                                                                                                   lizzieLet6_2_r,
                                                                                                                                   lizzieLet6_1_r}));
  assign readPointer_QTree_Intq4a8u_1_argbuf_rwb_r = (& readPointer_QTree_Intq4a8u_1_argbuf_rwb_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Intq4a8u_1_argbuf_rwb_emitted <= 6'd0;
    else
      readPointer_QTree_Intq4a8u_1_argbuf_rwb_emitted <= (readPointer_QTree_Intq4a8u_1_argbuf_rwb_r ? 6'd0 :
                                                          readPointer_QTree_Intq4a8u_1_argbuf_rwb_done);
  
  /* buf (Ty QTree_Int) : (readPointer_QTree_IntwsiX_1_1_argbuf,QTree_Int) > (readPointer_QTree_IntwsiX_1_1_argbuf_rwb,QTree_Int) */
  QTree_Int_t readPointer_QTree_IntwsiX_1_1_argbuf_bufchan_d;
  logic readPointer_QTree_IntwsiX_1_1_argbuf_bufchan_r;
  assign readPointer_QTree_IntwsiX_1_1_argbuf_r = ((! readPointer_QTree_IntwsiX_1_1_argbuf_bufchan_d[0]) || readPointer_QTree_IntwsiX_1_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_IntwsiX_1_1_argbuf_bufchan_d <= {66'd0, 1'd0};
    else
      if (readPointer_QTree_IntwsiX_1_1_argbuf_r)
        readPointer_QTree_IntwsiX_1_1_argbuf_bufchan_d <= readPointer_QTree_IntwsiX_1_1_argbuf_d;
  QTree_Int_t readPointer_QTree_IntwsiX_1_1_argbuf_bufchan_buf;
  assign readPointer_QTree_IntwsiX_1_1_argbuf_bufchan_r = (! readPointer_QTree_IntwsiX_1_1_argbuf_bufchan_buf[0]);
  assign readPointer_QTree_IntwsiX_1_1_argbuf_rwb_d = (readPointer_QTree_IntwsiX_1_1_argbuf_bufchan_buf[0] ? readPointer_QTree_IntwsiX_1_1_argbuf_bufchan_buf :
                                                       readPointer_QTree_IntwsiX_1_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_IntwsiX_1_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((readPointer_QTree_IntwsiX_1_1_argbuf_rwb_r && readPointer_QTree_IntwsiX_1_1_argbuf_bufchan_buf[0]))
        readPointer_QTree_IntwsiX_1_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
      else if (((! readPointer_QTree_IntwsiX_1_1_argbuf_rwb_r) && (! readPointer_QTree_IntwsiX_1_1_argbuf_bufchan_buf[0])))
        readPointer_QTree_IntwsiX_1_1_argbuf_bufchan_buf <= readPointer_QTree_IntwsiX_1_1_argbuf_bufchan_d;
  
  /* fork (Ty QTree_Int) : (readPointer_QTree_IntwsiX_1_1_argbuf_rwb,QTree_Int) > [(lizzieLet4_1,QTree_Int),
                                                                              (lizzieLet4_2,QTree_Int),
                                                                              (lizzieLet4_3,QTree_Int),
                                                                              (lizzieLet4_4,QTree_Int)] */
  logic [3:0] readPointer_QTree_IntwsiX_1_1_argbuf_rwb_emitted;
  logic [3:0] readPointer_QTree_IntwsiX_1_1_argbuf_rwb_done;
  assign lizzieLet4_1_d = {readPointer_QTree_IntwsiX_1_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_IntwsiX_1_1_argbuf_rwb_d[0] && (! readPointer_QTree_IntwsiX_1_1_argbuf_rwb_emitted[0]))};
  assign lizzieLet4_2_d = {readPointer_QTree_IntwsiX_1_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_IntwsiX_1_1_argbuf_rwb_d[0] && (! readPointer_QTree_IntwsiX_1_1_argbuf_rwb_emitted[1]))};
  assign lizzieLet4_3_d = {readPointer_QTree_IntwsiX_1_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_IntwsiX_1_1_argbuf_rwb_d[0] && (! readPointer_QTree_IntwsiX_1_1_argbuf_rwb_emitted[2]))};
  assign lizzieLet4_4_d = {readPointer_QTree_IntwsiX_1_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_IntwsiX_1_1_argbuf_rwb_d[0] && (! readPointer_QTree_IntwsiX_1_1_argbuf_rwb_emitted[3]))};
  assign readPointer_QTree_IntwsiX_1_1_argbuf_rwb_done = (readPointer_QTree_IntwsiX_1_1_argbuf_rwb_emitted | ({lizzieLet4_4_d[0],
                                                                                                               lizzieLet4_3_d[0],
                                                                                                               lizzieLet4_2_d[0],
                                                                                                               lizzieLet4_1_d[0]} & {lizzieLet4_4_r,
                                                                                                                                     lizzieLet4_3_r,
                                                                                                                                     lizzieLet4_2_r,
                                                                                                                                     lizzieLet4_1_r}));
  assign readPointer_QTree_IntwsiX_1_1_argbuf_rwb_r = (& readPointer_QTree_IntwsiX_1_1_argbuf_rwb_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_IntwsiX_1_1_argbuf_rwb_emitted <= 4'd0;
    else
      readPointer_QTree_IntwsiX_1_1_argbuf_rwb_emitted <= (readPointer_QTree_IntwsiX_1_1_argbuf_rwb_r ? 4'd0 :
                                                           readPointer_QTree_IntwsiX_1_1_argbuf_rwb_done);
  
  /* buf (Ty Pointer_CTf''''''''_f''''''''_Int_Int) : (sc_0_10_destruct,Pointer_CTf''''''''_f''''''''_Int_Int) > (sc_0_10_1_argbuf,Pointer_CTf''''''''_f''''''''_Int_Int) */
  \Pointer_CTf''''''''_f''''''''_Int_Int_t  sc_0_10_destruct_bufchan_d;
  logic sc_0_10_destruct_bufchan_r;
  assign sc_0_10_destruct_r = ((! sc_0_10_destruct_bufchan_d[0]) || sc_0_10_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) sc_0_10_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (sc_0_10_destruct_r)
        sc_0_10_destruct_bufchan_d <= sc_0_10_destruct_d;
  \Pointer_CTf''''''''_f''''''''_Int_Int_t  sc_0_10_destruct_bufchan_buf;
  assign sc_0_10_destruct_bufchan_r = (! sc_0_10_destruct_bufchan_buf[0]);
  assign sc_0_10_1_argbuf_d = (sc_0_10_destruct_bufchan_buf[0] ? sc_0_10_destruct_bufchan_buf :
                               sc_0_10_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) sc_0_10_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((sc_0_10_1_argbuf_r && sc_0_10_destruct_bufchan_buf[0]))
        sc_0_10_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! sc_0_10_1_argbuf_r) && (! sc_0_10_destruct_bufchan_buf[0])))
        sc_0_10_destruct_bufchan_buf <= sc_0_10_destruct_bufchan_d;
  
  /* buf (Ty Pointer_CTf_f_Int_Int) : (sc_0_14_destruct,Pointer_CTf_f_Int_Int) > (sc_0_14_1_argbuf,Pointer_CTf_f_Int_Int) */
  Pointer_CTf_f_Int_Int_t sc_0_14_destruct_bufchan_d;
  logic sc_0_14_destruct_bufchan_r;
  assign sc_0_14_destruct_r = ((! sc_0_14_destruct_bufchan_d[0]) || sc_0_14_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) sc_0_14_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (sc_0_14_destruct_r)
        sc_0_14_destruct_bufchan_d <= sc_0_14_destruct_d;
  Pointer_CTf_f_Int_Int_t sc_0_14_destruct_bufchan_buf;
  assign sc_0_14_destruct_bufchan_r = (! sc_0_14_destruct_bufchan_buf[0]);
  assign sc_0_14_1_argbuf_d = (sc_0_14_destruct_bufchan_buf[0] ? sc_0_14_destruct_bufchan_buf :
                               sc_0_14_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) sc_0_14_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((sc_0_14_1_argbuf_r && sc_0_14_destruct_bufchan_buf[0]))
        sc_0_14_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! sc_0_14_1_argbuf_r) && (! sc_0_14_destruct_bufchan_buf[0])))
        sc_0_14_destruct_bufchan_buf <= sc_0_14_destruct_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz) : (sc_0_6_destruct,Pointer_CT$wnnz) > (sc_0_6_1_argbuf,Pointer_CT$wnnz) */
  Pointer_CT$wnnz_t sc_0_6_destruct_bufchan_d;
  logic sc_0_6_destruct_bufchan_r;
  assign sc_0_6_destruct_r = ((! sc_0_6_destruct_bufchan_d[0]) || sc_0_6_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) sc_0_6_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (sc_0_6_destruct_r)
        sc_0_6_destruct_bufchan_d <= sc_0_6_destruct_d;
  Pointer_CT$wnnz_t sc_0_6_destruct_bufchan_buf;
  assign sc_0_6_destruct_bufchan_r = (! sc_0_6_destruct_bufchan_buf[0]);
  assign sc_0_6_1_argbuf_d = (sc_0_6_destruct_bufchan_buf[0] ? sc_0_6_destruct_bufchan_buf :
                              sc_0_6_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) sc_0_6_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((sc_0_6_1_argbuf_r && sc_0_6_destruct_bufchan_buf[0]))
        sc_0_6_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! sc_0_6_1_argbuf_r) && (! sc_0_6_destruct_bufchan_buf[0])))
        sc_0_6_destruct_bufchan_buf <= sc_0_6_destruct_bufchan_d;
  
  /* buf (Ty Pointer_CTf''''''''_f''''''''_Int_Int) : (scfarg_0_1_goMux_mux,Pointer_CTf''''''''_f''''''''_Int_Int) > (scfarg_0_1_1_argbuf,Pointer_CTf''''''''_f''''''''_Int_Int) */
  \Pointer_CTf''''''''_f''''''''_Int_Int_t  scfarg_0_1_goMux_mux_bufchan_d;
  logic scfarg_0_1_goMux_mux_bufchan_r;
  assign scfarg_0_1_goMux_mux_r = ((! scfarg_0_1_goMux_mux_bufchan_d[0]) || scfarg_0_1_goMux_mux_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      scfarg_0_1_goMux_mux_bufchan_d <= {16'd0, 1'd0};
    else
      if (scfarg_0_1_goMux_mux_r)
        scfarg_0_1_goMux_mux_bufchan_d <= scfarg_0_1_goMux_mux_d;
  \Pointer_CTf''''''''_f''''''''_Int_Int_t  scfarg_0_1_goMux_mux_bufchan_buf;
  assign scfarg_0_1_goMux_mux_bufchan_r = (! scfarg_0_1_goMux_mux_bufchan_buf[0]);
  assign scfarg_0_1_1_argbuf_d = (scfarg_0_1_goMux_mux_bufchan_buf[0] ? scfarg_0_1_goMux_mux_bufchan_buf :
                                  scfarg_0_1_goMux_mux_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      scfarg_0_1_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((scfarg_0_1_1_argbuf_r && scfarg_0_1_goMux_mux_bufchan_buf[0]))
        scfarg_0_1_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
      else if (((! scfarg_0_1_1_argbuf_r) && (! scfarg_0_1_goMux_mux_bufchan_buf[0])))
        scfarg_0_1_goMux_mux_bufchan_buf <= scfarg_0_1_goMux_mux_bufchan_d;
  
  /* buf (Ty Pointer_CTf_f_Int_Int) : (scfarg_0_2_goMux_mux,Pointer_CTf_f_Int_Int) > (scfarg_0_2_1_argbuf,Pointer_CTf_f_Int_Int) */
  Pointer_CTf_f_Int_Int_t scfarg_0_2_goMux_mux_bufchan_d;
  logic scfarg_0_2_goMux_mux_bufchan_r;
  assign scfarg_0_2_goMux_mux_r = ((! scfarg_0_2_goMux_mux_bufchan_d[0]) || scfarg_0_2_goMux_mux_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      scfarg_0_2_goMux_mux_bufchan_d <= {16'd0, 1'd0};
    else
      if (scfarg_0_2_goMux_mux_r)
        scfarg_0_2_goMux_mux_bufchan_d <= scfarg_0_2_goMux_mux_d;
  Pointer_CTf_f_Int_Int_t scfarg_0_2_goMux_mux_bufchan_buf;
  assign scfarg_0_2_goMux_mux_bufchan_r = (! scfarg_0_2_goMux_mux_bufchan_buf[0]);
  assign scfarg_0_2_1_argbuf_d = (scfarg_0_2_goMux_mux_bufchan_buf[0] ? scfarg_0_2_goMux_mux_bufchan_buf :
                                  scfarg_0_2_goMux_mux_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      scfarg_0_2_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((scfarg_0_2_1_argbuf_r && scfarg_0_2_goMux_mux_bufchan_buf[0]))
        scfarg_0_2_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
      else if (((! scfarg_0_2_1_argbuf_r) && (! scfarg_0_2_goMux_mux_bufchan_buf[0])))
        scfarg_0_2_goMux_mux_bufchan_buf <= scfarg_0_2_goMux_mux_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz) : (scfarg_0_goMux_mux,Pointer_CT$wnnz) > (scfarg_0_1_argbuf,Pointer_CT$wnnz) */
  Pointer_CT$wnnz_t scfarg_0_goMux_mux_bufchan_d;
  logic scfarg_0_goMux_mux_bufchan_r;
  assign scfarg_0_goMux_mux_r = ((! scfarg_0_goMux_mux_bufchan_d[0]) || scfarg_0_goMux_mux_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) scfarg_0_goMux_mux_bufchan_d <= {16'd0, 1'd0};
    else
      if (scfarg_0_goMux_mux_r)
        scfarg_0_goMux_mux_bufchan_d <= scfarg_0_goMux_mux_d;
  Pointer_CT$wnnz_t scfarg_0_goMux_mux_bufchan_buf;
  assign scfarg_0_goMux_mux_bufchan_r = (! scfarg_0_goMux_mux_bufchan_buf[0]);
  assign scfarg_0_1_argbuf_d = (scfarg_0_goMux_mux_bufchan_buf[0] ? scfarg_0_goMux_mux_bufchan_buf :
                                scfarg_0_goMux_mux_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      scfarg_0_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((scfarg_0_1_argbuf_r && scfarg_0_goMux_mux_bufchan_buf[0]))
        scfarg_0_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
      else if (((! scfarg_0_1_argbuf_r) && (! scfarg_0_goMux_mux_bufchan_buf[0])))
        scfarg_0_goMux_mux_bufchan_buf <= scfarg_0_goMux_mux_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (t1a8Y_3_destruct,Pointer_QTree_Int) > (t1a8Y_3_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t t1a8Y_3_destruct_bufchan_d;
  logic t1a8Y_3_destruct_bufchan_r;
  assign t1a8Y_3_destruct_r = ((! t1a8Y_3_destruct_bufchan_d[0]) || t1a8Y_3_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t1a8Y_3_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (t1a8Y_3_destruct_r)
        t1a8Y_3_destruct_bufchan_d <= t1a8Y_3_destruct_d;
  Pointer_QTree_Int_t t1a8Y_3_destruct_bufchan_buf;
  assign t1a8Y_3_destruct_bufchan_r = (! t1a8Y_3_destruct_bufchan_buf[0]);
  assign t1a8Y_3_1_argbuf_d = (t1a8Y_3_destruct_bufchan_buf[0] ? t1a8Y_3_destruct_bufchan_buf :
                               t1a8Y_3_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t1a8Y_3_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((t1a8Y_3_1_argbuf_r && t1a8Y_3_destruct_bufchan_buf[0]))
        t1a8Y_3_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! t1a8Y_3_1_argbuf_r) && (! t1a8Y_3_destruct_bufchan_buf[0])))
        t1a8Y_3_destruct_bufchan_buf <= t1a8Y_3_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (t2a8Z_2_destruct,Pointer_QTree_Int) > (t2a8Z_2_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t t2a8Z_2_destruct_bufchan_d;
  logic t2a8Z_2_destruct_bufchan_r;
  assign t2a8Z_2_destruct_r = ((! t2a8Z_2_destruct_bufchan_d[0]) || t2a8Z_2_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t2a8Z_2_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (t2a8Z_2_destruct_r)
        t2a8Z_2_destruct_bufchan_d <= t2a8Z_2_destruct_d;
  Pointer_QTree_Int_t t2a8Z_2_destruct_bufchan_buf;
  assign t2a8Z_2_destruct_bufchan_r = (! t2a8Z_2_destruct_bufchan_buf[0]);
  assign t2a8Z_2_1_argbuf_d = (t2a8Z_2_destruct_bufchan_buf[0] ? t2a8Z_2_destruct_bufchan_buf :
                               t2a8Z_2_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t2a8Z_2_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((t2a8Z_2_1_argbuf_r && t2a8Z_2_destruct_bufchan_buf[0]))
        t2a8Z_2_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! t2a8Z_2_1_argbuf_r) && (! t2a8Z_2_destruct_bufchan_buf[0])))
        t2a8Z_2_destruct_bufchan_buf <= t2a8Z_2_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (t3a90_1_destruct,Pointer_QTree_Int) > (t3a90_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t t3a90_1_destruct_bufchan_d;
  logic t3a90_1_destruct_bufchan_r;
  assign t3a90_1_destruct_r = ((! t3a90_1_destruct_bufchan_d[0]) || t3a90_1_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t3a90_1_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (t3a90_1_destruct_r)
        t3a90_1_destruct_bufchan_d <= t3a90_1_destruct_d;
  Pointer_QTree_Int_t t3a90_1_destruct_bufchan_buf;
  assign t3a90_1_destruct_bufchan_r = (! t3a90_1_destruct_bufchan_buf[0]);
  assign t3a90_1_1_argbuf_d = (t3a90_1_destruct_bufchan_buf[0] ? t3a90_1_destruct_bufchan_buf :
                               t3a90_1_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t3a90_1_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((t3a90_1_1_argbuf_r && t3a90_1_destruct_bufchan_buf[0]))
        t3a90_1_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! t3a90_1_1_argbuf_r) && (! t3a90_1_destruct_bufchan_buf[0])))
        t3a90_1_destruct_bufchan_buf <= t3a90_1_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (t4a91_destruct,Pointer_QTree_Int) > (t4a91_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t t4a91_destruct_bufchan_d;
  logic t4a91_destruct_bufchan_r;
  assign t4a91_destruct_r = ((! t4a91_destruct_bufchan_d[0]) || t4a91_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t4a91_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (t4a91_destruct_r) t4a91_destruct_bufchan_d <= t4a91_destruct_d;
  Pointer_QTree_Int_t t4a91_destruct_bufchan_buf;
  assign t4a91_destruct_bufchan_r = (! t4a91_destruct_bufchan_buf[0]);
  assign t4a91_1_argbuf_d = (t4a91_destruct_bufchan_buf[0] ? t4a91_destruct_bufchan_buf :
                             t4a91_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t4a91_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((t4a91_1_argbuf_r && t4a91_destruct_bufchan_buf[0]))
        t4a91_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! t4a91_1_argbuf_r) && (! t4a91_destruct_bufchan_buf[0])))
        t4a91_destruct_bufchan_buf <= t4a91_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (tla8J_destruct,Pointer_QTree_Int) > (tla8J_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t tla8J_destruct_bufchan_d;
  logic tla8J_destruct_bufchan_r;
  assign tla8J_destruct_r = ((! tla8J_destruct_bufchan_d[0]) || tla8J_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) tla8J_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (tla8J_destruct_r) tla8J_destruct_bufchan_d <= tla8J_destruct_d;
  Pointer_QTree_Int_t tla8J_destruct_bufchan_buf;
  assign tla8J_destruct_bufchan_r = (! tla8J_destruct_bufchan_buf[0]);
  assign tla8J_1_argbuf_d = (tla8J_destruct_bufchan_buf[0] ? tla8J_destruct_bufchan_buf :
                             tla8J_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) tla8J_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((tla8J_1_argbuf_r && tla8J_destruct_bufchan_buf[0]))
        tla8J_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! tla8J_1_argbuf_r) && (! tla8J_destruct_bufchan_buf[0])))
        tla8J_destruct_bufchan_buf <= tla8J_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (tla8y_3_destruct,Pointer_QTree_Int) > (tla8y_3_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t tla8y_3_destruct_bufchan_d;
  logic tla8y_3_destruct_bufchan_r;
  assign tla8y_3_destruct_r = ((! tla8y_3_destruct_bufchan_d[0]) || tla8y_3_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) tla8y_3_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (tla8y_3_destruct_r)
        tla8y_3_destruct_bufchan_d <= tla8y_3_destruct_d;
  Pointer_QTree_Int_t tla8y_3_destruct_bufchan_buf;
  assign tla8y_3_destruct_bufchan_r = (! tla8y_3_destruct_bufchan_buf[0]);
  assign tla8y_3_1_argbuf_d = (tla8y_3_destruct_bufchan_buf[0] ? tla8y_3_destruct_bufchan_buf :
                               tla8y_3_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) tla8y_3_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((tla8y_3_1_argbuf_r && tla8y_3_destruct_bufchan_buf[0]))
        tla8y_3_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! tla8y_3_1_argbuf_r) && (! tla8y_3_destruct_bufchan_buf[0])))
        tla8y_3_destruct_bufchan_buf <= tla8y_3_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (tra8K_destruct,Pointer_QTree_Int) > (tra8K_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t tra8K_destruct_bufchan_d;
  logic tra8K_destruct_bufchan_r;
  assign tra8K_destruct_r = ((! tra8K_destruct_bufchan_d[0]) || tra8K_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) tra8K_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (tra8K_destruct_r) tra8K_destruct_bufchan_d <= tra8K_destruct_d;
  Pointer_QTree_Int_t tra8K_destruct_bufchan_buf;
  assign tra8K_destruct_bufchan_r = (! tra8K_destruct_bufchan_buf[0]);
  assign tra8K_1_argbuf_d = (tra8K_destruct_bufchan_buf[0] ? tra8K_destruct_bufchan_buf :
                             tra8K_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) tra8K_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((tra8K_1_argbuf_r && tra8K_destruct_bufchan_buf[0]))
        tra8K_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! tra8K_1_argbuf_r) && (! tra8K_destruct_bufchan_buf[0])))
        tra8K_destruct_bufchan_buf <= tra8K_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (tra8z_2_destruct,Pointer_QTree_Int) > (tra8z_2_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t tra8z_2_destruct_bufchan_d;
  logic tra8z_2_destruct_bufchan_r;
  assign tra8z_2_destruct_r = ((! tra8z_2_destruct_bufchan_d[0]) || tra8z_2_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) tra8z_2_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (tra8z_2_destruct_r)
        tra8z_2_destruct_bufchan_d <= tra8z_2_destruct_d;
  Pointer_QTree_Int_t tra8z_2_destruct_bufchan_buf;
  assign tra8z_2_destruct_bufchan_r = (! tra8z_2_destruct_bufchan_buf[0]);
  assign tra8z_2_1_argbuf_d = (tra8z_2_destruct_bufchan_buf[0] ? tra8z_2_destruct_bufchan_buf :
                               tra8z_2_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) tra8z_2_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((tra8z_2_1_argbuf_r && tra8z_2_destruct_bufchan_buf[0]))
        tra8z_2_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! tra8z_2_1_argbuf_r) && (! tra8z_2_destruct_bufchan_buf[0])))
        tra8z_2_destruct_bufchan_buf <= tra8z_2_destruct_bufchan_d;
  
  /* buf (Ty Int) : (va8I_1,Int) > (va8I_1_argbuf,Int) */
  Int_t va8I_1_bufchan_d;
  logic va8I_1_bufchan_r;
  assign va8I_1_r = ((! va8I_1_bufchan_d[0]) || va8I_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) va8I_1_bufchan_d <= {32'd0, 1'd0};
    else if (va8I_1_r) va8I_1_bufchan_d <= va8I_1_d;
  Int_t va8I_1_bufchan_buf;
  assign va8I_1_bufchan_r = (! va8I_1_bufchan_buf[0]);
  assign va8I_1_argbuf_d = (va8I_1_bufchan_buf[0] ? va8I_1_bufchan_buf :
                            va8I_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) va8I_1_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((va8I_1_argbuf_r && va8I_1_bufchan_buf[0]))
        va8I_1_bufchan_buf <= {32'd0, 1'd0};
      else if (((! va8I_1_argbuf_r) && (! va8I_1_bufchan_buf[0])))
        va8I_1_bufchan_buf <= va8I_1_bufchan_d;
  
  /* fork (Ty Int) : (va8I_destruct,Int) > [(va8I_1,Int),(va8I_2,Int)] */
  logic [1:0] va8I_destruct_emitted;
  logic [1:0] va8I_destruct_done;
  assign va8I_1_d = {va8I_destruct_d[32:1],
                     (va8I_destruct_d[0] && (! va8I_destruct_emitted[0]))};
  assign va8I_2_d = {va8I_destruct_d[32:1],
                     (va8I_destruct_d[0] && (! va8I_destruct_emitted[1]))};
  assign va8I_destruct_done = (va8I_destruct_emitted | ({va8I_2_d[0],
                                                         va8I_1_d[0]} & {va8I_2_r, va8I_1_r}));
  assign va8I_destruct_r = (& va8I_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) va8I_destruct_emitted <= 2'd0;
    else
      va8I_destruct_emitted <= (va8I_destruct_r ? 2'd0 :
                                va8I_destruct_done);
  
  /* buf (Ty Int) : (va8O_1,Int) > (va8O_1_argbuf,Int) */
  Int_t va8O_1_bufchan_d;
  logic va8O_1_bufchan_r;
  assign va8O_1_r = ((! va8O_1_bufchan_d[0]) || va8O_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) va8O_1_bufchan_d <= {32'd0, 1'd0};
    else if (va8O_1_r) va8O_1_bufchan_d <= va8O_1_d;
  Int_t va8O_1_bufchan_buf;
  assign va8O_1_bufchan_r = (! va8O_1_bufchan_buf[0]);
  assign va8O_1_argbuf_d = (va8O_1_bufchan_buf[0] ? va8O_1_bufchan_buf :
                            va8O_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) va8O_1_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((va8O_1_argbuf_r && va8O_1_bufchan_buf[0]))
        va8O_1_bufchan_buf <= {32'd0, 1'd0};
      else if (((! va8O_1_argbuf_r) && (! va8O_1_bufchan_buf[0])))
        va8O_1_bufchan_buf <= va8O_1_bufchan_d;
  
  /* fork (Ty Int) : (va8O_destruct,Int) > [(va8O_1,Int),(va8O_2,Int)] */
  logic [1:0] va8O_destruct_emitted;
  logic [1:0] va8O_destruct_done;
  assign va8O_1_d = {va8O_destruct_d[32:1],
                     (va8O_destruct_d[0] && (! va8O_destruct_emitted[0]))};
  assign va8O_2_d = {va8O_destruct_d[32:1],
                     (va8O_destruct_d[0] && (! va8O_destruct_emitted[1]))};
  assign va8O_destruct_done = (va8O_destruct_emitted | ({va8O_2_d[0],
                                                         va8O_1_d[0]} & {va8O_2_r, va8O_1_r}));
  assign va8O_destruct_r = (& va8O_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) va8O_destruct_emitted <= 2'd0;
    else
      va8O_destruct_emitted <= (va8O_destruct_r ? 2'd0 :
                                va8O_destruct_done);
  
  /* buf (Ty Int) : (va8x_1,Int) > (va8x_1_argbuf,Int) */
  Int_t va8x_1_bufchan_d;
  logic va8x_1_bufchan_r;
  assign va8x_1_r = ((! va8x_1_bufchan_d[0]) || va8x_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) va8x_1_bufchan_d <= {32'd0, 1'd0};
    else if (va8x_1_r) va8x_1_bufchan_d <= va8x_1_d;
  Int_t va8x_1_bufchan_buf;
  assign va8x_1_bufchan_r = (! va8x_1_bufchan_buf[0]);
  assign va8x_1_argbuf_d = (va8x_1_bufchan_buf[0] ? va8x_1_bufchan_buf :
                            va8x_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) va8x_1_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((va8x_1_argbuf_r && va8x_1_bufchan_buf[0]))
        va8x_1_bufchan_buf <= {32'd0, 1'd0};
      else if (((! va8x_1_argbuf_r) && (! va8x_1_bufchan_buf[0])))
        va8x_1_bufchan_buf <= va8x_1_bufchan_d;
  
  /* fork (Ty Int) : (va8x_destruct,Int) > [(va8x_1,Int),(va8x_2,Int)] */
  logic [1:0] va8x_destruct_emitted;
  logic [1:0] va8x_destruct_done;
  assign va8x_1_d = {va8x_destruct_d[32:1],
                     (va8x_destruct_d[0] && (! va8x_destruct_emitted[0]))};
  assign va8x_2_d = {va8x_destruct_d[32:1],
                     (va8x_destruct_d[0] && (! va8x_destruct_emitted[1]))};
  assign va8x_destruct_done = (va8x_destruct_emitted | ({va8x_2_d[0],
                                                         va8x_1_d[0]} & {va8x_2_r, va8x_1_r}));
  assign va8x_destruct_r = (& va8x_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) va8x_destruct_emitted <= 2'd0;
    else
      va8x_destruct_emitted <= (va8x_destruct_r ? 2'd0 :
                                va8x_destruct_done);
  
  /* buf (Ty Pointer_CT$wnnz) : (writeCT$wnnzlizzieLet0_1_argbuf,Pointer_CT$wnnz) > (writeCT$wnnzlizzieLet0_1_argbuf_rwb,Pointer_CT$wnnz) */
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet0_1_argbuf_bufchan_d;
  logic writeCT$wnnzlizzieLet0_1_argbuf_bufchan_r;
  assign writeCT$wnnzlizzieLet0_1_argbuf_r = ((! writeCT$wnnzlizzieLet0_1_argbuf_bufchan_d[0]) || writeCT$wnnzlizzieLet0_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnzlizzieLet0_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCT$wnnzlizzieLet0_1_argbuf_r)
        writeCT$wnnzlizzieLet0_1_argbuf_bufchan_d <= writeCT$wnnzlizzieLet0_1_argbuf_d;
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet0_1_argbuf_bufchan_buf;
  assign writeCT$wnnzlizzieLet0_1_argbuf_bufchan_r = (! writeCT$wnnzlizzieLet0_1_argbuf_bufchan_buf[0]);
  assign writeCT$wnnzlizzieLet0_1_argbuf_rwb_d = (writeCT$wnnzlizzieLet0_1_argbuf_bufchan_buf[0] ? writeCT$wnnzlizzieLet0_1_argbuf_bufchan_buf :
                                                  writeCT$wnnzlizzieLet0_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnzlizzieLet0_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeCT$wnnzlizzieLet0_1_argbuf_rwb_r && writeCT$wnnzlizzieLet0_1_argbuf_bufchan_buf[0]))
        writeCT$wnnzlizzieLet0_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeCT$wnnzlizzieLet0_1_argbuf_rwb_r) && (! writeCT$wnnzlizzieLet0_1_argbuf_bufchan_buf[0])))
        writeCT$wnnzlizzieLet0_1_argbuf_bufchan_buf <= writeCT$wnnzlizzieLet0_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz) : (writeCT$wnnzlizzieLet0_1_argbuf_rwb,Pointer_CT$wnnz) > (lizzieLet25_1_argbuf,Pointer_CT$wnnz) */
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet0_1_argbuf_rwb_bufchan_d;
  logic writeCT$wnnzlizzieLet0_1_argbuf_rwb_bufchan_r;
  assign writeCT$wnnzlizzieLet0_1_argbuf_rwb_r = ((! writeCT$wnnzlizzieLet0_1_argbuf_rwb_bufchan_d[0]) || writeCT$wnnzlizzieLet0_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnzlizzieLet0_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCT$wnnzlizzieLet0_1_argbuf_rwb_r)
        writeCT$wnnzlizzieLet0_1_argbuf_rwb_bufchan_d <= writeCT$wnnzlizzieLet0_1_argbuf_rwb_d;
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet0_1_argbuf_rwb_bufchan_buf;
  assign writeCT$wnnzlizzieLet0_1_argbuf_rwb_bufchan_r = (! writeCT$wnnzlizzieLet0_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet25_1_argbuf_d = (writeCT$wnnzlizzieLet0_1_argbuf_rwb_bufchan_buf[0] ? writeCT$wnnzlizzieLet0_1_argbuf_rwb_bufchan_buf :
                                   writeCT$wnnzlizzieLet0_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnzlizzieLet0_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet25_1_argbuf_r && writeCT$wnnzlizzieLet0_1_argbuf_rwb_bufchan_buf[0]))
        writeCT$wnnzlizzieLet0_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet25_1_argbuf_r) && (! writeCT$wnnzlizzieLet0_1_argbuf_rwb_bufchan_buf[0])))
        writeCT$wnnzlizzieLet0_1_argbuf_rwb_bufchan_buf <= writeCT$wnnzlizzieLet0_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz) : (writeCT$wnnzlizzieLet36_1_argbuf,Pointer_CT$wnnz) > (writeCT$wnnzlizzieLet36_1_argbuf_rwb,Pointer_CT$wnnz) */
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet36_1_argbuf_bufchan_d;
  logic writeCT$wnnzlizzieLet36_1_argbuf_bufchan_r;
  assign writeCT$wnnzlizzieLet36_1_argbuf_r = ((! writeCT$wnnzlizzieLet36_1_argbuf_bufchan_d[0]) || writeCT$wnnzlizzieLet36_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnzlizzieLet36_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCT$wnnzlizzieLet36_1_argbuf_r)
        writeCT$wnnzlizzieLet36_1_argbuf_bufchan_d <= writeCT$wnnzlizzieLet36_1_argbuf_d;
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet36_1_argbuf_bufchan_buf;
  assign writeCT$wnnzlizzieLet36_1_argbuf_bufchan_r = (! writeCT$wnnzlizzieLet36_1_argbuf_bufchan_buf[0]);
  assign writeCT$wnnzlizzieLet36_1_argbuf_rwb_d = (writeCT$wnnzlizzieLet36_1_argbuf_bufchan_buf[0] ? writeCT$wnnzlizzieLet36_1_argbuf_bufchan_buf :
                                                   writeCT$wnnzlizzieLet36_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnzlizzieLet36_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeCT$wnnzlizzieLet36_1_argbuf_rwb_r && writeCT$wnnzlizzieLet36_1_argbuf_bufchan_buf[0]))
        writeCT$wnnzlizzieLet36_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeCT$wnnzlizzieLet36_1_argbuf_rwb_r) && (! writeCT$wnnzlizzieLet36_1_argbuf_bufchan_buf[0])))
        writeCT$wnnzlizzieLet36_1_argbuf_bufchan_buf <= writeCT$wnnzlizzieLet36_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz) : (writeCT$wnnzlizzieLet36_1_argbuf_rwb,Pointer_CT$wnnz) > (sca2_1_argbuf,Pointer_CT$wnnz) */
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet36_1_argbuf_rwb_bufchan_d;
  logic writeCT$wnnzlizzieLet36_1_argbuf_rwb_bufchan_r;
  assign writeCT$wnnzlizzieLet36_1_argbuf_rwb_r = ((! writeCT$wnnzlizzieLet36_1_argbuf_rwb_bufchan_d[0]) || writeCT$wnnzlizzieLet36_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnzlizzieLet36_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCT$wnnzlizzieLet36_1_argbuf_rwb_r)
        writeCT$wnnzlizzieLet36_1_argbuf_rwb_bufchan_d <= writeCT$wnnzlizzieLet36_1_argbuf_rwb_d;
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet36_1_argbuf_rwb_bufchan_buf;
  assign writeCT$wnnzlizzieLet36_1_argbuf_rwb_bufchan_r = (! writeCT$wnnzlizzieLet36_1_argbuf_rwb_bufchan_buf[0]);
  assign sca2_1_argbuf_d = (writeCT$wnnzlizzieLet36_1_argbuf_rwb_bufchan_buf[0] ? writeCT$wnnzlizzieLet36_1_argbuf_rwb_bufchan_buf :
                            writeCT$wnnzlizzieLet36_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnzlizzieLet36_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((sca2_1_argbuf_r && writeCT$wnnzlizzieLet36_1_argbuf_rwb_bufchan_buf[0]))
        writeCT$wnnzlizzieLet36_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
      else if (((! sca2_1_argbuf_r) && (! writeCT$wnnzlizzieLet36_1_argbuf_rwb_bufchan_buf[0])))
        writeCT$wnnzlizzieLet36_1_argbuf_rwb_bufchan_buf <= writeCT$wnnzlizzieLet36_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz) : (writeCT$wnnzlizzieLet37_1_argbuf,Pointer_CT$wnnz) > (writeCT$wnnzlizzieLet37_1_argbuf_rwb,Pointer_CT$wnnz) */
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet37_1_argbuf_bufchan_d;
  logic writeCT$wnnzlizzieLet37_1_argbuf_bufchan_r;
  assign writeCT$wnnzlizzieLet37_1_argbuf_r = ((! writeCT$wnnzlizzieLet37_1_argbuf_bufchan_d[0]) || writeCT$wnnzlizzieLet37_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnzlizzieLet37_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCT$wnnzlizzieLet37_1_argbuf_r)
        writeCT$wnnzlizzieLet37_1_argbuf_bufchan_d <= writeCT$wnnzlizzieLet37_1_argbuf_d;
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet37_1_argbuf_bufchan_buf;
  assign writeCT$wnnzlizzieLet37_1_argbuf_bufchan_r = (! writeCT$wnnzlizzieLet37_1_argbuf_bufchan_buf[0]);
  assign writeCT$wnnzlizzieLet37_1_argbuf_rwb_d = (writeCT$wnnzlizzieLet37_1_argbuf_bufchan_buf[0] ? writeCT$wnnzlizzieLet37_1_argbuf_bufchan_buf :
                                                   writeCT$wnnzlizzieLet37_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnzlizzieLet37_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeCT$wnnzlizzieLet37_1_argbuf_rwb_r && writeCT$wnnzlizzieLet37_1_argbuf_bufchan_buf[0]))
        writeCT$wnnzlizzieLet37_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeCT$wnnzlizzieLet37_1_argbuf_rwb_r) && (! writeCT$wnnzlizzieLet37_1_argbuf_bufchan_buf[0])))
        writeCT$wnnzlizzieLet37_1_argbuf_bufchan_buf <= writeCT$wnnzlizzieLet37_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz) : (writeCT$wnnzlizzieLet37_1_argbuf_rwb,Pointer_CT$wnnz) > (sca1_1_argbuf,Pointer_CT$wnnz) */
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet37_1_argbuf_rwb_bufchan_d;
  logic writeCT$wnnzlizzieLet37_1_argbuf_rwb_bufchan_r;
  assign writeCT$wnnzlizzieLet37_1_argbuf_rwb_r = ((! writeCT$wnnzlizzieLet37_1_argbuf_rwb_bufchan_d[0]) || writeCT$wnnzlizzieLet37_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnzlizzieLet37_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCT$wnnzlizzieLet37_1_argbuf_rwb_r)
        writeCT$wnnzlizzieLet37_1_argbuf_rwb_bufchan_d <= writeCT$wnnzlizzieLet37_1_argbuf_rwb_d;
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet37_1_argbuf_rwb_bufchan_buf;
  assign writeCT$wnnzlizzieLet37_1_argbuf_rwb_bufchan_r = (! writeCT$wnnzlizzieLet37_1_argbuf_rwb_bufchan_buf[0]);
  assign sca1_1_argbuf_d = (writeCT$wnnzlizzieLet37_1_argbuf_rwb_bufchan_buf[0] ? writeCT$wnnzlizzieLet37_1_argbuf_rwb_bufchan_buf :
                            writeCT$wnnzlizzieLet37_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnzlizzieLet37_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((sca1_1_argbuf_r && writeCT$wnnzlizzieLet37_1_argbuf_rwb_bufchan_buf[0]))
        writeCT$wnnzlizzieLet37_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
      else if (((! sca1_1_argbuf_r) && (! writeCT$wnnzlizzieLet37_1_argbuf_rwb_bufchan_buf[0])))
        writeCT$wnnzlizzieLet37_1_argbuf_rwb_bufchan_buf <= writeCT$wnnzlizzieLet37_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz) : (writeCT$wnnzlizzieLet38_1_argbuf,Pointer_CT$wnnz) > (writeCT$wnnzlizzieLet38_1_argbuf_rwb,Pointer_CT$wnnz) */
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet38_1_argbuf_bufchan_d;
  logic writeCT$wnnzlizzieLet38_1_argbuf_bufchan_r;
  assign writeCT$wnnzlizzieLet38_1_argbuf_r = ((! writeCT$wnnzlizzieLet38_1_argbuf_bufchan_d[0]) || writeCT$wnnzlizzieLet38_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnzlizzieLet38_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCT$wnnzlizzieLet38_1_argbuf_r)
        writeCT$wnnzlizzieLet38_1_argbuf_bufchan_d <= writeCT$wnnzlizzieLet38_1_argbuf_d;
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet38_1_argbuf_bufchan_buf;
  assign writeCT$wnnzlizzieLet38_1_argbuf_bufchan_r = (! writeCT$wnnzlizzieLet38_1_argbuf_bufchan_buf[0]);
  assign writeCT$wnnzlizzieLet38_1_argbuf_rwb_d = (writeCT$wnnzlizzieLet38_1_argbuf_bufchan_buf[0] ? writeCT$wnnzlizzieLet38_1_argbuf_bufchan_buf :
                                                   writeCT$wnnzlizzieLet38_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnzlizzieLet38_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeCT$wnnzlizzieLet38_1_argbuf_rwb_r && writeCT$wnnzlizzieLet38_1_argbuf_bufchan_buf[0]))
        writeCT$wnnzlizzieLet38_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeCT$wnnzlizzieLet38_1_argbuf_rwb_r) && (! writeCT$wnnzlizzieLet38_1_argbuf_bufchan_buf[0])))
        writeCT$wnnzlizzieLet38_1_argbuf_bufchan_buf <= writeCT$wnnzlizzieLet38_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz) : (writeCT$wnnzlizzieLet38_1_argbuf_rwb,Pointer_CT$wnnz) > (sca0_1_argbuf,Pointer_CT$wnnz) */
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet38_1_argbuf_rwb_bufchan_d;
  logic writeCT$wnnzlizzieLet38_1_argbuf_rwb_bufchan_r;
  assign writeCT$wnnzlizzieLet38_1_argbuf_rwb_r = ((! writeCT$wnnzlizzieLet38_1_argbuf_rwb_bufchan_d[0]) || writeCT$wnnzlizzieLet38_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnzlizzieLet38_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCT$wnnzlizzieLet38_1_argbuf_rwb_r)
        writeCT$wnnzlizzieLet38_1_argbuf_rwb_bufchan_d <= writeCT$wnnzlizzieLet38_1_argbuf_rwb_d;
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet38_1_argbuf_rwb_bufchan_buf;
  assign writeCT$wnnzlizzieLet38_1_argbuf_rwb_bufchan_r = (! writeCT$wnnzlizzieLet38_1_argbuf_rwb_bufchan_buf[0]);
  assign sca0_1_argbuf_d = (writeCT$wnnzlizzieLet38_1_argbuf_rwb_bufchan_buf[0] ? writeCT$wnnzlizzieLet38_1_argbuf_rwb_bufchan_buf :
                            writeCT$wnnzlizzieLet38_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnzlizzieLet38_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((sca0_1_argbuf_r && writeCT$wnnzlizzieLet38_1_argbuf_rwb_bufchan_buf[0]))
        writeCT$wnnzlizzieLet38_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
      else if (((! sca0_1_argbuf_r) && (! writeCT$wnnzlizzieLet38_1_argbuf_rwb_bufchan_buf[0])))
        writeCT$wnnzlizzieLet38_1_argbuf_rwb_bufchan_buf <= writeCT$wnnzlizzieLet38_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz) : (writeCT$wnnzlizzieLet5_1_argbuf,Pointer_CT$wnnz) > (writeCT$wnnzlizzieLet5_1_argbuf_rwb,Pointer_CT$wnnz) */
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet5_1_argbuf_bufchan_d;
  logic writeCT$wnnzlizzieLet5_1_argbuf_bufchan_r;
  assign writeCT$wnnzlizzieLet5_1_argbuf_r = ((! writeCT$wnnzlizzieLet5_1_argbuf_bufchan_d[0]) || writeCT$wnnzlizzieLet5_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnzlizzieLet5_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCT$wnnzlizzieLet5_1_argbuf_r)
        writeCT$wnnzlizzieLet5_1_argbuf_bufchan_d <= writeCT$wnnzlizzieLet5_1_argbuf_d;
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet5_1_argbuf_bufchan_buf;
  assign writeCT$wnnzlizzieLet5_1_argbuf_bufchan_r = (! writeCT$wnnzlizzieLet5_1_argbuf_bufchan_buf[0]);
  assign writeCT$wnnzlizzieLet5_1_argbuf_rwb_d = (writeCT$wnnzlizzieLet5_1_argbuf_bufchan_buf[0] ? writeCT$wnnzlizzieLet5_1_argbuf_bufchan_buf :
                                                  writeCT$wnnzlizzieLet5_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnzlizzieLet5_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeCT$wnnzlizzieLet5_1_argbuf_rwb_r && writeCT$wnnzlizzieLet5_1_argbuf_bufchan_buf[0]))
        writeCT$wnnzlizzieLet5_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeCT$wnnzlizzieLet5_1_argbuf_rwb_r) && (! writeCT$wnnzlizzieLet5_1_argbuf_bufchan_buf[0])))
        writeCT$wnnzlizzieLet5_1_argbuf_bufchan_buf <= writeCT$wnnzlizzieLet5_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz) : (writeCT$wnnzlizzieLet5_1_argbuf_rwb,Pointer_CT$wnnz) > (sca3_1_argbuf,Pointer_CT$wnnz) */
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet5_1_argbuf_rwb_bufchan_d;
  logic writeCT$wnnzlizzieLet5_1_argbuf_rwb_bufchan_r;
  assign writeCT$wnnzlizzieLet5_1_argbuf_rwb_r = ((! writeCT$wnnzlizzieLet5_1_argbuf_rwb_bufchan_d[0]) || writeCT$wnnzlizzieLet5_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnzlizzieLet5_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCT$wnnzlizzieLet5_1_argbuf_rwb_r)
        writeCT$wnnzlizzieLet5_1_argbuf_rwb_bufchan_d <= writeCT$wnnzlizzieLet5_1_argbuf_rwb_d;
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet5_1_argbuf_rwb_bufchan_buf;
  assign writeCT$wnnzlizzieLet5_1_argbuf_rwb_bufchan_r = (! writeCT$wnnzlizzieLet5_1_argbuf_rwb_bufchan_buf[0]);
  assign sca3_1_argbuf_d = (writeCT$wnnzlizzieLet5_1_argbuf_rwb_bufchan_buf[0] ? writeCT$wnnzlizzieLet5_1_argbuf_rwb_bufchan_buf :
                            writeCT$wnnzlizzieLet5_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnzlizzieLet5_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((sca3_1_argbuf_r && writeCT$wnnzlizzieLet5_1_argbuf_rwb_bufchan_buf[0]))
        writeCT$wnnzlizzieLet5_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
      else if (((! sca3_1_argbuf_r) && (! writeCT$wnnzlizzieLet5_1_argbuf_rwb_bufchan_buf[0])))
        writeCT$wnnzlizzieLet5_1_argbuf_rwb_bufchan_buf <= writeCT$wnnzlizzieLet5_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CTf''''''''_f''''''''_Int_Int) : (writeCTf''''''''_f''''''''_Int_IntlizzieLet10_1_argbuf,Pointer_CTf''''''''_f''''''''_Int_Int) > (writeCTf''''''''_f''''''''_Int_IntlizzieLet10_1_argbuf_rwb,Pointer_CTf''''''''_f''''''''_Int_Int) */
  \Pointer_CTf''''''''_f''''''''_Int_Int_t  \writeCTf''''''''_f''''''''_Int_IntlizzieLet10_1_argbuf_bufchan_d ;
  logic \writeCTf''''''''_f''''''''_Int_IntlizzieLet10_1_argbuf_bufchan_r ;
  assign \writeCTf''''''''_f''''''''_Int_IntlizzieLet10_1_argbuf_r  = ((! \writeCTf''''''''_f''''''''_Int_IntlizzieLet10_1_argbuf_bufchan_d [0]) || \writeCTf''''''''_f''''''''_Int_IntlizzieLet10_1_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf''''''''_f''''''''_Int_IntlizzieLet10_1_argbuf_bufchan_d  <= {16'd0,
                                                                             1'd0};
    else
      if (\writeCTf''''''''_f''''''''_Int_IntlizzieLet10_1_argbuf_r )
        \writeCTf''''''''_f''''''''_Int_IntlizzieLet10_1_argbuf_bufchan_d  <= \writeCTf''''''''_f''''''''_Int_IntlizzieLet10_1_argbuf_d ;
  \Pointer_CTf''''''''_f''''''''_Int_Int_t  \writeCTf''''''''_f''''''''_Int_IntlizzieLet10_1_argbuf_bufchan_buf ;
  assign \writeCTf''''''''_f''''''''_Int_IntlizzieLet10_1_argbuf_bufchan_r  = (! \writeCTf''''''''_f''''''''_Int_IntlizzieLet10_1_argbuf_bufchan_buf [0]);
  assign \writeCTf''''''''_f''''''''_Int_IntlizzieLet10_1_argbuf_rwb_d  = (\writeCTf''''''''_f''''''''_Int_IntlizzieLet10_1_argbuf_bufchan_buf [0] ? \writeCTf''''''''_f''''''''_Int_IntlizzieLet10_1_argbuf_bufchan_buf  :
                                                                           \writeCTf''''''''_f''''''''_Int_IntlizzieLet10_1_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf''''''''_f''''''''_Int_IntlizzieLet10_1_argbuf_bufchan_buf  <= {16'd0,
                                                                               1'd0};
    else
      if ((\writeCTf''''''''_f''''''''_Int_IntlizzieLet10_1_argbuf_rwb_r  && \writeCTf''''''''_f''''''''_Int_IntlizzieLet10_1_argbuf_bufchan_buf [0]))
        \writeCTf''''''''_f''''''''_Int_IntlizzieLet10_1_argbuf_bufchan_buf  <= {16'd0,
                                                                                 1'd0};
      else if (((! \writeCTf''''''''_f''''''''_Int_IntlizzieLet10_1_argbuf_rwb_r ) && (! \writeCTf''''''''_f''''''''_Int_IntlizzieLet10_1_argbuf_bufchan_buf [0])))
        \writeCTf''''''''_f''''''''_Int_IntlizzieLet10_1_argbuf_bufchan_buf  <= \writeCTf''''''''_f''''''''_Int_IntlizzieLet10_1_argbuf_bufchan_d ;
  
  /* buf (Ty Pointer_CTf''''''''_f''''''''_Int_Int) : (writeCTf''''''''_f''''''''_Int_IntlizzieLet10_1_argbuf_rwb,Pointer_CTf''''''''_f''''''''_Int_Int) > (sca3_1_1_argbuf,Pointer_CTf''''''''_f''''''''_Int_Int) */
  \Pointer_CTf''''''''_f''''''''_Int_Int_t  \writeCTf''''''''_f''''''''_Int_IntlizzieLet10_1_argbuf_rwb_bufchan_d ;
  logic \writeCTf''''''''_f''''''''_Int_IntlizzieLet10_1_argbuf_rwb_bufchan_r ;
  assign \writeCTf''''''''_f''''''''_Int_IntlizzieLet10_1_argbuf_rwb_r  = ((! \writeCTf''''''''_f''''''''_Int_IntlizzieLet10_1_argbuf_rwb_bufchan_d [0]) || \writeCTf''''''''_f''''''''_Int_IntlizzieLet10_1_argbuf_rwb_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf''''''''_f''''''''_Int_IntlizzieLet10_1_argbuf_rwb_bufchan_d  <= {16'd0,
                                                                                 1'd0};
    else
      if (\writeCTf''''''''_f''''''''_Int_IntlizzieLet10_1_argbuf_rwb_r )
        \writeCTf''''''''_f''''''''_Int_IntlizzieLet10_1_argbuf_rwb_bufchan_d  <= \writeCTf''''''''_f''''''''_Int_IntlizzieLet10_1_argbuf_rwb_d ;
  \Pointer_CTf''''''''_f''''''''_Int_Int_t  \writeCTf''''''''_f''''''''_Int_IntlizzieLet10_1_argbuf_rwb_bufchan_buf ;
  assign \writeCTf''''''''_f''''''''_Int_IntlizzieLet10_1_argbuf_rwb_bufchan_r  = (! \writeCTf''''''''_f''''''''_Int_IntlizzieLet10_1_argbuf_rwb_bufchan_buf [0]);
  assign sca3_1_1_argbuf_d = (\writeCTf''''''''_f''''''''_Int_IntlizzieLet10_1_argbuf_rwb_bufchan_buf [0] ? \writeCTf''''''''_f''''''''_Int_IntlizzieLet10_1_argbuf_rwb_bufchan_buf  :
                              \writeCTf''''''''_f''''''''_Int_IntlizzieLet10_1_argbuf_rwb_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf''''''''_f''''''''_Int_IntlizzieLet10_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                                   1'd0};
    else
      if ((sca3_1_1_argbuf_r && \writeCTf''''''''_f''''''''_Int_IntlizzieLet10_1_argbuf_rwb_bufchan_buf [0]))
        \writeCTf''''''''_f''''''''_Int_IntlizzieLet10_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                                     1'd0};
      else if (((! sca3_1_1_argbuf_r) && (! \writeCTf''''''''_f''''''''_Int_IntlizzieLet10_1_argbuf_rwb_bufchan_buf [0])))
        \writeCTf''''''''_f''''''''_Int_IntlizzieLet10_1_argbuf_rwb_bufchan_buf  <= \writeCTf''''''''_f''''''''_Int_IntlizzieLet10_1_argbuf_rwb_bufchan_d ;
  
  /* buf (Ty Pointer_CTf''''''''_f''''''''_Int_Int) : (writeCTf''''''''_f''''''''_Int_IntlizzieLet33_1_argbuf,Pointer_CTf''''''''_f''''''''_Int_Int) > (writeCTf''''''''_f''''''''_Int_IntlizzieLet33_1_argbuf_rwb,Pointer_CTf''''''''_f''''''''_Int_Int) */
  \Pointer_CTf''''''''_f''''''''_Int_Int_t  \writeCTf''''''''_f''''''''_Int_IntlizzieLet33_1_argbuf_bufchan_d ;
  logic \writeCTf''''''''_f''''''''_Int_IntlizzieLet33_1_argbuf_bufchan_r ;
  assign \writeCTf''''''''_f''''''''_Int_IntlizzieLet33_1_argbuf_r  = ((! \writeCTf''''''''_f''''''''_Int_IntlizzieLet33_1_argbuf_bufchan_d [0]) || \writeCTf''''''''_f''''''''_Int_IntlizzieLet33_1_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf''''''''_f''''''''_Int_IntlizzieLet33_1_argbuf_bufchan_d  <= {16'd0,
                                                                             1'd0};
    else
      if (\writeCTf''''''''_f''''''''_Int_IntlizzieLet33_1_argbuf_r )
        \writeCTf''''''''_f''''''''_Int_IntlizzieLet33_1_argbuf_bufchan_d  <= \writeCTf''''''''_f''''''''_Int_IntlizzieLet33_1_argbuf_d ;
  \Pointer_CTf''''''''_f''''''''_Int_Int_t  \writeCTf''''''''_f''''''''_Int_IntlizzieLet33_1_argbuf_bufchan_buf ;
  assign \writeCTf''''''''_f''''''''_Int_IntlizzieLet33_1_argbuf_bufchan_r  = (! \writeCTf''''''''_f''''''''_Int_IntlizzieLet33_1_argbuf_bufchan_buf [0]);
  assign \writeCTf''''''''_f''''''''_Int_IntlizzieLet33_1_argbuf_rwb_d  = (\writeCTf''''''''_f''''''''_Int_IntlizzieLet33_1_argbuf_bufchan_buf [0] ? \writeCTf''''''''_f''''''''_Int_IntlizzieLet33_1_argbuf_bufchan_buf  :
                                                                           \writeCTf''''''''_f''''''''_Int_IntlizzieLet33_1_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf''''''''_f''''''''_Int_IntlizzieLet33_1_argbuf_bufchan_buf  <= {16'd0,
                                                                               1'd0};
    else
      if ((\writeCTf''''''''_f''''''''_Int_IntlizzieLet33_1_argbuf_rwb_r  && \writeCTf''''''''_f''''''''_Int_IntlizzieLet33_1_argbuf_bufchan_buf [0]))
        \writeCTf''''''''_f''''''''_Int_IntlizzieLet33_1_argbuf_bufchan_buf  <= {16'd0,
                                                                                 1'd0};
      else if (((! \writeCTf''''''''_f''''''''_Int_IntlizzieLet33_1_argbuf_rwb_r ) && (! \writeCTf''''''''_f''''''''_Int_IntlizzieLet33_1_argbuf_bufchan_buf [0])))
        \writeCTf''''''''_f''''''''_Int_IntlizzieLet33_1_argbuf_bufchan_buf  <= \writeCTf''''''''_f''''''''_Int_IntlizzieLet33_1_argbuf_bufchan_d ;
  
  /* buf (Ty Pointer_CTf''''''''_f''''''''_Int_Int) : (writeCTf''''''''_f''''''''_Int_IntlizzieLet33_1_argbuf_rwb,Pointer_CTf''''''''_f''''''''_Int_Int) > (lizzieLet5_1_1_argbuf,Pointer_CTf''''''''_f''''''''_Int_Int) */
  \Pointer_CTf''''''''_f''''''''_Int_Int_t  \writeCTf''''''''_f''''''''_Int_IntlizzieLet33_1_argbuf_rwb_bufchan_d ;
  logic \writeCTf''''''''_f''''''''_Int_IntlizzieLet33_1_argbuf_rwb_bufchan_r ;
  assign \writeCTf''''''''_f''''''''_Int_IntlizzieLet33_1_argbuf_rwb_r  = ((! \writeCTf''''''''_f''''''''_Int_IntlizzieLet33_1_argbuf_rwb_bufchan_d [0]) || \writeCTf''''''''_f''''''''_Int_IntlizzieLet33_1_argbuf_rwb_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf''''''''_f''''''''_Int_IntlizzieLet33_1_argbuf_rwb_bufchan_d  <= {16'd0,
                                                                                 1'd0};
    else
      if (\writeCTf''''''''_f''''''''_Int_IntlizzieLet33_1_argbuf_rwb_r )
        \writeCTf''''''''_f''''''''_Int_IntlizzieLet33_1_argbuf_rwb_bufchan_d  <= \writeCTf''''''''_f''''''''_Int_IntlizzieLet33_1_argbuf_rwb_d ;
  \Pointer_CTf''''''''_f''''''''_Int_Int_t  \writeCTf''''''''_f''''''''_Int_IntlizzieLet33_1_argbuf_rwb_bufchan_buf ;
  assign \writeCTf''''''''_f''''''''_Int_IntlizzieLet33_1_argbuf_rwb_bufchan_r  = (! \writeCTf''''''''_f''''''''_Int_IntlizzieLet33_1_argbuf_rwb_bufchan_buf [0]);
  assign lizzieLet5_1_1_argbuf_d = (\writeCTf''''''''_f''''''''_Int_IntlizzieLet33_1_argbuf_rwb_bufchan_buf [0] ? \writeCTf''''''''_f''''''''_Int_IntlizzieLet33_1_argbuf_rwb_bufchan_buf  :
                                    \writeCTf''''''''_f''''''''_Int_IntlizzieLet33_1_argbuf_rwb_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf''''''''_f''''''''_Int_IntlizzieLet33_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                                   1'd0};
    else
      if ((lizzieLet5_1_1_argbuf_r && \writeCTf''''''''_f''''''''_Int_IntlizzieLet33_1_argbuf_rwb_bufchan_buf [0]))
        \writeCTf''''''''_f''''''''_Int_IntlizzieLet33_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                                     1'd0};
      else if (((! lizzieLet5_1_1_argbuf_r) && (! \writeCTf''''''''_f''''''''_Int_IntlizzieLet33_1_argbuf_rwb_bufchan_buf [0])))
        \writeCTf''''''''_f''''''''_Int_IntlizzieLet33_1_argbuf_rwb_bufchan_buf  <= \writeCTf''''''''_f''''''''_Int_IntlizzieLet33_1_argbuf_rwb_bufchan_d ;
  
  /* buf (Ty Pointer_CTf''''''''_f''''''''_Int_Int) : (writeCTf''''''''_f''''''''_Int_IntlizzieLet40_1_argbuf,Pointer_CTf''''''''_f''''''''_Int_Int) > (writeCTf''''''''_f''''''''_Int_IntlizzieLet40_1_argbuf_rwb,Pointer_CTf''''''''_f''''''''_Int_Int) */
  \Pointer_CTf''''''''_f''''''''_Int_Int_t  \writeCTf''''''''_f''''''''_Int_IntlizzieLet40_1_argbuf_bufchan_d ;
  logic \writeCTf''''''''_f''''''''_Int_IntlizzieLet40_1_argbuf_bufchan_r ;
  assign \writeCTf''''''''_f''''''''_Int_IntlizzieLet40_1_argbuf_r  = ((! \writeCTf''''''''_f''''''''_Int_IntlizzieLet40_1_argbuf_bufchan_d [0]) || \writeCTf''''''''_f''''''''_Int_IntlizzieLet40_1_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf''''''''_f''''''''_Int_IntlizzieLet40_1_argbuf_bufchan_d  <= {16'd0,
                                                                             1'd0};
    else
      if (\writeCTf''''''''_f''''''''_Int_IntlizzieLet40_1_argbuf_r )
        \writeCTf''''''''_f''''''''_Int_IntlizzieLet40_1_argbuf_bufchan_d  <= \writeCTf''''''''_f''''''''_Int_IntlizzieLet40_1_argbuf_d ;
  \Pointer_CTf''''''''_f''''''''_Int_Int_t  \writeCTf''''''''_f''''''''_Int_IntlizzieLet40_1_argbuf_bufchan_buf ;
  assign \writeCTf''''''''_f''''''''_Int_IntlizzieLet40_1_argbuf_bufchan_r  = (! \writeCTf''''''''_f''''''''_Int_IntlizzieLet40_1_argbuf_bufchan_buf [0]);
  assign \writeCTf''''''''_f''''''''_Int_IntlizzieLet40_1_argbuf_rwb_d  = (\writeCTf''''''''_f''''''''_Int_IntlizzieLet40_1_argbuf_bufchan_buf [0] ? \writeCTf''''''''_f''''''''_Int_IntlizzieLet40_1_argbuf_bufchan_buf  :
                                                                           \writeCTf''''''''_f''''''''_Int_IntlizzieLet40_1_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf''''''''_f''''''''_Int_IntlizzieLet40_1_argbuf_bufchan_buf  <= {16'd0,
                                                                               1'd0};
    else
      if ((\writeCTf''''''''_f''''''''_Int_IntlizzieLet40_1_argbuf_rwb_r  && \writeCTf''''''''_f''''''''_Int_IntlizzieLet40_1_argbuf_bufchan_buf [0]))
        \writeCTf''''''''_f''''''''_Int_IntlizzieLet40_1_argbuf_bufchan_buf  <= {16'd0,
                                                                                 1'd0};
      else if (((! \writeCTf''''''''_f''''''''_Int_IntlizzieLet40_1_argbuf_rwb_r ) && (! \writeCTf''''''''_f''''''''_Int_IntlizzieLet40_1_argbuf_bufchan_buf [0])))
        \writeCTf''''''''_f''''''''_Int_IntlizzieLet40_1_argbuf_bufchan_buf  <= \writeCTf''''''''_f''''''''_Int_IntlizzieLet40_1_argbuf_bufchan_d ;
  
  /* buf (Ty Pointer_CTf''''''''_f''''''''_Int_Int) : (writeCTf''''''''_f''''''''_Int_IntlizzieLet40_1_argbuf_rwb,Pointer_CTf''''''''_f''''''''_Int_Int) > (sca2_1_1_argbuf,Pointer_CTf''''''''_f''''''''_Int_Int) */
  \Pointer_CTf''''''''_f''''''''_Int_Int_t  \writeCTf''''''''_f''''''''_Int_IntlizzieLet40_1_argbuf_rwb_bufchan_d ;
  logic \writeCTf''''''''_f''''''''_Int_IntlizzieLet40_1_argbuf_rwb_bufchan_r ;
  assign \writeCTf''''''''_f''''''''_Int_IntlizzieLet40_1_argbuf_rwb_r  = ((! \writeCTf''''''''_f''''''''_Int_IntlizzieLet40_1_argbuf_rwb_bufchan_d [0]) || \writeCTf''''''''_f''''''''_Int_IntlizzieLet40_1_argbuf_rwb_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf''''''''_f''''''''_Int_IntlizzieLet40_1_argbuf_rwb_bufchan_d  <= {16'd0,
                                                                                 1'd0};
    else
      if (\writeCTf''''''''_f''''''''_Int_IntlizzieLet40_1_argbuf_rwb_r )
        \writeCTf''''''''_f''''''''_Int_IntlizzieLet40_1_argbuf_rwb_bufchan_d  <= \writeCTf''''''''_f''''''''_Int_IntlizzieLet40_1_argbuf_rwb_d ;
  \Pointer_CTf''''''''_f''''''''_Int_Int_t  \writeCTf''''''''_f''''''''_Int_IntlizzieLet40_1_argbuf_rwb_bufchan_buf ;
  assign \writeCTf''''''''_f''''''''_Int_IntlizzieLet40_1_argbuf_rwb_bufchan_r  = (! \writeCTf''''''''_f''''''''_Int_IntlizzieLet40_1_argbuf_rwb_bufchan_buf [0]);
  assign sca2_1_1_argbuf_d = (\writeCTf''''''''_f''''''''_Int_IntlizzieLet40_1_argbuf_rwb_bufchan_buf [0] ? \writeCTf''''''''_f''''''''_Int_IntlizzieLet40_1_argbuf_rwb_bufchan_buf  :
                              \writeCTf''''''''_f''''''''_Int_IntlizzieLet40_1_argbuf_rwb_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf''''''''_f''''''''_Int_IntlizzieLet40_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                                   1'd0};
    else
      if ((sca2_1_1_argbuf_r && \writeCTf''''''''_f''''''''_Int_IntlizzieLet40_1_argbuf_rwb_bufchan_buf [0]))
        \writeCTf''''''''_f''''''''_Int_IntlizzieLet40_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                                     1'd0};
      else if (((! sca2_1_1_argbuf_r) && (! \writeCTf''''''''_f''''''''_Int_IntlizzieLet40_1_argbuf_rwb_bufchan_buf [0])))
        \writeCTf''''''''_f''''''''_Int_IntlizzieLet40_1_argbuf_rwb_bufchan_buf  <= \writeCTf''''''''_f''''''''_Int_IntlizzieLet40_1_argbuf_rwb_bufchan_d ;
  
  /* buf (Ty Pointer_CTf''''''''_f''''''''_Int_Int) : (writeCTf''''''''_f''''''''_Int_IntlizzieLet41_1_argbuf,Pointer_CTf''''''''_f''''''''_Int_Int) > (writeCTf''''''''_f''''''''_Int_IntlizzieLet41_1_argbuf_rwb,Pointer_CTf''''''''_f''''''''_Int_Int) */
  \Pointer_CTf''''''''_f''''''''_Int_Int_t  \writeCTf''''''''_f''''''''_Int_IntlizzieLet41_1_argbuf_bufchan_d ;
  logic \writeCTf''''''''_f''''''''_Int_IntlizzieLet41_1_argbuf_bufchan_r ;
  assign \writeCTf''''''''_f''''''''_Int_IntlizzieLet41_1_argbuf_r  = ((! \writeCTf''''''''_f''''''''_Int_IntlizzieLet41_1_argbuf_bufchan_d [0]) || \writeCTf''''''''_f''''''''_Int_IntlizzieLet41_1_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf''''''''_f''''''''_Int_IntlizzieLet41_1_argbuf_bufchan_d  <= {16'd0,
                                                                             1'd0};
    else
      if (\writeCTf''''''''_f''''''''_Int_IntlizzieLet41_1_argbuf_r )
        \writeCTf''''''''_f''''''''_Int_IntlizzieLet41_1_argbuf_bufchan_d  <= \writeCTf''''''''_f''''''''_Int_IntlizzieLet41_1_argbuf_d ;
  \Pointer_CTf''''''''_f''''''''_Int_Int_t  \writeCTf''''''''_f''''''''_Int_IntlizzieLet41_1_argbuf_bufchan_buf ;
  assign \writeCTf''''''''_f''''''''_Int_IntlizzieLet41_1_argbuf_bufchan_r  = (! \writeCTf''''''''_f''''''''_Int_IntlizzieLet41_1_argbuf_bufchan_buf [0]);
  assign \writeCTf''''''''_f''''''''_Int_IntlizzieLet41_1_argbuf_rwb_d  = (\writeCTf''''''''_f''''''''_Int_IntlizzieLet41_1_argbuf_bufchan_buf [0] ? \writeCTf''''''''_f''''''''_Int_IntlizzieLet41_1_argbuf_bufchan_buf  :
                                                                           \writeCTf''''''''_f''''''''_Int_IntlizzieLet41_1_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf''''''''_f''''''''_Int_IntlizzieLet41_1_argbuf_bufchan_buf  <= {16'd0,
                                                                               1'd0};
    else
      if ((\writeCTf''''''''_f''''''''_Int_IntlizzieLet41_1_argbuf_rwb_r  && \writeCTf''''''''_f''''''''_Int_IntlizzieLet41_1_argbuf_bufchan_buf [0]))
        \writeCTf''''''''_f''''''''_Int_IntlizzieLet41_1_argbuf_bufchan_buf  <= {16'd0,
                                                                                 1'd0};
      else if (((! \writeCTf''''''''_f''''''''_Int_IntlizzieLet41_1_argbuf_rwb_r ) && (! \writeCTf''''''''_f''''''''_Int_IntlizzieLet41_1_argbuf_bufchan_buf [0])))
        \writeCTf''''''''_f''''''''_Int_IntlizzieLet41_1_argbuf_bufchan_buf  <= \writeCTf''''''''_f''''''''_Int_IntlizzieLet41_1_argbuf_bufchan_d ;
  
  /* buf (Ty Pointer_CTf''''''''_f''''''''_Int_Int) : (writeCTf''''''''_f''''''''_Int_IntlizzieLet41_1_argbuf_rwb,Pointer_CTf''''''''_f''''''''_Int_Int) > (sca1_1_1_argbuf,Pointer_CTf''''''''_f''''''''_Int_Int) */
  \Pointer_CTf''''''''_f''''''''_Int_Int_t  \writeCTf''''''''_f''''''''_Int_IntlizzieLet41_1_argbuf_rwb_bufchan_d ;
  logic \writeCTf''''''''_f''''''''_Int_IntlizzieLet41_1_argbuf_rwb_bufchan_r ;
  assign \writeCTf''''''''_f''''''''_Int_IntlizzieLet41_1_argbuf_rwb_r  = ((! \writeCTf''''''''_f''''''''_Int_IntlizzieLet41_1_argbuf_rwb_bufchan_d [0]) || \writeCTf''''''''_f''''''''_Int_IntlizzieLet41_1_argbuf_rwb_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf''''''''_f''''''''_Int_IntlizzieLet41_1_argbuf_rwb_bufchan_d  <= {16'd0,
                                                                                 1'd0};
    else
      if (\writeCTf''''''''_f''''''''_Int_IntlizzieLet41_1_argbuf_rwb_r )
        \writeCTf''''''''_f''''''''_Int_IntlizzieLet41_1_argbuf_rwb_bufchan_d  <= \writeCTf''''''''_f''''''''_Int_IntlizzieLet41_1_argbuf_rwb_d ;
  \Pointer_CTf''''''''_f''''''''_Int_Int_t  \writeCTf''''''''_f''''''''_Int_IntlizzieLet41_1_argbuf_rwb_bufchan_buf ;
  assign \writeCTf''''''''_f''''''''_Int_IntlizzieLet41_1_argbuf_rwb_bufchan_r  = (! \writeCTf''''''''_f''''''''_Int_IntlizzieLet41_1_argbuf_rwb_bufchan_buf [0]);
  assign sca1_1_1_argbuf_d = (\writeCTf''''''''_f''''''''_Int_IntlizzieLet41_1_argbuf_rwb_bufchan_buf [0] ? \writeCTf''''''''_f''''''''_Int_IntlizzieLet41_1_argbuf_rwb_bufchan_buf  :
                              \writeCTf''''''''_f''''''''_Int_IntlizzieLet41_1_argbuf_rwb_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf''''''''_f''''''''_Int_IntlizzieLet41_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                                   1'd0};
    else
      if ((sca1_1_1_argbuf_r && \writeCTf''''''''_f''''''''_Int_IntlizzieLet41_1_argbuf_rwb_bufchan_buf [0]))
        \writeCTf''''''''_f''''''''_Int_IntlizzieLet41_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                                     1'd0};
      else if (((! sca1_1_1_argbuf_r) && (! \writeCTf''''''''_f''''''''_Int_IntlizzieLet41_1_argbuf_rwb_bufchan_buf [0])))
        \writeCTf''''''''_f''''''''_Int_IntlizzieLet41_1_argbuf_rwb_bufchan_buf  <= \writeCTf''''''''_f''''''''_Int_IntlizzieLet41_1_argbuf_rwb_bufchan_d ;
  
  /* buf (Ty Pointer_CTf''''''''_f''''''''_Int_Int) : (writeCTf''''''''_f''''''''_Int_IntlizzieLet42_1_argbuf,Pointer_CTf''''''''_f''''''''_Int_Int) > (writeCTf''''''''_f''''''''_Int_IntlizzieLet42_1_argbuf_rwb,Pointer_CTf''''''''_f''''''''_Int_Int) */
  \Pointer_CTf''''''''_f''''''''_Int_Int_t  \writeCTf''''''''_f''''''''_Int_IntlizzieLet42_1_argbuf_bufchan_d ;
  logic \writeCTf''''''''_f''''''''_Int_IntlizzieLet42_1_argbuf_bufchan_r ;
  assign \writeCTf''''''''_f''''''''_Int_IntlizzieLet42_1_argbuf_r  = ((! \writeCTf''''''''_f''''''''_Int_IntlizzieLet42_1_argbuf_bufchan_d [0]) || \writeCTf''''''''_f''''''''_Int_IntlizzieLet42_1_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf''''''''_f''''''''_Int_IntlizzieLet42_1_argbuf_bufchan_d  <= {16'd0,
                                                                             1'd0};
    else
      if (\writeCTf''''''''_f''''''''_Int_IntlizzieLet42_1_argbuf_r )
        \writeCTf''''''''_f''''''''_Int_IntlizzieLet42_1_argbuf_bufchan_d  <= \writeCTf''''''''_f''''''''_Int_IntlizzieLet42_1_argbuf_d ;
  \Pointer_CTf''''''''_f''''''''_Int_Int_t  \writeCTf''''''''_f''''''''_Int_IntlizzieLet42_1_argbuf_bufchan_buf ;
  assign \writeCTf''''''''_f''''''''_Int_IntlizzieLet42_1_argbuf_bufchan_r  = (! \writeCTf''''''''_f''''''''_Int_IntlizzieLet42_1_argbuf_bufchan_buf [0]);
  assign \writeCTf''''''''_f''''''''_Int_IntlizzieLet42_1_argbuf_rwb_d  = (\writeCTf''''''''_f''''''''_Int_IntlizzieLet42_1_argbuf_bufchan_buf [0] ? \writeCTf''''''''_f''''''''_Int_IntlizzieLet42_1_argbuf_bufchan_buf  :
                                                                           \writeCTf''''''''_f''''''''_Int_IntlizzieLet42_1_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf''''''''_f''''''''_Int_IntlizzieLet42_1_argbuf_bufchan_buf  <= {16'd0,
                                                                               1'd0};
    else
      if ((\writeCTf''''''''_f''''''''_Int_IntlizzieLet42_1_argbuf_rwb_r  && \writeCTf''''''''_f''''''''_Int_IntlizzieLet42_1_argbuf_bufchan_buf [0]))
        \writeCTf''''''''_f''''''''_Int_IntlizzieLet42_1_argbuf_bufchan_buf  <= {16'd0,
                                                                                 1'd0};
      else if (((! \writeCTf''''''''_f''''''''_Int_IntlizzieLet42_1_argbuf_rwb_r ) && (! \writeCTf''''''''_f''''''''_Int_IntlizzieLet42_1_argbuf_bufchan_buf [0])))
        \writeCTf''''''''_f''''''''_Int_IntlizzieLet42_1_argbuf_bufchan_buf  <= \writeCTf''''''''_f''''''''_Int_IntlizzieLet42_1_argbuf_bufchan_d ;
  
  /* buf (Ty Pointer_CTf''''''''_f''''''''_Int_Int) : (writeCTf''''''''_f''''''''_Int_IntlizzieLet42_1_argbuf_rwb,Pointer_CTf''''''''_f''''''''_Int_Int) > (sca0_1_1_argbuf,Pointer_CTf''''''''_f''''''''_Int_Int) */
  \Pointer_CTf''''''''_f''''''''_Int_Int_t  \writeCTf''''''''_f''''''''_Int_IntlizzieLet42_1_argbuf_rwb_bufchan_d ;
  logic \writeCTf''''''''_f''''''''_Int_IntlizzieLet42_1_argbuf_rwb_bufchan_r ;
  assign \writeCTf''''''''_f''''''''_Int_IntlizzieLet42_1_argbuf_rwb_r  = ((! \writeCTf''''''''_f''''''''_Int_IntlizzieLet42_1_argbuf_rwb_bufchan_d [0]) || \writeCTf''''''''_f''''''''_Int_IntlizzieLet42_1_argbuf_rwb_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf''''''''_f''''''''_Int_IntlizzieLet42_1_argbuf_rwb_bufchan_d  <= {16'd0,
                                                                                 1'd0};
    else
      if (\writeCTf''''''''_f''''''''_Int_IntlizzieLet42_1_argbuf_rwb_r )
        \writeCTf''''''''_f''''''''_Int_IntlizzieLet42_1_argbuf_rwb_bufchan_d  <= \writeCTf''''''''_f''''''''_Int_IntlizzieLet42_1_argbuf_rwb_d ;
  \Pointer_CTf''''''''_f''''''''_Int_Int_t  \writeCTf''''''''_f''''''''_Int_IntlizzieLet42_1_argbuf_rwb_bufchan_buf ;
  assign \writeCTf''''''''_f''''''''_Int_IntlizzieLet42_1_argbuf_rwb_bufchan_r  = (! \writeCTf''''''''_f''''''''_Int_IntlizzieLet42_1_argbuf_rwb_bufchan_buf [0]);
  assign sca0_1_1_argbuf_d = (\writeCTf''''''''_f''''''''_Int_IntlizzieLet42_1_argbuf_rwb_bufchan_buf [0] ? \writeCTf''''''''_f''''''''_Int_IntlizzieLet42_1_argbuf_rwb_bufchan_buf  :
                              \writeCTf''''''''_f''''''''_Int_IntlizzieLet42_1_argbuf_rwb_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf''''''''_f''''''''_Int_IntlizzieLet42_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                                   1'd0};
    else
      if ((sca0_1_1_argbuf_r && \writeCTf''''''''_f''''''''_Int_IntlizzieLet42_1_argbuf_rwb_bufchan_buf [0]))
        \writeCTf''''''''_f''''''''_Int_IntlizzieLet42_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                                     1'd0};
      else if (((! sca0_1_1_argbuf_r) && (! \writeCTf''''''''_f''''''''_Int_IntlizzieLet42_1_argbuf_rwb_bufchan_buf [0])))
        \writeCTf''''''''_f''''''''_Int_IntlizzieLet42_1_argbuf_rwb_bufchan_buf  <= \writeCTf''''''''_f''''''''_Int_IntlizzieLet42_1_argbuf_rwb_bufchan_d ;
  
  /* buf (Ty Pointer_CTf_f_Int_Int) : (writeCTf_f_Int_IntlizzieLet30_1_argbuf,Pointer_CTf_f_Int_Int) > (writeCTf_f_Int_IntlizzieLet30_1_argbuf_rwb,Pointer_CTf_f_Int_Int) */
  Pointer_CTf_f_Int_Int_t writeCTf_f_Int_IntlizzieLet30_1_argbuf_bufchan_d;
  logic writeCTf_f_Int_IntlizzieLet30_1_argbuf_bufchan_r;
  assign writeCTf_f_Int_IntlizzieLet30_1_argbuf_r = ((! writeCTf_f_Int_IntlizzieLet30_1_argbuf_bufchan_d[0]) || writeCTf_f_Int_IntlizzieLet30_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTf_f_Int_IntlizzieLet30_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCTf_f_Int_IntlizzieLet30_1_argbuf_r)
        writeCTf_f_Int_IntlizzieLet30_1_argbuf_bufchan_d <= writeCTf_f_Int_IntlizzieLet30_1_argbuf_d;
  Pointer_CTf_f_Int_Int_t writeCTf_f_Int_IntlizzieLet30_1_argbuf_bufchan_buf;
  assign writeCTf_f_Int_IntlizzieLet30_1_argbuf_bufchan_r = (! writeCTf_f_Int_IntlizzieLet30_1_argbuf_bufchan_buf[0]);
  assign writeCTf_f_Int_IntlizzieLet30_1_argbuf_rwb_d = (writeCTf_f_Int_IntlizzieLet30_1_argbuf_bufchan_buf[0] ? writeCTf_f_Int_IntlizzieLet30_1_argbuf_bufchan_buf :
                                                         writeCTf_f_Int_IntlizzieLet30_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTf_f_Int_IntlizzieLet30_1_argbuf_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((writeCTf_f_Int_IntlizzieLet30_1_argbuf_rwb_r && writeCTf_f_Int_IntlizzieLet30_1_argbuf_bufchan_buf[0]))
        writeCTf_f_Int_IntlizzieLet30_1_argbuf_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! writeCTf_f_Int_IntlizzieLet30_1_argbuf_rwb_r) && (! writeCTf_f_Int_IntlizzieLet30_1_argbuf_bufchan_buf[0])))
        writeCTf_f_Int_IntlizzieLet30_1_argbuf_bufchan_buf <= writeCTf_f_Int_IntlizzieLet30_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CTf_f_Int_Int) : (writeCTf_f_Int_IntlizzieLet30_1_argbuf_rwb,Pointer_CTf_f_Int_Int) > (sca3_2_1_argbuf,Pointer_CTf_f_Int_Int) */
  Pointer_CTf_f_Int_Int_t writeCTf_f_Int_IntlizzieLet30_1_argbuf_rwb_bufchan_d;
  logic writeCTf_f_Int_IntlizzieLet30_1_argbuf_rwb_bufchan_r;
  assign writeCTf_f_Int_IntlizzieLet30_1_argbuf_rwb_r = ((! writeCTf_f_Int_IntlizzieLet30_1_argbuf_rwb_bufchan_d[0]) || writeCTf_f_Int_IntlizzieLet30_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTf_f_Int_IntlizzieLet30_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                               1'd0};
    else
      if (writeCTf_f_Int_IntlizzieLet30_1_argbuf_rwb_r)
        writeCTf_f_Int_IntlizzieLet30_1_argbuf_rwb_bufchan_d <= writeCTf_f_Int_IntlizzieLet30_1_argbuf_rwb_d;
  Pointer_CTf_f_Int_Int_t writeCTf_f_Int_IntlizzieLet30_1_argbuf_rwb_bufchan_buf;
  assign writeCTf_f_Int_IntlizzieLet30_1_argbuf_rwb_bufchan_r = (! writeCTf_f_Int_IntlizzieLet30_1_argbuf_rwb_bufchan_buf[0]);
  assign sca3_2_1_argbuf_d = (writeCTf_f_Int_IntlizzieLet30_1_argbuf_rwb_bufchan_buf[0] ? writeCTf_f_Int_IntlizzieLet30_1_argbuf_rwb_bufchan_buf :
                              writeCTf_f_Int_IntlizzieLet30_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTf_f_Int_IntlizzieLet30_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                 1'd0};
    else
      if ((sca3_2_1_argbuf_r && writeCTf_f_Int_IntlizzieLet30_1_argbuf_rwb_bufchan_buf[0]))
        writeCTf_f_Int_IntlizzieLet30_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                   1'd0};
      else if (((! sca3_2_1_argbuf_r) && (! writeCTf_f_Int_IntlizzieLet30_1_argbuf_rwb_bufchan_buf[0])))
        writeCTf_f_Int_IntlizzieLet30_1_argbuf_rwb_bufchan_buf <= writeCTf_f_Int_IntlizzieLet30_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CTf_f_Int_Int) : (writeCTf_f_Int_IntlizzieLet34_1_argbuf,Pointer_CTf_f_Int_Int) > (writeCTf_f_Int_IntlizzieLet34_1_argbuf_rwb,Pointer_CTf_f_Int_Int) */
  Pointer_CTf_f_Int_Int_t writeCTf_f_Int_IntlizzieLet34_1_argbuf_bufchan_d;
  logic writeCTf_f_Int_IntlizzieLet34_1_argbuf_bufchan_r;
  assign writeCTf_f_Int_IntlizzieLet34_1_argbuf_r = ((! writeCTf_f_Int_IntlizzieLet34_1_argbuf_bufchan_d[0]) || writeCTf_f_Int_IntlizzieLet34_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTf_f_Int_IntlizzieLet34_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCTf_f_Int_IntlizzieLet34_1_argbuf_r)
        writeCTf_f_Int_IntlizzieLet34_1_argbuf_bufchan_d <= writeCTf_f_Int_IntlizzieLet34_1_argbuf_d;
  Pointer_CTf_f_Int_Int_t writeCTf_f_Int_IntlizzieLet34_1_argbuf_bufchan_buf;
  assign writeCTf_f_Int_IntlizzieLet34_1_argbuf_bufchan_r = (! writeCTf_f_Int_IntlizzieLet34_1_argbuf_bufchan_buf[0]);
  assign writeCTf_f_Int_IntlizzieLet34_1_argbuf_rwb_d = (writeCTf_f_Int_IntlizzieLet34_1_argbuf_bufchan_buf[0] ? writeCTf_f_Int_IntlizzieLet34_1_argbuf_bufchan_buf :
                                                         writeCTf_f_Int_IntlizzieLet34_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTf_f_Int_IntlizzieLet34_1_argbuf_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((writeCTf_f_Int_IntlizzieLet34_1_argbuf_rwb_r && writeCTf_f_Int_IntlizzieLet34_1_argbuf_bufchan_buf[0]))
        writeCTf_f_Int_IntlizzieLet34_1_argbuf_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! writeCTf_f_Int_IntlizzieLet34_1_argbuf_rwb_r) && (! writeCTf_f_Int_IntlizzieLet34_1_argbuf_bufchan_buf[0])))
        writeCTf_f_Int_IntlizzieLet34_1_argbuf_bufchan_buf <= writeCTf_f_Int_IntlizzieLet34_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CTf_f_Int_Int) : (writeCTf_f_Int_IntlizzieLet34_1_argbuf_rwb,Pointer_CTf_f_Int_Int) > (lizzieLet22_1_1_argbuf,Pointer_CTf_f_Int_Int) */
  Pointer_CTf_f_Int_Int_t writeCTf_f_Int_IntlizzieLet34_1_argbuf_rwb_bufchan_d;
  logic writeCTf_f_Int_IntlizzieLet34_1_argbuf_rwb_bufchan_r;
  assign writeCTf_f_Int_IntlizzieLet34_1_argbuf_rwb_r = ((! writeCTf_f_Int_IntlizzieLet34_1_argbuf_rwb_bufchan_d[0]) || writeCTf_f_Int_IntlizzieLet34_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTf_f_Int_IntlizzieLet34_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                               1'd0};
    else
      if (writeCTf_f_Int_IntlizzieLet34_1_argbuf_rwb_r)
        writeCTf_f_Int_IntlizzieLet34_1_argbuf_rwb_bufchan_d <= writeCTf_f_Int_IntlizzieLet34_1_argbuf_rwb_d;
  Pointer_CTf_f_Int_Int_t writeCTf_f_Int_IntlizzieLet34_1_argbuf_rwb_bufchan_buf;
  assign writeCTf_f_Int_IntlizzieLet34_1_argbuf_rwb_bufchan_r = (! writeCTf_f_Int_IntlizzieLet34_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet22_1_1_argbuf_d = (writeCTf_f_Int_IntlizzieLet34_1_argbuf_rwb_bufchan_buf[0] ? writeCTf_f_Int_IntlizzieLet34_1_argbuf_rwb_bufchan_buf :
                                     writeCTf_f_Int_IntlizzieLet34_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTf_f_Int_IntlizzieLet34_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                 1'd0};
    else
      if ((lizzieLet22_1_1_argbuf_r && writeCTf_f_Int_IntlizzieLet34_1_argbuf_rwb_bufchan_buf[0]))
        writeCTf_f_Int_IntlizzieLet34_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                   1'd0};
      else if (((! lizzieLet22_1_1_argbuf_r) && (! writeCTf_f_Int_IntlizzieLet34_1_argbuf_rwb_bufchan_buf[0])))
        writeCTf_f_Int_IntlizzieLet34_1_argbuf_rwb_bufchan_buf <= writeCTf_f_Int_IntlizzieLet34_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CTf_f_Int_Int) : (writeCTf_f_Int_IntlizzieLet45_1_argbuf,Pointer_CTf_f_Int_Int) > (writeCTf_f_Int_IntlizzieLet45_1_argbuf_rwb,Pointer_CTf_f_Int_Int) */
  Pointer_CTf_f_Int_Int_t writeCTf_f_Int_IntlizzieLet45_1_argbuf_bufchan_d;
  logic writeCTf_f_Int_IntlizzieLet45_1_argbuf_bufchan_r;
  assign writeCTf_f_Int_IntlizzieLet45_1_argbuf_r = ((! writeCTf_f_Int_IntlizzieLet45_1_argbuf_bufchan_d[0]) || writeCTf_f_Int_IntlizzieLet45_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTf_f_Int_IntlizzieLet45_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCTf_f_Int_IntlizzieLet45_1_argbuf_r)
        writeCTf_f_Int_IntlizzieLet45_1_argbuf_bufchan_d <= writeCTf_f_Int_IntlizzieLet45_1_argbuf_d;
  Pointer_CTf_f_Int_Int_t writeCTf_f_Int_IntlizzieLet45_1_argbuf_bufchan_buf;
  assign writeCTf_f_Int_IntlizzieLet45_1_argbuf_bufchan_r = (! writeCTf_f_Int_IntlizzieLet45_1_argbuf_bufchan_buf[0]);
  assign writeCTf_f_Int_IntlizzieLet45_1_argbuf_rwb_d = (writeCTf_f_Int_IntlizzieLet45_1_argbuf_bufchan_buf[0] ? writeCTf_f_Int_IntlizzieLet45_1_argbuf_bufchan_buf :
                                                         writeCTf_f_Int_IntlizzieLet45_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTf_f_Int_IntlizzieLet45_1_argbuf_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((writeCTf_f_Int_IntlizzieLet45_1_argbuf_rwb_r && writeCTf_f_Int_IntlizzieLet45_1_argbuf_bufchan_buf[0]))
        writeCTf_f_Int_IntlizzieLet45_1_argbuf_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! writeCTf_f_Int_IntlizzieLet45_1_argbuf_rwb_r) && (! writeCTf_f_Int_IntlizzieLet45_1_argbuf_bufchan_buf[0])))
        writeCTf_f_Int_IntlizzieLet45_1_argbuf_bufchan_buf <= writeCTf_f_Int_IntlizzieLet45_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CTf_f_Int_Int) : (writeCTf_f_Int_IntlizzieLet45_1_argbuf_rwb,Pointer_CTf_f_Int_Int) > (sca2_2_1_argbuf,Pointer_CTf_f_Int_Int) */
  Pointer_CTf_f_Int_Int_t writeCTf_f_Int_IntlizzieLet45_1_argbuf_rwb_bufchan_d;
  logic writeCTf_f_Int_IntlizzieLet45_1_argbuf_rwb_bufchan_r;
  assign writeCTf_f_Int_IntlizzieLet45_1_argbuf_rwb_r = ((! writeCTf_f_Int_IntlizzieLet45_1_argbuf_rwb_bufchan_d[0]) || writeCTf_f_Int_IntlizzieLet45_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTf_f_Int_IntlizzieLet45_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                               1'd0};
    else
      if (writeCTf_f_Int_IntlizzieLet45_1_argbuf_rwb_r)
        writeCTf_f_Int_IntlizzieLet45_1_argbuf_rwb_bufchan_d <= writeCTf_f_Int_IntlizzieLet45_1_argbuf_rwb_d;
  Pointer_CTf_f_Int_Int_t writeCTf_f_Int_IntlizzieLet45_1_argbuf_rwb_bufchan_buf;
  assign writeCTf_f_Int_IntlizzieLet45_1_argbuf_rwb_bufchan_r = (! writeCTf_f_Int_IntlizzieLet45_1_argbuf_rwb_bufchan_buf[0]);
  assign sca2_2_1_argbuf_d = (writeCTf_f_Int_IntlizzieLet45_1_argbuf_rwb_bufchan_buf[0] ? writeCTf_f_Int_IntlizzieLet45_1_argbuf_rwb_bufchan_buf :
                              writeCTf_f_Int_IntlizzieLet45_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTf_f_Int_IntlizzieLet45_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                 1'd0};
    else
      if ((sca2_2_1_argbuf_r && writeCTf_f_Int_IntlizzieLet45_1_argbuf_rwb_bufchan_buf[0]))
        writeCTf_f_Int_IntlizzieLet45_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                   1'd0};
      else if (((! sca2_2_1_argbuf_r) && (! writeCTf_f_Int_IntlizzieLet45_1_argbuf_rwb_bufchan_buf[0])))
        writeCTf_f_Int_IntlizzieLet45_1_argbuf_rwb_bufchan_buf <= writeCTf_f_Int_IntlizzieLet45_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CTf_f_Int_Int) : (writeCTf_f_Int_IntlizzieLet46_1_argbuf,Pointer_CTf_f_Int_Int) > (writeCTf_f_Int_IntlizzieLet46_1_argbuf_rwb,Pointer_CTf_f_Int_Int) */
  Pointer_CTf_f_Int_Int_t writeCTf_f_Int_IntlizzieLet46_1_argbuf_bufchan_d;
  logic writeCTf_f_Int_IntlizzieLet46_1_argbuf_bufchan_r;
  assign writeCTf_f_Int_IntlizzieLet46_1_argbuf_r = ((! writeCTf_f_Int_IntlizzieLet46_1_argbuf_bufchan_d[0]) || writeCTf_f_Int_IntlizzieLet46_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTf_f_Int_IntlizzieLet46_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCTf_f_Int_IntlizzieLet46_1_argbuf_r)
        writeCTf_f_Int_IntlizzieLet46_1_argbuf_bufchan_d <= writeCTf_f_Int_IntlizzieLet46_1_argbuf_d;
  Pointer_CTf_f_Int_Int_t writeCTf_f_Int_IntlizzieLet46_1_argbuf_bufchan_buf;
  assign writeCTf_f_Int_IntlizzieLet46_1_argbuf_bufchan_r = (! writeCTf_f_Int_IntlizzieLet46_1_argbuf_bufchan_buf[0]);
  assign writeCTf_f_Int_IntlizzieLet46_1_argbuf_rwb_d = (writeCTf_f_Int_IntlizzieLet46_1_argbuf_bufchan_buf[0] ? writeCTf_f_Int_IntlizzieLet46_1_argbuf_bufchan_buf :
                                                         writeCTf_f_Int_IntlizzieLet46_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTf_f_Int_IntlizzieLet46_1_argbuf_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((writeCTf_f_Int_IntlizzieLet46_1_argbuf_rwb_r && writeCTf_f_Int_IntlizzieLet46_1_argbuf_bufchan_buf[0]))
        writeCTf_f_Int_IntlizzieLet46_1_argbuf_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! writeCTf_f_Int_IntlizzieLet46_1_argbuf_rwb_r) && (! writeCTf_f_Int_IntlizzieLet46_1_argbuf_bufchan_buf[0])))
        writeCTf_f_Int_IntlizzieLet46_1_argbuf_bufchan_buf <= writeCTf_f_Int_IntlizzieLet46_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CTf_f_Int_Int) : (writeCTf_f_Int_IntlizzieLet46_1_argbuf_rwb,Pointer_CTf_f_Int_Int) > (sca1_2_1_argbuf,Pointer_CTf_f_Int_Int) */
  Pointer_CTf_f_Int_Int_t writeCTf_f_Int_IntlizzieLet46_1_argbuf_rwb_bufchan_d;
  logic writeCTf_f_Int_IntlizzieLet46_1_argbuf_rwb_bufchan_r;
  assign writeCTf_f_Int_IntlizzieLet46_1_argbuf_rwb_r = ((! writeCTf_f_Int_IntlizzieLet46_1_argbuf_rwb_bufchan_d[0]) || writeCTf_f_Int_IntlizzieLet46_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTf_f_Int_IntlizzieLet46_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                               1'd0};
    else
      if (writeCTf_f_Int_IntlizzieLet46_1_argbuf_rwb_r)
        writeCTf_f_Int_IntlizzieLet46_1_argbuf_rwb_bufchan_d <= writeCTf_f_Int_IntlizzieLet46_1_argbuf_rwb_d;
  Pointer_CTf_f_Int_Int_t writeCTf_f_Int_IntlizzieLet46_1_argbuf_rwb_bufchan_buf;
  assign writeCTf_f_Int_IntlizzieLet46_1_argbuf_rwb_bufchan_r = (! writeCTf_f_Int_IntlizzieLet46_1_argbuf_rwb_bufchan_buf[0]);
  assign sca1_2_1_argbuf_d = (writeCTf_f_Int_IntlizzieLet46_1_argbuf_rwb_bufchan_buf[0] ? writeCTf_f_Int_IntlizzieLet46_1_argbuf_rwb_bufchan_buf :
                              writeCTf_f_Int_IntlizzieLet46_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTf_f_Int_IntlizzieLet46_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                 1'd0};
    else
      if ((sca1_2_1_argbuf_r && writeCTf_f_Int_IntlizzieLet46_1_argbuf_rwb_bufchan_buf[0]))
        writeCTf_f_Int_IntlizzieLet46_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                   1'd0};
      else if (((! sca1_2_1_argbuf_r) && (! writeCTf_f_Int_IntlizzieLet46_1_argbuf_rwb_bufchan_buf[0])))
        writeCTf_f_Int_IntlizzieLet46_1_argbuf_rwb_bufchan_buf <= writeCTf_f_Int_IntlizzieLet46_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CTf_f_Int_Int) : (writeCTf_f_Int_IntlizzieLet47_1_argbuf,Pointer_CTf_f_Int_Int) > (writeCTf_f_Int_IntlizzieLet47_1_argbuf_rwb,Pointer_CTf_f_Int_Int) */
  Pointer_CTf_f_Int_Int_t writeCTf_f_Int_IntlizzieLet47_1_argbuf_bufchan_d;
  logic writeCTf_f_Int_IntlizzieLet47_1_argbuf_bufchan_r;
  assign writeCTf_f_Int_IntlizzieLet47_1_argbuf_r = ((! writeCTf_f_Int_IntlizzieLet47_1_argbuf_bufchan_d[0]) || writeCTf_f_Int_IntlizzieLet47_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTf_f_Int_IntlizzieLet47_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCTf_f_Int_IntlizzieLet47_1_argbuf_r)
        writeCTf_f_Int_IntlizzieLet47_1_argbuf_bufchan_d <= writeCTf_f_Int_IntlizzieLet47_1_argbuf_d;
  Pointer_CTf_f_Int_Int_t writeCTf_f_Int_IntlizzieLet47_1_argbuf_bufchan_buf;
  assign writeCTf_f_Int_IntlizzieLet47_1_argbuf_bufchan_r = (! writeCTf_f_Int_IntlizzieLet47_1_argbuf_bufchan_buf[0]);
  assign writeCTf_f_Int_IntlizzieLet47_1_argbuf_rwb_d = (writeCTf_f_Int_IntlizzieLet47_1_argbuf_bufchan_buf[0] ? writeCTf_f_Int_IntlizzieLet47_1_argbuf_bufchan_buf :
                                                         writeCTf_f_Int_IntlizzieLet47_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTf_f_Int_IntlizzieLet47_1_argbuf_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((writeCTf_f_Int_IntlizzieLet47_1_argbuf_rwb_r && writeCTf_f_Int_IntlizzieLet47_1_argbuf_bufchan_buf[0]))
        writeCTf_f_Int_IntlizzieLet47_1_argbuf_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! writeCTf_f_Int_IntlizzieLet47_1_argbuf_rwb_r) && (! writeCTf_f_Int_IntlizzieLet47_1_argbuf_bufchan_buf[0])))
        writeCTf_f_Int_IntlizzieLet47_1_argbuf_bufchan_buf <= writeCTf_f_Int_IntlizzieLet47_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CTf_f_Int_Int) : (writeCTf_f_Int_IntlizzieLet47_1_argbuf_rwb,Pointer_CTf_f_Int_Int) > (sca0_2_1_argbuf,Pointer_CTf_f_Int_Int) */
  Pointer_CTf_f_Int_Int_t writeCTf_f_Int_IntlizzieLet47_1_argbuf_rwb_bufchan_d;
  logic writeCTf_f_Int_IntlizzieLet47_1_argbuf_rwb_bufchan_r;
  assign writeCTf_f_Int_IntlizzieLet47_1_argbuf_rwb_r = ((! writeCTf_f_Int_IntlizzieLet47_1_argbuf_rwb_bufchan_d[0]) || writeCTf_f_Int_IntlizzieLet47_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTf_f_Int_IntlizzieLet47_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                               1'd0};
    else
      if (writeCTf_f_Int_IntlizzieLet47_1_argbuf_rwb_r)
        writeCTf_f_Int_IntlizzieLet47_1_argbuf_rwb_bufchan_d <= writeCTf_f_Int_IntlizzieLet47_1_argbuf_rwb_d;
  Pointer_CTf_f_Int_Int_t writeCTf_f_Int_IntlizzieLet47_1_argbuf_rwb_bufchan_buf;
  assign writeCTf_f_Int_IntlizzieLet47_1_argbuf_rwb_bufchan_r = (! writeCTf_f_Int_IntlizzieLet47_1_argbuf_rwb_bufchan_buf[0]);
  assign sca0_2_1_argbuf_d = (writeCTf_f_Int_IntlizzieLet47_1_argbuf_rwb_bufchan_buf[0] ? writeCTf_f_Int_IntlizzieLet47_1_argbuf_rwb_bufchan_buf :
                              writeCTf_f_Int_IntlizzieLet47_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTf_f_Int_IntlizzieLet47_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                 1'd0};
    else
      if ((sca0_2_1_argbuf_r && writeCTf_f_Int_IntlizzieLet47_1_argbuf_rwb_bufchan_buf[0]))
        writeCTf_f_Int_IntlizzieLet47_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                   1'd0};
      else if (((! sca0_2_1_argbuf_r) && (! writeCTf_f_Int_IntlizzieLet47_1_argbuf_rwb_bufchan_buf[0])))
        writeCTf_f_Int_IntlizzieLet47_1_argbuf_rwb_bufchan_buf <= writeCTf_f_Int_IntlizzieLet47_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet11_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet11_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet11_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet11_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet11_1_argbuf_r = ((! writeQTree_IntlizzieLet11_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet11_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet11_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet11_1_argbuf_r)
        writeQTree_IntlizzieLet11_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet11_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet11_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet11_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet11_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet11_1_argbuf_rwb_d = (writeQTree_IntlizzieLet11_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet11_1_argbuf_bufchan_buf :
                                                     writeQTree_IntlizzieLet11_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet11_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet11_1_argbuf_rwb_r && writeQTree_IntlizzieLet11_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet11_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet11_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet11_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet11_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet11_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet11_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet4_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet11_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet11_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet11_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet11_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet11_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet11_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet11_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet11_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet11_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet11_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet11_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet11_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet4_1_1_argbuf_d = (writeQTree_IntlizzieLet11_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet11_1_argbuf_rwb_bufchan_buf :
                                    writeQTree_IntlizzieLet11_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet11_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((lizzieLet4_1_1_argbuf_r && writeQTree_IntlizzieLet11_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet11_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! lizzieLet4_1_1_argbuf_r) && (! writeQTree_IntlizzieLet11_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet11_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet11_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet14_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet14_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet14_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet14_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet14_1_argbuf_r = ((! writeQTree_IntlizzieLet14_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet14_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet14_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet14_1_argbuf_r)
        writeQTree_IntlizzieLet14_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet14_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet14_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet14_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet14_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet14_1_argbuf_rwb_d = (writeQTree_IntlizzieLet14_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet14_1_argbuf_bufchan_buf :
                                                     writeQTree_IntlizzieLet14_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet14_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet14_1_argbuf_rwb_r && writeQTree_IntlizzieLet14_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet14_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet14_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet14_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet14_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet14_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet14_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet6_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet14_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet14_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet14_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet14_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet14_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet14_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet14_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet14_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet14_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet14_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet14_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet14_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet6_1_1_argbuf_d = (writeQTree_IntlizzieLet14_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet14_1_argbuf_rwb_bufchan_buf :
                                    writeQTree_IntlizzieLet14_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet14_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((lizzieLet6_1_1_argbuf_r && writeQTree_IntlizzieLet14_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet14_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! lizzieLet6_1_1_argbuf_r) && (! writeQTree_IntlizzieLet14_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet14_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet14_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet15_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet15_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet15_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet15_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet15_1_argbuf_r = ((! writeQTree_IntlizzieLet15_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet15_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet15_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet15_1_argbuf_r)
        writeQTree_IntlizzieLet15_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet15_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet15_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet15_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet15_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet15_1_argbuf_rwb_d = (writeQTree_IntlizzieLet15_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet15_1_argbuf_bufchan_buf :
                                                     writeQTree_IntlizzieLet15_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet15_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet15_1_argbuf_rwb_r && writeQTree_IntlizzieLet15_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet15_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet15_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet15_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet15_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet15_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet15_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet7_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet15_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet15_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet15_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet15_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet15_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet15_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet15_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet15_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet15_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet15_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet15_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet15_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet7_1_1_argbuf_d = (writeQTree_IntlizzieLet15_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet15_1_argbuf_rwb_bufchan_buf :
                                    writeQTree_IntlizzieLet15_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet15_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((lizzieLet7_1_1_argbuf_r && writeQTree_IntlizzieLet15_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet15_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! lizzieLet7_1_1_argbuf_r) && (! writeQTree_IntlizzieLet15_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet15_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet15_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet16_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet16_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet16_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet16_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet16_1_argbuf_r = ((! writeQTree_IntlizzieLet16_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet16_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet16_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet16_1_argbuf_r)
        writeQTree_IntlizzieLet16_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet16_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet16_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet16_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet16_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet16_1_argbuf_rwb_d = (writeQTree_IntlizzieLet16_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet16_1_argbuf_bufchan_buf :
                                                     writeQTree_IntlizzieLet16_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet16_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet16_1_argbuf_rwb_r && writeQTree_IntlizzieLet16_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet16_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet16_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet16_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet16_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet16_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet16_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet8_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet16_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet16_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet16_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet16_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet16_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet16_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet16_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet16_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet16_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet16_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet16_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet16_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet8_1_1_argbuf_d = (writeQTree_IntlizzieLet16_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet16_1_argbuf_rwb_bufchan_buf :
                                    writeQTree_IntlizzieLet16_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet16_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((lizzieLet8_1_1_argbuf_r && writeQTree_IntlizzieLet16_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet16_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! lizzieLet8_1_1_argbuf_r) && (! writeQTree_IntlizzieLet16_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet16_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet16_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet17_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet17_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet17_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet17_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet17_1_argbuf_r = ((! writeQTree_IntlizzieLet17_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet17_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet17_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet17_1_argbuf_r)
        writeQTree_IntlizzieLet17_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet17_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet17_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet17_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet17_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet17_1_argbuf_rwb_d = (writeQTree_IntlizzieLet17_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet17_1_argbuf_bufchan_buf :
                                                     writeQTree_IntlizzieLet17_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet17_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet17_1_argbuf_rwb_r && writeQTree_IntlizzieLet17_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet17_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet17_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet17_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet17_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet17_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet17_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet9_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet17_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet17_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet17_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet17_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet17_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet17_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet17_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet17_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet17_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet17_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet17_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet17_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet9_1_1_argbuf_d = (writeQTree_IntlizzieLet17_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet17_1_argbuf_rwb_bufchan_buf :
                                    writeQTree_IntlizzieLet17_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet17_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((lizzieLet9_1_1_argbuf_r && writeQTree_IntlizzieLet17_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet17_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! lizzieLet9_1_1_argbuf_r) && (! writeQTree_IntlizzieLet17_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet17_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet17_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet18_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet18_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet18_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet18_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet18_1_argbuf_r = ((! writeQTree_IntlizzieLet18_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet18_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet18_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet18_1_argbuf_r)
        writeQTree_IntlizzieLet18_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet18_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet18_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet18_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet18_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet18_1_argbuf_rwb_d = (writeQTree_IntlizzieLet18_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet18_1_argbuf_bufchan_buf :
                                                     writeQTree_IntlizzieLet18_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet18_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet18_1_argbuf_rwb_r && writeQTree_IntlizzieLet18_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet18_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet18_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet18_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet18_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet18_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet18_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet10_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet18_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet18_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet18_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet18_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet18_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet18_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet18_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet18_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet18_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet18_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet18_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet18_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet10_1_1_argbuf_d = (writeQTree_IntlizzieLet18_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet18_1_argbuf_rwb_bufchan_buf :
                                     writeQTree_IntlizzieLet18_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet18_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((lizzieLet10_1_1_argbuf_r && writeQTree_IntlizzieLet18_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet18_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! lizzieLet10_1_1_argbuf_r) && (! writeQTree_IntlizzieLet18_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet18_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet18_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet20_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet20_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet20_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet20_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet20_1_argbuf_r = ((! writeQTree_IntlizzieLet20_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet20_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet20_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet20_1_argbuf_r)
        writeQTree_IntlizzieLet20_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet20_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet20_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet20_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet20_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet20_1_argbuf_rwb_d = (writeQTree_IntlizzieLet20_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet20_1_argbuf_bufchan_buf :
                                                     writeQTree_IntlizzieLet20_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet20_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet20_1_argbuf_rwb_r && writeQTree_IntlizzieLet20_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet20_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet20_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet20_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet20_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet20_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet20_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet11_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet20_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet20_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet20_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet20_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet20_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet20_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet20_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet20_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet20_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet20_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet20_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet20_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet11_1_1_argbuf_d = (writeQTree_IntlizzieLet20_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet20_1_argbuf_rwb_bufchan_buf :
                                     writeQTree_IntlizzieLet20_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet20_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((lizzieLet11_1_1_argbuf_r && writeQTree_IntlizzieLet20_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet20_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! lizzieLet11_1_1_argbuf_r) && (! writeQTree_IntlizzieLet20_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet20_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet20_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet21_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet21_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet21_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet21_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet21_1_argbuf_r = ((! writeQTree_IntlizzieLet21_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet21_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet21_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet21_1_argbuf_r)
        writeQTree_IntlizzieLet21_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet21_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet21_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet21_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet21_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet21_1_argbuf_rwb_d = (writeQTree_IntlizzieLet21_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet21_1_argbuf_bufchan_buf :
                                                     writeQTree_IntlizzieLet21_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet21_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet21_1_argbuf_rwb_r && writeQTree_IntlizzieLet21_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet21_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet21_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet21_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet21_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet21_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet21_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet12_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet21_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet21_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet21_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet21_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet21_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet21_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet21_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet21_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet21_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet21_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet21_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet21_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet12_1_1_argbuf_d = (writeQTree_IntlizzieLet21_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet21_1_argbuf_rwb_bufchan_buf :
                                     writeQTree_IntlizzieLet21_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet21_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((lizzieLet12_1_1_argbuf_r && writeQTree_IntlizzieLet21_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet21_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! lizzieLet12_1_1_argbuf_r) && (! writeQTree_IntlizzieLet21_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet21_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet21_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet22_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet22_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet22_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet22_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet22_1_argbuf_r = ((! writeQTree_IntlizzieLet22_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet22_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet22_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet22_1_argbuf_r)
        writeQTree_IntlizzieLet22_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet22_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet22_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet22_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet22_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet22_1_argbuf_rwb_d = (writeQTree_IntlizzieLet22_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet22_1_argbuf_bufchan_buf :
                                                     writeQTree_IntlizzieLet22_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet22_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet22_1_argbuf_rwb_r && writeQTree_IntlizzieLet22_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet22_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet22_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet22_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet22_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet22_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet22_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet13_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet22_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet22_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet22_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet22_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet22_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet22_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet22_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet22_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet22_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet22_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet22_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet22_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet13_1_1_argbuf_d = (writeQTree_IntlizzieLet22_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet22_1_argbuf_rwb_bufchan_buf :
                                     writeQTree_IntlizzieLet22_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet22_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((lizzieLet13_1_1_argbuf_r && writeQTree_IntlizzieLet22_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet22_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! lizzieLet13_1_1_argbuf_r) && (! writeQTree_IntlizzieLet22_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet22_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet22_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet23_2_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet23_2_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet23_2_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet23_2_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet23_2_1_argbuf_r = ((! writeQTree_IntlizzieLet23_2_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet23_2_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet23_2_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet23_2_1_argbuf_r)
        writeQTree_IntlizzieLet23_2_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet23_2_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet23_2_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet23_2_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet23_2_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet23_2_1_argbuf_rwb_d = (writeQTree_IntlizzieLet23_2_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet23_2_1_argbuf_bufchan_buf :
                                                       writeQTree_IntlizzieLet23_2_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet23_2_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet23_2_1_argbuf_rwb_r && writeQTree_IntlizzieLet23_2_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet23_2_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet23_2_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet23_2_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet23_2_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet23_2_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet23_2_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet14_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet23_2_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet23_2_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet23_2_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet23_2_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet23_2_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet23_2_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                             1'd0};
    else
      if (writeQTree_IntlizzieLet23_2_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet23_2_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet23_2_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet23_2_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet23_2_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet23_2_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet14_1_1_argbuf_d = (writeQTree_IntlizzieLet23_2_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet23_2_1_argbuf_rwb_bufchan_buf :
                                     writeQTree_IntlizzieLet23_2_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet23_2_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
    else
      if ((lizzieLet14_1_1_argbuf_r && writeQTree_IntlizzieLet23_2_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet23_2_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                 1'd0};
      else if (((! lizzieLet14_1_1_argbuf_r) && (! writeQTree_IntlizzieLet23_2_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet23_2_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet23_2_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet24_1_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet24_1_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet24_1_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet24_1_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet24_1_1_argbuf_r = ((! writeQTree_IntlizzieLet24_1_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet24_1_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet24_1_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet24_1_1_argbuf_r)
        writeQTree_IntlizzieLet24_1_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet24_1_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet24_1_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet24_1_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet24_1_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet24_1_1_argbuf_rwb_d = (writeQTree_IntlizzieLet24_1_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet24_1_1_argbuf_bufchan_buf :
                                                       writeQTree_IntlizzieLet24_1_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet24_1_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet24_1_1_argbuf_rwb_r && writeQTree_IntlizzieLet24_1_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet24_1_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet24_1_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet24_1_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet24_1_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet24_1_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet24_1_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet15_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet24_1_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet24_1_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet24_1_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet24_1_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet24_1_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet24_1_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                             1'd0};
    else
      if (writeQTree_IntlizzieLet24_1_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet24_1_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet24_1_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet24_1_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet24_1_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet24_1_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet15_1_1_argbuf_d = (writeQTree_IntlizzieLet24_1_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet24_1_1_argbuf_rwb_bufchan_buf :
                                     writeQTree_IntlizzieLet24_1_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet24_1_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
    else
      if ((lizzieLet15_1_1_argbuf_r && writeQTree_IntlizzieLet24_1_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet24_1_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                 1'd0};
      else if (((! lizzieLet15_1_1_argbuf_r) && (! writeQTree_IntlizzieLet24_1_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet24_1_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet24_1_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet25_1_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet25_1_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet25_1_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet25_1_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet25_1_1_argbuf_r = ((! writeQTree_IntlizzieLet25_1_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet25_1_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet25_1_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet25_1_1_argbuf_r)
        writeQTree_IntlizzieLet25_1_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet25_1_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet25_1_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet25_1_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet25_1_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet25_1_1_argbuf_rwb_d = (writeQTree_IntlizzieLet25_1_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet25_1_1_argbuf_bufchan_buf :
                                                       writeQTree_IntlizzieLet25_1_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet25_1_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet25_1_1_argbuf_rwb_r && writeQTree_IntlizzieLet25_1_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet25_1_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet25_1_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet25_1_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet25_1_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet25_1_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet25_1_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet16_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet25_1_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet25_1_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet25_1_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet25_1_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet25_1_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet25_1_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                             1'd0};
    else
      if (writeQTree_IntlizzieLet25_1_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet25_1_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet25_1_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet25_1_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet25_1_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet25_1_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet16_1_1_argbuf_d = (writeQTree_IntlizzieLet25_1_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet25_1_1_argbuf_rwb_bufchan_buf :
                                     writeQTree_IntlizzieLet25_1_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet25_1_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
    else
      if ((lizzieLet16_1_1_argbuf_r && writeQTree_IntlizzieLet25_1_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet25_1_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                 1'd0};
      else if (((! lizzieLet16_1_1_argbuf_r) && (! writeQTree_IntlizzieLet25_1_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet25_1_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet25_1_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet26_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet26_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet26_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet26_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet26_1_argbuf_r = ((! writeQTree_IntlizzieLet26_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet26_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet26_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet26_1_argbuf_r)
        writeQTree_IntlizzieLet26_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet26_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet26_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet26_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet26_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet26_1_argbuf_rwb_d = (writeQTree_IntlizzieLet26_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet26_1_argbuf_bufchan_buf :
                                                     writeQTree_IntlizzieLet26_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet26_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet26_1_argbuf_rwb_r && writeQTree_IntlizzieLet26_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet26_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet26_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet26_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet26_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet26_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet26_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet17_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet26_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet26_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet26_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet26_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet26_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet26_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet26_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet26_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet26_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet26_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet26_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet26_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet17_1_1_argbuf_d = (writeQTree_IntlizzieLet26_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet26_1_argbuf_rwb_bufchan_buf :
                                     writeQTree_IntlizzieLet26_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet26_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((lizzieLet17_1_1_argbuf_r && writeQTree_IntlizzieLet26_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet26_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! lizzieLet17_1_1_argbuf_r) && (! writeQTree_IntlizzieLet26_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet26_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet26_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet28_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet28_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet28_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet28_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet28_1_argbuf_r = ((! writeQTree_IntlizzieLet28_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet28_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet28_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet28_1_argbuf_r)
        writeQTree_IntlizzieLet28_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet28_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet28_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet28_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet28_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet28_1_argbuf_rwb_d = (writeQTree_IntlizzieLet28_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet28_1_argbuf_bufchan_buf :
                                                     writeQTree_IntlizzieLet28_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet28_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet28_1_argbuf_rwb_r && writeQTree_IntlizzieLet28_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet28_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet28_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet28_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet28_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet28_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet28_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet18_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet28_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet28_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet28_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet28_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet28_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet28_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet28_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet28_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet28_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet28_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet28_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet28_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet18_1_1_argbuf_d = (writeQTree_IntlizzieLet28_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet28_1_argbuf_rwb_bufchan_buf :
                                     writeQTree_IntlizzieLet28_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet28_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((lizzieLet18_1_1_argbuf_r && writeQTree_IntlizzieLet28_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet28_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! lizzieLet18_1_1_argbuf_r) && (! writeQTree_IntlizzieLet28_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet28_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet28_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet29_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet29_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet29_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet29_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet29_1_argbuf_r = ((! writeQTree_IntlizzieLet29_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet29_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet29_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet29_1_argbuf_r)
        writeQTree_IntlizzieLet29_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet29_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet29_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet29_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet29_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet29_1_argbuf_rwb_d = (writeQTree_IntlizzieLet29_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet29_1_argbuf_bufchan_buf :
                                                     writeQTree_IntlizzieLet29_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet29_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet29_1_argbuf_rwb_r && writeQTree_IntlizzieLet29_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet29_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet29_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet29_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet29_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet29_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet29_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet19_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet29_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet29_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet29_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet29_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet29_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet29_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet29_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet29_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet29_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet29_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet29_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet29_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet19_1_argbuf_d = (writeQTree_IntlizzieLet29_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet29_1_argbuf_rwb_bufchan_buf :
                                   writeQTree_IntlizzieLet29_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet29_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((lizzieLet19_1_argbuf_r && writeQTree_IntlizzieLet29_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet29_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! lizzieLet19_1_argbuf_r) && (! writeQTree_IntlizzieLet29_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet29_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet29_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet31_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet31_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet31_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet31_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet31_1_argbuf_r = ((! writeQTree_IntlizzieLet31_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet31_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet31_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet31_1_argbuf_r)
        writeQTree_IntlizzieLet31_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet31_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet31_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet31_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet31_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet31_1_argbuf_rwb_d = (writeQTree_IntlizzieLet31_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet31_1_argbuf_bufchan_buf :
                                                     writeQTree_IntlizzieLet31_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet31_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet31_1_argbuf_rwb_r && writeQTree_IntlizzieLet31_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet31_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet31_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet31_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet31_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet31_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet31_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet20_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet31_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet31_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet31_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet31_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet31_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet31_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet31_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet31_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet31_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet31_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet31_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet31_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet20_1_1_argbuf_d = (writeQTree_IntlizzieLet31_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet31_1_argbuf_rwb_bufchan_buf :
                                     writeQTree_IntlizzieLet31_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet31_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((lizzieLet20_1_1_argbuf_r && writeQTree_IntlizzieLet31_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet31_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! lizzieLet20_1_1_argbuf_r) && (! writeQTree_IntlizzieLet31_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet31_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet31_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet32_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet32_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet32_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet32_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet32_1_argbuf_r = ((! writeQTree_IntlizzieLet32_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet32_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet32_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet32_1_argbuf_r)
        writeQTree_IntlizzieLet32_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet32_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet32_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet32_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet32_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet32_1_argbuf_rwb_d = (writeQTree_IntlizzieLet32_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet32_1_argbuf_bufchan_buf :
                                                     writeQTree_IntlizzieLet32_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet32_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet32_1_argbuf_rwb_r && writeQTree_IntlizzieLet32_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet32_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet32_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet32_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet32_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet32_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet32_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet21_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet32_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet32_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet32_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet32_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet32_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet32_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet32_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet32_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet32_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet32_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet32_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet32_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet21_1_1_argbuf_d = (writeQTree_IntlizzieLet32_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet32_1_argbuf_rwb_bufchan_buf :
                                     writeQTree_IntlizzieLet32_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet32_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((lizzieLet21_1_1_argbuf_r && writeQTree_IntlizzieLet32_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet32_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! lizzieLet21_1_1_argbuf_r) && (! writeQTree_IntlizzieLet32_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet32_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet32_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet43_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet43_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet43_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet43_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet43_1_argbuf_r = ((! writeQTree_IntlizzieLet43_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet43_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet43_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet43_1_argbuf_r)
        writeQTree_IntlizzieLet43_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet43_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet43_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet43_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet43_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet43_1_argbuf_rwb_d = (writeQTree_IntlizzieLet43_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet43_1_argbuf_bufchan_buf :
                                                     writeQTree_IntlizzieLet43_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet43_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet43_1_argbuf_rwb_r && writeQTree_IntlizzieLet43_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet43_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet43_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet43_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet43_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet43_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet43_1_argbuf_rwb,Pointer_QTree_Int) > (contRet_0_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet43_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet43_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet43_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet43_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet43_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet43_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet43_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet43_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet43_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet43_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet43_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet43_1_argbuf_rwb_bufchan_buf[0]);
  assign contRet_0_1_1_argbuf_d = (writeQTree_IntlizzieLet43_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet43_1_argbuf_rwb_bufchan_buf :
                                   writeQTree_IntlizzieLet43_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet43_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((contRet_0_1_1_argbuf_r && writeQTree_IntlizzieLet43_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet43_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! contRet_0_1_1_argbuf_r) && (! writeQTree_IntlizzieLet43_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet43_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet43_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet48_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet48_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet48_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet48_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet48_1_argbuf_r = ((! writeQTree_IntlizzieLet48_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet48_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet48_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet48_1_argbuf_r)
        writeQTree_IntlizzieLet48_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet48_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet48_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet48_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet48_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet48_1_argbuf_rwb_d = (writeQTree_IntlizzieLet48_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet48_1_argbuf_bufchan_buf :
                                                     writeQTree_IntlizzieLet48_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet48_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet48_1_argbuf_rwb_r && writeQTree_IntlizzieLet48_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet48_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet48_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet48_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet48_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet48_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet48_1_argbuf_rwb,Pointer_QTree_Int) > (contRet_0_2_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet48_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet48_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet48_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet48_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet48_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet48_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet48_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet48_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet48_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet48_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet48_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet48_1_argbuf_rwb_bufchan_buf[0]);
  assign contRet_0_2_1_argbuf_d = (writeQTree_IntlizzieLet48_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet48_1_argbuf_rwb_bufchan_buf :
                                   writeQTree_IntlizzieLet48_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet48_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((contRet_0_2_1_argbuf_r && writeQTree_IntlizzieLet48_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet48_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! contRet_0_2_1_argbuf_r) && (! writeQTree_IntlizzieLet48_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet48_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet48_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet7_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet7_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet7_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet7_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet7_1_argbuf_r = ((! writeQTree_IntlizzieLet7_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet7_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet7_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet7_1_argbuf_r)
        writeQTree_IntlizzieLet7_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet7_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet7_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet7_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet7_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet7_1_argbuf_rwb_d = (writeQTree_IntlizzieLet7_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet7_1_argbuf_bufchan_buf :
                                                    writeQTree_IntlizzieLet7_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet7_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet7_1_argbuf_rwb_r && writeQTree_IntlizzieLet7_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet7_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet7_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet7_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet7_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet7_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet7_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet1_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet7_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet7_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet7_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet7_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet7_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet7_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet7_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet7_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet7_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet7_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet7_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet7_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet1_1_1_argbuf_d = (writeQTree_IntlizzieLet7_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet7_1_argbuf_rwb_bufchan_buf :
                                    writeQTree_IntlizzieLet7_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet7_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet1_1_1_argbuf_r && writeQTree_IntlizzieLet7_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet7_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet1_1_1_argbuf_r) && (! writeQTree_IntlizzieLet7_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet7_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet7_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet8_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet8_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet8_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet8_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet8_1_argbuf_r = ((! writeQTree_IntlizzieLet8_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet8_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet8_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet8_1_argbuf_r)
        writeQTree_IntlizzieLet8_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet8_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet8_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet8_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet8_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet8_1_argbuf_rwb_d = (writeQTree_IntlizzieLet8_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet8_1_argbuf_bufchan_buf :
                                                    writeQTree_IntlizzieLet8_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet8_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet8_1_argbuf_rwb_r && writeQTree_IntlizzieLet8_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet8_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet8_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet8_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet8_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet8_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet8_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet2_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet8_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet8_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet8_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet8_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet8_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet8_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet8_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet8_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet8_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet8_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet8_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet8_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet2_1_1_argbuf_d = (writeQTree_IntlizzieLet8_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet8_1_argbuf_rwb_bufchan_buf :
                                    writeQTree_IntlizzieLet8_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet8_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet2_1_1_argbuf_r && writeQTree_IntlizzieLet8_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet8_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet2_1_1_argbuf_r) && (! writeQTree_IntlizzieLet8_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet8_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet8_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet9_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet9_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet9_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet9_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet9_1_argbuf_r = ((! writeQTree_IntlizzieLet9_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet9_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet9_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet9_1_argbuf_r)
        writeQTree_IntlizzieLet9_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet9_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet9_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet9_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet9_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet9_1_argbuf_rwb_d = (writeQTree_IntlizzieLet9_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet9_1_argbuf_bufchan_buf :
                                                    writeQTree_IntlizzieLet9_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet9_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet9_1_argbuf_rwb_r && writeQTree_IntlizzieLet9_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet9_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet9_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet9_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet9_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet9_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet9_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet3_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet9_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet9_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet9_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet9_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet9_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet9_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet9_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet9_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet9_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet9_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet9_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet9_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet3_1_1_argbuf_d = (writeQTree_IntlizzieLet9_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet9_1_argbuf_rwb_bufchan_buf :
                                    writeQTree_IntlizzieLet9_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet9_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet3_1_1_argbuf_r && writeQTree_IntlizzieLet9_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet9_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet3_1_1_argbuf_r) && (! writeQTree_IntlizzieLet9_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet9_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet9_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (wsiX_1_goMux_mux,Pointer_QTree_Int) > (wsiX_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t wsiX_1_goMux_mux_bufchan_d;
  logic wsiX_1_goMux_mux_bufchan_r;
  assign wsiX_1_goMux_mux_r = ((! wsiX_1_goMux_mux_bufchan_d[0]) || wsiX_1_goMux_mux_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) wsiX_1_goMux_mux_bufchan_d <= {16'd0, 1'd0};
    else
      if (wsiX_1_goMux_mux_r)
        wsiX_1_goMux_mux_bufchan_d <= wsiX_1_goMux_mux_d;
  Pointer_QTree_Int_t wsiX_1_goMux_mux_bufchan_buf;
  assign wsiX_1_goMux_mux_bufchan_r = (! wsiX_1_goMux_mux_bufchan_buf[0]);
  assign wsiX_1_1_argbuf_d = (wsiX_1_goMux_mux_bufchan_buf[0] ? wsiX_1_goMux_mux_bufchan_buf :
                              wsiX_1_goMux_mux_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) wsiX_1_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((wsiX_1_1_argbuf_r && wsiX_1_goMux_mux_bufchan_buf[0]))
        wsiX_1_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
      else if (((! wsiX_1_1_argbuf_r) && (! wsiX_1_goMux_mux_bufchan_buf[0])))
        wsiX_1_goMux_mux_bufchan_buf <= wsiX_1_goMux_mux_bufchan_d;
  
  /* buf (Ty CT$wnnz) : (wwsj0_2_1lizzieLet35_4Lcall_$wnnz2_1sc_0_4_1q4a87_2_1Lcall_$wnnz1,CT$wnnz) > (lizzieLet37_1_argbuf,CT$wnnz) */
  CT$wnnz_t wwsj0_2_1lizzieLet35_4Lcall_$wnnz2_1sc_0_4_1q4a87_2_1Lcall_$wnnz1_bufchan_d;
  logic wwsj0_2_1lizzieLet35_4Lcall_$wnnz2_1sc_0_4_1q4a87_2_1Lcall_$wnnz1_bufchan_r;
  assign wwsj0_2_1lizzieLet35_4Lcall_$wnnz2_1sc_0_4_1q4a87_2_1Lcall_$wnnz1_r = ((! wwsj0_2_1lizzieLet35_4Lcall_$wnnz2_1sc_0_4_1q4a87_2_1Lcall_$wnnz1_bufchan_d[0]) || wwsj0_2_1lizzieLet35_4Lcall_$wnnz2_1sc_0_4_1q4a87_2_1Lcall_$wnnz1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      wwsj0_2_1lizzieLet35_4Lcall_$wnnz2_1sc_0_4_1q4a87_2_1Lcall_$wnnz1_bufchan_d <= {115'd0,
                                                                                      1'd0};
    else
      if (wwsj0_2_1lizzieLet35_4Lcall_$wnnz2_1sc_0_4_1q4a87_2_1Lcall_$wnnz1_r)
        wwsj0_2_1lizzieLet35_4Lcall_$wnnz2_1sc_0_4_1q4a87_2_1Lcall_$wnnz1_bufchan_d <= wwsj0_2_1lizzieLet35_4Lcall_$wnnz2_1sc_0_4_1q4a87_2_1Lcall_$wnnz1_d;
  CT$wnnz_t wwsj0_2_1lizzieLet35_4Lcall_$wnnz2_1sc_0_4_1q4a87_2_1Lcall_$wnnz1_bufchan_buf;
  assign wwsj0_2_1lizzieLet35_4Lcall_$wnnz2_1sc_0_4_1q4a87_2_1Lcall_$wnnz1_bufchan_r = (! wwsj0_2_1lizzieLet35_4Lcall_$wnnz2_1sc_0_4_1q4a87_2_1Lcall_$wnnz1_bufchan_buf[0]);
  assign lizzieLet37_1_argbuf_d = (wwsj0_2_1lizzieLet35_4Lcall_$wnnz2_1sc_0_4_1q4a87_2_1Lcall_$wnnz1_bufchan_buf[0] ? wwsj0_2_1lizzieLet35_4Lcall_$wnnz2_1sc_0_4_1q4a87_2_1Lcall_$wnnz1_bufchan_buf :
                                   wwsj0_2_1lizzieLet35_4Lcall_$wnnz2_1sc_0_4_1q4a87_2_1Lcall_$wnnz1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      wwsj0_2_1lizzieLet35_4Lcall_$wnnz2_1sc_0_4_1q4a87_2_1Lcall_$wnnz1_bufchan_buf <= {115'd0,
                                                                                        1'd0};
    else
      if ((lizzieLet37_1_argbuf_r && wwsj0_2_1lizzieLet35_4Lcall_$wnnz2_1sc_0_4_1q4a87_2_1Lcall_$wnnz1_bufchan_buf[0]))
        wwsj0_2_1lizzieLet35_4Lcall_$wnnz2_1sc_0_4_1q4a87_2_1Lcall_$wnnz1_bufchan_buf <= {115'd0,
                                                                                          1'd0};
      else if (((! lizzieLet37_1_argbuf_r) && (! wwsj0_2_1lizzieLet35_4Lcall_$wnnz2_1sc_0_4_1q4a87_2_1Lcall_$wnnz1_bufchan_buf[0])))
        wwsj0_2_1lizzieLet35_4Lcall_$wnnz2_1sc_0_4_1q4a87_2_1Lcall_$wnnz1_bufchan_buf <= wwsj0_2_1lizzieLet35_4Lcall_$wnnz2_1sc_0_4_1q4a87_2_1Lcall_$wnnz1_bufchan_d;
  
  /* dcon (Ty CT$wnnz,Dcon Lcall_$wnnz1) : [(wwsj0_2_destruct,Int#),
                                       (lizzieLet35_4Lcall_$wnnz2,Int#),
                                       (sc_0_4_destruct,Pointer_CT$wnnz),
                                       (q4a87_2_destruct,Pointer_QTree_Int)] > (wwsj0_2_1lizzieLet35_4Lcall_$wnnz2_1sc_0_4_1q4a87_2_1Lcall_$wnnz1,CT$wnnz) */
  assign wwsj0_2_1lizzieLet35_4Lcall_$wnnz2_1sc_0_4_1q4a87_2_1Lcall_$wnnz1_d = Lcall_$wnnz1_dc((& {wwsj0_2_destruct_d[0],
                                                                                                   lizzieLet35_4Lcall_$wnnz2_d[0],
                                                                                                   sc_0_4_destruct_d[0],
                                                                                                   q4a87_2_destruct_d[0]}), wwsj0_2_destruct_d, lizzieLet35_4Lcall_$wnnz2_d, sc_0_4_destruct_d, q4a87_2_destruct_d);
  assign {wwsj0_2_destruct_r,
          lizzieLet35_4Lcall_$wnnz2_r,
          sc_0_4_destruct_r,
          q4a87_2_destruct_r} = {4 {(wwsj0_2_1lizzieLet35_4Lcall_$wnnz2_1sc_0_4_1q4a87_2_1Lcall_$wnnz1_r && wwsj0_2_1lizzieLet35_4Lcall_$wnnz2_1sc_0_4_1q4a87_2_1Lcall_$wnnz1_d[0])}};
  
  /* buf (Ty CT$wnnz) : (wwsj0_3_1ww1Xju_1_1lizzieLet35_4Lcall_$wnnz1_1sc_0_5_1Lcall_$wnnz0,CT$wnnz) > (lizzieLet38_1_argbuf,CT$wnnz) */
  CT$wnnz_t wwsj0_3_1ww1Xju_1_1lizzieLet35_4Lcall_$wnnz1_1sc_0_5_1Lcall_$wnnz0_bufchan_d;
  logic wwsj0_3_1ww1Xju_1_1lizzieLet35_4Lcall_$wnnz1_1sc_0_5_1Lcall_$wnnz0_bufchan_r;
  assign wwsj0_3_1ww1Xju_1_1lizzieLet35_4Lcall_$wnnz1_1sc_0_5_1Lcall_$wnnz0_r = ((! wwsj0_3_1ww1Xju_1_1lizzieLet35_4Lcall_$wnnz1_1sc_0_5_1Lcall_$wnnz0_bufchan_d[0]) || wwsj0_3_1ww1Xju_1_1lizzieLet35_4Lcall_$wnnz1_1sc_0_5_1Lcall_$wnnz0_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      wwsj0_3_1ww1Xju_1_1lizzieLet35_4Lcall_$wnnz1_1sc_0_5_1Lcall_$wnnz0_bufchan_d <= {115'd0,
                                                                                       1'd0};
    else
      if (wwsj0_3_1ww1Xju_1_1lizzieLet35_4Lcall_$wnnz1_1sc_0_5_1Lcall_$wnnz0_r)
        wwsj0_3_1ww1Xju_1_1lizzieLet35_4Lcall_$wnnz1_1sc_0_5_1Lcall_$wnnz0_bufchan_d <= wwsj0_3_1ww1Xju_1_1lizzieLet35_4Lcall_$wnnz1_1sc_0_5_1Lcall_$wnnz0_d;
  CT$wnnz_t wwsj0_3_1ww1Xju_1_1lizzieLet35_4Lcall_$wnnz1_1sc_0_5_1Lcall_$wnnz0_bufchan_buf;
  assign wwsj0_3_1ww1Xju_1_1lizzieLet35_4Lcall_$wnnz1_1sc_0_5_1Lcall_$wnnz0_bufchan_r = (! wwsj0_3_1ww1Xju_1_1lizzieLet35_4Lcall_$wnnz1_1sc_0_5_1Lcall_$wnnz0_bufchan_buf[0]);
  assign lizzieLet38_1_argbuf_d = (wwsj0_3_1ww1Xju_1_1lizzieLet35_4Lcall_$wnnz1_1sc_0_5_1Lcall_$wnnz0_bufchan_buf[0] ? wwsj0_3_1ww1Xju_1_1lizzieLet35_4Lcall_$wnnz1_1sc_0_5_1Lcall_$wnnz0_bufchan_buf :
                                   wwsj0_3_1ww1Xju_1_1lizzieLet35_4Lcall_$wnnz1_1sc_0_5_1Lcall_$wnnz0_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      wwsj0_3_1ww1Xju_1_1lizzieLet35_4Lcall_$wnnz1_1sc_0_5_1Lcall_$wnnz0_bufchan_buf <= {115'd0,
                                                                                         1'd0};
    else
      if ((lizzieLet38_1_argbuf_r && wwsj0_3_1ww1Xju_1_1lizzieLet35_4Lcall_$wnnz1_1sc_0_5_1Lcall_$wnnz0_bufchan_buf[0]))
        wwsj0_3_1ww1Xju_1_1lizzieLet35_4Lcall_$wnnz1_1sc_0_5_1Lcall_$wnnz0_bufchan_buf <= {115'd0,
                                                                                           1'd0};
      else if (((! lizzieLet38_1_argbuf_r) && (! wwsj0_3_1ww1Xju_1_1lizzieLet35_4Lcall_$wnnz1_1sc_0_5_1Lcall_$wnnz0_bufchan_buf[0])))
        wwsj0_3_1ww1Xju_1_1lizzieLet35_4Lcall_$wnnz1_1sc_0_5_1Lcall_$wnnz0_bufchan_buf <= wwsj0_3_1ww1Xju_1_1lizzieLet35_4Lcall_$wnnz1_1sc_0_5_1Lcall_$wnnz0_bufchan_d;
  
  /* dcon (Ty CT$wnnz,Dcon Lcall_$wnnz0) : [(wwsj0_3_destruct,Int#),
                                       (ww1Xju_1_destruct,Int#),
                                       (lizzieLet35_4Lcall_$wnnz1,Int#),
                                       (sc_0_5_destruct,Pointer_CT$wnnz)] > (wwsj0_3_1ww1Xju_1_1lizzieLet35_4Lcall_$wnnz1_1sc_0_5_1Lcall_$wnnz0,CT$wnnz) */
  assign wwsj0_3_1ww1Xju_1_1lizzieLet35_4Lcall_$wnnz1_1sc_0_5_1Lcall_$wnnz0_d = Lcall_$wnnz0_dc((& {wwsj0_3_destruct_d[0],
                                                                                                    ww1Xju_1_destruct_d[0],
                                                                                                    lizzieLet35_4Lcall_$wnnz1_d[0],
                                                                                                    sc_0_5_destruct_d[0]}), wwsj0_3_destruct_d, ww1Xju_1_destruct_d, lizzieLet35_4Lcall_$wnnz1_d, sc_0_5_destruct_d);
  assign {wwsj0_3_destruct_r,
          ww1Xju_1_destruct_r,
          lizzieLet35_4Lcall_$wnnz1_r,
          sc_0_5_destruct_r} = {4 {(wwsj0_3_1ww1Xju_1_1lizzieLet35_4Lcall_$wnnz1_1sc_0_5_1Lcall_$wnnz0_r && wwsj0_3_1ww1Xju_1_1lizzieLet35_4Lcall_$wnnz1_1sc_0_5_1Lcall_$wnnz0_d[0])}};
  
  /* op_add (Ty Int#) : (wwsj0_4_1ww1Xju_2_1_Add32,Int#) (ww2Xjx_1_destruct,Int#) > (es_6_2_1ww2Xjx_1_1_Add32,Int#) */
  assign es_6_2_1ww2Xjx_1_1_Add32_d = {(wwsj0_4_1ww1Xju_2_1_Add32_d[32:1] + ww2Xjx_1_destruct_d[32:1]),
                                       (wwsj0_4_1ww1Xju_2_1_Add32_d[0] && ww2Xjx_1_destruct_d[0])};
  assign {wwsj0_4_1ww1Xju_2_1_Add32_r,
          ww2Xjx_1_destruct_r} = {2 {(es_6_2_1ww2Xjx_1_1_Add32_r && es_6_2_1ww2Xjx_1_1_Add32_d[0])}};
  
  /* op_add (Ty Int#) : (wwsj0_4_destruct,Int#) (ww1Xju_2_destruct,Int#) > (wwsj0_4_1ww1Xju_2_1_Add32,Int#) */
  assign wwsj0_4_1ww1Xju_2_1_Add32_d = {(wwsj0_4_destruct_d[32:1] + ww1Xju_2_destruct_d[32:1]),
                                        (wwsj0_4_destruct_d[0] && ww1Xju_2_destruct_d[0])};
  assign {wwsj0_4_destruct_r,
          ww1Xju_2_destruct_r} = {2 {(wwsj0_4_1ww1Xju_2_1_Add32_r && wwsj0_4_1ww1Xju_2_1_Add32_d[0])}};
  
  /* dcon (Ty Int,
      Dcon I#) : [(x1agS_1lizzieLet0_1_1_Add32,Int#)] > (es_0_1_1I#,Int) */
  assign \es_0_1_1I#_d  = \I#_dc ((& {x1agS_1lizzieLet0_1_1_Add32_d[0]}), x1agS_1lizzieLet0_1_1_Add32_d);
  assign {x1agS_1lizzieLet0_1_1_Add32_r} = {1 {(\es_0_1_1I#_r  && \es_0_1_1I#_d [0])}};
  
  /* op_add (Ty Int#) : (x1agS_destruct,Int#) (arg0_2_1Dcon_main1_3I#_1_argbuf_2,Int#) > (x1agS_1lizzieLet0_1_1_Add32,Int#) */
  assign x1agS_1lizzieLet0_1_1_Add32_d = {(x1agS_destruct_d[32:1] + \arg0_2_1Dcon_main1_3I#_1_argbuf_2_d [32:1]),
                                          (x1agS_destruct_d[0] && \arg0_2_1Dcon_main1_3I#_1_argbuf_2_d [0])};
  assign {x1agS_destruct_r,
          \arg0_2_1Dcon_main1_3I#_1_argbuf_2_r } = {2 {(x1agS_1lizzieLet0_1_1_Add32_r && x1agS_1lizzieLet0_1_1_Add32_d[0])}};
endmodule