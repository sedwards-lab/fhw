`timescale 1ns/1ns
import mMaskKron_package::*;

module mMaskKron(
  input logic clk,
  input logic reset,
  input Go_t \\QTree_Int_src_d ,
  output logic \\QTree_Int_src_r ,
  input QTree_Int_t dummy_write_QTree_Int_d,
  output logic dummy_write_QTree_Int_r,
  input Go_t sourceGo_d,
  output logic sourceGo_r,
  input Pointer_QTree_Int_t w1svB_1_1_d,
  output logic w1svB_1_1_r,
  input Pointer_QTree_Int_t wsvA_1_0_d,
  output logic wsvA_1_0_r,
  output \Word16#_t  forkHP1_QTree_Int_snk_dout,
  input logic forkHP1_QTree_Int_snk_rout,
  output Pointer_QTree_Int_t dummy_write_QTree_Int_sink_dout,
  input logic dummy_write_QTree_Int_sink_rout,
  output Int_t \es_0_1I#_dout ,
  input logic \es_0_1I#_rout 
  );
  /* --define=INPUTS=((__05CQTree_Int_src, 0, 1, Go), (dummy_write_QTree_Int, 66, 73786976294838206464, QTree_Int), (sourceGo, 0, 1, Go), (w1svB_1_1, 16, 65536, Pointer_QTree_Int), (wsvA_1_0, 16, 65536, Pointer_QTree_Int)) */
  /* --define=TAPS=() */
  /* --define=OUTPUTS=((forkHP1_QTree_Int_snk, 16, 65536, Word16__023), (dummy_write_QTree_Int_sink, 16, 65536, Pointer_QTree_Int), (es_0_1I__023, 32, 4294967296, Int)) */
  /* TYPE_START
CT__024wnnz_Int 16 3 (0,[0]) (1,[16p,16p,16p,16p]) (2,[32,16p,16p,16p]) (3,[32,32,16p,16p]) (4,[32,32,32,16p])
QTree_Int 16 2 (0,[0]) (1,[32]) (2,[16p,16p,16p,16p]) (3,[0])
CTmain_map__027_Int_Int 16 3 (0,[0]) (1,[16p,0,0,16p,16p,16p]) (2,[16p,16p,0,0,16p,16p]) (3,[16p,16p,16p,0,0,16p]) (4,[16p,16p,16p,16p])
CTmap__027__027_map__027__027_Int_Int_Int 16 3 (0,[0]) (1,[16p,0,0,32,16p,16p,16p]) (2,[16p,16p,0,0,32,16p,16p]) (3,[16p,16p,16p,0,0,32,16p]) (4,[16p,16p,16p,16p])
CTkron_kron_Int_Int_Int 16 3 (0,[0]) (1,[16p,0,0,16p,16p,16p,16p]) (2,[16p,16p,0,0,16p,16p,16p]) (3,[16p,16p,16p,0,0,16p,16p]) (4,[16p,16p,16p,16p])
TupGo___Pointer_QTree_Int___Pointer_QTree_Int 16 0 (0,[0,16p,16p])
TupGo___Pointer_QTree_Int 16 0 (0,[0,16p])
TupGo___Pointer_QTree_Int___Pointer_CT__024wnnz_Int 16 0 (0,[0,16p,16p])
TupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Int 16 0 (0,[0,0,0,16p,16p,16p])
TupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int___Pointer_CTmain_map__027_Int_Int 16 0 (0,[0,0,0,16p,16p])
TupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap__027__027_map__027__027_Int_Int_Int 16 0 (0,[0,0,0,32,16p,16p])
TupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int 16 0 (0,[0,0,0,16p,16p])
TupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int 16 0 (0,[0,0,0,16p])
TupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int 16 0 (0,[0,0,0,32,16p])
TYPE_END */
  /*  */
  /*  */
  Go_t goFork_d;
  logic goFork_r;
  Go_t goFor_2_d;
  logic goFor_2_r;
  Go_t goFor_3_d;
  logic goFor_3_r;
  Go_t goFor_4_d;
  logic goFor_4_r;
  Go_t goFor_5_d;
  logic goFor_5_r;
  Go_t goFor_6_d;
  logic goFor_6_r;
  Go_t goFor_7_d;
  logic goFor_7_r;
  Go_t goFor_8_d;
  logic goFor_8_r;
  Go_t goFor_9_d;
  logic goFor_9_r;
  \Word16#_t  initHP_CT$wnnz_Int_d;
  logic initHP_CT$wnnz_Int_r;
  \Word16#_t  incrHP_CT$wnnz_Int_d;
  logic incrHP_CT$wnnz_Int_r;
  Go_t incrHP_mergeCT$wnnz_Int_d;
  logic incrHP_mergeCT$wnnz_Int_r;
  Go_t incrHP_CT$wnnz_Int1_d;
  logic incrHP_CT$wnnz_Int1_r;
  Go_t incrHP_CT$wnnz_Int2_d;
  logic incrHP_CT$wnnz_Int2_r;
  \Word16#_t  addHP_CT$wnnz_Int_d;
  logic addHP_CT$wnnz_Int_r;
  \Word16#_t  mergeHP_CT$wnnz_Int_d;
  logic mergeHP_CT$wnnz_Int_r;
  Go_t incrHP_mergeCT$wnnz_Int_buf_d;
  logic incrHP_mergeCT$wnnz_Int_buf_r;
  \Word16#_t  mergeHP_CT$wnnz_Int_buf_d;
  logic mergeHP_CT$wnnz_Int_buf_r;
  \Word16#_t  forkHP1_CT$wnnz_Int_d;
  logic forkHP1_CT$wnnz_Int_r;
  \Word16#_t  forkHP1_CT$wnnz_In2_d;
  logic forkHP1_CT$wnnz_In2_r;
  \Word16#_t  forkHP1_CT$wnnz_In3_d;
  logic forkHP1_CT$wnnz_In3_r;
  C2_t memMergeChoice_CT$wnnz_Int_d;
  logic memMergeChoice_CT$wnnz_Int_r;
  MemIn_CT$wnnz_Int_t memMergeIn_CT$wnnz_Int_d;
  logic memMergeIn_CT$wnnz_Int_r;
  MemOut_CT$wnnz_Int_t memOut_CT$wnnz_Int_d;
  logic memOut_CT$wnnz_Int_r;
  MemOut_CT$wnnz_Int_t memReadOut_CT$wnnz_Int_d;
  logic memReadOut_CT$wnnz_Int_r;
  MemOut_CT$wnnz_Int_t memWriteOut_CT$wnnz_Int_d;
  logic memWriteOut_CT$wnnz_Int_r;
  MemIn_CT$wnnz_Int_t memMergeIn_CT$wnnz_Int_dbuf_d;
  logic memMergeIn_CT$wnnz_Int_dbuf_r;
  MemIn_CT$wnnz_Int_t memMergeIn_CT$wnnz_Int_rbuf_d;
  logic memMergeIn_CT$wnnz_Int_rbuf_r;
  MemOut_CT$wnnz_Int_t memOut_CT$wnnz_Int_dbuf_d;
  logic memOut_CT$wnnz_Int_dbuf_r;
  MemOut_CT$wnnz_Int_t memOut_CT$wnnz_Int_rbuf_d;
  logic memOut_CT$wnnz_Int_rbuf_r;
  \Word16#_t  destructReadIn_CT$wnnz_Int_d;
  logic destructReadIn_CT$wnnz_Int_r;
  MemIn_CT$wnnz_Int_t dconReadIn_CT$wnnz_Int_d;
  logic dconReadIn_CT$wnnz_Int_r;
  CT$wnnz_Int_t readPointer_CT$wnnz_Intscfarg_0_1_argbuf_d;
  logic readPointer_CT$wnnz_Intscfarg_0_1_argbuf_r;
  C5_t writeMerge_choice_CT$wnnz_Int_d;
  logic writeMerge_choice_CT$wnnz_Int_r;
  CT$wnnz_Int_t writeMerge_data_CT$wnnz_Int_d;
  logic writeMerge_data_CT$wnnz_Int_r;
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet0_1_argbuf_d;
  logic writeCT$wnnz_IntlizzieLet0_1_argbuf_r;
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet26_1_argbuf_d;
  logic writeCT$wnnz_IntlizzieLet26_1_argbuf_r;
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet27_1_argbuf_d;
  logic writeCT$wnnz_IntlizzieLet27_1_argbuf_r;
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet28_1_argbuf_d;
  logic writeCT$wnnz_IntlizzieLet28_1_argbuf_r;
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet5_1_argbuf_d;
  logic writeCT$wnnz_IntlizzieLet5_1_argbuf_r;
  MemIn_CT$wnnz_Int_t dconWriteIn_CT$wnnz_Int_d;
  logic dconWriteIn_CT$wnnz_Int_r;
  Pointer_CT$wnnz_Int_t dconPtr_CT$wnnz_Int_d;
  logic dconPtr_CT$wnnz_Int_r;
  Pointer_CT$wnnz_Int_t _39_d;
  logic _39_r;
  assign _39_r = 1'd1;
  Pointer_CT$wnnz_Int_t demuxWriteResult_CT$wnnz_Int_d;
  logic demuxWriteResult_CT$wnnz_Int_r;
  \Word16#_t  initHP_QTree_Int_d;
  logic initHP_QTree_Int_r;
  \Word16#_t  incrHP_QTree_Int_d;
  logic incrHP_QTree_Int_r;
  Go_t incrHP_mergeQTree_Int_d;
  logic incrHP_mergeQTree_Int_r;
  Go_t incrHP_QTree_Int1_d;
  logic incrHP_QTree_Int1_r;
  Go_t incrHP_QTree_Int2_d;
  logic incrHP_QTree_Int2_r;
  \Word16#_t  addHP_QTree_Int_d;
  logic addHP_QTree_Int_r;
  \Word16#_t  mergeHP_QTree_Int_d;
  logic mergeHP_QTree_Int_r;
  Go_t incrHP_mergeQTree_Int_buf_d;
  logic incrHP_mergeQTree_Int_buf_r;
  \Word16#_t  mergeHP_QTree_Int_buf_d;
  logic mergeHP_QTree_Int_buf_r;
  Go_t go_1_dummy_write_QTree_Int_d;
  logic go_1_dummy_write_QTree_Int_r;
  Go_t go_2_dummy_write_QTree_Int_d;
  logic go_2_dummy_write_QTree_Int_r;
  \Word16#_t  forkHP1_QTree_Int_d;
  logic forkHP1_QTree_Int_r;
  \Word16#_t  forkHP1_QTree_Int_snk_d;
  logic forkHP1_QTree_Int_snk_r;
  \Word16#_t  forkHP1_QTree_In3_d;
  logic forkHP1_QTree_In3_r;
  \Word16#_t  forkHP1_QTree_In4_d;
  logic forkHP1_QTree_In4_r;
  C2_t memMergeChoice_QTree_Int_d;
  logic memMergeChoice_QTree_Int_r;
  MemIn_QTree_Int_t memMergeIn_QTree_Int_d;
  logic memMergeIn_QTree_Int_r;
  MemOut_QTree_Int_t memOut_QTree_Int_d;
  logic memOut_QTree_Int_r;
  MemOut_QTree_Int_t memReadOut_QTree_Int_d;
  logic memReadOut_QTree_Int_r;
  MemOut_QTree_Int_t memWriteOut_QTree_Int_d;
  logic memWriteOut_QTree_Int_r;
  MemIn_QTree_Int_t memMergeIn_QTree_Int_dbuf_d;
  logic memMergeIn_QTree_Int_dbuf_r;
  MemIn_QTree_Int_t memMergeIn_QTree_Int_rbuf_d;
  logic memMergeIn_QTree_Int_rbuf_r;
  MemOut_QTree_Int_t memOut_QTree_Int_dbuf_d;
  logic memOut_QTree_Int_dbuf_r;
  MemOut_QTree_Int_t memOut_QTree_Int_rbuf_d;
  logic memOut_QTree_Int_rbuf_r;
  C4_t readMerge_choice_QTree_Int_d;
  logic readMerge_choice_QTree_Int_r;
  Pointer_QTree_Int_t readMerge_data_QTree_Int_d;
  logic readMerge_data_QTree_Int_r;
  QTree_Int_t readPointer_QTree_Intm1ad4_1_argbuf_d;
  logic readPointer_QTree_Intm1ad4_1_argbuf_r;
  QTree_Int_t readPointer_QTree_IntmacN_1_argbuf_d;
  logic readPointer_QTree_IntmacN_1_argbuf_r;
  QTree_Int_t readPointer_QTree_IntmacW_1_argbuf_d;
  logic readPointer_QTree_IntmacW_1_argbuf_r;
  QTree_Int_t readPointer_QTree_Intwsvt_1_1_argbuf_d;
  logic readPointer_QTree_Intwsvt_1_1_argbuf_r;
  \Word16#_t  destructReadIn_QTree_Int_d;
  logic destructReadIn_QTree_Int_r;
  MemIn_QTree_Int_t dconReadIn_QTree_Int_d;
  logic dconReadIn_QTree_Int_r;
  QTree_Int_t destructReadOut_QTree_Int_d;
  logic destructReadOut_QTree_Int_r;
  C14_t writeMerge_choice_QTree_Int_d;
  logic writeMerge_choice_QTree_Int_r;
  QTree_Int_t writeMerge_data_QTree_Int_d;
  logic writeMerge_data_QTree_Int_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet11_1_1_argbuf_d;
  logic writeQTree_IntlizzieLet11_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet12_1_1_argbuf_d;
  logic writeQTree_IntlizzieLet12_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet13_1_1_argbuf_d;
  logic writeQTree_IntlizzieLet13_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet15_2_1_argbuf_d;
  logic writeQTree_IntlizzieLet15_2_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet17_1_1_argbuf_d;
  logic writeQTree_IntlizzieLet17_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet18_1_argbuf_d;
  logic writeQTree_IntlizzieLet18_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet19_1_argbuf_d;
  logic writeQTree_IntlizzieLet19_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet21_1_argbuf_d;
  logic writeQTree_IntlizzieLet21_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet33_1_argbuf_d;
  logic writeQTree_IntlizzieLet33_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet38_1_argbuf_d;
  logic writeQTree_IntlizzieLet38_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet43_1_argbuf_d;
  logic writeQTree_IntlizzieLet43_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet7_1_argbuf_d;
  logic writeQTree_IntlizzieLet7_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet9_1_argbuf_d;
  logic writeQTree_IntlizzieLet9_1_argbuf_r;
  Pointer_QTree_Int_t dummy_write_QTree_Int_sink_d;
  logic dummy_write_QTree_Int_sink_r;
  MemIn_QTree_Int_t dconWriteIn_QTree_Int_d;
  logic dconWriteIn_QTree_Int_r;
  Pointer_QTree_Int_t dconPtr_QTree_Int_d;
  logic dconPtr_QTree_Int_r;
  Pointer_QTree_Int_t _38_d;
  logic _38_r;
  assign _38_r = 1'd1;
  Pointer_QTree_Int_t demuxWriteResult_QTree_Int_d;
  logic demuxWriteResult_QTree_Int_r;
  \Word16#_t  \initHP_CTmain_map'_Int_Int_d ;
  logic \initHP_CTmain_map'_Int_Int_r ;
  \Word16#_t  \incrHP_CTmain_map'_Int_Int_d ;
  logic \incrHP_CTmain_map'_Int_Int_r ;
  Go_t \incrHP_mergeCTmain_map'_Int_Int_d ;
  logic \incrHP_mergeCTmain_map'_Int_Int_r ;
  Go_t \incrHP_CTmain_map'_Int_Int1_d ;
  logic \incrHP_CTmain_map'_Int_Int1_r ;
  Go_t \incrHP_CTmain_map'_Int_Int2_d ;
  logic \incrHP_CTmain_map'_Int_Int2_r ;
  \Word16#_t  \addHP_CTmain_map'_Int_Int_d ;
  logic \addHP_CTmain_map'_Int_Int_r ;
  \Word16#_t  \mergeHP_CTmain_map'_Int_Int_d ;
  logic \mergeHP_CTmain_map'_Int_Int_r ;
  Go_t \incrHP_mergeCTmain_map'_Int_Int_buf_d ;
  logic \incrHP_mergeCTmain_map'_Int_Int_buf_r ;
  \Word16#_t  \mergeHP_CTmain_map'_Int_Int_buf_d ;
  logic \mergeHP_CTmain_map'_Int_Int_buf_r ;
  \Word16#_t  \forkHP1_CTmain_map'_Int_Int_d ;
  logic \forkHP1_CTmain_map'_Int_Int_r ;
  \Word16#_t  \forkHP1_CTmain_map'_Int_In2_d ;
  logic \forkHP1_CTmain_map'_Int_In2_r ;
  \Word16#_t  \forkHP1_CTmain_map'_Int_In3_d ;
  logic \forkHP1_CTmain_map'_Int_In3_r ;
  C2_t \memMergeChoice_CTmain_map'_Int_Int_d ;
  logic \memMergeChoice_CTmain_map'_Int_Int_r ;
  \MemIn_CTmain_map'_Int_Int_t  \memMergeIn_CTmain_map'_Int_Int_d ;
  logic \memMergeIn_CTmain_map'_Int_Int_r ;
  \MemOut_CTmain_map'_Int_Int_t  \memOut_CTmain_map'_Int_Int_d ;
  logic \memOut_CTmain_map'_Int_Int_r ;
  \MemOut_CTmain_map'_Int_Int_t  \memReadOut_CTmain_map'_Int_Int_d ;
  logic \memReadOut_CTmain_map'_Int_Int_r ;
  \MemOut_CTmain_map'_Int_Int_t  \memWriteOut_CTmain_map'_Int_Int_d ;
  logic \memWriteOut_CTmain_map'_Int_Int_r ;
  \MemIn_CTmain_map'_Int_Int_t  \memMergeIn_CTmain_map'_Int_Int_dbuf_d ;
  logic \memMergeIn_CTmain_map'_Int_Int_dbuf_r ;
  \MemIn_CTmain_map'_Int_Int_t  \memMergeIn_CTmain_map'_Int_Int_rbuf_d ;
  logic \memMergeIn_CTmain_map'_Int_Int_rbuf_r ;
  \MemOut_CTmain_map'_Int_Int_t  \memOut_CTmain_map'_Int_Int_dbuf_d ;
  logic \memOut_CTmain_map'_Int_Int_dbuf_r ;
  \MemOut_CTmain_map'_Int_Int_t  \memOut_CTmain_map'_Int_Int_rbuf_d ;
  logic \memOut_CTmain_map'_Int_Int_rbuf_r ;
  \Word16#_t  \destructReadIn_CTmain_map'_Int_Int_d ;
  logic \destructReadIn_CTmain_map'_Int_Int_r ;
  \MemIn_CTmain_map'_Int_Int_t  \dconReadIn_CTmain_map'_Int_Int_d ;
  logic \dconReadIn_CTmain_map'_Int_Int_r ;
  \CTmain_map'_Int_Int_t  \readPointer_CTmain_map'_Int_Intscfarg_0_2_1_argbuf_d ;
  logic \readPointer_CTmain_map'_Int_Intscfarg_0_2_1_argbuf_r ;
  C5_t \writeMerge_choice_CTmain_map'_Int_Int_d ;
  logic \writeMerge_choice_CTmain_map'_Int_Int_r ;
  \CTmain_map'_Int_Int_t  \writeMerge_data_CTmain_map'_Int_Int_d ;
  logic \writeMerge_data_CTmain_map'_Int_Int_r ;
  \Pointer_CTmain_map'_Int_Int_t  \writeCTmain_map'_Int_IntlizzieLet14_1_argbuf_d ;
  logic \writeCTmain_map'_Int_IntlizzieLet14_1_argbuf_r ;
  \Pointer_CTmain_map'_Int_Int_t  \writeCTmain_map'_Int_IntlizzieLet23_1_argbuf_d ;
  logic \writeCTmain_map'_Int_IntlizzieLet23_1_argbuf_r ;
  \Pointer_CTmain_map'_Int_Int_t  \writeCTmain_map'_Int_IntlizzieLet35_1_argbuf_d ;
  logic \writeCTmain_map'_Int_IntlizzieLet35_1_argbuf_r ;
  \Pointer_CTmain_map'_Int_Int_t  \writeCTmain_map'_Int_IntlizzieLet36_1_argbuf_d ;
  logic \writeCTmain_map'_Int_IntlizzieLet36_1_argbuf_r ;
  \Pointer_CTmain_map'_Int_Int_t  \writeCTmain_map'_Int_IntlizzieLet37_1_argbuf_d ;
  logic \writeCTmain_map'_Int_IntlizzieLet37_1_argbuf_r ;
  \MemIn_CTmain_map'_Int_Int_t  \dconWriteIn_CTmain_map'_Int_Int_d ;
  logic \dconWriteIn_CTmain_map'_Int_Int_r ;
  \Pointer_CTmain_map'_Int_Int_t  \dconPtr_CTmain_map'_Int_Int_d ;
  logic \dconPtr_CTmain_map'_Int_Int_r ;
  \Pointer_CTmain_map'_Int_Int_t  _37_d;
  logic _37_r;
  assign _37_r = 1'd1;
  \Pointer_CTmain_map'_Int_Int_t  \demuxWriteResult_CTmain_map'_Int_Int_d ;
  logic \demuxWriteResult_CTmain_map'_Int_Int_r ;
  \Word16#_t  \initHP_CTmap''_map''_Int_Int_Int_d ;
  logic \initHP_CTmap''_map''_Int_Int_Int_r ;
  \Word16#_t  \incrHP_CTmap''_map''_Int_Int_Int_d ;
  logic \incrHP_CTmap''_map''_Int_Int_Int_r ;
  Go_t \incrHP_mergeCTmap''_map''_Int_Int_Int_d ;
  logic \incrHP_mergeCTmap''_map''_Int_Int_Int_r ;
  Go_t \incrHP_CTmap''_map''_Int_Int_Int1_d ;
  logic \incrHP_CTmap''_map''_Int_Int_Int1_r ;
  Go_t \incrHP_CTmap''_map''_Int_Int_Int2_d ;
  logic \incrHP_CTmap''_map''_Int_Int_Int2_r ;
  \Word16#_t  \addHP_CTmap''_map''_Int_Int_Int_d ;
  logic \addHP_CTmap''_map''_Int_Int_Int_r ;
  \Word16#_t  \mergeHP_CTmap''_map''_Int_Int_Int_d ;
  logic \mergeHP_CTmap''_map''_Int_Int_Int_r ;
  Go_t \incrHP_mergeCTmap''_map''_Int_Int_Int_buf_d ;
  logic \incrHP_mergeCTmap''_map''_Int_Int_Int_buf_r ;
  \Word16#_t  \mergeHP_CTmap''_map''_Int_Int_Int_buf_d ;
  logic \mergeHP_CTmap''_map''_Int_Int_Int_buf_r ;
  \Word16#_t  \forkHP1_CTmap''_map''_Int_Int_Int_d ;
  logic \forkHP1_CTmap''_map''_Int_Int_Int_r ;
  \Word16#_t  \forkHP1_CTmap''_map''_Int_Int_In2_d ;
  logic \forkHP1_CTmap''_map''_Int_Int_In2_r ;
  \Word16#_t  \forkHP1_CTmap''_map''_Int_Int_In3_d ;
  logic \forkHP1_CTmap''_map''_Int_Int_In3_r ;
  C2_t \memMergeChoice_CTmap''_map''_Int_Int_Int_d ;
  logic \memMergeChoice_CTmap''_map''_Int_Int_Int_r ;
  \MemIn_CTmap''_map''_Int_Int_Int_t  \memMergeIn_CTmap''_map''_Int_Int_Int_d ;
  logic \memMergeIn_CTmap''_map''_Int_Int_Int_r ;
  \MemOut_CTmap''_map''_Int_Int_Int_t  \memOut_CTmap''_map''_Int_Int_Int_d ;
  logic \memOut_CTmap''_map''_Int_Int_Int_r ;
  \MemOut_CTmap''_map''_Int_Int_Int_t  \memReadOut_CTmap''_map''_Int_Int_Int_d ;
  logic \memReadOut_CTmap''_map''_Int_Int_Int_r ;
  \MemOut_CTmap''_map''_Int_Int_Int_t  \memWriteOut_CTmap''_map''_Int_Int_Int_d ;
  logic \memWriteOut_CTmap''_map''_Int_Int_Int_r ;
  \MemIn_CTmap''_map''_Int_Int_Int_t  \memMergeIn_CTmap''_map''_Int_Int_Int_dbuf_d ;
  logic \memMergeIn_CTmap''_map''_Int_Int_Int_dbuf_r ;
  \MemIn_CTmap''_map''_Int_Int_Int_t  \memMergeIn_CTmap''_map''_Int_Int_Int_rbuf_d ;
  logic \memMergeIn_CTmap''_map''_Int_Int_Int_rbuf_r ;
  \MemOut_CTmap''_map''_Int_Int_Int_t  \memOut_CTmap''_map''_Int_Int_Int_dbuf_d ;
  logic \memOut_CTmap''_map''_Int_Int_Int_dbuf_r ;
  \MemOut_CTmap''_map''_Int_Int_Int_t  \memOut_CTmap''_map''_Int_Int_Int_rbuf_d ;
  logic \memOut_CTmap''_map''_Int_Int_Int_rbuf_r ;
  \Word16#_t  \destructReadIn_CTmap''_map''_Int_Int_Int_d ;
  logic \destructReadIn_CTmap''_map''_Int_Int_Int_r ;
  \MemIn_CTmap''_map''_Int_Int_Int_t  \dconReadIn_CTmap''_map''_Int_Int_Int_d ;
  logic \dconReadIn_CTmap''_map''_Int_Int_Int_r ;
  \CTmap''_map''_Int_Int_Int_t  \readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf_d ;
  logic \readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf_r ;
  C5_t \writeMerge_choice_CTmap''_map''_Int_Int_Int_d ;
  logic \writeMerge_choice_CTmap''_map''_Int_Int_Int_r ;
  \CTmap''_map''_Int_Int_Int_t  \writeMerge_data_CTmap''_map''_Int_Int_Int_d ;
  logic \writeMerge_data_CTmap''_map''_Int_Int_Int_r ;
  \Pointer_CTmap''_map''_Int_Int_Int_t  \writeCTmap''_map''_Int_Int_IntlizzieLet20_1_argbuf_d ;
  logic \writeCTmap''_map''_Int_Int_IntlizzieLet20_1_argbuf_r ;
  \Pointer_CTmap''_map''_Int_Int_Int_t  \writeCTmap''_map''_Int_Int_IntlizzieLet24_1_argbuf_d ;
  logic \writeCTmap''_map''_Int_Int_IntlizzieLet24_1_argbuf_r ;
  \Pointer_CTmap''_map''_Int_Int_Int_t  \writeCTmap''_map''_Int_Int_IntlizzieLet40_1_argbuf_d ;
  logic \writeCTmap''_map''_Int_Int_IntlizzieLet40_1_argbuf_r ;
  \Pointer_CTmap''_map''_Int_Int_Int_t  \writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf_d ;
  logic \writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf_r ;
  \Pointer_CTmap''_map''_Int_Int_Int_t  \writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf_d ;
  logic \writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf_r ;
  \MemIn_CTmap''_map''_Int_Int_Int_t  \dconWriteIn_CTmap''_map''_Int_Int_Int_d ;
  logic \dconWriteIn_CTmap''_map''_Int_Int_Int_r ;
  \Pointer_CTmap''_map''_Int_Int_Int_t  \dconPtr_CTmap''_map''_Int_Int_Int_d ;
  logic \dconPtr_CTmap''_map''_Int_Int_Int_r ;
  \Pointer_CTmap''_map''_Int_Int_Int_t  _36_d;
  logic _36_r;
  assign _36_r = 1'd1;
  \Pointer_CTmap''_map''_Int_Int_Int_t  \demuxWriteResult_CTmap''_map''_Int_Int_Int_d ;
  logic \demuxWriteResult_CTmap''_map''_Int_Int_Int_r ;
  \Word16#_t  initHP_CTkron_kron_Int_Int_Int_d;
  logic initHP_CTkron_kron_Int_Int_Int_r;
  \Word16#_t  incrHP_CTkron_kron_Int_Int_Int_d;
  logic incrHP_CTkron_kron_Int_Int_Int_r;
  Go_t incrHP_mergeCTkron_kron_Int_Int_Int_d;
  logic incrHP_mergeCTkron_kron_Int_Int_Int_r;
  Go_t incrHP_CTkron_kron_Int_Int_Int1_d;
  logic incrHP_CTkron_kron_Int_Int_Int1_r;
  Go_t incrHP_CTkron_kron_Int_Int_Int2_d;
  logic incrHP_CTkron_kron_Int_Int_Int2_r;
  \Word16#_t  addHP_CTkron_kron_Int_Int_Int_d;
  logic addHP_CTkron_kron_Int_Int_Int_r;
  \Word16#_t  mergeHP_CTkron_kron_Int_Int_Int_d;
  logic mergeHP_CTkron_kron_Int_Int_Int_r;
  Go_t incrHP_mergeCTkron_kron_Int_Int_Int_buf_d;
  logic incrHP_mergeCTkron_kron_Int_Int_Int_buf_r;
  \Word16#_t  mergeHP_CTkron_kron_Int_Int_Int_buf_d;
  logic mergeHP_CTkron_kron_Int_Int_Int_buf_r;
  \Word16#_t  forkHP1_CTkron_kron_Int_Int_Int_d;
  logic forkHP1_CTkron_kron_Int_Int_Int_r;
  \Word16#_t  forkHP1_CTkron_kron_Int_Int_In2_d;
  logic forkHP1_CTkron_kron_Int_Int_In2_r;
  \Word16#_t  forkHP1_CTkron_kron_Int_Int_In3_d;
  logic forkHP1_CTkron_kron_Int_Int_In3_r;
  C2_t memMergeChoice_CTkron_kron_Int_Int_Int_d;
  logic memMergeChoice_CTkron_kron_Int_Int_Int_r;
  MemIn_CTkron_kron_Int_Int_Int_t memMergeIn_CTkron_kron_Int_Int_Int_d;
  logic memMergeIn_CTkron_kron_Int_Int_Int_r;
  MemOut_CTkron_kron_Int_Int_Int_t memOut_CTkron_kron_Int_Int_Int_d;
  logic memOut_CTkron_kron_Int_Int_Int_r;
  MemOut_CTkron_kron_Int_Int_Int_t memReadOut_CTkron_kron_Int_Int_Int_d;
  logic memReadOut_CTkron_kron_Int_Int_Int_r;
  MemOut_CTkron_kron_Int_Int_Int_t memWriteOut_CTkron_kron_Int_Int_Int_d;
  logic memWriteOut_CTkron_kron_Int_Int_Int_r;
  MemIn_CTkron_kron_Int_Int_Int_t memMergeIn_CTkron_kron_Int_Int_Int_dbuf_d;
  logic memMergeIn_CTkron_kron_Int_Int_Int_dbuf_r;
  MemIn_CTkron_kron_Int_Int_Int_t memMergeIn_CTkron_kron_Int_Int_Int_rbuf_d;
  logic memMergeIn_CTkron_kron_Int_Int_Int_rbuf_r;
  MemOut_CTkron_kron_Int_Int_Int_t memOut_CTkron_kron_Int_Int_Int_dbuf_d;
  logic memOut_CTkron_kron_Int_Int_Int_dbuf_r;
  MemOut_CTkron_kron_Int_Int_Int_t memOut_CTkron_kron_Int_Int_Int_rbuf_d;
  logic memOut_CTkron_kron_Int_Int_Int_rbuf_r;
  \Word16#_t  destructReadIn_CTkron_kron_Int_Int_Int_d;
  logic destructReadIn_CTkron_kron_Int_Int_Int_r;
  MemIn_CTkron_kron_Int_Int_Int_t dconReadIn_CTkron_kron_Int_Int_Int_d;
  logic dconReadIn_CTkron_kron_Int_Int_Int_r;
  CTkron_kron_Int_Int_Int_t readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf_d;
  logic readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf_r;
  C5_t writeMerge_choice_CTkron_kron_Int_Int_Int_d;
  logic writeMerge_choice_CTkron_kron_Int_Int_Int_r;
  CTkron_kron_Int_Int_Int_t writeMerge_data_CTkron_kron_Int_Int_Int_d;
  logic writeMerge_data_CTkron_kron_Int_Int_Int_r;
  Pointer_CTkron_kron_Int_Int_Int_t writeCTkron_kron_Int_Int_IntlizzieLet22_1_argbuf_d;
  logic writeCTkron_kron_Int_Int_IntlizzieLet22_1_argbuf_r;
  Pointer_CTkron_kron_Int_Int_Int_t writeCTkron_kron_Int_Int_IntlizzieLet30_1_argbuf_d;
  logic writeCTkron_kron_Int_Int_IntlizzieLet30_1_argbuf_r;
  Pointer_CTkron_kron_Int_Int_Int_t writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf_d;
  logic writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf_r;
  Pointer_CTkron_kron_Int_Int_Int_t writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf_d;
  logic writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf_r;
  Pointer_CTkron_kron_Int_Int_Int_t writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf_d;
  logic writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf_r;
  MemIn_CTkron_kron_Int_Int_Int_t dconWriteIn_CTkron_kron_Int_Int_Int_d;
  logic dconWriteIn_CTkron_kron_Int_Int_Int_r;
  Pointer_CTkron_kron_Int_Int_Int_t dconPtr_CTkron_kron_Int_Int_Int_d;
  logic dconPtr_CTkron_kron_Int_Int_Int_r;
  Pointer_CTkron_kron_Int_Int_Int_t _35_d;
  logic _35_r;
  assign _35_r = 1'd1;
  Pointer_CTkron_kron_Int_Int_Int_t demuxWriteResult_CTkron_kron_Int_Int_Int_d;
  logic demuxWriteResult_CTkron_kron_Int_Int_Int_r;
  Go_t go_1_argbuf_d;
  logic go_1_argbuf_r;
  Go_t \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intgo_7_d ;
  logic \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intgo_7_r ;
  Pointer_QTree_Int_t \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_IntwsvA_d ;
  logic \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_IntwsvA_r ;
  Pointer_QTree_Int_t \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intw1svB_d ;
  logic \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intw1svB_r ;
  Go_t go_7_1_d;
  logic go_7_1_r;
  Go_t go_7_2_d;
  logic go_7_2_r;
  Go_t go_7_3_d;
  logic go_7_3_r;
  Go_t go_7_4_d;
  logic go_7_4_r;
  Go_t go_7_5_d;
  logic go_7_5_r;
  Go_t go_7_6_d;
  logic go_7_6_r;
  Go_t go_7_7_d;
  logic go_7_7_r;
  Pointer_QTree_Int_t w1svB_1_argbuf_d;
  logic w1svB_1_argbuf_r;
  Pointer_QTree_Int_t wsvA_1_argbuf_d;
  logic wsvA_1_argbuf_r;
  Int_t \es_0_1I#_d ;
  logic \es_0_1I#_r ;
  Go_t \$wnnz_IntTupGo___Pointer_QTree_Intgo_8_d ;
  logic \$wnnz_IntTupGo___Pointer_QTree_Intgo_8_r ;
  Pointer_QTree_Int_t \$wnnz_IntTupGo___Pointer_QTree_Intwsvt_d ;
  logic \$wnnz_IntTupGo___Pointer_QTree_Intwsvt_r ;
  Go_t go_8_1_d;
  logic go_8_1_r;
  Go_t go_8_2_d;
  logic go_8_2_r;
  Pointer_QTree_Int_t wsvt_1_argbuf_d;
  logic wsvt_1_argbuf_r;
  \Int#_t  \$wmain_resbuf_d ;
  logic \$wmain_resbuf_r ;
  C2_t applyfnInt_Bool_5_choice_d;
  logic applyfnInt_Bool_5_choice_r;
  TupGo___MyDTInt_Bool___Int_t applyfnInt_Bool_5_data_d;
  logic applyfnInt_Bool_5_data_r;
  MyDTInt_Bool_t arg0_1_d;
  logic arg0_1_r;
  MyDTInt_Bool_t arg0_2_d;
  logic arg0_2_r;
  MyDTInt_Bool_t arg0_3_d;
  logic arg0_3_r;
  MyBool_t applyfnInt_Bool_5_resbuf_d;
  logic applyfnInt_Bool_5_resbuf_r;
  MyBool_t applyfnInt_Bool_5_2_argbuf_d;
  logic applyfnInt_Bool_5_2_argbuf_r;
  MyBool_t es_0_4_1_d;
  logic es_0_4_1_r;
  MyBool_t es_0_4_2_d;
  logic es_0_4_2_r;
  MyBool_t es_0_4_3_d;
  logic es_0_4_3_r;
  MyBool_t applyfnInt_Bool_5_1_d;
  logic applyfnInt_Bool_5_1_r;
  MyBool_t applyfnInt_Bool_5_2_d;
  logic applyfnInt_Bool_5_2_r;
  Go_t applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intgo_9_d;
  logic applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intgo_9_r;
  MyDTInt_Bool_t applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_d;
  logic applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_r;
  Int_t applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg1_d;
  logic applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg1_r;
  MyBool_t es_0_5_1_d;
  logic es_0_5_1_r;
  MyBool_t es_0_5_2_d;
  logic es_0_5_2_r;
  MyBool_t es_0_5_3_d;
  logic es_0_5_3_r;
  Go_t applyfnInt_Int_5TupGo___MyDTInt_Int___Intgo_10_d;
  logic applyfnInt_Int_5TupGo___MyDTInt_Int___Intgo_10_r;
  MyDTInt_Int_t applyfnInt_Int_5TupGo___MyDTInt_Int___Intarg0_2_d;
  logic applyfnInt_Int_5TupGo___MyDTInt_Int___Intarg0_2_r;
  Int_t applyfnInt_Int_5TupGo___MyDTInt_Int___Intarg1_1_d;
  logic applyfnInt_Int_5TupGo___MyDTInt_Int___Intarg1_1_r;
  MyDTInt_Int_t arg0_2_1_d;
  logic arg0_2_1_r;
  MyDTInt_Int_t arg0_2_2_d;
  logic arg0_2_2_r;
  MyDTInt_Int_t arg0_2_3_d;
  logic arg0_2_3_r;
  Int_t xacr_1_d;
  logic xacr_1_r;
  Int_t xacr_2_d;
  logic xacr_2_r;
  MyDTInt_Int_Int_t applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_4_d;
  logic applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_4_r;
  Int_t applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg2_d;
  logic applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg2_r;
  Int_t applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg1_2_d;
  logic applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg1_2_r;
  MyDTInt_Int_Int_t arg0_4_1_d;
  logic arg0_4_1_r;
  MyDTInt_Int_Int_t arg0_4_2_d;
  logic arg0_4_2_r;
  MyDTInt_Int_Int_t arg0_4_3_d;
  logic arg0_4_3_r;
  Int_t xacr_1_1_d;
  logic xacr_1_1_r;
  Int_t xacr_1_2_d;
  logic xacr_1_2_r;
  Int_t arg0_1Dcon_eqZero_d;
  logic arg0_1Dcon_eqZero_r;
  Int_t arg0_1Dcon_eqZero_1_d;
  logic arg0_1Dcon_eqZero_1_r;
  Int_t arg0_1Dcon_eqZero_2_d;
  logic arg0_1Dcon_eqZero_2_r;
  Int_t arg0_1Dcon_eqZero_3_d;
  logic arg0_1Dcon_eqZero_3_r;
  Int_t arg0_1Dcon_eqZero_4_d;
  logic arg0_1Dcon_eqZero_4_r;
  \Int#_t  x1aqk_destruct_d;
  logic x1aqk_destruct_r;
  Int_t \arg0_1Dcon_eqZero_1I#_d ;
  logic \arg0_1Dcon_eqZero_1I#_r ;
  Go_t \arg0_1Dcon_eqZero_3I#_d ;
  logic \arg0_1Dcon_eqZero_3I#_r ;
  Go_t \arg0_1Dcon_eqZero_3I#_1_d ;
  logic \arg0_1Dcon_eqZero_3I#_1_r ;
  Go_t \arg0_1Dcon_eqZero_3I#_2_d ;
  logic \arg0_1Dcon_eqZero_3I#_2_r ;
  Go_t \arg0_1Dcon_eqZero_3I#_3_d ;
  logic \arg0_1Dcon_eqZero_3I#_3_r ;
  Go_t \arg0_1Dcon_eqZero_3I#_1_argbuf_d ;
  logic \arg0_1Dcon_eqZero_3I#_1_argbuf_r ;
  \Int#_t  \arg0_1Dcon_eqZero_3I#_1_argbuf_0_d ;
  logic \arg0_1Dcon_eqZero_3I#_1_argbuf_0_r ;
  Bool_t lizzieLet1_1wild1X1h_1_Eq_d;
  logic lizzieLet1_1wild1X1h_1_Eq_r;
  Go_t \arg0_1Dcon_eqZero_3I#_2_argbuf_d ;
  logic \arg0_1Dcon_eqZero_3I#_2_argbuf_r ;
  TupGo___Bool_t boolConvert_1TupGo___Bool_1_d;
  logic boolConvert_1TupGo___Bool_1_r;
  MyBool_t lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_d;
  logic lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_r;
  Go_t arg0_2Dcon_eqZero_d;
  logic arg0_2Dcon_eqZero_r;
  Int_t arg0_2_1Dcon_main1_d;
  logic arg0_2_1Dcon_main1_r;
  Int_t arg0_2_1Dcon_main1_1_d;
  logic arg0_2_1Dcon_main1_1_r;
  Int_t arg0_2_1Dcon_main1_2_d;
  logic arg0_2_1Dcon_main1_2_r;
  Int_t arg0_2_1Dcon_main1_3_d;
  logic arg0_2_1Dcon_main1_3_r;
  Int_t arg0_2_1Dcon_main1_4_d;
  logic arg0_2_1Dcon_main1_4_r;
  \Int#_t  xaqa_destruct_d;
  logic xaqa_destruct_r;
  Int_t \arg0_2_1Dcon_main1_1I#_d ;
  logic \arg0_2_1Dcon_main1_1I#_r ;
  Go_t \arg0_2_1Dcon_main1_3I#_d ;
  logic \arg0_2_1Dcon_main1_3I#_r ;
  Go_t \arg0_2_1Dcon_main1_3I#_1_argbuf_d ;
  logic \arg0_2_1Dcon_main1_3I#_1_argbuf_r ;
  \Int#_t  \arg0_2_1Dcon_main1_3I#_1_argbuf_2_d ;
  logic \arg0_2_1Dcon_main1_3I#_1_argbuf_2_r ;
  Int_t \es_0_2_1I#_mux_d ;
  logic \es_0_2_1I#_mux_r ;
  Go_t arg0_2_2Dcon_main1_d;
  logic arg0_2_2Dcon_main1_r;
  Int_t \es_0_2_1I#_mux_mux_d ;
  logic \es_0_2_1I#_mux_mux_r ;
  MyBool_t lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_d;
  logic lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_r;
  Int_t \arg0_4_1Dcon_$fNumInt_$ctimes_d ;
  logic \arg0_4_1Dcon_$fNumInt_$ctimes_r ;
  Int_t \arg0_4_2Dcon_$fNumInt_$ctimes_d ;
  logic \arg0_4_2Dcon_$fNumInt_$ctimes_r ;
  Int_t \arg0_4_2Dcon_$fNumInt_$ctimes_1_d ;
  logic \arg0_4_2Dcon_$fNumInt_$ctimes_1_r ;
  Int_t \arg0_4_2Dcon_$fNumInt_$ctimes_2_d ;
  logic \arg0_4_2Dcon_$fNumInt_$ctimes_2_r ;
  Int_t \arg0_4_2Dcon_$fNumInt_$ctimes_3_d ;
  logic \arg0_4_2Dcon_$fNumInt_$ctimes_3_r ;
  Int_t \arg0_4_2Dcon_$fNumInt_$ctimes_4_d ;
  logic \arg0_4_2Dcon_$fNumInt_$ctimes_4_r ;
  \Int#_t  xa1m0_destruct_d;
  logic xa1m0_destruct_r;
  Int_t \arg0_4_2Dcon_$fNumInt_$ctimes_1I#_d ;
  logic \arg0_4_2Dcon_$fNumInt_$ctimes_1I#_r ;
  Int_t \arg0_4_2Dcon_$fNumInt_$ctimes_3I#_d ;
  logic \arg0_4_2Dcon_$fNumInt_$ctimes_3I#_r ;
  Int_t \arg0_4_2Dcon_$fNumInt_$ctimes_3I#_1_d ;
  logic \arg0_4_2Dcon_$fNumInt_$ctimes_3I#_1_r ;
  Int_t \arg0_4_2Dcon_$fNumInt_$ctimes_3I#_2_d ;
  logic \arg0_4_2Dcon_$fNumInt_$ctimes_3I#_2_r ;
  Int_t \arg0_4_2Dcon_$fNumInt_$ctimes_3I#_3_d ;
  logic \arg0_4_2Dcon_$fNumInt_$ctimes_3I#_3_r ;
  Int_t \arg0_4_2Dcon_$fNumInt_$ctimes_3I#_4_d ;
  logic \arg0_4_2Dcon_$fNumInt_$ctimes_3I#_4_r ;
  \Int#_t  ya1m1_destruct_d;
  logic ya1m1_destruct_r;
  Int_t \arg0_4_2Dcon_$fNumInt_$ctimes_3I#_1I#_d ;
  logic \arg0_4_2Dcon_$fNumInt_$ctimes_3I#_1I#_r ;
  \Int#_t  \arg0_4_2Dcon_$fNumInt_$ctimes_3I#_3I#_d ;
  logic \arg0_4_2Dcon_$fNumInt_$ctimes_3I#_3I#_r ;
  \Int#_t  \arg0_4_2Dcon_$fNumInt_$ctimes_3I#_3I#_1ya1m1_1_Mul32_d ;
  logic \arg0_4_2Dcon_$fNumInt_$ctimes_3I#_3I#_1ya1m1_1_Mul32_r ;
  Int_t \es_0_3_1I#_d ;
  logic \es_0_3_1I#_r ;
  Int_t \es_0_3_1I#_mux_d ;
  logic \es_0_3_1I#_mux_r ;
  Int_t \es_0_3_1I#_mux_mux_d ;
  logic \es_0_3_1I#_mux_mux_r ;
  Int_t \es_0_3_1I#_mux_mux_mux_d ;
  logic \es_0_3_1I#_mux_mux_mux_r ;
  Go_t boolConvert_1TupGo___Boolgo_1_d;
  logic boolConvert_1TupGo___Boolgo_1_r;
  Bool_t boolConvert_1TupGo___Boolbool_d;
  logic boolConvert_1TupGo___Boolbool_r;
  Bool_t bool_1_d;
  logic bool_1_r;
  Bool_t bool_2_d;
  logic bool_2_r;
  MyBool_t lizzieLet3_1_d;
  logic lizzieLet3_1_r;
  MyBool_t lizzieLet3_2_d;
  logic lizzieLet3_2_r;
  Go_t bool_1False_d;
  logic bool_1False_r;
  Go_t bool_1True_d;
  logic bool_1True_r;
  MyBool_t bool_1False_1MyFalse_d;
  logic bool_1False_1MyFalse_r;
  MyBool_t boolConvert_1_resbuf_d;
  logic boolConvert_1_resbuf_r;
  MyBool_t bool_1True_1MyTrue_d;
  logic bool_1True_1MyTrue_r;
  MyBool_t bool_1False_1MyFalsebool_1True_1MyTrue_mux_d;
  logic bool_1False_1MyFalsebool_1True_1MyTrue_mux_r;
  Go_t call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intgo_11_d;
  logic call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intgo_11_r;
  Pointer_QTree_Int_t call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intwsvt_1_d;
  logic call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intwsvt_1_r;
  Pointer_CT$wnnz_Int_t call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intsc_0_d;
  logic call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intsc_0_r;
  Go_t call_$wnnz_Int_initBufi_d;
  logic call_$wnnz_Int_initBufi_r;
  C5_t go_11_goMux_choice_d;
  logic go_11_goMux_choice_r;
  Go_t go_11_goMux_data_d;
  logic go_11_goMux_data_r;
  Go_t call_$wnnz_Int_unlockFork1_d;
  logic call_$wnnz_Int_unlockFork1_r;
  Go_t call_$wnnz_Int_unlockFork2_d;
  logic call_$wnnz_Int_unlockFork2_r;
  Go_t call_$wnnz_Int_unlockFork3_d;
  logic call_$wnnz_Int_unlockFork3_r;
  Go_t call_$wnnz_Int_initBuf_d;
  logic call_$wnnz_Int_initBuf_r;
  Go_t call_$wnnz_Int_goMux1_d;
  logic call_$wnnz_Int_goMux1_r;
  Pointer_QTree_Int_t call_$wnnz_Int_goMux2_d;
  logic call_$wnnz_Int_goMux2_r;
  Pointer_CT$wnnz_Int_t call_$wnnz_Int_goMux3_d;
  logic call_$wnnz_Int_goMux3_r;
  Go_t call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Intgo_12_d;
  logic call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Intgo_12_r;
  MyDTInt_Bool_t call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_IntisZad2_d;
  logic call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_IntisZad2_r;
  MyDTInt_Int_Int_t call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Intgad3_d;
  logic call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Intgad3_r;
  Pointer_QTree_Int_t call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Intm1ad4_d;
  logic call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Intm1ad4_r;
  Pointer_QTree_Int_t call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Intm2ad5_d;
  logic call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Intm2ad5_r;
  Pointer_CTkron_kron_Int_Int_Int_t call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Intsc_0_1_d;
  logic call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Intsc_0_1_r;
  Go_t call_kron_kron_Int_Int_Int_initBufi_d;
  logic call_kron_kron_Int_Int_Int_initBufi_r;
  C5_t go_12_goMux_choice_d;
  logic go_12_goMux_choice_r;
  Go_t go_12_goMux_data_d;
  logic go_12_goMux_data_r;
  Go_t call_kron_kron_Int_Int_Int_unlockFork1_d;
  logic call_kron_kron_Int_Int_Int_unlockFork1_r;
  Go_t call_kron_kron_Int_Int_Int_unlockFork2_d;
  logic call_kron_kron_Int_Int_Int_unlockFork2_r;
  Go_t call_kron_kron_Int_Int_Int_unlockFork3_d;
  logic call_kron_kron_Int_Int_Int_unlockFork3_r;
  Go_t call_kron_kron_Int_Int_Int_unlockFork4_d;
  logic call_kron_kron_Int_Int_Int_unlockFork4_r;
  Go_t call_kron_kron_Int_Int_Int_unlockFork5_d;
  logic call_kron_kron_Int_Int_Int_unlockFork5_r;
  Go_t call_kron_kron_Int_Int_Int_unlockFork6_d;
  logic call_kron_kron_Int_Int_Int_unlockFork6_r;
  Go_t call_kron_kron_Int_Int_Int_initBuf_d;
  logic call_kron_kron_Int_Int_Int_initBuf_r;
  Go_t call_kron_kron_Int_Int_Int_goMux1_d;
  logic call_kron_kron_Int_Int_Int_goMux1_r;
  MyDTInt_Bool_t call_kron_kron_Int_Int_Int_goMux2_d;
  logic call_kron_kron_Int_Int_Int_goMux2_r;
  MyDTInt_Int_Int_t call_kron_kron_Int_Int_Int_goMux3_d;
  logic call_kron_kron_Int_Int_Int_goMux3_r;
  Pointer_QTree_Int_t call_kron_kron_Int_Int_Int_goMux4_d;
  logic call_kron_kron_Int_Int_Int_goMux4_r;
  Pointer_QTree_Int_t call_kron_kron_Int_Int_Int_goMux5_d;
  logic call_kron_kron_Int_Int_Int_goMux5_r;
  Pointer_CTkron_kron_Int_Int_Int_t call_kron_kron_Int_Int_Int_goMux6_d;
  logic call_kron_kron_Int_Int_Int_goMux6_r;
  Go_t \call_main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Intgo_13_d ;
  logic \call_main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Intgo_13_r ;
  MyDTInt_Bool_t \call_main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int___Pointer_CTmain_map'_Int_IntisZacL_d ;
  logic \call_main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int___Pointer_CTmain_map'_Int_IntisZacL_r ;
  MyDTInt_Int_t \call_main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int___Pointer_CTmain_map'_Int_IntgacM_d ;
  logic \call_main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int___Pointer_CTmain_map'_Int_IntgacM_r ;
  Pointer_QTree_Int_t \call_main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int___Pointer_CTmain_map'_Int_IntmacN_d ;
  logic \call_main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int___Pointer_CTmain_map'_Int_IntmacN_r ;
  \Pointer_CTmain_map'_Int_Int_t  \call_main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Intsc_0_2_d ;
  logic \call_main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Intsc_0_2_r ;
  Go_t \call_main_map'_Int_Int_initBufi_d ;
  logic \call_main_map'_Int_Int_initBufi_r ;
  C5_t go_13_goMux_choice_d;
  logic go_13_goMux_choice_r;
  Go_t go_13_goMux_data_d;
  logic go_13_goMux_data_r;
  Go_t \call_main_map'_Int_Int_unlockFork1_d ;
  logic \call_main_map'_Int_Int_unlockFork1_r ;
  Go_t \call_main_map'_Int_Int_unlockFork2_d ;
  logic \call_main_map'_Int_Int_unlockFork2_r ;
  Go_t \call_main_map'_Int_Int_unlockFork3_d ;
  logic \call_main_map'_Int_Int_unlockFork3_r ;
  Go_t \call_main_map'_Int_Int_unlockFork4_d ;
  logic \call_main_map'_Int_Int_unlockFork4_r ;
  Go_t \call_main_map'_Int_Int_unlockFork5_d ;
  logic \call_main_map'_Int_Int_unlockFork5_r ;
  Go_t \call_main_map'_Int_Int_initBuf_d ;
  logic \call_main_map'_Int_Int_initBuf_r ;
  Go_t \call_main_map'_Int_Int_goMux1_d ;
  logic \call_main_map'_Int_Int_goMux1_r ;
  MyDTInt_Bool_t \call_main_map'_Int_Int_goMux2_d ;
  logic \call_main_map'_Int_Int_goMux2_r ;
  MyDTInt_Int_t \call_main_map'_Int_Int_goMux3_d ;
  logic \call_main_map'_Int_Int_goMux3_r ;
  Pointer_QTree_Int_t \call_main_map'_Int_Int_goMux4_d ;
  logic \call_main_map'_Int_Int_goMux4_r ;
  \Pointer_CTmain_map'_Int_Int_t  \call_main_map'_Int_Int_goMux5_d ;
  logic \call_main_map'_Int_Int_goMux5_r ;
  Go_t \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Intgo_14_d ;
  logic \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Intgo_14_r ;
  MyDTInt_Bool_t \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_IntisZacT_d ;
  logic \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_IntisZacT_r ;
  MyDTInt_Int_Int_t \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_IntgacU_d ;
  logic \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_IntgacU_r ;
  Int_t \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Intv'acV_d ;
  logic \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Intv'acV_r ;
  Pointer_QTree_Int_t \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_IntmacW_d ;
  logic \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_IntmacW_r ;
  \Pointer_CTmap''_map''_Int_Int_Int_t  \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Intsc_0_3_d ;
  logic \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Intsc_0_3_r ;
  Go_t \call_map''_map''_Int_Int_Int_initBufi_d ;
  logic \call_map''_map''_Int_Int_Int_initBufi_r ;
  C5_t go_14_goMux_choice_d;
  logic go_14_goMux_choice_r;
  Go_t go_14_goMux_data_d;
  logic go_14_goMux_data_r;
  Go_t \call_map''_map''_Int_Int_Int_unlockFork1_d ;
  logic \call_map''_map''_Int_Int_Int_unlockFork1_r ;
  Go_t \call_map''_map''_Int_Int_Int_unlockFork2_d ;
  logic \call_map''_map''_Int_Int_Int_unlockFork2_r ;
  Go_t \call_map''_map''_Int_Int_Int_unlockFork3_d ;
  logic \call_map''_map''_Int_Int_Int_unlockFork3_r ;
  Go_t \call_map''_map''_Int_Int_Int_unlockFork4_d ;
  logic \call_map''_map''_Int_Int_Int_unlockFork4_r ;
  Go_t \call_map''_map''_Int_Int_Int_unlockFork5_d ;
  logic \call_map''_map''_Int_Int_Int_unlockFork5_r ;
  Go_t \call_map''_map''_Int_Int_Int_unlockFork6_d ;
  logic \call_map''_map''_Int_Int_Int_unlockFork6_r ;
  Go_t \call_map''_map''_Int_Int_Int_initBuf_d ;
  logic \call_map''_map''_Int_Int_Int_initBuf_r ;
  Go_t \call_map''_map''_Int_Int_Int_goMux1_d ;
  logic \call_map''_map''_Int_Int_Int_goMux1_r ;
  MyDTInt_Bool_t \call_map''_map''_Int_Int_Int_goMux2_d ;
  logic \call_map''_map''_Int_Int_Int_goMux2_r ;
  MyDTInt_Int_Int_t \call_map''_map''_Int_Int_Int_goMux3_d ;
  logic \call_map''_map''_Int_Int_Int_goMux3_r ;
  Int_t \call_map''_map''_Int_Int_Int_goMux4_d ;
  logic \call_map''_map''_Int_Int_Int_goMux4_r ;
  Pointer_QTree_Int_t \call_map''_map''_Int_Int_Int_goMux5_d ;
  logic \call_map''_map''_Int_Int_Int_goMux5_r ;
  \Pointer_CTmap''_map''_Int_Int_Int_t  \call_map''_map''_Int_Int_Int_goMux6_d ;
  logic \call_map''_map''_Int_Int_Int_goMux6_r ;
  Int_t applyfnInt_Int_5_resbuf_d;
  logic applyfnInt_Int_5_resbuf_r;
  Int_t applyfnInt_Int_Int_5_resbuf_d;
  logic applyfnInt_Int_Int_5_resbuf_r;
  Go_t es_0_4_1MyFalse_d;
  logic es_0_4_1MyFalse_r;
  Go_t es_0_4_1MyTrue_d;
  logic es_0_4_1MyTrue_r;
  Go_t es_0_4_1MyFalse_1_argbuf_d;
  logic es_0_4_1MyFalse_1_argbuf_r;
  Go_t es_0_4_1MyTrue_1_d;
  logic es_0_4_1MyTrue_1_r;
  Go_t es_0_4_1MyTrue_2_d;
  logic es_0_4_1MyTrue_2_r;
  QTree_Int_t es_0_4_1MyTrue_1QNone_Int_d;
  logic es_0_4_1MyTrue_1QNone_Int_r;
  QTree_Int_t lizzieLet13_1_1_argbuf_d;
  logic lizzieLet13_1_1_argbuf_r;
  Go_t es_0_4_1MyTrue_2_argbuf_d;
  logic es_0_4_1MyTrue_2_argbuf_r;
  \Pointer_CTmain_map'_Int_Int_t  es_0_4_2MyFalse_d;
  logic es_0_4_2MyFalse_r;
  \Pointer_CTmain_map'_Int_Int_t  es_0_4_2MyTrue_d;
  logic es_0_4_2MyTrue_r;
  \Pointer_CTmain_map'_Int_Int_t  es_0_4_2MyFalse_1_argbuf_d;
  logic es_0_4_2MyFalse_1_argbuf_r;
  \Pointer_CTmain_map'_Int_Int_t  es_0_4_2MyTrue_1_argbuf_d;
  logic es_0_4_2MyTrue_1_argbuf_r;
  Int_t es_0_4_3MyFalse_d;
  logic es_0_4_3MyFalse_r;
  Int_t _34_d;
  logic _34_r;
  assign _34_r = 1'd1;
  QTree_Int_t es_0_4_3MyFalse_1QVal_Int_d;
  logic es_0_4_3MyFalse_1QVal_Int_r;
  QTree_Int_t lizzieLet12_1_1_argbuf_d;
  logic lizzieLet12_1_1_argbuf_r;
  Go_t es_0_5_1MyFalse_d;
  logic es_0_5_1MyFalse_r;
  Go_t es_0_5_1MyTrue_d;
  logic es_0_5_1MyTrue_r;
  Go_t es_0_5_1MyFalse_1_argbuf_d;
  logic es_0_5_1MyFalse_1_argbuf_r;
  Go_t es_0_5_1MyTrue_1_d;
  logic es_0_5_1MyTrue_1_r;
  Go_t es_0_5_1MyTrue_2_d;
  logic es_0_5_1MyTrue_2_r;
  QTree_Int_t es_0_5_1MyTrue_1QNone_Int_d;
  logic es_0_5_1MyTrue_1QNone_Int_r;
  QTree_Int_t lizzieLet19_1_argbuf_d;
  logic lizzieLet19_1_argbuf_r;
  Go_t es_0_5_1MyTrue_2_argbuf_d;
  logic es_0_5_1MyTrue_2_argbuf_r;
  \Pointer_CTmap''_map''_Int_Int_Int_t  es_0_5_2MyFalse_d;
  logic es_0_5_2MyFalse_r;
  \Pointer_CTmap''_map''_Int_Int_Int_t  es_0_5_2MyTrue_d;
  logic es_0_5_2MyTrue_r;
  \Pointer_CTmap''_map''_Int_Int_Int_t  es_0_5_2MyFalse_1_argbuf_d;
  logic es_0_5_2MyFalse_1_argbuf_r;
  \Pointer_CTmap''_map''_Int_Int_Int_t  es_0_5_2MyTrue_1_argbuf_d;
  logic es_0_5_2MyTrue_1_argbuf_r;
  Int_t es_0_5_3MyFalse_d;
  logic es_0_5_3MyFalse_r;
  Int_t _33_d;
  logic _33_r;
  assign _33_r = 1'd1;
  QTree_Int_t es_0_5_3MyFalse_1QVal_Int_d;
  logic es_0_5_3MyFalse_1QVal_Int_r;
  QTree_Int_t lizzieLet18_1_argbuf_d;
  logic lizzieLet18_1_argbuf_r;
  \Int#_t  contRet_0_1_argbuf_d;
  logic contRet_0_1_argbuf_r;
  \Int#_t  es_4_1_1lizzieLet25_4Lcall_$wnnz_Int0_1_Add32_d;
  logic es_4_1_1lizzieLet25_4Lcall_$wnnz_Int0_1_Add32_r;
  MyDTInt_Int_t gacM_2_2_argbuf_d;
  logic gacM_2_2_argbuf_r;
  MyDTInt_Int_t gacM_2_1_d;
  logic gacM_2_1_r;
  MyDTInt_Int_t gacM_2_2_d;
  logic gacM_2_2_r;
  MyDTInt_Int_t gacM_3_2_argbuf_d;
  logic gacM_3_2_argbuf_r;
  MyDTInt_Int_t gacM_3_1_d;
  logic gacM_3_1_r;
  MyDTInt_Int_t gacM_3_2_d;
  logic gacM_3_2_r;
  MyDTInt_Int_t gacM_4_1_argbuf_d;
  logic gacM_4_1_argbuf_r;
  MyDTInt_Int_Int_t gacU_2_2_argbuf_d;
  logic gacU_2_2_argbuf_r;
  MyDTInt_Int_Int_t gacU_2_1_d;
  logic gacU_2_1_r;
  MyDTInt_Int_Int_t gacU_2_2_d;
  logic gacU_2_2_r;
  MyDTInt_Int_Int_t gacU_3_2_argbuf_d;
  logic gacU_3_2_argbuf_r;
  MyDTInt_Int_Int_t gacU_3_1_d;
  logic gacU_3_1_r;
  MyDTInt_Int_Int_t gacU_3_2_d;
  logic gacU_3_2_r;
  MyDTInt_Int_Int_t gacU_4_1_argbuf_d;
  logic gacU_4_1_argbuf_r;
  MyDTInt_Int_Int_t gad3_2_2_argbuf_d;
  logic gad3_2_2_argbuf_r;
  MyDTInt_Int_Int_t gad3_2_1_d;
  logic gad3_2_1_r;
  MyDTInt_Int_Int_t gad3_2_2_d;
  logic gad3_2_2_r;
  MyDTInt_Int_Int_t gad3_3_2_argbuf_d;
  logic gad3_3_2_argbuf_r;
  MyDTInt_Int_Int_t gad3_3_1_d;
  logic gad3_3_1_r;
  MyDTInt_Int_Int_t gad3_3_2_d;
  logic gad3_3_2_r;
  MyDTInt_Int_Int_t gad3_4_1_argbuf_d;
  logic gad3_4_1_argbuf_r;
  C5_t go_11_goMux_choice_1_d;
  logic go_11_goMux_choice_1_r;
  C5_t go_11_goMux_choice_2_d;
  logic go_11_goMux_choice_2_r;
  Pointer_QTree_Int_t wsvt_1_goMux_mux_d;
  logic wsvt_1_goMux_mux_r;
  Pointer_CT$wnnz_Int_t sc_0_goMux_mux_d;
  logic sc_0_goMux_mux_r;
  C5_t go_12_goMux_choice_1_d;
  logic go_12_goMux_choice_1_r;
  C5_t go_12_goMux_choice_2_d;
  logic go_12_goMux_choice_2_r;
  C5_t go_12_goMux_choice_3_d;
  logic go_12_goMux_choice_3_r;
  C5_t go_12_goMux_choice_4_d;
  logic go_12_goMux_choice_4_r;
  C5_t go_12_goMux_choice_5_d;
  logic go_12_goMux_choice_5_r;
  MyDTInt_Bool_t isZad2_goMux_mux_d;
  logic isZad2_goMux_mux_r;
  MyDTInt_Int_Int_t gad3_goMux_mux_d;
  logic gad3_goMux_mux_r;
  Pointer_QTree_Int_t m1ad4_goMux_mux_d;
  logic m1ad4_goMux_mux_r;
  Pointer_QTree_Int_t m2ad5_goMux_mux_d;
  logic m2ad5_goMux_mux_r;
  Pointer_CTkron_kron_Int_Int_Int_t sc_0_1_goMux_mux_d;
  logic sc_0_1_goMux_mux_r;
  C5_t go_13_goMux_choice_1_d;
  logic go_13_goMux_choice_1_r;
  C5_t go_13_goMux_choice_2_d;
  logic go_13_goMux_choice_2_r;
  C5_t go_13_goMux_choice_3_d;
  logic go_13_goMux_choice_3_r;
  C5_t go_13_goMux_choice_4_d;
  logic go_13_goMux_choice_4_r;
  MyDTInt_Bool_t isZacL_goMux_mux_d;
  logic isZacL_goMux_mux_r;
  MyDTInt_Int_t gacM_goMux_mux_d;
  logic gacM_goMux_mux_r;
  Pointer_QTree_Int_t macN_goMux_mux_d;
  logic macN_goMux_mux_r;
  \Pointer_CTmain_map'_Int_Int_t  sc_0_2_goMux_mux_d;
  logic sc_0_2_goMux_mux_r;
  C5_t go_14_goMux_choice_1_d;
  logic go_14_goMux_choice_1_r;
  C5_t go_14_goMux_choice_2_d;
  logic go_14_goMux_choice_2_r;
  C5_t go_14_goMux_choice_3_d;
  logic go_14_goMux_choice_3_r;
  C5_t go_14_goMux_choice_4_d;
  logic go_14_goMux_choice_4_r;
  C5_t go_14_goMux_choice_5_d;
  logic go_14_goMux_choice_5_r;
  MyDTInt_Bool_t isZacT_goMux_mux_d;
  logic isZacT_goMux_mux_r;
  MyDTInt_Int_Int_t gacU_goMux_mux_d;
  logic gacU_goMux_mux_r;
  Int_t \v'acV_goMux_mux_d ;
  logic \v'acV_goMux_mux_r ;
  Pointer_QTree_Int_t macW_goMux_mux_d;
  logic macW_goMux_mux_r;
  \Pointer_CTmap''_map''_Int_Int_Int_t  sc_0_3_goMux_mux_d;
  logic sc_0_3_goMux_mux_r;
  CTkron_kron_Int_Int_Int_t go_15_1Lkron_kron_Int_Int_Intsbos_d;
  logic go_15_1Lkron_kron_Int_Int_Intsbos_r;
  CTkron_kron_Int_Int_Int_t lizzieLet22_1_argbuf_d;
  logic lizzieLet22_1_argbuf_r;
  Go_t go_15_2_argbuf_d;
  logic go_15_2_argbuf_r;
  TupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Int_t call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Int_1_d;
  logic call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Int_1_r;
  \CTmain_map'_Int_Int_t  \go_16_1Lmain_map'_Int_Intsbos_d ;
  logic \go_16_1Lmain_map'_Int_Intsbos_r ;
  \CTmain_map'_Int_Int_t  lizzieLet23_1_argbuf_d;
  logic lizzieLet23_1_argbuf_r;
  Go_t go_16_2_argbuf_d;
  logic go_16_2_argbuf_r;
  \TupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Int_t  \call_main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Int_1_d ;
  logic \call_main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Int_1_r ;
  \CTmap''_map''_Int_Int_Int_t  \go_17_1Lmap''_map''_Int_Int_Intsbos_d ;
  logic \go_17_1Lmap''_map''_Int_Int_Intsbos_r ;
  \CTmap''_map''_Int_Int_Int_t  lizzieLet24_1_argbuf_d;
  logic lizzieLet24_1_argbuf_r;
  Go_t go_17_2_argbuf_d;
  logic go_17_2_argbuf_r;
  \TupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Int_t  \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Int_1_d ;
  logic \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Int_1_r ;
  C4_t go_18_goMux_choice_1_d;
  logic go_18_goMux_choice_1_r;
  C4_t go_18_goMux_choice_2_d;
  logic go_18_goMux_choice_2_r;
  \Int#_t  srtarg_0_goMux_mux_d;
  logic srtarg_0_goMux_mux_r;
  Pointer_CT$wnnz_Int_t scfarg_0_goMux_mux_d;
  logic scfarg_0_goMux_mux_r;
  C4_t go_19_goMux_choice_1_d;
  logic go_19_goMux_choice_1_r;
  C4_t go_19_goMux_choice_2_d;
  logic go_19_goMux_choice_2_r;
  Pointer_QTree_Int_t srtarg_0_1_goMux_mux_d;
  logic srtarg_0_1_goMux_mux_r;
  Pointer_CTkron_kron_Int_Int_Int_t scfarg_0_1_goMux_mux_d;
  logic scfarg_0_1_goMux_mux_r;
  TupGo___Pointer_QTree_Int___Pointer_QTree_Int_t \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Int_1_d ;
  logic \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Int_1_r ;
  C5_t go_20_goMux_choice_1_d;
  logic go_20_goMux_choice_1_r;
  C5_t go_20_goMux_choice_2_d;
  logic go_20_goMux_choice_2_r;
  Pointer_QTree_Int_t srtarg_0_2_goMux_mux_d;
  logic srtarg_0_2_goMux_mux_r;
  \Pointer_CTmain_map'_Int_Int_t  scfarg_0_2_goMux_mux_d;
  logic scfarg_0_2_goMux_mux_r;
  C5_t go_21_goMux_choice_1_d;
  logic go_21_goMux_choice_1_r;
  C5_t go_21_goMux_choice_2_d;
  logic go_21_goMux_choice_2_r;
  Pointer_QTree_Int_t srtarg_0_3_goMux_mux_d;
  logic srtarg_0_3_goMux_mux_r;
  \Pointer_CTmap''_map''_Int_Int_Int_t  scfarg_0_3_goMux_mux_d;
  logic scfarg_0_3_goMux_mux_r;
  MyDTInt_Int_t go_7_1Dcon_main1_d;
  logic go_7_1Dcon_main1_r;
  MyDTInt_Int_t es_2_1_argbuf_d;
  logic es_2_1_argbuf_r;
  MyDTInt_Bool_t go_7_2Dcon_eqZero_d;
  logic go_7_2Dcon_eqZero_r;
  MyDTInt_Bool_t es_1_1_argbuf_d;
  logic es_1_1_argbuf_r;
  MyDTInt_Int_Int_t \go_7_3Dcon_$fNumInt_$ctimes_d ;
  logic \go_7_3Dcon_$fNumInt_$ctimes_r ;
  MyDTInt_Int_Int_t es_5_1_argbuf_d;
  logic es_5_1_argbuf_r;
  MyDTInt_Bool_t go_7_4Dcon_eqZero_d;
  logic go_7_4Dcon_eqZero_r;
  MyDTInt_Bool_t es_4_1_argbuf_d;
  logic es_4_1_argbuf_r;
  Go_t go_7_5_argbuf_d;
  logic go_7_5_argbuf_r;
  TupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_t kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1_d;
  logic kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1_r;
  Go_t go_7_6_argbuf_d;
  logic go_7_6_argbuf_r;
  TupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int_t \main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int_1_d ;
  logic \main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int_1_r ;
  Go_t go_7_7_argbuf_d;
  logic go_7_7_argbuf_r;
  TupGo___Pointer_QTree_Int_t \$wnnz_IntTupGo___Pointer_QTree_Int_1_d ;
  logic \$wnnz_IntTupGo___Pointer_QTree_Int_1_r ;
  CT$wnnz_Int_t go_8_1L$wnnz_Intsbos_d;
  logic go_8_1L$wnnz_Intsbos_r;
  CT$wnnz_Int_t lizzieLet0_1_argbuf_d;
  logic lizzieLet0_1_argbuf_r;
  Go_t go_8_2_argbuf_d;
  logic go_8_2_argbuf_r;
  TupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_t call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_d;
  logic call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_r;
  MyDTInt_Bool_t isZacL_2_2_argbuf_d;
  logic isZacL_2_2_argbuf_r;
  MyDTInt_Bool_t isZacL_2_1_d;
  logic isZacL_2_1_r;
  MyDTInt_Bool_t isZacL_2_2_d;
  logic isZacL_2_2_r;
  MyDTInt_Bool_t isZacL_3_2_argbuf_d;
  logic isZacL_3_2_argbuf_r;
  MyDTInt_Bool_t isZacL_3_1_d;
  logic isZacL_3_1_r;
  MyDTInt_Bool_t isZacL_3_2_d;
  logic isZacL_3_2_r;
  MyDTInt_Bool_t isZacL_4_1_argbuf_d;
  logic isZacL_4_1_argbuf_r;
  MyDTInt_Bool_t isZacT_2_2_argbuf_d;
  logic isZacT_2_2_argbuf_r;
  MyDTInt_Bool_t isZacT_2_1_d;
  logic isZacT_2_1_r;
  MyDTInt_Bool_t isZacT_2_2_d;
  logic isZacT_2_2_r;
  MyDTInt_Bool_t isZacT_3_2_argbuf_d;
  logic isZacT_3_2_argbuf_r;
  MyDTInt_Bool_t isZacT_3_1_d;
  logic isZacT_3_1_r;
  MyDTInt_Bool_t isZacT_3_2_d;
  logic isZacT_3_2_r;
  MyDTInt_Bool_t isZacT_4_1_argbuf_d;
  logic isZacT_4_1_argbuf_r;
  MyDTInt_Bool_t isZad2_2_2_argbuf_d;
  logic isZad2_2_2_argbuf_r;
  MyDTInt_Bool_t isZad2_2_1_d;
  logic isZad2_2_1_r;
  MyDTInt_Bool_t isZad2_2_2_d;
  logic isZad2_2_2_r;
  MyDTInt_Bool_t isZad2_3_2_argbuf_d;
  logic isZad2_3_2_argbuf_r;
  MyDTInt_Bool_t isZad2_3_1_d;
  logic isZad2_3_1_r;
  MyDTInt_Bool_t isZad2_3_2_d;
  logic isZad2_3_2_r;
  MyDTInt_Bool_t isZad2_4_1_argbuf_d;
  logic isZad2_4_1_argbuf_r;
  Go_t kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgo_15_d;
  logic kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgo_15_r;
  MyDTInt_Bool_t kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntisZad2_1_d;
  logic kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntisZad2_1_r;
  MyDTInt_Int_Int_t kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgad3_1_d;
  logic kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgad3_1_r;
  Pointer_QTree_Int_t kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm1ad4_1_d;
  logic kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm1ad4_1_r;
  Pointer_QTree_Int_t kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm2ad5_1_d;
  logic kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm2ad5_1_r;
  MyDTInt_Int_Int_t gad3_1_1_argbuf_d;
  logic gad3_1_1_argbuf_r;
  Go_t go_15_1_d;
  logic go_15_1_r;
  Go_t go_15_2_d;
  logic go_15_2_r;
  MyDTInt_Bool_t isZad2_1_1_argbuf_d;
  logic isZad2_1_1_argbuf_r;
  Pointer_QTree_Int_t m1ad4_1_1_argbuf_d;
  logic m1ad4_1_1_argbuf_r;
  Pointer_QTree_Int_t m2ad5_1_1_argbuf_d;
  logic m2ad5_1_1_argbuf_r;
  Pointer_QTree_Int_t es_3_1_argbuf_d;
  logic es_3_1_argbuf_r;
  Pointer_QTree_Int_t q1acP_destruct_d;
  logic q1acP_destruct_r;
  Pointer_QTree_Int_t q2acQ_destruct_d;
  logic q2acQ_destruct_r;
  Pointer_QTree_Int_t q3acR_destruct_d;
  logic q3acR_destruct_r;
  Pointer_QTree_Int_t q4acS_destruct_d;
  logic q4acS_destruct_r;
  Int_t vacO_destruct_d;
  logic vacO_destruct_r;
  QTree_Int_t _32_d;
  logic _32_r;
  assign _32_r = 1'd1;
  QTree_Int_t lizzieLet10_1QVal_Int_d;
  logic lizzieLet10_1QVal_Int_r;
  QTree_Int_t lizzieLet10_1QNode_Int_d;
  logic lizzieLet10_1QNode_Int_r;
  QTree_Int_t _31_d;
  logic _31_r;
  assign _31_r = 1'd1;
  MyDTInt_Int_t _30_d;
  logic _30_r;
  assign _30_r = 1'd1;
  MyDTInt_Int_t lizzieLet10_3QVal_Int_d;
  logic lizzieLet10_3QVal_Int_r;
  MyDTInt_Int_t lizzieLet10_3QNode_Int_d;
  logic lizzieLet10_3QNode_Int_r;
  MyDTInt_Int_t _29_d;
  logic _29_r;
  assign _29_r = 1'd1;
  MyDTInt_Int_t lizzieLet10_3QNode_Int_1_d;
  logic lizzieLet10_3QNode_Int_1_r;
  MyDTInt_Int_t lizzieLet10_3QNode_Int_2_d;
  logic lizzieLet10_3QNode_Int_2_r;
  MyDTInt_Int_t lizzieLet10_3QNode_Int_2_argbuf_d;
  logic lizzieLet10_3QNode_Int_2_argbuf_r;
  MyDTInt_Int_t lizzieLet10_3QVal_Int_1_argbuf_d;
  logic lizzieLet10_3QVal_Int_1_argbuf_r;
  Go_t lizzieLet10_4QNone_Int_d;
  logic lizzieLet10_4QNone_Int_r;
  Go_t lizzieLet10_4QVal_Int_d;
  logic lizzieLet10_4QVal_Int_r;
  Go_t lizzieLet10_4QNode_Int_d;
  logic lizzieLet10_4QNode_Int_r;
  Go_t lizzieLet10_4QError_Int_d;
  logic lizzieLet10_4QError_Int_r;
  Go_t lizzieLet10_4QError_Int_1_d;
  logic lizzieLet10_4QError_Int_1_r;
  Go_t lizzieLet10_4QError_Int_2_d;
  logic lizzieLet10_4QError_Int_2_r;
  QTree_Int_t lizzieLet10_4QError_Int_1QError_Int_d;
  logic lizzieLet10_4QError_Int_1QError_Int_r;
  QTree_Int_t lizzieLet15_2_1_argbuf_d;
  logic lizzieLet15_2_1_argbuf_r;
  Go_t lizzieLet10_4QError_Int_2_argbuf_d;
  logic lizzieLet10_4QError_Int_2_argbuf_r;
  Go_t lizzieLet10_4QNode_Int_1_argbuf_d;
  logic lizzieLet10_4QNode_Int_1_argbuf_r;
  Go_t lizzieLet10_4QNone_Int_1_d;
  logic lizzieLet10_4QNone_Int_1_r;
  Go_t lizzieLet10_4QNone_Int_2_d;
  logic lizzieLet10_4QNone_Int_2_r;
  QTree_Int_t lizzieLet10_4QNone_Int_1QNone_Int_d;
  logic lizzieLet10_4QNone_Int_1QNone_Int_r;
  QTree_Int_t lizzieLet11_1_1_argbuf_d;
  logic lizzieLet11_1_1_argbuf_r;
  Go_t lizzieLet10_4QNone_Int_2_argbuf_d;
  logic lizzieLet10_4QNone_Int_2_argbuf_r;
  C5_t go_20_goMux_choice_d;
  logic go_20_goMux_choice_r;
  Go_t go_20_goMux_data_d;
  logic go_20_goMux_data_r;
  Go_t lizzieLet10_4QVal_Int_1_d;
  logic lizzieLet10_4QVal_Int_1_r;
  Go_t lizzieLet10_4QVal_Int_2_d;
  logic lizzieLet10_4QVal_Int_2_r;
  Go_t lizzieLet10_4QVal_Int_3_d;
  logic lizzieLet10_4QVal_Int_3_r;
  Go_t lizzieLet10_4QVal_Int_1_argbuf_d;
  logic lizzieLet10_4QVal_Int_1_argbuf_r;
  TupGo___MyDTInt_Int___Int_t applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_d;
  logic applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_r;
  Go_t lizzieLet10_4QVal_Int_2_argbuf_d;
  logic lizzieLet10_4QVal_Int_2_argbuf_r;
  TupGo___MyDTInt_Bool___Int_t applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int2_d;
  logic applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int2_r;
  MyDTInt_Bool_t _28_d;
  logic _28_r;
  assign _28_r = 1'd1;
  MyDTInt_Bool_t lizzieLet10_5QVal_Int_d;
  logic lizzieLet10_5QVal_Int_r;
  MyDTInt_Bool_t lizzieLet10_5QNode_Int_d;
  logic lizzieLet10_5QNode_Int_r;
  MyDTInt_Bool_t _27_d;
  logic _27_r;
  assign _27_r = 1'd1;
  MyDTInt_Bool_t lizzieLet10_5QNode_Int_1_d;
  logic lizzieLet10_5QNode_Int_1_r;
  MyDTInt_Bool_t lizzieLet10_5QNode_Int_2_d;
  logic lizzieLet10_5QNode_Int_2_r;
  MyDTInt_Bool_t lizzieLet10_5QNode_Int_2_argbuf_d;
  logic lizzieLet10_5QNode_Int_2_argbuf_r;
  MyDTInt_Bool_t lizzieLet10_5QVal_Int_1_argbuf_d;
  logic lizzieLet10_5QVal_Int_1_argbuf_r;
  \Pointer_CTmain_map'_Int_Int_t  lizzieLet10_6QNone_Int_d;
  logic lizzieLet10_6QNone_Int_r;
  \Pointer_CTmain_map'_Int_Int_t  lizzieLet10_6QVal_Int_d;
  logic lizzieLet10_6QVal_Int_r;
  \Pointer_CTmain_map'_Int_Int_t  lizzieLet10_6QNode_Int_d;
  logic lizzieLet10_6QNode_Int_r;
  \Pointer_CTmain_map'_Int_Int_t  lizzieLet10_6QError_Int_d;
  logic lizzieLet10_6QError_Int_r;
  \Pointer_CTmain_map'_Int_Int_t  lizzieLet10_6QError_Int_1_argbuf_d;
  logic lizzieLet10_6QError_Int_1_argbuf_r;
  \CTmain_map'_Int_Int_t  \lizzieLet10_6QNode_Int_1lizzieLet10_5QNode_Int_1lizzieLet10_3QNode_Int_1q1acP_1q2acQ_1q3acR_1Lcall_main_map'_Int_Int3_d ;
  logic \lizzieLet10_6QNode_Int_1lizzieLet10_5QNode_Int_1lizzieLet10_3QNode_Int_1q1acP_1q2acQ_1q3acR_1Lcall_main_map'_Int_Int3_r ;
  \CTmain_map'_Int_Int_t  lizzieLet14_1_argbuf_d;
  logic lizzieLet14_1_argbuf_r;
  \Pointer_CTmain_map'_Int_Int_t  lizzieLet10_6QNone_Int_1_argbuf_d;
  logic lizzieLet10_6QNone_Int_1_argbuf_r;
  Pointer_QTree_Int_t q1acY_destruct_d;
  logic q1acY_destruct_r;
  Pointer_QTree_Int_t q2acZ_destruct_d;
  logic q2acZ_destruct_r;
  Pointer_QTree_Int_t q3ad0_destruct_d;
  logic q3ad0_destruct_r;
  Pointer_QTree_Int_t q4ad1_destruct_d;
  logic q4ad1_destruct_r;
  Int_t vacX_destruct_d;
  logic vacX_destruct_r;
  QTree_Int_t _26_d;
  logic _26_r;
  assign _26_r = 1'd1;
  QTree_Int_t lizzieLet16_1_1QVal_Int_d;
  logic lizzieLet16_1_1QVal_Int_r;
  QTree_Int_t lizzieLet16_1_1QNode_Int_d;
  logic lizzieLet16_1_1QNode_Int_r;
  QTree_Int_t _25_d;
  logic _25_r;
  assign _25_r = 1'd1;
  MyDTInt_Int_Int_t _24_d;
  logic _24_r;
  assign _24_r = 1'd1;
  MyDTInt_Int_Int_t lizzieLet16_1_3QVal_Int_d;
  logic lizzieLet16_1_3QVal_Int_r;
  MyDTInt_Int_Int_t lizzieLet16_1_3QNode_Int_d;
  logic lizzieLet16_1_3QNode_Int_r;
  MyDTInt_Int_Int_t _23_d;
  logic _23_r;
  assign _23_r = 1'd1;
  MyDTInt_Int_Int_t lizzieLet16_1_3QNode_Int_1_d;
  logic lizzieLet16_1_3QNode_Int_1_r;
  MyDTInt_Int_Int_t lizzieLet16_1_3QNode_Int_2_d;
  logic lizzieLet16_1_3QNode_Int_2_r;
  MyDTInt_Int_Int_t lizzieLet16_1_3QNode_Int_2_argbuf_d;
  logic lizzieLet16_1_3QNode_Int_2_argbuf_r;
  MyDTInt_Int_Int_t lizzieLet16_1_3QVal_Int_1_argbuf_d;
  logic lizzieLet16_1_3QVal_Int_1_argbuf_r;
  TupMyDTInt_Int_Int___Int___Int_t applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_d;
  logic applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_r;
  Go_t lizzieLet16_1_4QNone_Int_d;
  logic lizzieLet16_1_4QNone_Int_r;
  Go_t lizzieLet16_1_4QVal_Int_d;
  logic lizzieLet16_1_4QVal_Int_r;
  Go_t lizzieLet16_1_4QNode_Int_d;
  logic lizzieLet16_1_4QNode_Int_r;
  Go_t lizzieLet16_1_4QError_Int_d;
  logic lizzieLet16_1_4QError_Int_r;
  Go_t lizzieLet16_1_4QError_Int_1_d;
  logic lizzieLet16_1_4QError_Int_1_r;
  Go_t lizzieLet16_1_4QError_Int_2_d;
  logic lizzieLet16_1_4QError_Int_2_r;
  QTree_Int_t lizzieLet16_1_4QError_Int_1QError_Int_d;
  logic lizzieLet16_1_4QError_Int_1QError_Int_r;
  QTree_Int_t lizzieLet21_1_argbuf_d;
  logic lizzieLet21_1_argbuf_r;
  Go_t lizzieLet16_1_4QError_Int_2_argbuf_d;
  logic lizzieLet16_1_4QError_Int_2_argbuf_r;
  Go_t lizzieLet16_1_4QNode_Int_1_argbuf_d;
  logic lizzieLet16_1_4QNode_Int_1_argbuf_r;
  Go_t lizzieLet16_1_4QNone_Int_1_d;
  logic lizzieLet16_1_4QNone_Int_1_r;
  Go_t lizzieLet16_1_4QNone_Int_2_d;
  logic lizzieLet16_1_4QNone_Int_2_r;
  QTree_Int_t lizzieLet16_1_4QNone_Int_1QNone_Int_d;
  logic lizzieLet16_1_4QNone_Int_1QNone_Int_r;
  QTree_Int_t lizzieLet17_1_1_argbuf_d;
  logic lizzieLet17_1_1_argbuf_r;
  Go_t lizzieLet16_1_4QNone_Int_2_argbuf_d;
  logic lizzieLet16_1_4QNone_Int_2_argbuf_r;
  C5_t go_21_goMux_choice_d;
  logic go_21_goMux_choice_r;
  Go_t go_21_goMux_data_d;
  logic go_21_goMux_data_r;
  Go_t lizzieLet16_1_4QVal_Int_1_d;
  logic lizzieLet16_1_4QVal_Int_1_r;
  Go_t lizzieLet16_1_4QVal_Int_2_d;
  logic lizzieLet16_1_4QVal_Int_2_r;
  Go_t lizzieLet16_1_4QVal_Int_1_argbuf_d;
  logic lizzieLet16_1_4QVal_Int_1_argbuf_r;
  TupGo___MyDTInt_Bool___Int_t applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_d;
  logic applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_r;
  MyDTInt_Bool_t _22_d;
  logic _22_r;
  assign _22_r = 1'd1;
  MyDTInt_Bool_t lizzieLet16_1_5QVal_Int_d;
  logic lizzieLet16_1_5QVal_Int_r;
  MyDTInt_Bool_t lizzieLet16_1_5QNode_Int_d;
  logic lizzieLet16_1_5QNode_Int_r;
  MyDTInt_Bool_t _21_d;
  logic _21_r;
  assign _21_r = 1'd1;
  MyDTInt_Bool_t lizzieLet16_1_5QNode_Int_1_d;
  logic lizzieLet16_1_5QNode_Int_1_r;
  MyDTInt_Bool_t lizzieLet16_1_5QNode_Int_2_d;
  logic lizzieLet16_1_5QNode_Int_2_r;
  MyDTInt_Bool_t lizzieLet16_1_5QNode_Int_2_argbuf_d;
  logic lizzieLet16_1_5QNode_Int_2_argbuf_r;
  MyDTInt_Bool_t lizzieLet16_1_5QVal_Int_1_argbuf_d;
  logic lizzieLet16_1_5QVal_Int_1_argbuf_r;
  \Pointer_CTmap''_map''_Int_Int_Int_t  lizzieLet16_1_6QNone_Int_d;
  logic lizzieLet16_1_6QNone_Int_r;
  \Pointer_CTmap''_map''_Int_Int_Int_t  lizzieLet16_1_6QVal_Int_d;
  logic lizzieLet16_1_6QVal_Int_r;
  \Pointer_CTmap''_map''_Int_Int_Int_t  lizzieLet16_1_6QNode_Int_d;
  logic lizzieLet16_1_6QNode_Int_r;
  \Pointer_CTmap''_map''_Int_Int_Int_t  lizzieLet16_1_6QError_Int_d;
  logic lizzieLet16_1_6QError_Int_r;
  \Pointer_CTmap''_map''_Int_Int_Int_t  lizzieLet16_1_6QError_Int_1_argbuf_d;
  logic lizzieLet16_1_6QError_Int_1_argbuf_r;
  \CTmap''_map''_Int_Int_Int_t  \lizzieLet16_1_6QNode_Int_1lizzieLet16_1_5QNode_Int_1lizzieLet16_1_3QNode_Int_1lizzieLet16_1_7QNode_Int_1q1acY_1q2acZ_1q3ad0_1Lcall_map''_map''_Int_Int_Int3_d ;
  logic \lizzieLet16_1_6QNode_Int_1lizzieLet16_1_5QNode_Int_1lizzieLet16_1_3QNode_Int_1lizzieLet16_1_7QNode_Int_1q1acY_1q2acZ_1q3ad0_1Lcall_map''_map''_Int_Int_Int3_r ;
  \CTmap''_map''_Int_Int_Int_t  lizzieLet20_1_argbuf_d;
  logic lizzieLet20_1_argbuf_r;
  \Pointer_CTmap''_map''_Int_Int_Int_t  lizzieLet16_1_6QNone_Int_1_argbuf_d;
  logic lizzieLet16_1_6QNone_Int_1_argbuf_r;
  Int_t _20_d;
  logic _20_r;
  assign _20_r = 1'd1;
  Int_t lizzieLet16_1_7QVal_Int_d;
  logic lizzieLet16_1_7QVal_Int_r;
  Int_t lizzieLet16_1_7QNode_Int_d;
  logic lizzieLet16_1_7QNode_Int_r;
  Int_t _19_d;
  logic _19_r;
  assign _19_r = 1'd1;
  Int_t lizzieLet16_1_7QNode_Int_1_d;
  logic lizzieLet16_1_7QNode_Int_1_r;
  Int_t lizzieLet16_1_7QNode_Int_2_d;
  logic lizzieLet16_1_7QNode_Int_2_r;
  Int_t lizzieLet16_1_7QNode_Int_2_argbuf_d;
  logic lizzieLet16_1_7QNode_Int_2_argbuf_r;
  Int_t lizzieLet16_1_7QVal_Int_1_argbuf_d;
  logic lizzieLet16_1_7QVal_Int_1_argbuf_r;
  Bool_t lizzieLet2_1_argbuf_d;
  logic lizzieLet2_1_argbuf_r;
  \Int#_t  wwsvw_3_destruct_d;
  logic wwsvw_3_destruct_r;
  \Int#_t  ww1XwI_2_destruct_d;
  logic ww1XwI_2_destruct_r;
  \Int#_t  ww2XwL_1_destruct_d;
  logic ww2XwL_1_destruct_r;
  Pointer_CT$wnnz_Int_t sc_0_7_destruct_d;
  logic sc_0_7_destruct_r;
  \Int#_t  wwsvw_2_destruct_d;
  logic wwsvw_2_destruct_r;
  \Int#_t  ww1XwI_1_destruct_d;
  logic ww1XwI_1_destruct_r;
  Pointer_CT$wnnz_Int_t sc_0_6_destruct_d;
  logic sc_0_6_destruct_r;
  Pointer_QTree_Int_t q4ac3_3_destruct_d;
  logic q4ac3_3_destruct_r;
  \Int#_t  wwsvw_1_destruct_d;
  logic wwsvw_1_destruct_r;
  Pointer_CT$wnnz_Int_t sc_0_5_destruct_d;
  logic sc_0_5_destruct_r;
  Pointer_QTree_Int_t q4ac3_2_destruct_d;
  logic q4ac3_2_destruct_r;
  Pointer_QTree_Int_t q3ac2_2_destruct_d;
  logic q3ac2_2_destruct_r;
  Pointer_CT$wnnz_Int_t sc_0_4_destruct_d;
  logic sc_0_4_destruct_r;
  Pointer_QTree_Int_t q4ac3_1_destruct_d;
  logic q4ac3_1_destruct_r;
  Pointer_QTree_Int_t q3ac2_1_destruct_d;
  logic q3ac2_1_destruct_r;
  Pointer_QTree_Int_t q2ac1_1_destruct_d;
  logic q2ac1_1_destruct_r;
  CT$wnnz_Int_t _18_d;
  logic _18_r;
  assign _18_r = 1'd1;
  CT$wnnz_Int_t lizzieLet25_1Lcall_$wnnz_Int3_d;
  logic lizzieLet25_1Lcall_$wnnz_Int3_r;
  CT$wnnz_Int_t lizzieLet25_1Lcall_$wnnz_Int2_d;
  logic lizzieLet25_1Lcall_$wnnz_Int2_r;
  CT$wnnz_Int_t lizzieLet25_1Lcall_$wnnz_Int1_d;
  logic lizzieLet25_1Lcall_$wnnz_Int1_r;
  CT$wnnz_Int_t lizzieLet25_1Lcall_$wnnz_Int0_d;
  logic lizzieLet25_1Lcall_$wnnz_Int0_r;
  Go_t _17_d;
  logic _17_r;
  assign _17_r = 1'd1;
  Go_t lizzieLet25_3Lcall_$wnnz_Int3_d;
  logic lizzieLet25_3Lcall_$wnnz_Int3_r;
  Go_t lizzieLet25_3Lcall_$wnnz_Int2_d;
  logic lizzieLet25_3Lcall_$wnnz_Int2_r;
  Go_t lizzieLet25_3Lcall_$wnnz_Int1_d;
  logic lizzieLet25_3Lcall_$wnnz_Int1_r;
  Go_t lizzieLet25_3Lcall_$wnnz_Int0_d;
  logic lizzieLet25_3Lcall_$wnnz_Int0_r;
  Go_t lizzieLet25_3Lcall_$wnnz_Int0_1_argbuf_d;
  logic lizzieLet25_3Lcall_$wnnz_Int0_1_argbuf_r;
  Go_t lizzieLet25_3Lcall_$wnnz_Int1_1_argbuf_d;
  logic lizzieLet25_3Lcall_$wnnz_Int1_1_argbuf_r;
  Go_t lizzieLet25_3Lcall_$wnnz_Int2_1_argbuf_d;
  logic lizzieLet25_3Lcall_$wnnz_Int2_1_argbuf_r;
  Go_t lizzieLet25_3Lcall_$wnnz_Int3_1_argbuf_d;
  logic lizzieLet25_3Lcall_$wnnz_Int3_1_argbuf_r;
  \Int#_t  lizzieLet25_4L$wnnz_Intsbos_d;
  logic lizzieLet25_4L$wnnz_Intsbos_r;
  \Int#_t  lizzieLet25_4Lcall_$wnnz_Int3_d;
  logic lizzieLet25_4Lcall_$wnnz_Int3_r;
  \Int#_t  lizzieLet25_4Lcall_$wnnz_Int2_d;
  logic lizzieLet25_4Lcall_$wnnz_Int2_r;
  \Int#_t  lizzieLet25_4Lcall_$wnnz_Int1_d;
  logic lizzieLet25_4Lcall_$wnnz_Int1_r;
  \Int#_t  lizzieLet25_4Lcall_$wnnz_Int0_d;
  logic lizzieLet25_4Lcall_$wnnz_Int0_r;
  \Int#_t  lizzieLet25_4L$wnnz_Intsbos_1_merge_merge_fork_1_d;
  logic lizzieLet25_4L$wnnz_Intsbos_1_merge_merge_fork_1_r;
  \Int#_t  lizzieLet25_4L$wnnz_Intsbos_1_merge_merge_fork_2_d;
  logic lizzieLet25_4L$wnnz_Intsbos_1_merge_merge_fork_2_r;
  Go_t call_$wnnz_Int_goConst_d;
  logic call_$wnnz_Int_goConst_r;
  \Int#_t  \$wnnz_Int_resbuf_d ;
  logic \$wnnz_Int_resbuf_r ;
  CT$wnnz_Int_t lizzieLet25_4Lcall_$wnnz_Int3_1sc_0_4_1q4ac3_1_1q3ac2_1_1Lcall_$wnnz_Int2_d;
  logic lizzieLet25_4Lcall_$wnnz_Int3_1sc_0_4_1q4ac3_1_1q3ac2_1_1Lcall_$wnnz_Int2_r;
  CT$wnnz_Int_t lizzieLet26_1_argbuf_d;
  logic lizzieLet26_1_argbuf_r;
  Pointer_QTree_Int_t es_1_1_destruct_d;
  logic es_1_1_destruct_r;
  Pointer_QTree_Int_t es_2_2_destruct_d;
  logic es_2_2_destruct_r;
  Pointer_QTree_Int_t es_3_3_destruct_d;
  logic es_3_3_destruct_r;
  Pointer_CTkron_kron_Int_Int_Int_t sc_0_11_destruct_d;
  logic sc_0_11_destruct_r;
  Pointer_QTree_Int_t es_2_1_destruct_d;
  logic es_2_1_destruct_r;
  Pointer_QTree_Int_t es_3_2_destruct_d;
  logic es_3_2_destruct_r;
  Pointer_CTkron_kron_Int_Int_Int_t sc_0_10_destruct_d;
  logic sc_0_10_destruct_r;
  MyDTInt_Bool_t isZad2_4_destruct_d;
  logic isZad2_4_destruct_r;
  MyDTInt_Int_Int_t gad3_4_destruct_d;
  logic gad3_4_destruct_r;
  Pointer_QTree_Int_t q1ad7_3_destruct_d;
  logic q1ad7_3_destruct_r;
  Pointer_QTree_Int_t m2ad5_4_destruct_d;
  logic m2ad5_4_destruct_r;
  Pointer_QTree_Int_t es_3_1_destruct_d;
  logic es_3_1_destruct_r;
  Pointer_CTkron_kron_Int_Int_Int_t sc_0_9_destruct_d;
  logic sc_0_9_destruct_r;
  MyDTInt_Bool_t isZad2_3_destruct_d;
  logic isZad2_3_destruct_r;
  MyDTInt_Int_Int_t gad3_3_destruct_d;
  logic gad3_3_destruct_r;
  Pointer_QTree_Int_t q1ad7_2_destruct_d;
  logic q1ad7_2_destruct_r;
  Pointer_QTree_Int_t m2ad5_3_destruct_d;
  logic m2ad5_3_destruct_r;
  Pointer_QTree_Int_t q2ad8_2_destruct_d;
  logic q2ad8_2_destruct_r;
  Pointer_CTkron_kron_Int_Int_Int_t sc_0_8_destruct_d;
  logic sc_0_8_destruct_r;
  MyDTInt_Bool_t isZad2_2_destruct_d;
  logic isZad2_2_destruct_r;
  MyDTInt_Int_Int_t gad3_2_destruct_d;
  logic gad3_2_destruct_r;
  Pointer_QTree_Int_t q1ad7_1_destruct_d;
  logic q1ad7_1_destruct_r;
  Pointer_QTree_Int_t m2ad5_2_destruct_d;
  logic m2ad5_2_destruct_r;
  Pointer_QTree_Int_t q2ad8_1_destruct_d;
  logic q2ad8_1_destruct_r;
  Pointer_QTree_Int_t q3ad9_1_destruct_d;
  logic q3ad9_1_destruct_r;
  CTkron_kron_Int_Int_Int_t _16_d;
  logic _16_r;
  assign _16_r = 1'd1;
  CTkron_kron_Int_Int_Int_t lizzieLet29_1Lcall_kron_kron_Int_Int_Int3_d;
  logic lizzieLet29_1Lcall_kron_kron_Int_Int_Int3_r;
  CTkron_kron_Int_Int_Int_t lizzieLet29_1Lcall_kron_kron_Int_Int_Int2_d;
  logic lizzieLet29_1Lcall_kron_kron_Int_Int_Int2_r;
  CTkron_kron_Int_Int_Int_t lizzieLet29_1Lcall_kron_kron_Int_Int_Int1_d;
  logic lizzieLet29_1Lcall_kron_kron_Int_Int_Int1_r;
  CTkron_kron_Int_Int_Int_t lizzieLet29_1Lcall_kron_kron_Int_Int_Int0_d;
  logic lizzieLet29_1Lcall_kron_kron_Int_Int_Int0_r;
  Go_t _15_d;
  logic _15_r;
  assign _15_r = 1'd1;
  Go_t lizzieLet29_3Lcall_kron_kron_Int_Int_Int3_d;
  logic lizzieLet29_3Lcall_kron_kron_Int_Int_Int3_r;
  Go_t lizzieLet29_3Lcall_kron_kron_Int_Int_Int2_d;
  logic lizzieLet29_3Lcall_kron_kron_Int_Int_Int2_r;
  Go_t lizzieLet29_3Lcall_kron_kron_Int_Int_Int1_d;
  logic lizzieLet29_3Lcall_kron_kron_Int_Int_Int1_r;
  Go_t lizzieLet29_3Lcall_kron_kron_Int_Int_Int0_d;
  logic lizzieLet29_3Lcall_kron_kron_Int_Int_Int0_r;
  Go_t lizzieLet29_3Lcall_kron_kron_Int_Int_Int0_1_argbuf_d;
  logic lizzieLet29_3Lcall_kron_kron_Int_Int_Int0_1_argbuf_r;
  Go_t lizzieLet29_3Lcall_kron_kron_Int_Int_Int1_1_argbuf_d;
  logic lizzieLet29_3Lcall_kron_kron_Int_Int_Int1_1_argbuf_r;
  Go_t lizzieLet29_3Lcall_kron_kron_Int_Int_Int2_1_argbuf_d;
  logic lizzieLet29_3Lcall_kron_kron_Int_Int_Int2_1_argbuf_r;
  Go_t lizzieLet29_3Lcall_kron_kron_Int_Int_Int3_1_argbuf_d;
  logic lizzieLet29_3Lcall_kron_kron_Int_Int_Int3_1_argbuf_r;
  Pointer_QTree_Int_t lizzieLet29_4Lkron_kron_Int_Int_Intsbos_d;
  logic lizzieLet29_4Lkron_kron_Int_Int_Intsbos_r;
  Pointer_QTree_Int_t lizzieLet29_4Lcall_kron_kron_Int_Int_Int3_d;
  logic lizzieLet29_4Lcall_kron_kron_Int_Int_Int3_r;
  Pointer_QTree_Int_t lizzieLet29_4Lcall_kron_kron_Int_Int_Int2_d;
  logic lizzieLet29_4Lcall_kron_kron_Int_Int_Int2_r;
  Pointer_QTree_Int_t lizzieLet29_4Lcall_kron_kron_Int_Int_Int1_d;
  logic lizzieLet29_4Lcall_kron_kron_Int_Int_Int1_r;
  Pointer_QTree_Int_t lizzieLet29_4Lcall_kron_kron_Int_Int_Int0_d;
  logic lizzieLet29_4Lcall_kron_kron_Int_Int_Int0_r;
  QTree_Int_t lizzieLet29_4Lcall_kron_kron_Int_Int_Int0_1es_1_1_1es_2_2_1es_3_3_1QNode_Int_d;
  logic lizzieLet29_4Lcall_kron_kron_Int_Int_Int0_1es_1_1_1es_2_2_1es_3_3_1QNode_Int_r;
  QTree_Int_t lizzieLet33_1_argbuf_d;
  logic lizzieLet33_1_argbuf_r;
  CTkron_kron_Int_Int_Int_t lizzieLet29_4Lcall_kron_kron_Int_Int_Int1_1es_2_1_1es_3_2_1sc_0_10_1Lcall_kron_kron_Int_Int_Int0_d;
  logic lizzieLet29_4Lcall_kron_kron_Int_Int_Int1_1es_2_1_1es_3_2_1sc_0_10_1Lcall_kron_kron_Int_Int_Int0_r;
  CTkron_kron_Int_Int_Int_t lizzieLet32_1_argbuf_d;
  logic lizzieLet32_1_argbuf_r;
  CTkron_kron_Int_Int_Int_t lizzieLet29_4Lcall_kron_kron_Int_Int_Int2_1es_3_1_1sc_0_9_1isZad2_3_1gad3_3_1q1ad7_2_1m2ad5_3_1Lcall_kron_kron_Int_Int_Int1_d;
  logic lizzieLet29_4Lcall_kron_kron_Int_Int_Int2_1es_3_1_1sc_0_9_1isZad2_3_1gad3_3_1q1ad7_2_1m2ad5_3_1Lcall_kron_kron_Int_Int_Int1_r;
  CTkron_kron_Int_Int_Int_t lizzieLet31_1_argbuf_d;
  logic lizzieLet31_1_argbuf_r;
  CTkron_kron_Int_Int_Int_t lizzieLet29_4Lcall_kron_kron_Int_Int_Int3_1sc_0_8_1isZad2_2_1gad3_2_1q1ad7_1_1m2ad5_2_1q2ad8_1_1Lcall_kron_kron_Int_Int_Int2_d;
  logic lizzieLet29_4Lcall_kron_kron_Int_Int_Int3_1sc_0_8_1isZad2_2_1gad3_2_1q1ad7_1_1m2ad5_2_1q2ad8_1_1Lcall_kron_kron_Int_Int_Int2_r;
  CTkron_kron_Int_Int_Int_t lizzieLet30_1_argbuf_d;
  logic lizzieLet30_1_argbuf_r;
  Pointer_QTree_Int_t lizzieLet29_4Lkron_kron_Int_Int_Intsbos_1_merge_merge_fork_1_d;
  logic lizzieLet29_4Lkron_kron_Int_Int_Intsbos_1_merge_merge_fork_1_r;
  Pointer_QTree_Int_t lizzieLet29_4Lkron_kron_Int_Int_Intsbos_1_merge_merge_fork_2_d;
  logic lizzieLet29_4Lkron_kron_Int_Int_Intsbos_1_merge_merge_fork_2_r;
  Go_t call_kron_kron_Int_Int_Int_goConst_d;
  logic call_kron_kron_Int_Int_Int_goConst_r;
  Pointer_QTree_Int_t kron_kron_Int_Int_Int_resbuf_d;
  logic kron_kron_Int_Int_Int_resbuf_r;
  Pointer_QTree_Int_t es_2_3_destruct_d;
  logic es_2_3_destruct_r;
  Pointer_QTree_Int_t es_3_5_destruct_d;
  logic es_3_5_destruct_r;
  Pointer_QTree_Int_t es_4_4_destruct_d;
  logic es_4_4_destruct_r;
  \Pointer_CTmain_map'_Int_Int_t  sc_0_15_destruct_d;
  logic sc_0_15_destruct_r;
  Pointer_QTree_Int_t es_3_4_destruct_d;
  logic es_3_4_destruct_r;
  Pointer_QTree_Int_t es_4_3_destruct_d;
  logic es_4_3_destruct_r;
  \Pointer_CTmain_map'_Int_Int_t  sc_0_14_destruct_d;
  logic sc_0_14_destruct_r;
  MyDTInt_Bool_t isZacL_4_destruct_d;
  logic isZacL_4_destruct_r;
  MyDTInt_Int_t gacM_4_destruct_d;
  logic gacM_4_destruct_r;
  Pointer_QTree_Int_t q1acP_3_destruct_d;
  logic q1acP_3_destruct_r;
  Pointer_QTree_Int_t es_4_2_destruct_d;
  logic es_4_2_destruct_r;
  \Pointer_CTmain_map'_Int_Int_t  sc_0_13_destruct_d;
  logic sc_0_13_destruct_r;
  MyDTInt_Bool_t isZacL_3_destruct_d;
  logic isZacL_3_destruct_r;
  MyDTInt_Int_t gacM_3_destruct_d;
  logic gacM_3_destruct_r;
  Pointer_QTree_Int_t q1acP_2_destruct_d;
  logic q1acP_2_destruct_r;
  Pointer_QTree_Int_t q2acQ_2_destruct_d;
  logic q2acQ_2_destruct_r;
  \Pointer_CTmain_map'_Int_Int_t  sc_0_12_destruct_d;
  logic sc_0_12_destruct_r;
  MyDTInt_Bool_t isZacL_2_destruct_d;
  logic isZacL_2_destruct_r;
  MyDTInt_Int_t gacM_2_destruct_d;
  logic gacM_2_destruct_r;
  Pointer_QTree_Int_t q1acP_1_destruct_d;
  logic q1acP_1_destruct_r;
  Pointer_QTree_Int_t q2acQ_1_destruct_d;
  logic q2acQ_1_destruct_r;
  Pointer_QTree_Int_t q3acR_1_destruct_d;
  logic q3acR_1_destruct_r;
  \CTmain_map'_Int_Int_t  _14_d;
  logic _14_r;
  assign _14_r = 1'd1;
  \CTmain_map'_Int_Int_t  \lizzieLet34_1Lcall_main_map'_Int_Int3_d ;
  logic \lizzieLet34_1Lcall_main_map'_Int_Int3_r ;
  \CTmain_map'_Int_Int_t  \lizzieLet34_1Lcall_main_map'_Int_Int2_d ;
  logic \lizzieLet34_1Lcall_main_map'_Int_Int2_r ;
  \CTmain_map'_Int_Int_t  \lizzieLet34_1Lcall_main_map'_Int_Int1_d ;
  logic \lizzieLet34_1Lcall_main_map'_Int_Int1_r ;
  \CTmain_map'_Int_Int_t  \lizzieLet34_1Lcall_main_map'_Int_Int0_d ;
  logic \lizzieLet34_1Lcall_main_map'_Int_Int0_r ;
  Go_t _13_d;
  logic _13_r;
  assign _13_r = 1'd1;
  Go_t \lizzieLet34_3Lcall_main_map'_Int_Int3_d ;
  logic \lizzieLet34_3Lcall_main_map'_Int_Int3_r ;
  Go_t \lizzieLet34_3Lcall_main_map'_Int_Int2_d ;
  logic \lizzieLet34_3Lcall_main_map'_Int_Int2_r ;
  Go_t \lizzieLet34_3Lcall_main_map'_Int_Int1_d ;
  logic \lizzieLet34_3Lcall_main_map'_Int_Int1_r ;
  Go_t \lizzieLet34_3Lcall_main_map'_Int_Int0_d ;
  logic \lizzieLet34_3Lcall_main_map'_Int_Int0_r ;
  Go_t \lizzieLet34_3Lcall_main_map'_Int_Int0_1_argbuf_d ;
  logic \lizzieLet34_3Lcall_main_map'_Int_Int0_1_argbuf_r ;
  Go_t \lizzieLet34_3Lcall_main_map'_Int_Int1_1_argbuf_d ;
  logic \lizzieLet34_3Lcall_main_map'_Int_Int1_1_argbuf_r ;
  Go_t \lizzieLet34_3Lcall_main_map'_Int_Int2_1_argbuf_d ;
  logic \lizzieLet34_3Lcall_main_map'_Int_Int2_1_argbuf_r ;
  Go_t \lizzieLet34_3Lcall_main_map'_Int_Int3_1_argbuf_d ;
  logic \lizzieLet34_3Lcall_main_map'_Int_Int3_1_argbuf_r ;
  Pointer_QTree_Int_t \lizzieLet34_4Lmain_map'_Int_Intsbos_d ;
  logic \lizzieLet34_4Lmain_map'_Int_Intsbos_r ;
  Pointer_QTree_Int_t \lizzieLet34_4Lcall_main_map'_Int_Int3_d ;
  logic \lizzieLet34_4Lcall_main_map'_Int_Int3_r ;
  Pointer_QTree_Int_t \lizzieLet34_4Lcall_main_map'_Int_Int2_d ;
  logic \lizzieLet34_4Lcall_main_map'_Int_Int2_r ;
  Pointer_QTree_Int_t \lizzieLet34_4Lcall_main_map'_Int_Int1_d ;
  logic \lizzieLet34_4Lcall_main_map'_Int_Int1_r ;
  Pointer_QTree_Int_t \lizzieLet34_4Lcall_main_map'_Int_Int0_d ;
  logic \lizzieLet34_4Lcall_main_map'_Int_Int0_r ;
  QTree_Int_t \lizzieLet34_4Lcall_main_map'_Int_Int0_1es_2_3_1es_3_5_1es_4_4_1QNode_Int_d ;
  logic \lizzieLet34_4Lcall_main_map'_Int_Int0_1es_2_3_1es_3_5_1es_4_4_1QNode_Int_r ;
  QTree_Int_t lizzieLet38_1_argbuf_d;
  logic lizzieLet38_1_argbuf_r;
  \CTmain_map'_Int_Int_t  \lizzieLet34_4Lcall_main_map'_Int_Int1_1es_3_4_1es_4_3_1sc_0_14_1Lcall_main_map'_Int_Int0_d ;
  logic \lizzieLet34_4Lcall_main_map'_Int_Int1_1es_3_4_1es_4_3_1sc_0_14_1Lcall_main_map'_Int_Int0_r ;
  \CTmain_map'_Int_Int_t  lizzieLet37_1_argbuf_d;
  logic lizzieLet37_1_argbuf_r;
  \CTmain_map'_Int_Int_t  \lizzieLet34_4Lcall_main_map'_Int_Int2_1es_4_2_1sc_0_13_1isZacL_3_1gacM_3_1q1acP_2_1Lcall_main_map'_Int_Int1_d ;
  logic \lizzieLet34_4Lcall_main_map'_Int_Int2_1es_4_2_1sc_0_13_1isZacL_3_1gacM_3_1q1acP_2_1Lcall_main_map'_Int_Int1_r ;
  \CTmain_map'_Int_Int_t  lizzieLet36_1_argbuf_d;
  logic lizzieLet36_1_argbuf_r;
  \CTmain_map'_Int_Int_t  \lizzieLet34_4Lcall_main_map'_Int_Int3_1sc_0_12_1isZacL_2_1gacM_2_1q1acP_1_1q2acQ_1_1Lcall_main_map'_Int_Int2_d ;
  logic \lizzieLet34_4Lcall_main_map'_Int_Int3_1sc_0_12_1isZacL_2_1gacM_2_1q1acP_1_1q2acQ_1_1Lcall_main_map'_Int_Int2_r ;
  \CTmain_map'_Int_Int_t  lizzieLet35_1_argbuf_d;
  logic lizzieLet35_1_argbuf_r;
  Pointer_QTree_Int_t \lizzieLet34_4Lmain_map'_Int_Intsbos_1_merge_merge_fork_1_d ;
  logic \lizzieLet34_4Lmain_map'_Int_Intsbos_1_merge_merge_fork_1_r ;
  Pointer_QTree_Int_t \lizzieLet34_4Lmain_map'_Int_Intsbos_1_merge_merge_fork_2_d ;
  logic \lizzieLet34_4Lmain_map'_Int_Intsbos_1_merge_merge_fork_2_r ;
  Go_t \call_main_map'_Int_Int_goConst_d ;
  logic \call_main_map'_Int_Int_goConst_r ;
  Pointer_QTree_Int_t \main_map'_Int_Int_resbuf_d ;
  logic \main_map'_Int_Int_resbuf_r ;
  Pointer_QTree_Int_t es_2_4_destruct_d;
  logic es_2_4_destruct_r;
  Pointer_QTree_Int_t es_3_7_destruct_d;
  logic es_3_7_destruct_r;
  Pointer_QTree_Int_t es_4_7_destruct_d;
  logic es_4_7_destruct_r;
  \Pointer_CTmap''_map''_Int_Int_Int_t  sc_0_19_destruct_d;
  logic sc_0_19_destruct_r;
  Pointer_QTree_Int_t es_3_6_destruct_d;
  logic es_3_6_destruct_r;
  Pointer_QTree_Int_t es_4_6_destruct_d;
  logic es_4_6_destruct_r;
  \Pointer_CTmap''_map''_Int_Int_Int_t  sc_0_18_destruct_d;
  logic sc_0_18_destruct_r;
  MyDTInt_Bool_t isZacT_4_destruct_d;
  logic isZacT_4_destruct_r;
  MyDTInt_Int_Int_t gacU_4_destruct_d;
  logic gacU_4_destruct_r;
  Int_t \v'acV_4_destruct_d ;
  logic \v'acV_4_destruct_r ;
  Pointer_QTree_Int_t q1acY_3_destruct_d;
  logic q1acY_3_destruct_r;
  Pointer_QTree_Int_t es_4_5_destruct_d;
  logic es_4_5_destruct_r;
  \Pointer_CTmap''_map''_Int_Int_Int_t  sc_0_17_destruct_d;
  logic sc_0_17_destruct_r;
  MyDTInt_Bool_t isZacT_3_destruct_d;
  logic isZacT_3_destruct_r;
  MyDTInt_Int_Int_t gacU_3_destruct_d;
  logic gacU_3_destruct_r;
  Int_t \v'acV_3_destruct_d ;
  logic \v'acV_3_destruct_r ;
  Pointer_QTree_Int_t q1acY_2_destruct_d;
  logic q1acY_2_destruct_r;
  Pointer_QTree_Int_t q2acZ_2_destruct_d;
  logic q2acZ_2_destruct_r;
  \Pointer_CTmap''_map''_Int_Int_Int_t  sc_0_16_destruct_d;
  logic sc_0_16_destruct_r;
  MyDTInt_Bool_t isZacT_2_destruct_d;
  logic isZacT_2_destruct_r;
  MyDTInt_Int_Int_t gacU_2_destruct_d;
  logic gacU_2_destruct_r;
  Int_t \v'acV_2_destruct_d ;
  logic \v'acV_2_destruct_r ;
  Pointer_QTree_Int_t q1acY_1_destruct_d;
  logic q1acY_1_destruct_r;
  Pointer_QTree_Int_t q2acZ_1_destruct_d;
  logic q2acZ_1_destruct_r;
  Pointer_QTree_Int_t q3ad0_1_destruct_d;
  logic q3ad0_1_destruct_r;
  \CTmap''_map''_Int_Int_Int_t  _12_d;
  logic _12_r;
  assign _12_r = 1'd1;
  \CTmap''_map''_Int_Int_Int_t  \lizzieLet39_1Lcall_map''_map''_Int_Int_Int3_d ;
  logic \lizzieLet39_1Lcall_map''_map''_Int_Int_Int3_r ;
  \CTmap''_map''_Int_Int_Int_t  \lizzieLet39_1Lcall_map''_map''_Int_Int_Int2_d ;
  logic \lizzieLet39_1Lcall_map''_map''_Int_Int_Int2_r ;
  \CTmap''_map''_Int_Int_Int_t  \lizzieLet39_1Lcall_map''_map''_Int_Int_Int1_d ;
  logic \lizzieLet39_1Lcall_map''_map''_Int_Int_Int1_r ;
  \CTmap''_map''_Int_Int_Int_t  \lizzieLet39_1Lcall_map''_map''_Int_Int_Int0_d ;
  logic \lizzieLet39_1Lcall_map''_map''_Int_Int_Int0_r ;
  Go_t _11_d;
  logic _11_r;
  assign _11_r = 1'd1;
  Go_t \lizzieLet39_3Lcall_map''_map''_Int_Int_Int3_d ;
  logic \lizzieLet39_3Lcall_map''_map''_Int_Int_Int3_r ;
  Go_t \lizzieLet39_3Lcall_map''_map''_Int_Int_Int2_d ;
  logic \lizzieLet39_3Lcall_map''_map''_Int_Int_Int2_r ;
  Go_t \lizzieLet39_3Lcall_map''_map''_Int_Int_Int1_d ;
  logic \lizzieLet39_3Lcall_map''_map''_Int_Int_Int1_r ;
  Go_t \lizzieLet39_3Lcall_map''_map''_Int_Int_Int0_d ;
  logic \lizzieLet39_3Lcall_map''_map''_Int_Int_Int0_r ;
  Go_t \lizzieLet39_3Lcall_map''_map''_Int_Int_Int0_1_argbuf_d ;
  logic \lizzieLet39_3Lcall_map''_map''_Int_Int_Int0_1_argbuf_r ;
  Go_t \lizzieLet39_3Lcall_map''_map''_Int_Int_Int1_1_argbuf_d ;
  logic \lizzieLet39_3Lcall_map''_map''_Int_Int_Int1_1_argbuf_r ;
  Go_t \lizzieLet39_3Lcall_map''_map''_Int_Int_Int2_1_argbuf_d ;
  logic \lizzieLet39_3Lcall_map''_map''_Int_Int_Int2_1_argbuf_r ;
  Go_t \lizzieLet39_3Lcall_map''_map''_Int_Int_Int3_1_argbuf_d ;
  logic \lizzieLet39_3Lcall_map''_map''_Int_Int_Int3_1_argbuf_r ;
  Pointer_QTree_Int_t \lizzieLet39_4Lmap''_map''_Int_Int_Intsbos_d ;
  logic \lizzieLet39_4Lmap''_map''_Int_Int_Intsbos_r ;
  Pointer_QTree_Int_t \lizzieLet39_4Lcall_map''_map''_Int_Int_Int3_d ;
  logic \lizzieLet39_4Lcall_map''_map''_Int_Int_Int3_r ;
  Pointer_QTree_Int_t \lizzieLet39_4Lcall_map''_map''_Int_Int_Int2_d ;
  logic \lizzieLet39_4Lcall_map''_map''_Int_Int_Int2_r ;
  Pointer_QTree_Int_t \lizzieLet39_4Lcall_map''_map''_Int_Int_Int1_d ;
  logic \lizzieLet39_4Lcall_map''_map''_Int_Int_Int1_r ;
  Pointer_QTree_Int_t \lizzieLet39_4Lcall_map''_map''_Int_Int_Int0_d ;
  logic \lizzieLet39_4Lcall_map''_map''_Int_Int_Int0_r ;
  QTree_Int_t \lizzieLet39_4Lcall_map''_map''_Int_Int_Int0_1es_2_4_1es_3_7_1es_4_7_1QNode_Int_d ;
  logic \lizzieLet39_4Lcall_map''_map''_Int_Int_Int0_1es_2_4_1es_3_7_1es_4_7_1QNode_Int_r ;
  QTree_Int_t lizzieLet43_1_argbuf_d;
  logic lizzieLet43_1_argbuf_r;
  \CTmap''_map''_Int_Int_Int_t  \lizzieLet39_4Lcall_map''_map''_Int_Int_Int1_1es_3_6_1es_4_6_1sc_0_18_1Lcall_map''_map''_Int_Int_Int0_d ;
  logic \lizzieLet39_4Lcall_map''_map''_Int_Int_Int1_1es_3_6_1es_4_6_1sc_0_18_1Lcall_map''_map''_Int_Int_Int0_r ;
  \CTmap''_map''_Int_Int_Int_t  lizzieLet42_1_argbuf_d;
  logic lizzieLet42_1_argbuf_r;
  \CTmap''_map''_Int_Int_Int_t  \lizzieLet39_4Lcall_map''_map''_Int_Int_Int2_1es_4_5_1sc_0_17_1isZacT_3_1gacU_3_1v'acV_3_1q1acY_2_1Lcall_map''_map''_Int_Int_Int1_d ;
  logic \lizzieLet39_4Lcall_map''_map''_Int_Int_Int2_1es_4_5_1sc_0_17_1isZacT_3_1gacU_3_1v'acV_3_1q1acY_2_1Lcall_map''_map''_Int_Int_Int1_r ;
  \CTmap''_map''_Int_Int_Int_t  lizzieLet41_1_argbuf_d;
  logic lizzieLet41_1_argbuf_r;
  \CTmap''_map''_Int_Int_Int_t  \lizzieLet39_4Lcall_map''_map''_Int_Int_Int3_1sc_0_16_1isZacT_2_1gacU_2_1v'acV_2_1q1acY_1_1q2acZ_1_1Lcall_map''_map''_Int_Int_Int2_d ;
  logic \lizzieLet39_4Lcall_map''_map''_Int_Int_Int3_1sc_0_16_1isZacT_2_1gacU_2_1v'acV_2_1q1acY_1_1q2acZ_1_1Lcall_map''_map''_Int_Int_Int2_r ;
  \CTmap''_map''_Int_Int_Int_t  lizzieLet40_1_argbuf_d;
  logic lizzieLet40_1_argbuf_r;
  Pointer_QTree_Int_t \lizzieLet39_4Lmap''_map''_Int_Int_Intsbos_1_merge_merge_fork_1_d ;
  logic \lizzieLet39_4Lmap''_map''_Int_Int_Intsbos_1_merge_merge_fork_1_r ;
  Pointer_QTree_Int_t \lizzieLet39_4Lmap''_map''_Int_Int_Intsbos_1_merge_merge_fork_2_d ;
  logic \lizzieLet39_4Lmap''_map''_Int_Int_Intsbos_1_merge_merge_fork_2_r ;
  Go_t \call_map''_map''_Int_Int_Int_goConst_d ;
  logic \call_map''_map''_Int_Int_Int_goConst_r ;
  Pointer_QTree_Int_t \map''_map''_Int_Int_Int_resbuf_d ;
  logic \map''_map''_Int_Int_Int_resbuf_r ;
  Go_t lizzieLet3_1MyFalse_d;
  logic lizzieLet3_1MyFalse_r;
  Go_t lizzieLet3_1MyTrue_d;
  logic lizzieLet3_1MyTrue_r;
  MyBool_t lizzieLet3_1MyFalse_1MyFalse_d;
  logic lizzieLet3_1MyFalse_1MyFalse_r;
  MyBool_t lizzieLet3_1MyTrue_1MyTrue_d;
  logic lizzieLet3_1MyTrue_1MyTrue_r;
  MyBool_t lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_d;
  logic lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_r;
  Pointer_QTree_Int_t q1ac0_destruct_d;
  logic q1ac0_destruct_r;
  Pointer_QTree_Int_t q2ac1_destruct_d;
  logic q2ac1_destruct_r;
  Pointer_QTree_Int_t q3ac2_destruct_d;
  logic q3ac2_destruct_r;
  Pointer_QTree_Int_t q4ac3_destruct_d;
  logic q4ac3_destruct_r;
  QTree_Int_t _10_d;
  logic _10_r;
  assign _10_r = 1'd1;
  QTree_Int_t _9_d;
  logic _9_r;
  assign _9_r = 1'd1;
  QTree_Int_t lizzieLet4_1QNode_Int_d;
  logic lizzieLet4_1QNode_Int_r;
  QTree_Int_t _8_d;
  logic _8_r;
  assign _8_r = 1'd1;
  Go_t lizzieLet4_3QNone_Int_d;
  logic lizzieLet4_3QNone_Int_r;
  Go_t lizzieLet4_3QVal_Int_d;
  logic lizzieLet4_3QVal_Int_r;
  Go_t lizzieLet4_3QNode_Int_d;
  logic lizzieLet4_3QNode_Int_r;
  Go_t lizzieLet4_3QError_Int_d;
  logic lizzieLet4_3QError_Int_r;
  Go_t lizzieLet4_3QError_Int_1_d;
  logic lizzieLet4_3QError_Int_1_r;
  Go_t lizzieLet4_3QError_Int_2_d;
  logic lizzieLet4_3QError_Int_2_r;
  Go_t lizzieLet4_3QError_Int_1_argbuf_d;
  logic lizzieLet4_3QError_Int_1_argbuf_r;
  \Int#_t  lizzieLet4_3QError_Int_1_argbuf_0_d;
  logic lizzieLet4_3QError_Int_1_argbuf_0_r;
  \Int#_t  lizzieLet15_1_1_argbuf_d;
  logic lizzieLet15_1_1_argbuf_r;
  Go_t lizzieLet4_3QError_Int_2_argbuf_d;
  logic lizzieLet4_3QError_Int_2_argbuf_r;
  Go_t lizzieLet4_3QNode_Int_1_argbuf_d;
  logic lizzieLet4_3QNode_Int_1_argbuf_r;
  Go_t lizzieLet4_3QNone_Int_1_d;
  logic lizzieLet4_3QNone_Int_1_r;
  Go_t lizzieLet4_3QNone_Int_2_d;
  logic lizzieLet4_3QNone_Int_2_r;
  Go_t lizzieLet4_3QNone_Int_1_argbuf_d;
  logic lizzieLet4_3QNone_Int_1_argbuf_r;
  \Int#_t  lizzieLet4_3QNone_Int_1_argbuf_0_d;
  logic lizzieLet4_3QNone_Int_1_argbuf_0_r;
  \Int#_t  lizzieLet15_1_argbuf_d;
  logic lizzieLet15_1_argbuf_r;
  Go_t lizzieLet4_3QNone_Int_2_argbuf_d;
  logic lizzieLet4_3QNone_Int_2_argbuf_r;
  C4_t go_18_goMux_choice_d;
  logic go_18_goMux_choice_r;
  Go_t go_18_goMux_data_d;
  logic go_18_goMux_data_r;
  Go_t lizzieLet4_3QVal_Int_1_d;
  logic lizzieLet4_3QVal_Int_1_r;
  Go_t lizzieLet4_3QVal_Int_2_d;
  logic lizzieLet4_3QVal_Int_2_r;
  Go_t lizzieLet4_3QVal_Int_1_argbuf_d;
  logic lizzieLet4_3QVal_Int_1_argbuf_r;
  \Int#_t  lizzieLet4_3QVal_Int_1_argbuf_1_d;
  logic lizzieLet4_3QVal_Int_1_argbuf_1_r;
  \Int#_t  lizzieLet16_1_argbuf_d;
  logic lizzieLet16_1_argbuf_r;
  Go_t lizzieLet4_3QVal_Int_2_argbuf_d;
  logic lizzieLet4_3QVal_Int_2_argbuf_r;
  Pointer_CT$wnnz_Int_t lizzieLet4_4QNone_Int_d;
  logic lizzieLet4_4QNone_Int_r;
  Pointer_CT$wnnz_Int_t lizzieLet4_4QVal_Int_d;
  logic lizzieLet4_4QVal_Int_r;
  Pointer_CT$wnnz_Int_t lizzieLet4_4QNode_Int_d;
  logic lizzieLet4_4QNode_Int_r;
  Pointer_CT$wnnz_Int_t lizzieLet4_4QError_Int_d;
  logic lizzieLet4_4QError_Int_r;
  Pointer_CT$wnnz_Int_t lizzieLet4_4QError_Int_1_argbuf_d;
  logic lizzieLet4_4QError_Int_1_argbuf_r;
  CT$wnnz_Int_t lizzieLet4_4QNode_Int_1q4ac3_1q3ac2_1q2ac1_1Lcall_$wnnz_Int3_d;
  logic lizzieLet4_4QNode_Int_1q4ac3_1q3ac2_1q2ac1_1Lcall_$wnnz_Int3_r;
  CT$wnnz_Int_t lizzieLet5_1_argbuf_d;
  logic lizzieLet5_1_argbuf_r;
  Pointer_CT$wnnz_Int_t lizzieLet4_4QNone_Int_1_argbuf_d;
  logic lizzieLet4_4QNone_Int_1_argbuf_r;
  Pointer_CT$wnnz_Int_t lizzieLet4_4QVal_Int_1_argbuf_d;
  logic lizzieLet4_4QVal_Int_1_argbuf_r;
  Pointer_QTree_Int_t q1ad7_destruct_d;
  logic q1ad7_destruct_r;
  Pointer_QTree_Int_t q2ad8_destruct_d;
  logic q2ad8_destruct_r;
  Pointer_QTree_Int_t q3ad9_destruct_d;
  logic q3ad9_destruct_r;
  Pointer_QTree_Int_t q4ada_destruct_d;
  logic q4ada_destruct_r;
  Int_t vad6_destruct_d;
  logic vad6_destruct_r;
  QTree_Int_t _7_d;
  logic _7_r;
  assign _7_r = 1'd1;
  QTree_Int_t lizzieLet6_1QVal_Int_d;
  logic lizzieLet6_1QVal_Int_r;
  QTree_Int_t lizzieLet6_1QNode_Int_d;
  logic lizzieLet6_1QNode_Int_r;
  QTree_Int_t _6_d;
  logic _6_r;
  assign _6_r = 1'd1;
  MyDTInt_Int_Int_t _5_d;
  logic _5_r;
  assign _5_r = 1'd1;
  MyDTInt_Int_Int_t lizzieLet6_3QVal_Int_d;
  logic lizzieLet6_3QVal_Int_r;
  MyDTInt_Int_Int_t lizzieLet6_3QNode_Int_d;
  logic lizzieLet6_3QNode_Int_r;
  MyDTInt_Int_Int_t _4_d;
  logic _4_r;
  assign _4_r = 1'd1;
  MyDTInt_Int_Int_t lizzieLet6_3QNode_Int_1_d;
  logic lizzieLet6_3QNode_Int_1_r;
  MyDTInt_Int_Int_t lizzieLet6_3QNode_Int_2_d;
  logic lizzieLet6_3QNode_Int_2_r;
  MyDTInt_Int_Int_t lizzieLet6_3QNode_Int_2_argbuf_d;
  logic lizzieLet6_3QNode_Int_2_argbuf_r;
  MyDTInt_Int_Int_t lizzieLet6_3QVal_Int_1_argbuf_d;
  logic lizzieLet6_3QVal_Int_1_argbuf_r;
  Go_t lizzieLet6_4QNone_Int_d;
  logic lizzieLet6_4QNone_Int_r;
  Go_t lizzieLet6_4QVal_Int_d;
  logic lizzieLet6_4QVal_Int_r;
  Go_t lizzieLet6_4QNode_Int_d;
  logic lizzieLet6_4QNode_Int_r;
  Go_t lizzieLet6_4QError_Int_d;
  logic lizzieLet6_4QError_Int_r;
  Go_t lizzieLet6_4QError_Int_1_d;
  logic lizzieLet6_4QError_Int_1_r;
  Go_t lizzieLet6_4QError_Int_2_d;
  logic lizzieLet6_4QError_Int_2_r;
  QTree_Int_t lizzieLet6_4QError_Int_1QError_Int_d;
  logic lizzieLet6_4QError_Int_1QError_Int_r;
  QTree_Int_t lizzieLet9_1_argbuf_d;
  logic lizzieLet9_1_argbuf_r;
  Go_t lizzieLet6_4QError_Int_2_argbuf_d;
  logic lizzieLet6_4QError_Int_2_argbuf_r;
  Go_t lizzieLet6_4QNode_Int_1_argbuf_d;
  logic lizzieLet6_4QNode_Int_1_argbuf_r;
  Go_t lizzieLet6_4QNone_Int_1_d;
  logic lizzieLet6_4QNone_Int_1_r;
  Go_t lizzieLet6_4QNone_Int_2_d;
  logic lizzieLet6_4QNone_Int_2_r;
  QTree_Int_t lizzieLet6_4QNone_Int_1QNone_Int_d;
  logic lizzieLet6_4QNone_Int_1QNone_Int_r;
  QTree_Int_t lizzieLet7_1_argbuf_d;
  logic lizzieLet7_1_argbuf_r;
  Go_t lizzieLet6_4QNone_Int_2_argbuf_d;
  logic lizzieLet6_4QNone_Int_2_argbuf_r;
  C4_t go_19_goMux_choice_d;
  logic go_19_goMux_choice_r;
  Go_t go_19_goMux_data_d;
  logic go_19_goMux_data_r;
  Go_t lizzieLet6_4QVal_Int_1_d;
  logic lizzieLet6_4QVal_Int_1_r;
  Go_t lizzieLet6_4QVal_Int_2_d;
  logic lizzieLet6_4QVal_Int_2_r;
  Go_t lizzieLet6_4QVal_Int_1_argbuf_d;
  logic lizzieLet6_4QVal_Int_1_argbuf_r;
  TupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int_t \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int_1_d ;
  logic \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int_1_r ;
  Go_t lizzieLet6_4QVal_Int_2_argbuf_d;
  logic lizzieLet6_4QVal_Int_2_argbuf_r;
  MyDTInt_Bool_t _3_d;
  logic _3_r;
  assign _3_r = 1'd1;
  MyDTInt_Bool_t lizzieLet6_5QVal_Int_d;
  logic lizzieLet6_5QVal_Int_r;
  MyDTInt_Bool_t lizzieLet6_5QNode_Int_d;
  logic lizzieLet6_5QNode_Int_r;
  MyDTInt_Bool_t _2_d;
  logic _2_r;
  assign _2_r = 1'd1;
  MyDTInt_Bool_t lizzieLet6_5QNode_Int_1_d;
  logic lizzieLet6_5QNode_Int_1_r;
  MyDTInt_Bool_t lizzieLet6_5QNode_Int_2_d;
  logic lizzieLet6_5QNode_Int_2_r;
  MyDTInt_Bool_t lizzieLet6_5QNode_Int_2_argbuf_d;
  logic lizzieLet6_5QNode_Int_2_argbuf_r;
  MyDTInt_Bool_t lizzieLet6_5QVal_Int_1_argbuf_d;
  logic lizzieLet6_5QVal_Int_1_argbuf_r;
  Pointer_QTree_Int_t _1_d;
  logic _1_r;
  assign _1_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet6_6QVal_Int_d;
  logic lizzieLet6_6QVal_Int_r;
  Pointer_QTree_Int_t lizzieLet6_6QNode_Int_d;
  logic lizzieLet6_6QNode_Int_r;
  Pointer_QTree_Int_t _0_d;
  logic _0_r;
  assign _0_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet6_6QNode_Int_1_d;
  logic lizzieLet6_6QNode_Int_1_r;
  Pointer_QTree_Int_t lizzieLet6_6QNode_Int_2_d;
  logic lizzieLet6_6QNode_Int_2_r;
  Pointer_QTree_Int_t lizzieLet6_6QNode_Int_2_argbuf_d;
  logic lizzieLet6_6QNode_Int_2_argbuf_r;
  Pointer_QTree_Int_t lizzieLet6_6QVal_Int_1_argbuf_d;
  logic lizzieLet6_6QVal_Int_1_argbuf_r;
  Pointer_CTkron_kron_Int_Int_Int_t lizzieLet6_7QNone_Int_d;
  logic lizzieLet6_7QNone_Int_r;
  Pointer_CTkron_kron_Int_Int_Int_t lizzieLet6_7QVal_Int_d;
  logic lizzieLet6_7QVal_Int_r;
  Pointer_CTkron_kron_Int_Int_Int_t lizzieLet6_7QNode_Int_d;
  logic lizzieLet6_7QNode_Int_r;
  Pointer_CTkron_kron_Int_Int_Int_t lizzieLet6_7QError_Int_d;
  logic lizzieLet6_7QError_Int_r;
  Pointer_CTkron_kron_Int_Int_Int_t lizzieLet6_7QError_Int_1_argbuf_d;
  logic lizzieLet6_7QError_Int_1_argbuf_r;
  CTkron_kron_Int_Int_Int_t lizzieLet6_7QNode_Int_1lizzieLet6_5QNode_Int_1lizzieLet6_3QNode_Int_1q1ad7_1lizzieLet6_6QNode_Int_1q2ad8_1q3ad9_1Lcall_kron_kron_Int_Int_Int3_d;
  logic lizzieLet6_7QNode_Int_1lizzieLet6_5QNode_Int_1lizzieLet6_3QNode_Int_1q1ad7_1lizzieLet6_6QNode_Int_1q2ad8_1q3ad9_1Lcall_kron_kron_Int_Int_Int3_r;
  CTkron_kron_Int_Int_Int_t lizzieLet8_1_argbuf_d;
  logic lizzieLet8_1_argbuf_r;
  Pointer_CTkron_kron_Int_Int_Int_t lizzieLet6_7QNone_Int_1_argbuf_d;
  logic lizzieLet6_7QNone_Int_1_argbuf_r;
  Pointer_CTkron_kron_Int_Int_Int_t lizzieLet6_7QVal_Int_1_argbuf_d;
  logic lizzieLet6_7QVal_Int_1_argbuf_r;
  Pointer_QTree_Int_t m1ad4_1_argbuf_d;
  logic m1ad4_1_argbuf_r;
  Pointer_QTree_Int_t m2ad5_2_2_argbuf_d;
  logic m2ad5_2_2_argbuf_r;
  Pointer_QTree_Int_t m2ad5_2_1_d;
  logic m2ad5_2_1_r;
  Pointer_QTree_Int_t m2ad5_2_2_d;
  logic m2ad5_2_2_r;
  Pointer_QTree_Int_t m2ad5_3_2_argbuf_d;
  logic m2ad5_3_2_argbuf_r;
  Pointer_QTree_Int_t m2ad5_3_1_d;
  logic m2ad5_3_1_r;
  Pointer_QTree_Int_t m2ad5_3_2_d;
  logic m2ad5_3_2_r;
  Pointer_QTree_Int_t m2ad5_4_1_argbuf_d;
  logic m2ad5_4_1_argbuf_r;
  Pointer_QTree_Int_t macN_1_argbuf_d;
  logic macN_1_argbuf_r;
  Pointer_QTree_Int_t macW_1_argbuf_d;
  logic macW_1_argbuf_r;
  Go_t \main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Intgo_16_d ;
  logic \main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Intgo_16_r ;
  MyDTInt_Bool_t \main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_IntisZacL_1_d ;
  logic \main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_IntisZacL_1_r ;
  MyDTInt_Int_t \main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_IntgacM_1_d ;
  logic \main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_IntgacM_1_r ;
  Pointer_QTree_Int_t \main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_IntmacN_1_d ;
  logic \main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_IntmacN_1_r ;
  MyDTInt_Int_t gacM_1_1_argbuf_d;
  logic gacM_1_1_argbuf_r;
  Go_t go_16_1_d;
  logic go_16_1_r;
  Go_t go_16_2_d;
  logic go_16_2_r;
  MyDTInt_Bool_t isZacL_1_1_argbuf_d;
  logic isZacL_1_1_argbuf_r;
  Pointer_QTree_Int_t macN_1_1_argbuf_d;
  logic macN_1_1_argbuf_r;
  Pointer_QTree_Int_t es_0_1_1_argbuf_d;
  logic es_0_1_1_argbuf_r;
  Go_t \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Intgo_17_d ;
  logic \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Intgo_17_r ;
  MyDTInt_Bool_t \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntisZacT_1_d ;
  logic \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntisZacT_1_r ;
  MyDTInt_Int_Int_t \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntgacU_1_d ;
  logic \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntgacU_1_r ;
  Int_t \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Intv'acV_1_d ;
  logic \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Intv'acV_1_r ;
  Pointer_QTree_Int_t \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntmacW_1_d ;
  logic \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntmacW_1_r ;
  MyDTInt_Int_Int_t gacU_1_1_argbuf_d;
  logic gacU_1_1_argbuf_r;
  Go_t go_17_1_d;
  logic go_17_1_r;
  Go_t go_17_2_d;
  logic go_17_2_r;
  MyDTInt_Bool_t isZacT_1_1_argbuf_d;
  logic isZacT_1_1_argbuf_r;
  Pointer_QTree_Int_t macW_1_1_argbuf_d;
  logic macW_1_1_argbuf_r;
  Int_t \v'acV_1_1_argbuf_d ;
  logic \v'acV_1_1_argbuf_r ;
  Pointer_QTree_Int_t lizzieLet12_1_argbuf_d;
  logic lizzieLet12_1_argbuf_r;
  Pointer_QTree_Int_t q1ac0_1_argbuf_d;
  logic q1ac0_1_argbuf_r;
  Pointer_QTree_Int_t q1acP_3_1_argbuf_d;
  logic q1acP_3_1_argbuf_r;
  Pointer_QTree_Int_t q1acY_3_1_argbuf_d;
  logic q1acY_3_1_argbuf_r;
  Pointer_QTree_Int_t q1ad7_3_1_argbuf_d;
  logic q1ad7_3_1_argbuf_r;
  Pointer_QTree_Int_t q2ac1_1_1_argbuf_d;
  logic q2ac1_1_1_argbuf_r;
  Pointer_QTree_Int_t q2acQ_2_1_argbuf_d;
  logic q2acQ_2_1_argbuf_r;
  Pointer_QTree_Int_t q2acZ_2_1_argbuf_d;
  logic q2acZ_2_1_argbuf_r;
  Pointer_QTree_Int_t q2ad8_2_1_argbuf_d;
  logic q2ad8_2_1_argbuf_r;
  Pointer_QTree_Int_t q3ac2_2_1_argbuf_d;
  logic q3ac2_2_1_argbuf_r;
  Pointer_QTree_Int_t q3acR_1_1_argbuf_d;
  logic q3acR_1_1_argbuf_r;
  Pointer_QTree_Int_t q3ad0_1_1_argbuf_d;
  logic q3ad0_1_1_argbuf_r;
  Pointer_QTree_Int_t q3ad9_1_1_argbuf_d;
  logic q3ad9_1_1_argbuf_r;
  Pointer_QTree_Int_t q4ac3_3_1_argbuf_d;
  logic q4ac3_3_1_argbuf_r;
  Pointer_QTree_Int_t q4acS_1_argbuf_d;
  logic q4acS_1_argbuf_r;
  Pointer_QTree_Int_t q4ad1_1_argbuf_d;
  logic q4ad1_1_argbuf_r;
  Pointer_QTree_Int_t q4ada_1_argbuf_d;
  logic q4ada_1_argbuf_r;
  CT$wnnz_Int_t readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb_d;
  logic readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb_r;
  CT$wnnz_Int_t lizzieLet25_1_d;
  logic lizzieLet25_1_r;
  CT$wnnz_Int_t lizzieLet25_2_d;
  logic lizzieLet25_2_r;
  CT$wnnz_Int_t lizzieLet25_3_d;
  logic lizzieLet25_3_r;
  CT$wnnz_Int_t lizzieLet25_4_d;
  logic lizzieLet25_4_r;
  CTkron_kron_Int_Int_Int_t readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf_rwb_d;
  logic readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf_rwb_r;
  CTkron_kron_Int_Int_Int_t lizzieLet29_1_d;
  logic lizzieLet29_1_r;
  CTkron_kron_Int_Int_Int_t lizzieLet29_2_d;
  logic lizzieLet29_2_r;
  CTkron_kron_Int_Int_Int_t lizzieLet29_3_d;
  logic lizzieLet29_3_r;
  CTkron_kron_Int_Int_Int_t lizzieLet29_4_d;
  logic lizzieLet29_4_r;
  \CTmain_map'_Int_Int_t  \readPointer_CTmain_map'_Int_Intscfarg_0_2_1_argbuf_rwb_d ;
  logic \readPointer_CTmain_map'_Int_Intscfarg_0_2_1_argbuf_rwb_r ;
  \CTmain_map'_Int_Int_t  lizzieLet34_1_d;
  logic lizzieLet34_1_r;
  \CTmain_map'_Int_Int_t  lizzieLet34_2_d;
  logic lizzieLet34_2_r;
  \CTmain_map'_Int_Int_t  lizzieLet34_3_d;
  logic lizzieLet34_3_r;
  \CTmain_map'_Int_Int_t  lizzieLet34_4_d;
  logic lizzieLet34_4_r;
  \CTmap''_map''_Int_Int_Int_t  \readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf_rwb_d ;
  logic \readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf_rwb_r ;
  \CTmap''_map''_Int_Int_Int_t  lizzieLet39_1_d;
  logic lizzieLet39_1_r;
  \CTmap''_map''_Int_Int_Int_t  lizzieLet39_2_d;
  logic lizzieLet39_2_r;
  \CTmap''_map''_Int_Int_Int_t  lizzieLet39_3_d;
  logic lizzieLet39_3_r;
  \CTmap''_map''_Int_Int_Int_t  lizzieLet39_4_d;
  logic lizzieLet39_4_r;
  QTree_Int_t readPointer_QTree_Intm1ad4_1_argbuf_rwb_d;
  logic readPointer_QTree_Intm1ad4_1_argbuf_rwb_r;
  QTree_Int_t lizzieLet6_1_d;
  logic lizzieLet6_1_r;
  QTree_Int_t lizzieLet6_2_d;
  logic lizzieLet6_2_r;
  QTree_Int_t lizzieLet6_3_d;
  logic lizzieLet6_3_r;
  QTree_Int_t lizzieLet6_4_d;
  logic lizzieLet6_4_r;
  QTree_Int_t lizzieLet6_5_d;
  logic lizzieLet6_5_r;
  QTree_Int_t lizzieLet6_6_d;
  logic lizzieLet6_6_r;
  QTree_Int_t lizzieLet6_7_d;
  logic lizzieLet6_7_r;
  QTree_Int_t readPointer_QTree_IntmacN_1_argbuf_rwb_d;
  logic readPointer_QTree_IntmacN_1_argbuf_rwb_r;
  QTree_Int_t lizzieLet10_1_d;
  logic lizzieLet10_1_r;
  QTree_Int_t lizzieLet10_2_d;
  logic lizzieLet10_2_r;
  QTree_Int_t lizzieLet10_3_d;
  logic lizzieLet10_3_r;
  QTree_Int_t lizzieLet10_4_d;
  logic lizzieLet10_4_r;
  QTree_Int_t lizzieLet10_5_d;
  logic lizzieLet10_5_r;
  QTree_Int_t lizzieLet10_6_d;
  logic lizzieLet10_6_r;
  QTree_Int_t readPointer_QTree_IntmacW_1_argbuf_rwb_d;
  logic readPointer_QTree_IntmacW_1_argbuf_rwb_r;
  QTree_Int_t lizzieLet16_1_1_d;
  logic lizzieLet16_1_1_r;
  QTree_Int_t lizzieLet16_1_2_d;
  logic lizzieLet16_1_2_r;
  QTree_Int_t lizzieLet16_1_3_d;
  logic lizzieLet16_1_3_r;
  QTree_Int_t lizzieLet16_1_4_d;
  logic lizzieLet16_1_4_r;
  QTree_Int_t lizzieLet16_1_5_d;
  logic lizzieLet16_1_5_r;
  QTree_Int_t lizzieLet16_1_6_d;
  logic lizzieLet16_1_6_r;
  QTree_Int_t lizzieLet16_1_7_d;
  logic lizzieLet16_1_7_r;
  QTree_Int_t readPointer_QTree_Intwsvt_1_1_argbuf_rwb_d;
  logic readPointer_QTree_Intwsvt_1_1_argbuf_rwb_r;
  QTree_Int_t lizzieLet4_1_d;
  logic lizzieLet4_1_r;
  QTree_Int_t lizzieLet4_2_d;
  logic lizzieLet4_2_r;
  QTree_Int_t lizzieLet4_3_d;
  logic lizzieLet4_3_r;
  QTree_Int_t lizzieLet4_4_d;
  logic lizzieLet4_4_r;
  Pointer_CTkron_kron_Int_Int_Int_t sc_0_11_1_argbuf_d;
  logic sc_0_11_1_argbuf_r;
  \Pointer_CTmain_map'_Int_Int_t  sc_0_15_1_argbuf_d;
  logic sc_0_15_1_argbuf_r;
  \Pointer_CTmap''_map''_Int_Int_Int_t  sc_0_19_1_argbuf_d;
  logic sc_0_19_1_argbuf_r;
  Pointer_CT$wnnz_Int_t sc_0_7_1_argbuf_d;
  logic sc_0_7_1_argbuf_r;
  Pointer_CTkron_kron_Int_Int_Int_t scfarg_0_1_1_argbuf_d;
  logic scfarg_0_1_1_argbuf_r;
  \Pointer_CTmain_map'_Int_Int_t  scfarg_0_2_1_argbuf_d;
  logic scfarg_0_2_1_argbuf_r;
  \Pointer_CTmap''_map''_Int_Int_Int_t  scfarg_0_3_1_argbuf_d;
  logic scfarg_0_3_1_argbuf_r;
  Pointer_CT$wnnz_Int_t scfarg_0_1_argbuf_d;
  logic scfarg_0_1_argbuf_r;
  Int_t \v'acV_2_2_argbuf_d ;
  logic \v'acV_2_2_argbuf_r ;
  Int_t \v'acV_2_1_d ;
  logic \v'acV_2_1_r ;
  Int_t \v'acV_2_2_d ;
  logic \v'acV_2_2_r ;
  Int_t \v'acV_3_2_argbuf_d ;
  logic \v'acV_3_2_argbuf_r ;
  Int_t \v'acV_3_1_d ;
  logic \v'acV_3_1_r ;
  Int_t \v'acV_3_2_d ;
  logic \v'acV_3_2_r ;
  Int_t \v'acV_4_1_argbuf_d ;
  logic \v'acV_4_1_argbuf_r ;
  Int_t vacO_1_argbuf_d;
  logic vacO_1_argbuf_r;
  Int_t vacX_1_argbuf_d;
  logic vacX_1_argbuf_r;
  Int_t vad6_1_argbuf_d;
  logic vad6_1_argbuf_r;
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb_d;
  logic writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb_r;
  Pointer_CT$wnnz_Int_t lizzieLet17_1_argbuf_d;
  logic lizzieLet17_1_argbuf_r;
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet26_1_argbuf_rwb_d;
  logic writeCT$wnnz_IntlizzieLet26_1_argbuf_rwb_r;
  Pointer_CT$wnnz_Int_t sca2_1_argbuf_d;
  logic sca2_1_argbuf_r;
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet27_1_argbuf_rwb_d;
  logic writeCT$wnnz_IntlizzieLet27_1_argbuf_rwb_r;
  Pointer_CT$wnnz_Int_t sca1_1_argbuf_d;
  logic sca1_1_argbuf_r;
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet28_1_argbuf_rwb_d;
  logic writeCT$wnnz_IntlizzieLet28_1_argbuf_rwb_r;
  Pointer_CT$wnnz_Int_t sca0_1_argbuf_d;
  logic sca0_1_argbuf_r;
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb_d;
  logic writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb_r;
  Pointer_CT$wnnz_Int_t sca3_1_argbuf_d;
  logic sca3_1_argbuf_r;
  Pointer_CTkron_kron_Int_Int_Int_t writeCTkron_kron_Int_Int_IntlizzieLet22_1_argbuf_rwb_d;
  logic writeCTkron_kron_Int_Int_IntlizzieLet22_1_argbuf_rwb_r;
  Pointer_CTkron_kron_Int_Int_Int_t lizzieLet14_1_1_argbuf_d;
  logic lizzieLet14_1_1_argbuf_r;
  Pointer_CTkron_kron_Int_Int_Int_t writeCTkron_kron_Int_Int_IntlizzieLet30_1_argbuf_rwb_d;
  logic writeCTkron_kron_Int_Int_IntlizzieLet30_1_argbuf_rwb_r;
  Pointer_CTkron_kron_Int_Int_Int_t sca2_1_1_argbuf_d;
  logic sca2_1_1_argbuf_r;
  Pointer_CTkron_kron_Int_Int_Int_t writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf_rwb_d;
  logic writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf_rwb_r;
  Pointer_CTkron_kron_Int_Int_Int_t sca1_1_1_argbuf_d;
  logic sca1_1_1_argbuf_r;
  Pointer_CTkron_kron_Int_Int_Int_t writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf_rwb_d;
  logic writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf_rwb_r;
  Pointer_CTkron_kron_Int_Int_Int_t sca0_1_1_argbuf_d;
  logic sca0_1_1_argbuf_r;
  Pointer_CTkron_kron_Int_Int_Int_t writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf_rwb_d;
  logic writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf_rwb_r;
  Pointer_CTkron_kron_Int_Int_Int_t sca3_1_1_argbuf_d;
  logic sca3_1_1_argbuf_r;
  \Pointer_CTmain_map'_Int_Int_t  \writeCTmain_map'_Int_IntlizzieLet14_1_argbuf_rwb_d ;
  logic \writeCTmain_map'_Int_IntlizzieLet14_1_argbuf_rwb_r ;
  \Pointer_CTmain_map'_Int_Int_t  sca3_2_1_argbuf_d;
  logic sca3_2_1_argbuf_r;
  \Pointer_CTmain_map'_Int_Int_t  \writeCTmain_map'_Int_IntlizzieLet23_1_argbuf_rwb_d ;
  logic \writeCTmain_map'_Int_IntlizzieLet23_1_argbuf_rwb_r ;
  \Pointer_CTmain_map'_Int_Int_t  lizzieLet5_1_1_argbuf_d;
  logic lizzieLet5_1_1_argbuf_r;
  \Pointer_CTmain_map'_Int_Int_t  \writeCTmain_map'_Int_IntlizzieLet35_1_argbuf_rwb_d ;
  logic \writeCTmain_map'_Int_IntlizzieLet35_1_argbuf_rwb_r ;
  \Pointer_CTmain_map'_Int_Int_t  sca2_2_1_argbuf_d;
  logic sca2_2_1_argbuf_r;
  \Pointer_CTmain_map'_Int_Int_t  \writeCTmain_map'_Int_IntlizzieLet36_1_argbuf_rwb_d ;
  logic \writeCTmain_map'_Int_IntlizzieLet36_1_argbuf_rwb_r ;
  \Pointer_CTmain_map'_Int_Int_t  sca1_2_1_argbuf_d;
  logic sca1_2_1_argbuf_r;
  \Pointer_CTmain_map'_Int_Int_t  \writeCTmain_map'_Int_IntlizzieLet37_1_argbuf_rwb_d ;
  logic \writeCTmain_map'_Int_IntlizzieLet37_1_argbuf_rwb_r ;
  \Pointer_CTmain_map'_Int_Int_t  sca0_2_1_argbuf_d;
  logic sca0_2_1_argbuf_r;
  \Pointer_CTmap''_map''_Int_Int_Int_t  \writeCTmap''_map''_Int_Int_IntlizzieLet20_1_argbuf_rwb_d ;
  logic \writeCTmap''_map''_Int_Int_IntlizzieLet20_1_argbuf_rwb_r ;
  \Pointer_CTmap''_map''_Int_Int_Int_t  sca3_3_1_argbuf_d;
  logic sca3_3_1_argbuf_r;
  \Pointer_CTmap''_map''_Int_Int_Int_t  \writeCTmap''_map''_Int_Int_IntlizzieLet24_1_argbuf_rwb_d ;
  logic \writeCTmap''_map''_Int_Int_IntlizzieLet24_1_argbuf_rwb_r ;
  \Pointer_CTmap''_map''_Int_Int_Int_t  lizzieLet10_1_1_argbuf_d;
  logic lizzieLet10_1_1_argbuf_r;
  \Pointer_CTmap''_map''_Int_Int_Int_t  \writeCTmap''_map''_Int_Int_IntlizzieLet40_1_argbuf_rwb_d ;
  logic \writeCTmap''_map''_Int_Int_IntlizzieLet40_1_argbuf_rwb_r ;
  \Pointer_CTmap''_map''_Int_Int_Int_t  sca2_3_1_argbuf_d;
  logic sca2_3_1_argbuf_r;
  \Pointer_CTmap''_map''_Int_Int_Int_t  \writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf_rwb_d ;
  logic \writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf_rwb_r ;
  \Pointer_CTmap''_map''_Int_Int_Int_t  sca1_3_1_argbuf_d;
  logic sca1_3_1_argbuf_r;
  \Pointer_CTmap''_map''_Int_Int_Int_t  \writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf_rwb_d ;
  logic \writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf_rwb_r ;
  \Pointer_CTmap''_map''_Int_Int_Int_t  sca0_3_1_argbuf_d;
  logic sca0_3_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet11_1_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet11_1_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet1_1_1_argbuf_d;
  logic lizzieLet1_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet12_1_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet12_1_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet2_1_1_argbuf_d;
  logic lizzieLet2_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet13_1_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet13_1_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet3_1_1_argbuf_d;
  logic lizzieLet3_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet15_2_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet15_2_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet4_1_1_argbuf_d;
  logic lizzieLet4_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet17_1_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet17_1_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet6_1_1_argbuf_d;
  logic lizzieLet6_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet18_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet18_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet7_1_1_argbuf_d;
  logic lizzieLet7_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet19_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet19_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet8_1_1_argbuf_d;
  logic lizzieLet8_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet21_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet21_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet9_1_1_argbuf_d;
  logic lizzieLet9_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet33_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet33_1_argbuf_rwb_r;
  Pointer_QTree_Int_t contRet_0_1_1_argbuf_d;
  logic contRet_0_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet38_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet38_1_argbuf_rwb_r;
  Pointer_QTree_Int_t contRet_0_2_1_argbuf_d;
  logic contRet_0_2_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet43_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet43_1_argbuf_rwb_r;
  Pointer_QTree_Int_t contRet_0_3_1_argbuf_d;
  logic contRet_0_3_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet7_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet7_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet11_1_argbuf_d;
  logic lizzieLet11_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet9_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet9_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet13_1_argbuf_d;
  logic lizzieLet13_1_argbuf_r;
  Pointer_QTree_Int_t wsvt_1_1_argbuf_d;
  logic wsvt_1_1_argbuf_r;
  CT$wnnz_Int_t lizzieLet27_1_argbuf_d;
  logic lizzieLet27_1_argbuf_r;
  CT$wnnz_Int_t wwsvw_1_1lizzieLet25_4Lcall_$wnnz_Int2_1sc_0_5_1q4ac3_2_1Lcall_$wnnz_Int1_d;
  logic wwsvw_1_1lizzieLet25_4Lcall_$wnnz_Int2_1sc_0_5_1q4ac3_2_1Lcall_$wnnz_Int1_r;
  CT$wnnz_Int_t lizzieLet28_1_argbuf_d;
  logic lizzieLet28_1_argbuf_r;
  CT$wnnz_Int_t wwsvw_2_1ww1XwI_1_1lizzieLet25_4Lcall_$wnnz_Int1_1sc_0_6_1Lcall_$wnnz_Int0_d;
  logic wwsvw_2_1ww1XwI_1_1lizzieLet25_4Lcall_$wnnz_Int1_1sc_0_6_1Lcall_$wnnz_Int0_r;
  \Int#_t  es_6_1ww2XwL_1_1_Add32_d;
  logic es_6_1ww2XwL_1_1_Add32_r;
  \Int#_t  wwsvw_3_1ww1XwI_2_1_Add32_d;
  logic wwsvw_3_1ww1XwI_2_1_Add32_r;
  Int_t xacr_1_argbuf_d;
  logic xacr_1_argbuf_r;
  Int_t xacr_1_1_argbuf_d;
  logic xacr_1_1_argbuf_r;
  Int_t \es_0_2_1I#_d ;
  logic \es_0_2_1I#_r ;
  \Int#_t  xaqa_1lizzieLet0_1_1_Add32_d;
  logic xaqa_1lizzieLet0_1_1_Add32_r;
  
  /* fork (Ty Go) : (sourceGo,Go) > [(goFork,Go),
                                (goFor_2,Go),
                                (goFor_3,Go),
                                (goFor_4,Go),
                                (goFor_5,Go),
                                (goFor_6,Go),
                                (goFor_7,Go),
                                (goFor_8,Go),
                                (goFor_9,Go)] */
  logic [8:0] sourceGo_emitted;
  logic [8:0] sourceGo_done;
  assign goFork_d = (sourceGo_d[0] && (! sourceGo_emitted[0]));
  assign goFor_2_d = (sourceGo_d[0] && (! sourceGo_emitted[1]));
  assign goFor_3_d = (sourceGo_d[0] && (! sourceGo_emitted[2]));
  assign goFor_4_d = (sourceGo_d[0] && (! sourceGo_emitted[3]));
  assign goFor_5_d = (sourceGo_d[0] && (! sourceGo_emitted[4]));
  assign goFor_6_d = (sourceGo_d[0] && (! sourceGo_emitted[5]));
  assign goFor_7_d = (sourceGo_d[0] && (! sourceGo_emitted[6]));
  assign goFor_8_d = (sourceGo_d[0] && (! sourceGo_emitted[7]));
  assign goFor_9_d = (sourceGo_d[0] && (! sourceGo_emitted[8]));
  assign sourceGo_done = (sourceGo_emitted | ({goFor_9_d[0],
                                               goFor_8_d[0],
                                               goFor_7_d[0],
                                               goFor_6_d[0],
                                               goFor_5_d[0],
                                               goFor_4_d[0],
                                               goFor_3_d[0],
                                               goFor_2_d[0],
                                               goFork_d[0]} & {goFor_9_r,
                                                               goFor_8_r,
                                                               goFor_7_r,
                                                               goFor_6_r,
                                                               goFor_5_r,
                                                               goFor_4_r,
                                                               goFor_3_r,
                                                               goFor_2_r,
                                                               goFork_r}));
  assign sourceGo_r = (& sourceGo_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) sourceGo_emitted <= 9'd0;
    else
      sourceGo_emitted <= (sourceGo_r ? 9'd0 :
                           sourceGo_done);
  
  /* const (Ty Word16#,
       Lit 0) : (goFor_2,Go) > (initHP_CT$wnnz_Int,Word16#) */
  assign initHP_CT$wnnz_Int_d = {16'd0, goFor_2_d[0]};
  assign goFor_2_r = initHP_CT$wnnz_Int_r;
  
  /* const (Ty Word16#,
       Lit 1) : (incrHP_CT$wnnz_Int1,Go) > (incrHP_CT$wnnz_Int,Word16#) */
  assign incrHP_CT$wnnz_Int_d = {16'd1, incrHP_CT$wnnz_Int1_d[0]};
  assign incrHP_CT$wnnz_Int1_r = incrHP_CT$wnnz_Int_r;
  
  /* merge (Ty Go) : [(goFor_3,Go),
                 (incrHP_CT$wnnz_Int2,Go)] > (incrHP_mergeCT$wnnz_Int,Go) */
  logic [1:0] incrHP_mergeCT$wnnz_Int_selected;
  logic [1:0] incrHP_mergeCT$wnnz_Int_select;
  always_comb
    begin
      incrHP_mergeCT$wnnz_Int_selected = 2'd0;
      if ((| incrHP_mergeCT$wnnz_Int_select))
        incrHP_mergeCT$wnnz_Int_selected = incrHP_mergeCT$wnnz_Int_select;
      else
        if (goFor_3_d[0]) incrHP_mergeCT$wnnz_Int_selected[0] = 1'd1;
        else if (incrHP_CT$wnnz_Int2_d[0])
          incrHP_mergeCT$wnnz_Int_selected[1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeCT$wnnz_Int_select <= 2'd0;
    else
      incrHP_mergeCT$wnnz_Int_select <= (incrHP_mergeCT$wnnz_Int_r ? 2'd0 :
                                         incrHP_mergeCT$wnnz_Int_selected);
  always_comb
    if (incrHP_mergeCT$wnnz_Int_selected[0])
      incrHP_mergeCT$wnnz_Int_d = goFor_3_d;
    else if (incrHP_mergeCT$wnnz_Int_selected[1])
      incrHP_mergeCT$wnnz_Int_d = incrHP_CT$wnnz_Int2_d;
    else incrHP_mergeCT$wnnz_Int_d = 1'd0;
  assign {incrHP_CT$wnnz_Int2_r,
          goFor_3_r} = (incrHP_mergeCT$wnnz_Int_r ? incrHP_mergeCT$wnnz_Int_selected :
                        2'd0);
  
  /* fork (Ty Go) : (incrHP_mergeCT$wnnz_Int_buf,Go) > [(incrHP_CT$wnnz_Int1,Go),
                                                   (incrHP_CT$wnnz_Int2,Go)] */
  logic [1:0] incrHP_mergeCT$wnnz_Int_buf_emitted;
  logic [1:0] incrHP_mergeCT$wnnz_Int_buf_done;
  assign incrHP_CT$wnnz_Int1_d = (incrHP_mergeCT$wnnz_Int_buf_d[0] && (! incrHP_mergeCT$wnnz_Int_buf_emitted[0]));
  assign incrHP_CT$wnnz_Int2_d = (incrHP_mergeCT$wnnz_Int_buf_d[0] && (! incrHP_mergeCT$wnnz_Int_buf_emitted[1]));
  assign incrHP_mergeCT$wnnz_Int_buf_done = (incrHP_mergeCT$wnnz_Int_buf_emitted | ({incrHP_CT$wnnz_Int2_d[0],
                                                                                     incrHP_CT$wnnz_Int1_d[0]} & {incrHP_CT$wnnz_Int2_r,
                                                                                                                  incrHP_CT$wnnz_Int1_r}));
  assign incrHP_mergeCT$wnnz_Int_buf_r = (& incrHP_mergeCT$wnnz_Int_buf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeCT$wnnz_Int_buf_emitted <= 2'd0;
    else
      incrHP_mergeCT$wnnz_Int_buf_emitted <= (incrHP_mergeCT$wnnz_Int_buf_r ? 2'd0 :
                                              incrHP_mergeCT$wnnz_Int_buf_done);
  
  /* op_add (Ty Word16#) : (incrHP_CT$wnnz_Int,Word16#) (forkHP1_CT$wnnz_Int,Word16#) > (addHP_CT$wnnz_Int,Word16#) */
  assign addHP_CT$wnnz_Int_d = {(incrHP_CT$wnnz_Int_d[16:1] + forkHP1_CT$wnnz_Int_d[16:1]),
                                (incrHP_CT$wnnz_Int_d[0] && forkHP1_CT$wnnz_Int_d[0])};
  assign {incrHP_CT$wnnz_Int_r,
          forkHP1_CT$wnnz_Int_r} = {2 {(addHP_CT$wnnz_Int_r && addHP_CT$wnnz_Int_d[0])}};
  
  /* merge (Ty Word16#) : [(initHP_CT$wnnz_Int,Word16#),
                      (addHP_CT$wnnz_Int,Word16#)] > (mergeHP_CT$wnnz_Int,Word16#) */
  logic [1:0] mergeHP_CT$wnnz_Int_selected;
  logic [1:0] mergeHP_CT$wnnz_Int_select;
  always_comb
    begin
      mergeHP_CT$wnnz_Int_selected = 2'd0;
      if ((| mergeHP_CT$wnnz_Int_select))
        mergeHP_CT$wnnz_Int_selected = mergeHP_CT$wnnz_Int_select;
      else
        if (initHP_CT$wnnz_Int_d[0])
          mergeHP_CT$wnnz_Int_selected[0] = 1'd1;
        else if (addHP_CT$wnnz_Int_d[0])
          mergeHP_CT$wnnz_Int_selected[1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_CT$wnnz_Int_select <= 2'd0;
    else
      mergeHP_CT$wnnz_Int_select <= (mergeHP_CT$wnnz_Int_r ? 2'd0 :
                                     mergeHP_CT$wnnz_Int_selected);
  always_comb
    if (mergeHP_CT$wnnz_Int_selected[0])
      mergeHP_CT$wnnz_Int_d = initHP_CT$wnnz_Int_d;
    else if (mergeHP_CT$wnnz_Int_selected[1])
      mergeHP_CT$wnnz_Int_d = addHP_CT$wnnz_Int_d;
    else mergeHP_CT$wnnz_Int_d = {16'd0, 1'd0};
  assign {addHP_CT$wnnz_Int_r,
          initHP_CT$wnnz_Int_r} = (mergeHP_CT$wnnz_Int_r ? mergeHP_CT$wnnz_Int_selected :
                                   2'd0);
  
  /* buf (Ty Go) : (incrHP_mergeCT$wnnz_Int,Go) > (incrHP_mergeCT$wnnz_Int_buf,Go) */
  Go_t incrHP_mergeCT$wnnz_Int_bufchan_d;
  logic incrHP_mergeCT$wnnz_Int_bufchan_r;
  assign incrHP_mergeCT$wnnz_Int_r = ((! incrHP_mergeCT$wnnz_Int_bufchan_d[0]) || incrHP_mergeCT$wnnz_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeCT$wnnz_Int_bufchan_d <= 1'd0;
    else
      if (incrHP_mergeCT$wnnz_Int_r)
        incrHP_mergeCT$wnnz_Int_bufchan_d <= incrHP_mergeCT$wnnz_Int_d;
  Go_t incrHP_mergeCT$wnnz_Int_bufchan_buf;
  assign incrHP_mergeCT$wnnz_Int_bufchan_r = (! incrHP_mergeCT$wnnz_Int_bufchan_buf[0]);
  assign incrHP_mergeCT$wnnz_Int_buf_d = (incrHP_mergeCT$wnnz_Int_bufchan_buf[0] ? incrHP_mergeCT$wnnz_Int_bufchan_buf :
                                          incrHP_mergeCT$wnnz_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeCT$wnnz_Int_bufchan_buf <= 1'd0;
    else
      if ((incrHP_mergeCT$wnnz_Int_buf_r && incrHP_mergeCT$wnnz_Int_bufchan_buf[0]))
        incrHP_mergeCT$wnnz_Int_bufchan_buf <= 1'd0;
      else if (((! incrHP_mergeCT$wnnz_Int_buf_r) && (! incrHP_mergeCT$wnnz_Int_bufchan_buf[0])))
        incrHP_mergeCT$wnnz_Int_bufchan_buf <= incrHP_mergeCT$wnnz_Int_bufchan_d;
  
  /* buf (Ty Word16#) : (mergeHP_CT$wnnz_Int,Word16#) > (mergeHP_CT$wnnz_Int_buf,Word16#) */
  \Word16#_t  mergeHP_CT$wnnz_Int_bufchan_d;
  logic mergeHP_CT$wnnz_Int_bufchan_r;
  assign mergeHP_CT$wnnz_Int_r = ((! mergeHP_CT$wnnz_Int_bufchan_d[0]) || mergeHP_CT$wnnz_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      mergeHP_CT$wnnz_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (mergeHP_CT$wnnz_Int_r)
        mergeHP_CT$wnnz_Int_bufchan_d <= mergeHP_CT$wnnz_Int_d;
  \Word16#_t  mergeHP_CT$wnnz_Int_bufchan_buf;
  assign mergeHP_CT$wnnz_Int_bufchan_r = (! mergeHP_CT$wnnz_Int_bufchan_buf[0]);
  assign mergeHP_CT$wnnz_Int_buf_d = (mergeHP_CT$wnnz_Int_bufchan_buf[0] ? mergeHP_CT$wnnz_Int_bufchan_buf :
                                      mergeHP_CT$wnnz_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      mergeHP_CT$wnnz_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((mergeHP_CT$wnnz_Int_buf_r && mergeHP_CT$wnnz_Int_bufchan_buf[0]))
        mergeHP_CT$wnnz_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! mergeHP_CT$wnnz_Int_buf_r) && (! mergeHP_CT$wnnz_Int_bufchan_buf[0])))
        mergeHP_CT$wnnz_Int_bufchan_buf <= mergeHP_CT$wnnz_Int_bufchan_d;
  
  /* fork (Ty Word16#) : (mergeHP_CT$wnnz_Int_buf,Word16#) > [(forkHP1_CT$wnnz_Int,Word16#),
                                                         (forkHP1_CT$wnnz_In2,Word16#),
                                                         (forkHP1_CT$wnnz_In3,Word16#)] */
  logic [2:0] mergeHP_CT$wnnz_Int_buf_emitted;
  logic [2:0] mergeHP_CT$wnnz_Int_buf_done;
  assign forkHP1_CT$wnnz_Int_d = {mergeHP_CT$wnnz_Int_buf_d[16:1],
                                  (mergeHP_CT$wnnz_Int_buf_d[0] && (! mergeHP_CT$wnnz_Int_buf_emitted[0]))};
  assign forkHP1_CT$wnnz_In2_d = {mergeHP_CT$wnnz_Int_buf_d[16:1],
                                  (mergeHP_CT$wnnz_Int_buf_d[0] && (! mergeHP_CT$wnnz_Int_buf_emitted[1]))};
  assign forkHP1_CT$wnnz_In3_d = {mergeHP_CT$wnnz_Int_buf_d[16:1],
                                  (mergeHP_CT$wnnz_Int_buf_d[0] && (! mergeHP_CT$wnnz_Int_buf_emitted[2]))};
  assign mergeHP_CT$wnnz_Int_buf_done = (mergeHP_CT$wnnz_Int_buf_emitted | ({forkHP1_CT$wnnz_In3_d[0],
                                                                             forkHP1_CT$wnnz_In2_d[0],
                                                                             forkHP1_CT$wnnz_Int_d[0]} & {forkHP1_CT$wnnz_In3_r,
                                                                                                          forkHP1_CT$wnnz_In2_r,
                                                                                                          forkHP1_CT$wnnz_Int_r}));
  assign mergeHP_CT$wnnz_Int_buf_r = (& mergeHP_CT$wnnz_Int_buf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_CT$wnnz_Int_buf_emitted <= 3'd0;
    else
      mergeHP_CT$wnnz_Int_buf_emitted <= (mergeHP_CT$wnnz_Int_buf_r ? 3'd0 :
                                          mergeHP_CT$wnnz_Int_buf_done);
  
  /* mergectrl (Ty C2,
           Ty MemIn_CT$wnnz_Int) : [(dconReadIn_CT$wnnz_Int,MemIn_CT$wnnz_Int),
                                    (dconWriteIn_CT$wnnz_Int,MemIn_CT$wnnz_Int)] > (memMergeChoice_CT$wnnz_Int,C2) (memMergeIn_CT$wnnz_Int,MemIn_CT$wnnz_Int) */
  logic [1:0] dconReadIn_CT$wnnz_Int_select_d;
  assign dconReadIn_CT$wnnz_Int_select_d = ((| dconReadIn_CT$wnnz_Int_select_q) ? dconReadIn_CT$wnnz_Int_select_q :
                                            (dconReadIn_CT$wnnz_Int_d[0] ? 2'd1 :
                                             (dconWriteIn_CT$wnnz_Int_d[0] ? 2'd2 :
                                              2'd0)));
  logic [1:0] dconReadIn_CT$wnnz_Int_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) dconReadIn_CT$wnnz_Int_select_q <= 2'd0;
    else
      dconReadIn_CT$wnnz_Int_select_q <= (dconReadIn_CT$wnnz_Int_done ? 2'd0 :
                                          dconReadIn_CT$wnnz_Int_select_d);
  logic [1:0] dconReadIn_CT$wnnz_Int_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) dconReadIn_CT$wnnz_Int_emit_q <= 2'd0;
    else
      dconReadIn_CT$wnnz_Int_emit_q <= (dconReadIn_CT$wnnz_Int_done ? 2'd0 :
                                        dconReadIn_CT$wnnz_Int_emit_d);
  logic [1:0] dconReadIn_CT$wnnz_Int_emit_d;
  assign dconReadIn_CT$wnnz_Int_emit_d = (dconReadIn_CT$wnnz_Int_emit_q | ({memMergeChoice_CT$wnnz_Int_d[0],
                                                                            memMergeIn_CT$wnnz_Int_d[0]} & {memMergeChoice_CT$wnnz_Int_r,
                                                                                                            memMergeIn_CT$wnnz_Int_r}));
  logic dconReadIn_CT$wnnz_Int_done;
  assign dconReadIn_CT$wnnz_Int_done = (& dconReadIn_CT$wnnz_Int_emit_d);
  assign {dconWriteIn_CT$wnnz_Int_r,
          dconReadIn_CT$wnnz_Int_r} = (dconReadIn_CT$wnnz_Int_done ? dconReadIn_CT$wnnz_Int_select_d :
                                       2'd0);
  assign memMergeIn_CT$wnnz_Int_d = ((dconReadIn_CT$wnnz_Int_select_d[0] && (! dconReadIn_CT$wnnz_Int_emit_q[0])) ? dconReadIn_CT$wnnz_Int_d :
                                     ((dconReadIn_CT$wnnz_Int_select_d[1] && (! dconReadIn_CT$wnnz_Int_emit_q[0])) ? dconWriteIn_CT$wnnz_Int_d :
                                      {132'd0, 1'd0}));
  assign memMergeChoice_CT$wnnz_Int_d = ((dconReadIn_CT$wnnz_Int_select_d[0] && (! dconReadIn_CT$wnnz_Int_emit_q[1])) ? C1_2_dc(1'd1) :
                                         ((dconReadIn_CT$wnnz_Int_select_d[1] && (! dconReadIn_CT$wnnz_Int_emit_q[1])) ? C2_2_dc(1'd1) :
                                          {1'd0, 1'd0}));
  
  /* bram (Ty MemIn_CT$wnnz_Int,
      Ty MemOut_CT$wnnz_Int) : (memMergeIn_CT$wnnz_Int_dbuf,MemIn_CT$wnnz_Int) > (memOut_CT$wnnz_Int,MemOut_CT$wnnz_Int) */
  logic [114:0] memMergeIn_CT$wnnz_Int_dbuf_mem[65535:0];
  logic [15:0] memMergeIn_CT$wnnz_Int_dbuf_address;
  logic [114:0] memMergeIn_CT$wnnz_Int_dbuf_din;
  logic [114:0] memOut_CT$wnnz_Int_q;
  logic memOut_CT$wnnz_Int_valid;
  logic memMergeIn_CT$wnnz_Int_dbuf_we;
  logic memOut_CT$wnnz_Int_we;
  assign memMergeIn_CT$wnnz_Int_dbuf_din = memMergeIn_CT$wnnz_Int_dbuf_d[132:18];
  assign memMergeIn_CT$wnnz_Int_dbuf_address = memMergeIn_CT$wnnz_Int_dbuf_d[17:2];
  assign memMergeIn_CT$wnnz_Int_dbuf_we = (memMergeIn_CT$wnnz_Int_dbuf_d[1:1] && memMergeIn_CT$wnnz_Int_dbuf_d[0]);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        memOut_CT$wnnz_Int_we <= 1'd0;
        memOut_CT$wnnz_Int_valid <= 1'd0;
      end
    else
      begin
        memOut_CT$wnnz_Int_we <= memMergeIn_CT$wnnz_Int_dbuf_we;
        memOut_CT$wnnz_Int_valid <= memMergeIn_CT$wnnz_Int_dbuf_d[0];
        if (memMergeIn_CT$wnnz_Int_dbuf_we)
          begin
            memMergeIn_CT$wnnz_Int_dbuf_mem[memMergeIn_CT$wnnz_Int_dbuf_address] <= memMergeIn_CT$wnnz_Int_dbuf_din;
            memOut_CT$wnnz_Int_q <= memMergeIn_CT$wnnz_Int_dbuf_din;
          end
        else
          memOut_CT$wnnz_Int_q <= memMergeIn_CT$wnnz_Int_dbuf_mem[memMergeIn_CT$wnnz_Int_dbuf_address];
      end
  assign memOut_CT$wnnz_Int_d = {memOut_CT$wnnz_Int_q,
                                 memOut_CT$wnnz_Int_we,
                                 memOut_CT$wnnz_Int_valid};
  assign memMergeIn_CT$wnnz_Int_dbuf_r = ((! memOut_CT$wnnz_Int_valid) || memOut_CT$wnnz_Int_r);
  
  /* demux (Ty C2,
       Ty MemOut_CT$wnnz_Int) : (memMergeChoice_CT$wnnz_Int,C2) (memOut_CT$wnnz_Int_dbuf,MemOut_CT$wnnz_Int) > [(memReadOut_CT$wnnz_Int,MemOut_CT$wnnz_Int),
                                                                                                                (memWriteOut_CT$wnnz_Int,MemOut_CT$wnnz_Int)] */
  logic [1:0] memOut_CT$wnnz_Int_dbuf_onehotd;
  always_comb
    if ((memMergeChoice_CT$wnnz_Int_d[0] && memOut_CT$wnnz_Int_dbuf_d[0]))
      unique case (memMergeChoice_CT$wnnz_Int_d[1:1])
        1'd0: memOut_CT$wnnz_Int_dbuf_onehotd = 2'd1;
        1'd1: memOut_CT$wnnz_Int_dbuf_onehotd = 2'd2;
        default: memOut_CT$wnnz_Int_dbuf_onehotd = 2'd0;
      endcase
    else memOut_CT$wnnz_Int_dbuf_onehotd = 2'd0;
  assign memReadOut_CT$wnnz_Int_d = {memOut_CT$wnnz_Int_dbuf_d[116:1],
                                     memOut_CT$wnnz_Int_dbuf_onehotd[0]};
  assign memWriteOut_CT$wnnz_Int_d = {memOut_CT$wnnz_Int_dbuf_d[116:1],
                                      memOut_CT$wnnz_Int_dbuf_onehotd[1]};
  assign memOut_CT$wnnz_Int_dbuf_r = (| (memOut_CT$wnnz_Int_dbuf_onehotd & {memWriteOut_CT$wnnz_Int_r,
                                                                            memReadOut_CT$wnnz_Int_r}));
  assign memMergeChoice_CT$wnnz_Int_r = memOut_CT$wnnz_Int_dbuf_r;
  
  /* dbuf (Ty MemIn_CT$wnnz_Int) : (memMergeIn_CT$wnnz_Int_rbuf,MemIn_CT$wnnz_Int) > (memMergeIn_CT$wnnz_Int_dbuf,MemIn_CT$wnnz_Int) */
  assign memMergeIn_CT$wnnz_Int_rbuf_r = ((! memMergeIn_CT$wnnz_Int_dbuf_d[0]) || memMergeIn_CT$wnnz_Int_dbuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      memMergeIn_CT$wnnz_Int_dbuf_d <= {132'd0, 1'd0};
    else
      if (memMergeIn_CT$wnnz_Int_rbuf_r)
        memMergeIn_CT$wnnz_Int_dbuf_d <= memMergeIn_CT$wnnz_Int_rbuf_d;
  
  /* rbuf (Ty MemIn_CT$wnnz_Int) : (memMergeIn_CT$wnnz_Int,MemIn_CT$wnnz_Int) > (memMergeIn_CT$wnnz_Int_rbuf,MemIn_CT$wnnz_Int) */
  MemIn_CT$wnnz_Int_t memMergeIn_CT$wnnz_Int_buf;
  assign memMergeIn_CT$wnnz_Int_r = (! memMergeIn_CT$wnnz_Int_buf[0]);
  assign memMergeIn_CT$wnnz_Int_rbuf_d = (memMergeIn_CT$wnnz_Int_buf[0] ? memMergeIn_CT$wnnz_Int_buf :
                                          memMergeIn_CT$wnnz_Int_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memMergeIn_CT$wnnz_Int_buf <= {132'd0, 1'd0};
    else
      if ((memMergeIn_CT$wnnz_Int_rbuf_r && memMergeIn_CT$wnnz_Int_buf[0]))
        memMergeIn_CT$wnnz_Int_buf <= {132'd0, 1'd0};
      else if (((! memMergeIn_CT$wnnz_Int_rbuf_r) && (! memMergeIn_CT$wnnz_Int_buf[0])))
        memMergeIn_CT$wnnz_Int_buf <= memMergeIn_CT$wnnz_Int_d;
  
  /* dbuf (Ty MemOut_CT$wnnz_Int) : (memOut_CT$wnnz_Int_rbuf,MemOut_CT$wnnz_Int) > (memOut_CT$wnnz_Int_dbuf,MemOut_CT$wnnz_Int) */
  assign memOut_CT$wnnz_Int_rbuf_r = ((! memOut_CT$wnnz_Int_dbuf_d[0]) || memOut_CT$wnnz_Int_dbuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memOut_CT$wnnz_Int_dbuf_d <= {116'd0, 1'd0};
    else
      if (memOut_CT$wnnz_Int_rbuf_r)
        memOut_CT$wnnz_Int_dbuf_d <= memOut_CT$wnnz_Int_rbuf_d;
  
  /* rbuf (Ty MemOut_CT$wnnz_Int) : (memOut_CT$wnnz_Int,MemOut_CT$wnnz_Int) > (memOut_CT$wnnz_Int_rbuf,MemOut_CT$wnnz_Int) */
  MemOut_CT$wnnz_Int_t memOut_CT$wnnz_Int_buf;
  assign memOut_CT$wnnz_Int_r = (! memOut_CT$wnnz_Int_buf[0]);
  assign memOut_CT$wnnz_Int_rbuf_d = (memOut_CT$wnnz_Int_buf[0] ? memOut_CT$wnnz_Int_buf :
                                      memOut_CT$wnnz_Int_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memOut_CT$wnnz_Int_buf <= {116'd0, 1'd0};
    else
      if ((memOut_CT$wnnz_Int_rbuf_r && memOut_CT$wnnz_Int_buf[0]))
        memOut_CT$wnnz_Int_buf <= {116'd0, 1'd0};
      else if (((! memOut_CT$wnnz_Int_rbuf_r) && (! memOut_CT$wnnz_Int_buf[0])))
        memOut_CT$wnnz_Int_buf <= memOut_CT$wnnz_Int_d;
  
  /* destruct (Ty Pointer_CT$wnnz_Int,
          Dcon Pointer_CT$wnnz_Int) : (scfarg_0_1_argbuf,Pointer_CT$wnnz_Int) > [(destructReadIn_CT$wnnz_Int,Word16#)] */
  assign destructReadIn_CT$wnnz_Int_d = {scfarg_0_1_argbuf_d[16:1],
                                         scfarg_0_1_argbuf_d[0]};
  assign scfarg_0_1_argbuf_r = destructReadIn_CT$wnnz_Int_r;
  
  /* dcon (Ty MemIn_CT$wnnz_Int,
      Dcon ReadIn_CT$wnnz_Int) : [(destructReadIn_CT$wnnz_Int,Word16#)] > (dconReadIn_CT$wnnz_Int,MemIn_CT$wnnz_Int) */
  assign dconReadIn_CT$wnnz_Int_d = ReadIn_CT$wnnz_Int_dc((& {destructReadIn_CT$wnnz_Int_d[0]}), destructReadIn_CT$wnnz_Int_d);
  assign {destructReadIn_CT$wnnz_Int_r} = {1 {(dconReadIn_CT$wnnz_Int_r && dconReadIn_CT$wnnz_Int_d[0])}};
  
  /* destruct (Ty MemOut_CT$wnnz_Int,
          Dcon ReadOut_CT$wnnz_Int) : (memReadOut_CT$wnnz_Int,MemOut_CT$wnnz_Int) > [(readPointer_CT$wnnz_Intscfarg_0_1_argbuf,CT$wnnz_Int)] */
  assign readPointer_CT$wnnz_Intscfarg_0_1_argbuf_d = {memReadOut_CT$wnnz_Int_d[116:2],
                                                       memReadOut_CT$wnnz_Int_d[0]};
  assign memReadOut_CT$wnnz_Int_r = readPointer_CT$wnnz_Intscfarg_0_1_argbuf_r;
  
  /* mergectrl (Ty C5,
           Ty CT$wnnz_Int) : [(lizzieLet0_1_argbuf,CT$wnnz_Int),
                              (lizzieLet26_1_argbuf,CT$wnnz_Int),
                              (lizzieLet27_1_argbuf,CT$wnnz_Int),
                              (lizzieLet28_1_argbuf,CT$wnnz_Int),
                              (lizzieLet5_1_argbuf,CT$wnnz_Int)] > (writeMerge_choice_CT$wnnz_Int,C5) (writeMerge_data_CT$wnnz_Int,CT$wnnz_Int) */
  logic [4:0] lizzieLet0_1_argbuf_select_d;
  assign lizzieLet0_1_argbuf_select_d = ((| lizzieLet0_1_argbuf_select_q) ? lizzieLet0_1_argbuf_select_q :
                                         (lizzieLet0_1_argbuf_d[0] ? 5'd1 :
                                          (lizzieLet26_1_argbuf_d[0] ? 5'd2 :
                                           (lizzieLet27_1_argbuf_d[0] ? 5'd4 :
                                            (lizzieLet28_1_argbuf_d[0] ? 5'd8 :
                                             (lizzieLet5_1_argbuf_d[0] ? 5'd16 :
                                              5'd0))))));
  logic [4:0] lizzieLet0_1_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet0_1_argbuf_select_q <= 5'd0;
    else
      lizzieLet0_1_argbuf_select_q <= (lizzieLet0_1_argbuf_done ? 5'd0 :
                                       lizzieLet0_1_argbuf_select_d);
  logic [1:0] lizzieLet0_1_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet0_1_argbuf_emit_q <= 2'd0;
    else
      lizzieLet0_1_argbuf_emit_q <= (lizzieLet0_1_argbuf_done ? 2'd0 :
                                     lizzieLet0_1_argbuf_emit_d);
  logic [1:0] lizzieLet0_1_argbuf_emit_d;
  assign lizzieLet0_1_argbuf_emit_d = (lizzieLet0_1_argbuf_emit_q | ({writeMerge_choice_CT$wnnz_Int_d[0],
                                                                      writeMerge_data_CT$wnnz_Int_d[0]} & {writeMerge_choice_CT$wnnz_Int_r,
                                                                                                           writeMerge_data_CT$wnnz_Int_r}));
  logic lizzieLet0_1_argbuf_done;
  assign lizzieLet0_1_argbuf_done = (& lizzieLet0_1_argbuf_emit_d);
  assign {lizzieLet5_1_argbuf_r,
          lizzieLet28_1_argbuf_r,
          lizzieLet27_1_argbuf_r,
          lizzieLet26_1_argbuf_r,
          lizzieLet0_1_argbuf_r} = (lizzieLet0_1_argbuf_done ? lizzieLet0_1_argbuf_select_d :
                                    5'd0);
  assign writeMerge_data_CT$wnnz_Int_d = ((lizzieLet0_1_argbuf_select_d[0] && (! lizzieLet0_1_argbuf_emit_q[0])) ? lizzieLet0_1_argbuf_d :
                                          ((lizzieLet0_1_argbuf_select_d[1] && (! lizzieLet0_1_argbuf_emit_q[0])) ? lizzieLet26_1_argbuf_d :
                                           ((lizzieLet0_1_argbuf_select_d[2] && (! lizzieLet0_1_argbuf_emit_q[0])) ? lizzieLet27_1_argbuf_d :
                                            ((lizzieLet0_1_argbuf_select_d[3] && (! lizzieLet0_1_argbuf_emit_q[0])) ? lizzieLet28_1_argbuf_d :
                                             ((lizzieLet0_1_argbuf_select_d[4] && (! lizzieLet0_1_argbuf_emit_q[0])) ? lizzieLet5_1_argbuf_d :
                                              {115'd0, 1'd0})))));
  assign writeMerge_choice_CT$wnnz_Int_d = ((lizzieLet0_1_argbuf_select_d[0] && (! lizzieLet0_1_argbuf_emit_q[1])) ? C1_5_dc(1'd1) :
                                            ((lizzieLet0_1_argbuf_select_d[1] && (! lizzieLet0_1_argbuf_emit_q[1])) ? C2_5_dc(1'd1) :
                                             ((lizzieLet0_1_argbuf_select_d[2] && (! lizzieLet0_1_argbuf_emit_q[1])) ? C3_5_dc(1'd1) :
                                              ((lizzieLet0_1_argbuf_select_d[3] && (! lizzieLet0_1_argbuf_emit_q[1])) ? C4_5_dc(1'd1) :
                                               ((lizzieLet0_1_argbuf_select_d[4] && (! lizzieLet0_1_argbuf_emit_q[1])) ? C5_5_dc(1'd1) :
                                                {3'd0, 1'd0})))));
  
  /* demux (Ty C5,
       Ty Pointer_CT$wnnz_Int) : (writeMerge_choice_CT$wnnz_Int,C5) (demuxWriteResult_CT$wnnz_Int,Pointer_CT$wnnz_Int) > [(writeCT$wnnz_IntlizzieLet0_1_argbuf,Pointer_CT$wnnz_Int),
                                                                                                                          (writeCT$wnnz_IntlizzieLet26_1_argbuf,Pointer_CT$wnnz_Int),
                                                                                                                          (writeCT$wnnz_IntlizzieLet27_1_argbuf,Pointer_CT$wnnz_Int),
                                                                                                                          (writeCT$wnnz_IntlizzieLet28_1_argbuf,Pointer_CT$wnnz_Int),
                                                                                                                          (writeCT$wnnz_IntlizzieLet5_1_argbuf,Pointer_CT$wnnz_Int)] */
  logic [4:0] demuxWriteResult_CT$wnnz_Int_onehotd;
  always_comb
    if ((writeMerge_choice_CT$wnnz_Int_d[0] && demuxWriteResult_CT$wnnz_Int_d[0]))
      unique case (writeMerge_choice_CT$wnnz_Int_d[3:1])
        3'd0: demuxWriteResult_CT$wnnz_Int_onehotd = 5'd1;
        3'd1: demuxWriteResult_CT$wnnz_Int_onehotd = 5'd2;
        3'd2: demuxWriteResult_CT$wnnz_Int_onehotd = 5'd4;
        3'd3: demuxWriteResult_CT$wnnz_Int_onehotd = 5'd8;
        3'd4: demuxWriteResult_CT$wnnz_Int_onehotd = 5'd16;
        default: demuxWriteResult_CT$wnnz_Int_onehotd = 5'd0;
      endcase
    else demuxWriteResult_CT$wnnz_Int_onehotd = 5'd0;
  assign writeCT$wnnz_IntlizzieLet0_1_argbuf_d = {demuxWriteResult_CT$wnnz_Int_d[16:1],
                                                  demuxWriteResult_CT$wnnz_Int_onehotd[0]};
  assign writeCT$wnnz_IntlizzieLet26_1_argbuf_d = {demuxWriteResult_CT$wnnz_Int_d[16:1],
                                                   demuxWriteResult_CT$wnnz_Int_onehotd[1]};
  assign writeCT$wnnz_IntlizzieLet27_1_argbuf_d = {demuxWriteResult_CT$wnnz_Int_d[16:1],
                                                   demuxWriteResult_CT$wnnz_Int_onehotd[2]};
  assign writeCT$wnnz_IntlizzieLet28_1_argbuf_d = {demuxWriteResult_CT$wnnz_Int_d[16:1],
                                                   demuxWriteResult_CT$wnnz_Int_onehotd[3]};
  assign writeCT$wnnz_IntlizzieLet5_1_argbuf_d = {demuxWriteResult_CT$wnnz_Int_d[16:1],
                                                  demuxWriteResult_CT$wnnz_Int_onehotd[4]};
  assign demuxWriteResult_CT$wnnz_Int_r = (| (demuxWriteResult_CT$wnnz_Int_onehotd & {writeCT$wnnz_IntlizzieLet5_1_argbuf_r,
                                                                                      writeCT$wnnz_IntlizzieLet28_1_argbuf_r,
                                                                                      writeCT$wnnz_IntlizzieLet27_1_argbuf_r,
                                                                                      writeCT$wnnz_IntlizzieLet26_1_argbuf_r,
                                                                                      writeCT$wnnz_IntlizzieLet0_1_argbuf_r}));
  assign writeMerge_choice_CT$wnnz_Int_r = demuxWriteResult_CT$wnnz_Int_r;
  
  /* dcon (Ty MemIn_CT$wnnz_Int,
      Dcon WriteIn_CT$wnnz_Int) : [(forkHP1_CT$wnnz_In2,Word16#),
                                   (writeMerge_data_CT$wnnz_Int,CT$wnnz_Int)] > (dconWriteIn_CT$wnnz_Int,MemIn_CT$wnnz_Int) */
  assign dconWriteIn_CT$wnnz_Int_d = WriteIn_CT$wnnz_Int_dc((& {forkHP1_CT$wnnz_In2_d[0],
                                                                writeMerge_data_CT$wnnz_Int_d[0]}), forkHP1_CT$wnnz_In2_d, writeMerge_data_CT$wnnz_Int_d);
  assign {forkHP1_CT$wnnz_In2_r,
          writeMerge_data_CT$wnnz_Int_r} = {2 {(dconWriteIn_CT$wnnz_Int_r && dconWriteIn_CT$wnnz_Int_d[0])}};
  
  /* dcon (Ty Pointer_CT$wnnz_Int,
      Dcon Pointer_CT$wnnz_Int) : [(forkHP1_CT$wnnz_In3,Word16#)] > (dconPtr_CT$wnnz_Int,Pointer_CT$wnnz_Int) */
  assign dconPtr_CT$wnnz_Int_d = Pointer_CT$wnnz_Int_dc((& {forkHP1_CT$wnnz_In3_d[0]}), forkHP1_CT$wnnz_In3_d);
  assign {forkHP1_CT$wnnz_In3_r} = {1 {(dconPtr_CT$wnnz_Int_r && dconPtr_CT$wnnz_Int_d[0])}};
  
  /* demux (Ty MemOut_CT$wnnz_Int,
       Ty Pointer_CT$wnnz_Int) : (memWriteOut_CT$wnnz_Int,MemOut_CT$wnnz_Int) (dconPtr_CT$wnnz_Int,Pointer_CT$wnnz_Int) > [(_39,Pointer_CT$wnnz_Int),
                                                                                                                           (demuxWriteResult_CT$wnnz_Int,Pointer_CT$wnnz_Int)] */
  logic [1:0] dconPtr_CT$wnnz_Int_onehotd;
  always_comb
    if ((memWriteOut_CT$wnnz_Int_d[0] && dconPtr_CT$wnnz_Int_d[0]))
      unique case (memWriteOut_CT$wnnz_Int_d[1:1])
        1'd0: dconPtr_CT$wnnz_Int_onehotd = 2'd1;
        1'd1: dconPtr_CT$wnnz_Int_onehotd = 2'd2;
        default: dconPtr_CT$wnnz_Int_onehotd = 2'd0;
      endcase
    else dconPtr_CT$wnnz_Int_onehotd = 2'd0;
  assign _39_d = {dconPtr_CT$wnnz_Int_d[16:1],
                  dconPtr_CT$wnnz_Int_onehotd[0]};
  assign demuxWriteResult_CT$wnnz_Int_d = {dconPtr_CT$wnnz_Int_d[16:1],
                                           dconPtr_CT$wnnz_Int_onehotd[1]};
  assign dconPtr_CT$wnnz_Int_r = (| (dconPtr_CT$wnnz_Int_onehotd & {demuxWriteResult_CT$wnnz_Int_r,
                                                                    _39_r}));
  assign memWriteOut_CT$wnnz_Int_r = dconPtr_CT$wnnz_Int_r;
  
  /* const (Ty Word16#,
       Lit 0) : (go_1_dummy_write_QTree_Int,Go) > (initHP_QTree_Int,Word16#) */
  assign initHP_QTree_Int_d = {16'd0,
                               go_1_dummy_write_QTree_Int_d[0]};
  assign go_1_dummy_write_QTree_Int_r = initHP_QTree_Int_r;
  
  /* const (Ty Word16#,
       Lit 1) : (incrHP_QTree_Int1,Go) > (incrHP_QTree_Int,Word16#) */
  assign incrHP_QTree_Int_d = {16'd1, incrHP_QTree_Int1_d[0]};
  assign incrHP_QTree_Int1_r = incrHP_QTree_Int_r;
  
  /* merge (Ty Go) : [(go_2_dummy_write_QTree_Int,Go),
                 (incrHP_QTree_Int2,Go)] > (incrHP_mergeQTree_Int,Go) */
  logic [1:0] incrHP_mergeQTree_Int_selected;
  logic [1:0] incrHP_mergeQTree_Int_select;
  always_comb
    begin
      incrHP_mergeQTree_Int_selected = 2'd0;
      if ((| incrHP_mergeQTree_Int_select))
        incrHP_mergeQTree_Int_selected = incrHP_mergeQTree_Int_select;
      else
        if (go_2_dummy_write_QTree_Int_d[0])
          incrHP_mergeQTree_Int_selected[0] = 1'd1;
        else if (incrHP_QTree_Int2_d[0])
          incrHP_mergeQTree_Int_selected[1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeQTree_Int_select <= 2'd0;
    else
      incrHP_mergeQTree_Int_select <= (incrHP_mergeQTree_Int_r ? 2'd0 :
                                       incrHP_mergeQTree_Int_selected);
  always_comb
    if (incrHP_mergeQTree_Int_selected[0])
      incrHP_mergeQTree_Int_d = go_2_dummy_write_QTree_Int_d;
    else if (incrHP_mergeQTree_Int_selected[1])
      incrHP_mergeQTree_Int_d = incrHP_QTree_Int2_d;
    else incrHP_mergeQTree_Int_d = 1'd0;
  assign {incrHP_QTree_Int2_r,
          go_2_dummy_write_QTree_Int_r} = (incrHP_mergeQTree_Int_r ? incrHP_mergeQTree_Int_selected :
                                           2'd0);
  
  /* fork (Ty Go) : (incrHP_mergeQTree_Int_buf,Go) > [(incrHP_QTree_Int1,Go),
                                                 (incrHP_QTree_Int2,Go)] */
  logic [1:0] incrHP_mergeQTree_Int_buf_emitted;
  logic [1:0] incrHP_mergeQTree_Int_buf_done;
  assign incrHP_QTree_Int1_d = (incrHP_mergeQTree_Int_buf_d[0] && (! incrHP_mergeQTree_Int_buf_emitted[0]));
  assign incrHP_QTree_Int2_d = (incrHP_mergeQTree_Int_buf_d[0] && (! incrHP_mergeQTree_Int_buf_emitted[1]));
  assign incrHP_mergeQTree_Int_buf_done = (incrHP_mergeQTree_Int_buf_emitted | ({incrHP_QTree_Int2_d[0],
                                                                                 incrHP_QTree_Int1_d[0]} & {incrHP_QTree_Int2_r,
                                                                                                            incrHP_QTree_Int1_r}));
  assign incrHP_mergeQTree_Int_buf_r = (& incrHP_mergeQTree_Int_buf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeQTree_Int_buf_emitted <= 2'd0;
    else
      incrHP_mergeQTree_Int_buf_emitted <= (incrHP_mergeQTree_Int_buf_r ? 2'd0 :
                                            incrHP_mergeQTree_Int_buf_done);
  
  /* op_add (Ty Word16#) : (incrHP_QTree_Int,Word16#) (forkHP1_QTree_Int,Word16#) > (addHP_QTree_Int,Word16#) */
  assign addHP_QTree_Int_d = {(incrHP_QTree_Int_d[16:1] + forkHP1_QTree_Int_d[16:1]),
                              (incrHP_QTree_Int_d[0] && forkHP1_QTree_Int_d[0])};
  assign {incrHP_QTree_Int_r,
          forkHP1_QTree_Int_r} = {2 {(addHP_QTree_Int_r && addHP_QTree_Int_d[0])}};
  
  /* merge (Ty Word16#) : [(initHP_QTree_Int,Word16#),
                      (addHP_QTree_Int,Word16#)] > (mergeHP_QTree_Int,Word16#) */
  logic [1:0] mergeHP_QTree_Int_selected;
  logic [1:0] mergeHP_QTree_Int_select;
  always_comb
    begin
      mergeHP_QTree_Int_selected = 2'd0;
      if ((| mergeHP_QTree_Int_select))
        mergeHP_QTree_Int_selected = mergeHP_QTree_Int_select;
      else
        if (initHP_QTree_Int_d[0]) mergeHP_QTree_Int_selected[0] = 1'd1;
        else if (addHP_QTree_Int_d[0])
          mergeHP_QTree_Int_selected[1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_QTree_Int_select <= 2'd0;
    else
      mergeHP_QTree_Int_select <= (mergeHP_QTree_Int_r ? 2'd0 :
                                   mergeHP_QTree_Int_selected);
  always_comb
    if (mergeHP_QTree_Int_selected[0])
      mergeHP_QTree_Int_d = initHP_QTree_Int_d;
    else if (mergeHP_QTree_Int_selected[1])
      mergeHP_QTree_Int_d = addHP_QTree_Int_d;
    else mergeHP_QTree_Int_d = {16'd0, 1'd0};
  assign {addHP_QTree_Int_r,
          initHP_QTree_Int_r} = (mergeHP_QTree_Int_r ? mergeHP_QTree_Int_selected :
                                 2'd0);
  
  /* buf (Ty Go) : (incrHP_mergeQTree_Int,Go) > (incrHP_mergeQTree_Int_buf,Go) */
  Go_t incrHP_mergeQTree_Int_bufchan_d;
  logic incrHP_mergeQTree_Int_bufchan_r;
  assign incrHP_mergeQTree_Int_r = ((! incrHP_mergeQTree_Int_bufchan_d[0]) || incrHP_mergeQTree_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeQTree_Int_bufchan_d <= 1'd0;
    else
      if (incrHP_mergeQTree_Int_r)
        incrHP_mergeQTree_Int_bufchan_d <= incrHP_mergeQTree_Int_d;
  Go_t incrHP_mergeQTree_Int_bufchan_buf;
  assign incrHP_mergeQTree_Int_bufchan_r = (! incrHP_mergeQTree_Int_bufchan_buf[0]);
  assign incrHP_mergeQTree_Int_buf_d = (incrHP_mergeQTree_Int_bufchan_buf[0] ? incrHP_mergeQTree_Int_bufchan_buf :
                                        incrHP_mergeQTree_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeQTree_Int_bufchan_buf <= 1'd0;
    else
      if ((incrHP_mergeQTree_Int_buf_r && incrHP_mergeQTree_Int_bufchan_buf[0]))
        incrHP_mergeQTree_Int_bufchan_buf <= 1'd0;
      else if (((! incrHP_mergeQTree_Int_buf_r) && (! incrHP_mergeQTree_Int_bufchan_buf[0])))
        incrHP_mergeQTree_Int_bufchan_buf <= incrHP_mergeQTree_Int_bufchan_d;
  
  /* buf (Ty Word16#) : (mergeHP_QTree_Int,Word16#) > (mergeHP_QTree_Int_buf,Word16#) */
  \Word16#_t  mergeHP_QTree_Int_bufchan_d;
  logic mergeHP_QTree_Int_bufchan_r;
  assign mergeHP_QTree_Int_r = ((! mergeHP_QTree_Int_bufchan_d[0]) || mergeHP_QTree_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_QTree_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (mergeHP_QTree_Int_r)
        mergeHP_QTree_Int_bufchan_d <= mergeHP_QTree_Int_d;
  \Word16#_t  mergeHP_QTree_Int_bufchan_buf;
  assign mergeHP_QTree_Int_bufchan_r = (! mergeHP_QTree_Int_bufchan_buf[0]);
  assign mergeHP_QTree_Int_buf_d = (mergeHP_QTree_Int_bufchan_buf[0] ? mergeHP_QTree_Int_bufchan_buf :
                                    mergeHP_QTree_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      mergeHP_QTree_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((mergeHP_QTree_Int_buf_r && mergeHP_QTree_Int_bufchan_buf[0]))
        mergeHP_QTree_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! mergeHP_QTree_Int_buf_r) && (! mergeHP_QTree_Int_bufchan_buf[0])))
        mergeHP_QTree_Int_bufchan_buf <= mergeHP_QTree_Int_bufchan_d;
  
  /* sink (Ty Word16#) : (forkHP1_QTree_Int_snk,Word16#) > */
  assign {forkHP1_QTree_Int_snk_r,
          forkHP1_QTree_Int_snk_dout} = {forkHP1_QTree_Int_snk_rout,
                                         forkHP1_QTree_Int_snk_d};
  
  /* source (Ty Go) : > (\QTree_Int_src,Go) */
  
  /* fork (Ty Go) : (\QTree_Int_src,Go) > [(go_1_dummy_write_QTree_Int,Go),
                                      (go_2_dummy_write_QTree_Int,Go)] */
  logic [1:0] \\QTree_Int_src_emitted ;
  logic [1:0] \\QTree_Int_src_done ;
  assign go_1_dummy_write_QTree_Int_d = (\\QTree_Int_src_d [0] && (! \\QTree_Int_src_emitted [0]));
  assign go_2_dummy_write_QTree_Int_d = (\\QTree_Int_src_d [0] && (! \\QTree_Int_src_emitted [1]));
  assign \\QTree_Int_src_done  = (\\QTree_Int_src_emitted  | ({go_2_dummy_write_QTree_Int_d[0],
                                                               go_1_dummy_write_QTree_Int_d[0]} & {go_2_dummy_write_QTree_Int_r,
                                                                                                   go_1_dummy_write_QTree_Int_r}));
  assign \\QTree_Int_src_r  = (& \\QTree_Int_src_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \\QTree_Int_src_emitted  <= 2'd0;
    else
      \\QTree_Int_src_emitted  <= (\\QTree_Int_src_r  ? 2'd0 :
                                   \\QTree_Int_src_done );
  
  /* source (Ty QTree_Int) : > (dummy_write_QTree_Int,QTree_Int) */
  
  /* sink (Ty Pointer_QTree_Int) : (dummy_write_QTree_Int_sink,Pointer_QTree_Int) > */
  assign {dummy_write_QTree_Int_sink_r,
          dummy_write_QTree_Int_sink_dout} = {dummy_write_QTree_Int_sink_rout,
                                              dummy_write_QTree_Int_sink_d};
  
  /* fork (Ty Word16#) : (mergeHP_QTree_Int_buf,Word16#) > [(forkHP1_QTree_Int,Word16#),
                                                       (forkHP1_QTree_Int_snk,Word16#),
                                                       (forkHP1_QTree_In3,Word16#),
                                                       (forkHP1_QTree_In4,Word16#)] */
  logic [3:0] mergeHP_QTree_Int_buf_emitted;
  logic [3:0] mergeHP_QTree_Int_buf_done;
  assign forkHP1_QTree_Int_d = {mergeHP_QTree_Int_buf_d[16:1],
                                (mergeHP_QTree_Int_buf_d[0] && (! mergeHP_QTree_Int_buf_emitted[0]))};
  assign forkHP1_QTree_Int_snk_d = {mergeHP_QTree_Int_buf_d[16:1],
                                    (mergeHP_QTree_Int_buf_d[0] && (! mergeHP_QTree_Int_buf_emitted[1]))};
  assign forkHP1_QTree_In3_d = {mergeHP_QTree_Int_buf_d[16:1],
                                (mergeHP_QTree_Int_buf_d[0] && (! mergeHP_QTree_Int_buf_emitted[2]))};
  assign forkHP1_QTree_In4_d = {mergeHP_QTree_Int_buf_d[16:1],
                                (mergeHP_QTree_Int_buf_d[0] && (! mergeHP_QTree_Int_buf_emitted[3]))};
  assign mergeHP_QTree_Int_buf_done = (mergeHP_QTree_Int_buf_emitted | ({forkHP1_QTree_In4_d[0],
                                                                         forkHP1_QTree_In3_d[0],
                                                                         forkHP1_QTree_Int_snk_d[0],
                                                                         forkHP1_QTree_Int_d[0]} & {forkHP1_QTree_In4_r,
                                                                                                    forkHP1_QTree_In3_r,
                                                                                                    forkHP1_QTree_Int_snk_r,
                                                                                                    forkHP1_QTree_Int_r}));
  assign mergeHP_QTree_Int_buf_r = (& mergeHP_QTree_Int_buf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_QTree_Int_buf_emitted <= 4'd0;
    else
      mergeHP_QTree_Int_buf_emitted <= (mergeHP_QTree_Int_buf_r ? 4'd0 :
                                        mergeHP_QTree_Int_buf_done);
  
  /* mergectrl (Ty C2,
           Ty MemIn_QTree_Int) : [(dconReadIn_QTree_Int,MemIn_QTree_Int),
                                  (dconWriteIn_QTree_Int,MemIn_QTree_Int)] > (memMergeChoice_QTree_Int,C2) (memMergeIn_QTree_Int,MemIn_QTree_Int) */
  logic [1:0] dconReadIn_QTree_Int_select_d;
  assign dconReadIn_QTree_Int_select_d = ((| dconReadIn_QTree_Int_select_q) ? dconReadIn_QTree_Int_select_q :
                                          (dconReadIn_QTree_Int_d[0] ? 2'd1 :
                                           (dconWriteIn_QTree_Int_d[0] ? 2'd2 :
                                            2'd0)));
  logic [1:0] dconReadIn_QTree_Int_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) dconReadIn_QTree_Int_select_q <= 2'd0;
    else
      dconReadIn_QTree_Int_select_q <= (dconReadIn_QTree_Int_done ? 2'd0 :
                                        dconReadIn_QTree_Int_select_d);
  logic [1:0] dconReadIn_QTree_Int_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) dconReadIn_QTree_Int_emit_q <= 2'd0;
    else
      dconReadIn_QTree_Int_emit_q <= (dconReadIn_QTree_Int_done ? 2'd0 :
                                      dconReadIn_QTree_Int_emit_d);
  logic [1:0] dconReadIn_QTree_Int_emit_d;
  assign dconReadIn_QTree_Int_emit_d = (dconReadIn_QTree_Int_emit_q | ({memMergeChoice_QTree_Int_d[0],
                                                                        memMergeIn_QTree_Int_d[0]} & {memMergeChoice_QTree_Int_r,
                                                                                                      memMergeIn_QTree_Int_r}));
  logic dconReadIn_QTree_Int_done;
  assign dconReadIn_QTree_Int_done = (& dconReadIn_QTree_Int_emit_d);
  assign {dconWriteIn_QTree_Int_r,
          dconReadIn_QTree_Int_r} = (dconReadIn_QTree_Int_done ? dconReadIn_QTree_Int_select_d :
                                     2'd0);
  assign memMergeIn_QTree_Int_d = ((dconReadIn_QTree_Int_select_d[0] && (! dconReadIn_QTree_Int_emit_q[0])) ? dconReadIn_QTree_Int_d :
                                   ((dconReadIn_QTree_Int_select_d[1] && (! dconReadIn_QTree_Int_emit_q[0])) ? dconWriteIn_QTree_Int_d :
                                    {83'd0, 1'd0}));
  assign memMergeChoice_QTree_Int_d = ((dconReadIn_QTree_Int_select_d[0] && (! dconReadIn_QTree_Int_emit_q[1])) ? C1_2_dc(1'd1) :
                                       ((dconReadIn_QTree_Int_select_d[1] && (! dconReadIn_QTree_Int_emit_q[1])) ? C2_2_dc(1'd1) :
                                        {1'd0, 1'd0}));
  
  /* bram (Ty MemIn_QTree_Int,
      Ty MemOut_QTree_Int) : (memMergeIn_QTree_Int_dbuf,MemIn_QTree_Int) > (memOut_QTree_Int,MemOut_QTree_Int) */
  logic [65:0] memMergeIn_QTree_Int_dbuf_mem[65535:0];
  logic [15:0] memMergeIn_QTree_Int_dbuf_address;
  logic [65:0] memMergeIn_QTree_Int_dbuf_din;
  logic [65:0] memOut_QTree_Int_q;
  logic memOut_QTree_Int_valid;
  logic memMergeIn_QTree_Int_dbuf_we;
  logic memOut_QTree_Int_we;
  assign memMergeIn_QTree_Int_dbuf_din = memMergeIn_QTree_Int_dbuf_d[83:18];
  assign memMergeIn_QTree_Int_dbuf_address = memMergeIn_QTree_Int_dbuf_d[17:2];
  assign memMergeIn_QTree_Int_dbuf_we = (memMergeIn_QTree_Int_dbuf_d[1:1] && memMergeIn_QTree_Int_dbuf_d[0]);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        memOut_QTree_Int_we <= 1'd0;
        memOut_QTree_Int_valid <= 1'd0;
      end
    else
      begin
        memOut_QTree_Int_we <= memMergeIn_QTree_Int_dbuf_we;
        memOut_QTree_Int_valid <= memMergeIn_QTree_Int_dbuf_d[0];
        if (memMergeIn_QTree_Int_dbuf_we)
          begin
            memMergeIn_QTree_Int_dbuf_mem[memMergeIn_QTree_Int_dbuf_address] <= memMergeIn_QTree_Int_dbuf_din;
            memOut_QTree_Int_q <= memMergeIn_QTree_Int_dbuf_din;
          end
        else
          memOut_QTree_Int_q <= memMergeIn_QTree_Int_dbuf_mem[memMergeIn_QTree_Int_dbuf_address];
      end
  assign memOut_QTree_Int_d = {memOut_QTree_Int_q,
                               memOut_QTree_Int_we,
                               memOut_QTree_Int_valid};
  assign memMergeIn_QTree_Int_dbuf_r = ((! memOut_QTree_Int_valid) || memOut_QTree_Int_r);
  
  /* demux (Ty C2,
       Ty MemOut_QTree_Int) : (memMergeChoice_QTree_Int,C2) (memOut_QTree_Int_dbuf,MemOut_QTree_Int) > [(memReadOut_QTree_Int,MemOut_QTree_Int),
                                                                                                        (memWriteOut_QTree_Int,MemOut_QTree_Int)] */
  logic [1:0] memOut_QTree_Int_dbuf_onehotd;
  always_comb
    if ((memMergeChoice_QTree_Int_d[0] && memOut_QTree_Int_dbuf_d[0]))
      unique case (memMergeChoice_QTree_Int_d[1:1])
        1'd0: memOut_QTree_Int_dbuf_onehotd = 2'd1;
        1'd1: memOut_QTree_Int_dbuf_onehotd = 2'd2;
        default: memOut_QTree_Int_dbuf_onehotd = 2'd0;
      endcase
    else memOut_QTree_Int_dbuf_onehotd = 2'd0;
  assign memReadOut_QTree_Int_d = {memOut_QTree_Int_dbuf_d[67:1],
                                   memOut_QTree_Int_dbuf_onehotd[0]};
  assign memWriteOut_QTree_Int_d = {memOut_QTree_Int_dbuf_d[67:1],
                                    memOut_QTree_Int_dbuf_onehotd[1]};
  assign memOut_QTree_Int_dbuf_r = (| (memOut_QTree_Int_dbuf_onehotd & {memWriteOut_QTree_Int_r,
                                                                        memReadOut_QTree_Int_r}));
  assign memMergeChoice_QTree_Int_r = memOut_QTree_Int_dbuf_r;
  
  /* dbuf (Ty MemIn_QTree_Int) : (memMergeIn_QTree_Int_rbuf,MemIn_QTree_Int) > (memMergeIn_QTree_Int_dbuf,MemIn_QTree_Int) */
  assign memMergeIn_QTree_Int_rbuf_r = ((! memMergeIn_QTree_Int_dbuf_d[0]) || memMergeIn_QTree_Int_dbuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memMergeIn_QTree_Int_dbuf_d <= {83'd0, 1'd0};
    else
      if (memMergeIn_QTree_Int_rbuf_r)
        memMergeIn_QTree_Int_dbuf_d <= memMergeIn_QTree_Int_rbuf_d;
  
  /* rbuf (Ty MemIn_QTree_Int) : (memMergeIn_QTree_Int,MemIn_QTree_Int) > (memMergeIn_QTree_Int_rbuf,MemIn_QTree_Int) */
  MemIn_QTree_Int_t memMergeIn_QTree_Int_buf;
  assign memMergeIn_QTree_Int_r = (! memMergeIn_QTree_Int_buf[0]);
  assign memMergeIn_QTree_Int_rbuf_d = (memMergeIn_QTree_Int_buf[0] ? memMergeIn_QTree_Int_buf :
                                        memMergeIn_QTree_Int_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memMergeIn_QTree_Int_buf <= {83'd0, 1'd0};
    else
      if ((memMergeIn_QTree_Int_rbuf_r && memMergeIn_QTree_Int_buf[0]))
        memMergeIn_QTree_Int_buf <= {83'd0, 1'd0};
      else if (((! memMergeIn_QTree_Int_rbuf_r) && (! memMergeIn_QTree_Int_buf[0])))
        memMergeIn_QTree_Int_buf <= memMergeIn_QTree_Int_d;
  
  /* dbuf (Ty MemOut_QTree_Int) : (memOut_QTree_Int_rbuf,MemOut_QTree_Int) > (memOut_QTree_Int_dbuf,MemOut_QTree_Int) */
  assign memOut_QTree_Int_rbuf_r = ((! memOut_QTree_Int_dbuf_d[0]) || memOut_QTree_Int_dbuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memOut_QTree_Int_dbuf_d <= {67'd0, 1'd0};
    else
      if (memOut_QTree_Int_rbuf_r)
        memOut_QTree_Int_dbuf_d <= memOut_QTree_Int_rbuf_d;
  
  /* rbuf (Ty MemOut_QTree_Int) : (memOut_QTree_Int,MemOut_QTree_Int) > (memOut_QTree_Int_rbuf,MemOut_QTree_Int) */
  MemOut_QTree_Int_t memOut_QTree_Int_buf;
  assign memOut_QTree_Int_r = (! memOut_QTree_Int_buf[0]);
  assign memOut_QTree_Int_rbuf_d = (memOut_QTree_Int_buf[0] ? memOut_QTree_Int_buf :
                                    memOut_QTree_Int_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memOut_QTree_Int_buf <= {67'd0, 1'd0};
    else
      if ((memOut_QTree_Int_rbuf_r && memOut_QTree_Int_buf[0]))
        memOut_QTree_Int_buf <= {67'd0, 1'd0};
      else if (((! memOut_QTree_Int_rbuf_r) && (! memOut_QTree_Int_buf[0])))
        memOut_QTree_Int_buf <= memOut_QTree_Int_d;
  
  /* mergectrl (Ty C4,
           Ty Pointer_QTree_Int) : [(m1ad4_1_argbuf,Pointer_QTree_Int),
                                    (macN_1_argbuf,Pointer_QTree_Int),
                                    (macW_1_argbuf,Pointer_QTree_Int),
                                    (wsvt_1_1_argbuf,Pointer_QTree_Int)] > (readMerge_choice_QTree_Int,C4) (readMerge_data_QTree_Int,Pointer_QTree_Int) */
  logic [3:0] m1ad4_1_argbuf_select_d;
  assign m1ad4_1_argbuf_select_d = ((| m1ad4_1_argbuf_select_q) ? m1ad4_1_argbuf_select_q :
                                    (m1ad4_1_argbuf_d[0] ? 4'd1 :
                                     (macN_1_argbuf_d[0] ? 4'd2 :
                                      (macW_1_argbuf_d[0] ? 4'd4 :
                                       (wsvt_1_1_argbuf_d[0] ? 4'd8 :
                                        4'd0)))));
  logic [3:0] m1ad4_1_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m1ad4_1_argbuf_select_q <= 4'd0;
    else
      m1ad4_1_argbuf_select_q <= (m1ad4_1_argbuf_done ? 4'd0 :
                                  m1ad4_1_argbuf_select_d);
  logic [1:0] m1ad4_1_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m1ad4_1_argbuf_emit_q <= 2'd0;
    else
      m1ad4_1_argbuf_emit_q <= (m1ad4_1_argbuf_done ? 2'd0 :
                                m1ad4_1_argbuf_emit_d);
  logic [1:0] m1ad4_1_argbuf_emit_d;
  assign m1ad4_1_argbuf_emit_d = (m1ad4_1_argbuf_emit_q | ({readMerge_choice_QTree_Int_d[0],
                                                            readMerge_data_QTree_Int_d[0]} & {readMerge_choice_QTree_Int_r,
                                                                                              readMerge_data_QTree_Int_r}));
  logic m1ad4_1_argbuf_done;
  assign m1ad4_1_argbuf_done = (& m1ad4_1_argbuf_emit_d);
  assign {wsvt_1_1_argbuf_r,
          macW_1_argbuf_r,
          macN_1_argbuf_r,
          m1ad4_1_argbuf_r} = (m1ad4_1_argbuf_done ? m1ad4_1_argbuf_select_d :
                               4'd0);
  assign readMerge_data_QTree_Int_d = ((m1ad4_1_argbuf_select_d[0] && (! m1ad4_1_argbuf_emit_q[0])) ? m1ad4_1_argbuf_d :
                                       ((m1ad4_1_argbuf_select_d[1] && (! m1ad4_1_argbuf_emit_q[0])) ? macN_1_argbuf_d :
                                        ((m1ad4_1_argbuf_select_d[2] && (! m1ad4_1_argbuf_emit_q[0])) ? macW_1_argbuf_d :
                                         ((m1ad4_1_argbuf_select_d[3] && (! m1ad4_1_argbuf_emit_q[0])) ? wsvt_1_1_argbuf_d :
                                          {16'd0, 1'd0}))));
  assign readMerge_choice_QTree_Int_d = ((m1ad4_1_argbuf_select_d[0] && (! m1ad4_1_argbuf_emit_q[1])) ? C1_4_dc(1'd1) :
                                         ((m1ad4_1_argbuf_select_d[1] && (! m1ad4_1_argbuf_emit_q[1])) ? C2_4_dc(1'd1) :
                                          ((m1ad4_1_argbuf_select_d[2] && (! m1ad4_1_argbuf_emit_q[1])) ? C3_4_dc(1'd1) :
                                           ((m1ad4_1_argbuf_select_d[3] && (! m1ad4_1_argbuf_emit_q[1])) ? C4_4_dc(1'd1) :
                                            {2'd0, 1'd0}))));
  
  /* demux (Ty C4,
       Ty QTree_Int) : (readMerge_choice_QTree_Int,C4) (destructReadOut_QTree_Int,QTree_Int) > [(readPointer_QTree_Intm1ad4_1_argbuf,QTree_Int),
                                                                                                (readPointer_QTree_IntmacN_1_argbuf,QTree_Int),
                                                                                                (readPointer_QTree_IntmacW_1_argbuf,QTree_Int),
                                                                                                (readPointer_QTree_Intwsvt_1_1_argbuf,QTree_Int)] */
  logic [3:0] destructReadOut_QTree_Int_onehotd;
  always_comb
    if ((readMerge_choice_QTree_Int_d[0] && destructReadOut_QTree_Int_d[0]))
      unique case (readMerge_choice_QTree_Int_d[2:1])
        2'd0: destructReadOut_QTree_Int_onehotd = 4'd1;
        2'd1: destructReadOut_QTree_Int_onehotd = 4'd2;
        2'd2: destructReadOut_QTree_Int_onehotd = 4'd4;
        2'd3: destructReadOut_QTree_Int_onehotd = 4'd8;
        default: destructReadOut_QTree_Int_onehotd = 4'd0;
      endcase
    else destructReadOut_QTree_Int_onehotd = 4'd0;
  assign readPointer_QTree_Intm1ad4_1_argbuf_d = {destructReadOut_QTree_Int_d[66:1],
                                                  destructReadOut_QTree_Int_onehotd[0]};
  assign readPointer_QTree_IntmacN_1_argbuf_d = {destructReadOut_QTree_Int_d[66:1],
                                                 destructReadOut_QTree_Int_onehotd[1]};
  assign readPointer_QTree_IntmacW_1_argbuf_d = {destructReadOut_QTree_Int_d[66:1],
                                                 destructReadOut_QTree_Int_onehotd[2]};
  assign readPointer_QTree_Intwsvt_1_1_argbuf_d = {destructReadOut_QTree_Int_d[66:1],
                                                   destructReadOut_QTree_Int_onehotd[3]};
  assign destructReadOut_QTree_Int_r = (| (destructReadOut_QTree_Int_onehotd & {readPointer_QTree_Intwsvt_1_1_argbuf_r,
                                                                                readPointer_QTree_IntmacW_1_argbuf_r,
                                                                                readPointer_QTree_IntmacN_1_argbuf_r,
                                                                                readPointer_QTree_Intm1ad4_1_argbuf_r}));
  assign readMerge_choice_QTree_Int_r = destructReadOut_QTree_Int_r;
  
  /* destruct (Ty Pointer_QTree_Int,
          Dcon Pointer_QTree_Int) : (readMerge_data_QTree_Int,Pointer_QTree_Int) > [(destructReadIn_QTree_Int,Word16#)] */
  assign destructReadIn_QTree_Int_d = {readMerge_data_QTree_Int_d[16:1],
                                       readMerge_data_QTree_Int_d[0]};
  assign readMerge_data_QTree_Int_r = destructReadIn_QTree_Int_r;
  
  /* dcon (Ty MemIn_QTree_Int,
      Dcon ReadIn_QTree_Int) : [(destructReadIn_QTree_Int,Word16#)] > (dconReadIn_QTree_Int,MemIn_QTree_Int) */
  assign dconReadIn_QTree_Int_d = ReadIn_QTree_Int_dc((& {destructReadIn_QTree_Int_d[0]}), destructReadIn_QTree_Int_d);
  assign {destructReadIn_QTree_Int_r} = {1 {(dconReadIn_QTree_Int_r && dconReadIn_QTree_Int_d[0])}};
  
  /* destruct (Ty MemOut_QTree_Int,
          Dcon ReadOut_QTree_Int) : (memReadOut_QTree_Int,MemOut_QTree_Int) > [(destructReadOut_QTree_Int,QTree_Int)] */
  assign destructReadOut_QTree_Int_d = {memReadOut_QTree_Int_d[67:2],
                                        memReadOut_QTree_Int_d[0]};
  assign memReadOut_QTree_Int_r = destructReadOut_QTree_Int_r;
  
  /* mergectrl (Ty C14,
           Ty QTree_Int) : [(lizzieLet11_1_1_argbuf,QTree_Int),
                            (lizzieLet12_1_1_argbuf,QTree_Int),
                            (lizzieLet13_1_1_argbuf,QTree_Int),
                            (lizzieLet15_2_1_argbuf,QTree_Int),
                            (lizzieLet17_1_1_argbuf,QTree_Int),
                            (lizzieLet18_1_argbuf,QTree_Int),
                            (lizzieLet19_1_argbuf,QTree_Int),
                            (lizzieLet21_1_argbuf,QTree_Int),
                            (lizzieLet33_1_argbuf,QTree_Int),
                            (lizzieLet38_1_argbuf,QTree_Int),
                            (lizzieLet43_1_argbuf,QTree_Int),
                            (lizzieLet7_1_argbuf,QTree_Int),
                            (lizzieLet9_1_argbuf,QTree_Int),
                            (dummy_write_QTree_Int,QTree_Int)] > (writeMerge_choice_QTree_Int,C14) (writeMerge_data_QTree_Int,QTree_Int) */
  logic [13:0] lizzieLet11_1_1_argbuf_select_d;
  assign lizzieLet11_1_1_argbuf_select_d = ((| lizzieLet11_1_1_argbuf_select_q) ? lizzieLet11_1_1_argbuf_select_q :
                                            (lizzieLet11_1_1_argbuf_d[0] ? 14'd1 :
                                             (lizzieLet12_1_1_argbuf_d[0] ? 14'd2 :
                                              (lizzieLet13_1_1_argbuf_d[0] ? 14'd4 :
                                               (lizzieLet15_2_1_argbuf_d[0] ? 14'd8 :
                                                (lizzieLet17_1_1_argbuf_d[0] ? 14'd16 :
                                                 (lizzieLet18_1_argbuf_d[0] ? 14'd32 :
                                                  (lizzieLet19_1_argbuf_d[0] ? 14'd64 :
                                                   (lizzieLet21_1_argbuf_d[0] ? 14'd128 :
                                                    (lizzieLet33_1_argbuf_d[0] ? 14'd256 :
                                                     (lizzieLet38_1_argbuf_d[0] ? 14'd512 :
                                                      (lizzieLet43_1_argbuf_d[0] ? 14'd1024 :
                                                       (lizzieLet7_1_argbuf_d[0] ? 14'd2048 :
                                                        (lizzieLet9_1_argbuf_d[0] ? 14'd4096 :
                                                         (dummy_write_QTree_Int_d[0] ? 14'd8192 :
                                                          14'd0)))))))))))))));
  logic [13:0] lizzieLet11_1_1_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet11_1_1_argbuf_select_q <= 14'd0;
    else
      lizzieLet11_1_1_argbuf_select_q <= (lizzieLet11_1_1_argbuf_done ? 14'd0 :
                                          lizzieLet11_1_1_argbuf_select_d);
  logic [1:0] lizzieLet11_1_1_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet11_1_1_argbuf_emit_q <= 2'd0;
    else
      lizzieLet11_1_1_argbuf_emit_q <= (lizzieLet11_1_1_argbuf_done ? 2'd0 :
                                        lizzieLet11_1_1_argbuf_emit_d);
  logic [1:0] lizzieLet11_1_1_argbuf_emit_d;
  assign lizzieLet11_1_1_argbuf_emit_d = (lizzieLet11_1_1_argbuf_emit_q | ({writeMerge_choice_QTree_Int_d[0],
                                                                            writeMerge_data_QTree_Int_d[0]} & {writeMerge_choice_QTree_Int_r,
                                                                                                               writeMerge_data_QTree_Int_r}));
  logic lizzieLet11_1_1_argbuf_done;
  assign lizzieLet11_1_1_argbuf_done = (& lizzieLet11_1_1_argbuf_emit_d);
  assign {dummy_write_QTree_Int_r,
          lizzieLet9_1_argbuf_r,
          lizzieLet7_1_argbuf_r,
          lizzieLet43_1_argbuf_r,
          lizzieLet38_1_argbuf_r,
          lizzieLet33_1_argbuf_r,
          lizzieLet21_1_argbuf_r,
          lizzieLet19_1_argbuf_r,
          lizzieLet18_1_argbuf_r,
          lizzieLet17_1_1_argbuf_r,
          lizzieLet15_2_1_argbuf_r,
          lizzieLet13_1_1_argbuf_r,
          lizzieLet12_1_1_argbuf_r,
          lizzieLet11_1_1_argbuf_r} = (lizzieLet11_1_1_argbuf_done ? lizzieLet11_1_1_argbuf_select_d :
                                       14'd0);
  assign writeMerge_data_QTree_Int_d = ((lizzieLet11_1_1_argbuf_select_d[0] && (! lizzieLet11_1_1_argbuf_emit_q[0])) ? lizzieLet11_1_1_argbuf_d :
                                        ((lizzieLet11_1_1_argbuf_select_d[1] && (! lizzieLet11_1_1_argbuf_emit_q[0])) ? lizzieLet12_1_1_argbuf_d :
                                         ((lizzieLet11_1_1_argbuf_select_d[2] && (! lizzieLet11_1_1_argbuf_emit_q[0])) ? lizzieLet13_1_1_argbuf_d :
                                          ((lizzieLet11_1_1_argbuf_select_d[3] && (! lizzieLet11_1_1_argbuf_emit_q[0])) ? lizzieLet15_2_1_argbuf_d :
                                           ((lizzieLet11_1_1_argbuf_select_d[4] && (! lizzieLet11_1_1_argbuf_emit_q[0])) ? lizzieLet17_1_1_argbuf_d :
                                            ((lizzieLet11_1_1_argbuf_select_d[5] && (! lizzieLet11_1_1_argbuf_emit_q[0])) ? lizzieLet18_1_argbuf_d :
                                             ((lizzieLet11_1_1_argbuf_select_d[6] && (! lizzieLet11_1_1_argbuf_emit_q[0])) ? lizzieLet19_1_argbuf_d :
                                              ((lizzieLet11_1_1_argbuf_select_d[7] && (! lizzieLet11_1_1_argbuf_emit_q[0])) ? lizzieLet21_1_argbuf_d :
                                               ((lizzieLet11_1_1_argbuf_select_d[8] && (! lizzieLet11_1_1_argbuf_emit_q[0])) ? lizzieLet33_1_argbuf_d :
                                                ((lizzieLet11_1_1_argbuf_select_d[9] && (! lizzieLet11_1_1_argbuf_emit_q[0])) ? lizzieLet38_1_argbuf_d :
                                                 ((lizzieLet11_1_1_argbuf_select_d[10] && (! lizzieLet11_1_1_argbuf_emit_q[0])) ? lizzieLet43_1_argbuf_d :
                                                  ((lizzieLet11_1_1_argbuf_select_d[11] && (! lizzieLet11_1_1_argbuf_emit_q[0])) ? lizzieLet7_1_argbuf_d :
                                                   ((lizzieLet11_1_1_argbuf_select_d[12] && (! lizzieLet11_1_1_argbuf_emit_q[0])) ? lizzieLet9_1_argbuf_d :
                                                    ((lizzieLet11_1_1_argbuf_select_d[13] && (! lizzieLet11_1_1_argbuf_emit_q[0])) ? dummy_write_QTree_Int_d :
                                                     {66'd0, 1'd0}))))))))))))));
  assign writeMerge_choice_QTree_Int_d = ((lizzieLet11_1_1_argbuf_select_d[0] && (! lizzieLet11_1_1_argbuf_emit_q[1])) ? C1_14_dc(1'd1) :
                                          ((lizzieLet11_1_1_argbuf_select_d[1] && (! lizzieLet11_1_1_argbuf_emit_q[1])) ? C2_14_dc(1'd1) :
                                           ((lizzieLet11_1_1_argbuf_select_d[2] && (! lizzieLet11_1_1_argbuf_emit_q[1])) ? C3_14_dc(1'd1) :
                                            ((lizzieLet11_1_1_argbuf_select_d[3] && (! lizzieLet11_1_1_argbuf_emit_q[1])) ? C4_14_dc(1'd1) :
                                             ((lizzieLet11_1_1_argbuf_select_d[4] && (! lizzieLet11_1_1_argbuf_emit_q[1])) ? C5_14_dc(1'd1) :
                                              ((lizzieLet11_1_1_argbuf_select_d[5] && (! lizzieLet11_1_1_argbuf_emit_q[1])) ? C6_14_dc(1'd1) :
                                               ((lizzieLet11_1_1_argbuf_select_d[6] && (! lizzieLet11_1_1_argbuf_emit_q[1])) ? C7_14_dc(1'd1) :
                                                ((lizzieLet11_1_1_argbuf_select_d[7] && (! lizzieLet11_1_1_argbuf_emit_q[1])) ? C8_14_dc(1'd1) :
                                                 ((lizzieLet11_1_1_argbuf_select_d[8] && (! lizzieLet11_1_1_argbuf_emit_q[1])) ? C9_14_dc(1'd1) :
                                                  ((lizzieLet11_1_1_argbuf_select_d[9] && (! lizzieLet11_1_1_argbuf_emit_q[1])) ? C10_14_dc(1'd1) :
                                                   ((lizzieLet11_1_1_argbuf_select_d[10] && (! lizzieLet11_1_1_argbuf_emit_q[1])) ? C11_14_dc(1'd1) :
                                                    ((lizzieLet11_1_1_argbuf_select_d[11] && (! lizzieLet11_1_1_argbuf_emit_q[1])) ? C12_14_dc(1'd1) :
                                                     ((lizzieLet11_1_1_argbuf_select_d[12] && (! lizzieLet11_1_1_argbuf_emit_q[1])) ? C13_14_dc(1'd1) :
                                                      ((lizzieLet11_1_1_argbuf_select_d[13] && (! lizzieLet11_1_1_argbuf_emit_q[1])) ? C14_14_dc(1'd1) :
                                                       {4'd0, 1'd0}))))))))))))));
  
  /* demux (Ty C14,
       Ty Pointer_QTree_Int) : (writeMerge_choice_QTree_Int,C14) (demuxWriteResult_QTree_Int,Pointer_QTree_Int) > [(writeQTree_IntlizzieLet11_1_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet12_1_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet13_1_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet15_2_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet17_1_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet18_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet19_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet21_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet33_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet38_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet43_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet7_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet9_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (dummy_write_QTree_Int_sink,Pointer_QTree_Int)] */
  logic [13:0] demuxWriteResult_QTree_Int_onehotd;
  always_comb
    if ((writeMerge_choice_QTree_Int_d[0] && demuxWriteResult_QTree_Int_d[0]))
      unique case (writeMerge_choice_QTree_Int_d[4:1])
        4'd0: demuxWriteResult_QTree_Int_onehotd = 14'd1;
        4'd1: demuxWriteResult_QTree_Int_onehotd = 14'd2;
        4'd2: demuxWriteResult_QTree_Int_onehotd = 14'd4;
        4'd3: demuxWriteResult_QTree_Int_onehotd = 14'd8;
        4'd4: demuxWriteResult_QTree_Int_onehotd = 14'd16;
        4'd5: demuxWriteResult_QTree_Int_onehotd = 14'd32;
        4'd6: demuxWriteResult_QTree_Int_onehotd = 14'd64;
        4'd7: demuxWriteResult_QTree_Int_onehotd = 14'd128;
        4'd8: demuxWriteResult_QTree_Int_onehotd = 14'd256;
        4'd9: demuxWriteResult_QTree_Int_onehotd = 14'd512;
        4'd10: demuxWriteResult_QTree_Int_onehotd = 14'd1024;
        4'd11: demuxWriteResult_QTree_Int_onehotd = 14'd2048;
        4'd12: demuxWriteResult_QTree_Int_onehotd = 14'd4096;
        4'd13: demuxWriteResult_QTree_Int_onehotd = 14'd8192;
        default: demuxWriteResult_QTree_Int_onehotd = 14'd0;
      endcase
    else demuxWriteResult_QTree_Int_onehotd = 14'd0;
  assign writeQTree_IntlizzieLet11_1_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                   demuxWriteResult_QTree_Int_onehotd[0]};
  assign writeQTree_IntlizzieLet12_1_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                   demuxWriteResult_QTree_Int_onehotd[1]};
  assign writeQTree_IntlizzieLet13_1_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                   demuxWriteResult_QTree_Int_onehotd[2]};
  assign writeQTree_IntlizzieLet15_2_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                   demuxWriteResult_QTree_Int_onehotd[3]};
  assign writeQTree_IntlizzieLet17_1_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                   demuxWriteResult_QTree_Int_onehotd[4]};
  assign writeQTree_IntlizzieLet18_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                 demuxWriteResult_QTree_Int_onehotd[5]};
  assign writeQTree_IntlizzieLet19_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                 demuxWriteResult_QTree_Int_onehotd[6]};
  assign writeQTree_IntlizzieLet21_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                 demuxWriteResult_QTree_Int_onehotd[7]};
  assign writeQTree_IntlizzieLet33_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                 demuxWriteResult_QTree_Int_onehotd[8]};
  assign writeQTree_IntlizzieLet38_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                 demuxWriteResult_QTree_Int_onehotd[9]};
  assign writeQTree_IntlizzieLet43_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                 demuxWriteResult_QTree_Int_onehotd[10]};
  assign writeQTree_IntlizzieLet7_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                demuxWriteResult_QTree_Int_onehotd[11]};
  assign writeQTree_IntlizzieLet9_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                demuxWriteResult_QTree_Int_onehotd[12]};
  assign dummy_write_QTree_Int_sink_d = {demuxWriteResult_QTree_Int_d[16:1],
                                         demuxWriteResult_QTree_Int_onehotd[13]};
  assign demuxWriteResult_QTree_Int_r = (| (demuxWriteResult_QTree_Int_onehotd & {dummy_write_QTree_Int_sink_r,
                                                                                  writeQTree_IntlizzieLet9_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet7_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet43_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet38_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet33_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet21_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet19_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet18_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet17_1_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet15_2_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet13_1_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet12_1_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet11_1_1_argbuf_r}));
  assign writeMerge_choice_QTree_Int_r = demuxWriteResult_QTree_Int_r;
  
  /* dcon (Ty MemIn_QTree_Int,
      Dcon WriteIn_QTree_Int) : [(forkHP1_QTree_In3,Word16#),
                                 (writeMerge_data_QTree_Int,QTree_Int)] > (dconWriteIn_QTree_Int,MemIn_QTree_Int) */
  assign dconWriteIn_QTree_Int_d = WriteIn_QTree_Int_dc((& {forkHP1_QTree_In3_d[0],
                                                            writeMerge_data_QTree_Int_d[0]}), forkHP1_QTree_In3_d, writeMerge_data_QTree_Int_d);
  assign {forkHP1_QTree_In3_r,
          writeMerge_data_QTree_Int_r} = {2 {(dconWriteIn_QTree_Int_r && dconWriteIn_QTree_Int_d[0])}};
  
  /* dcon (Ty Pointer_QTree_Int,
      Dcon Pointer_QTree_Int) : [(forkHP1_QTree_In4,Word16#)] > (dconPtr_QTree_Int,Pointer_QTree_Int) */
  assign dconPtr_QTree_Int_d = Pointer_QTree_Int_dc((& {forkHP1_QTree_In4_d[0]}), forkHP1_QTree_In4_d);
  assign {forkHP1_QTree_In4_r} = {1 {(dconPtr_QTree_Int_r && dconPtr_QTree_Int_d[0])}};
  
  /* demux (Ty MemOut_QTree_Int,
       Ty Pointer_QTree_Int) : (memWriteOut_QTree_Int,MemOut_QTree_Int) (dconPtr_QTree_Int,Pointer_QTree_Int) > [(_38,Pointer_QTree_Int),
                                                                                                                 (demuxWriteResult_QTree_Int,Pointer_QTree_Int)] */
  logic [1:0] dconPtr_QTree_Int_onehotd;
  always_comb
    if ((memWriteOut_QTree_Int_d[0] && dconPtr_QTree_Int_d[0]))
      unique case (memWriteOut_QTree_Int_d[1:1])
        1'd0: dconPtr_QTree_Int_onehotd = 2'd1;
        1'd1: dconPtr_QTree_Int_onehotd = 2'd2;
        default: dconPtr_QTree_Int_onehotd = 2'd0;
      endcase
    else dconPtr_QTree_Int_onehotd = 2'd0;
  assign _38_d = {dconPtr_QTree_Int_d[16:1],
                  dconPtr_QTree_Int_onehotd[0]};
  assign demuxWriteResult_QTree_Int_d = {dconPtr_QTree_Int_d[16:1],
                                         dconPtr_QTree_Int_onehotd[1]};
  assign dconPtr_QTree_Int_r = (| (dconPtr_QTree_Int_onehotd & {demuxWriteResult_QTree_Int_r,
                                                                _38_r}));
  assign memWriteOut_QTree_Int_r = dconPtr_QTree_Int_r;
  
  /* const (Ty Word16#,
       Lit 0) : (goFor_4,Go) > (initHP_CTmain_map'_Int_Int,Word16#) */
  assign \initHP_CTmain_map'_Int_Int_d  = {16'd0, goFor_4_d[0]};
  assign goFor_4_r = \initHP_CTmain_map'_Int_Int_r ;
  
  /* const (Ty Word16#,
       Lit 1) : (incrHP_CTmain_map'_Int_Int1,Go) > (incrHP_CTmain_map'_Int_Int,Word16#) */
  assign \incrHP_CTmain_map'_Int_Int_d  = {16'd1,
                                           \incrHP_CTmain_map'_Int_Int1_d [0]};
  assign \incrHP_CTmain_map'_Int_Int1_r  = \incrHP_CTmain_map'_Int_Int_r ;
  
  /* merge (Ty Go) : [(goFor_5,Go),
                 (incrHP_CTmain_map'_Int_Int2,Go)] > (incrHP_mergeCTmain_map'_Int_Int,Go) */
  logic [1:0] \incrHP_mergeCTmain_map'_Int_Int_selected ;
  logic [1:0] \incrHP_mergeCTmain_map'_Int_Int_select ;
  always_comb
    begin
      \incrHP_mergeCTmain_map'_Int_Int_selected  = 2'd0;
      if ((| \incrHP_mergeCTmain_map'_Int_Int_select ))
        \incrHP_mergeCTmain_map'_Int_Int_selected  = \incrHP_mergeCTmain_map'_Int_Int_select ;
      else
        if (goFor_5_d[0])
          \incrHP_mergeCTmain_map'_Int_Int_selected [0] = 1'd1;
        else if (\incrHP_CTmain_map'_Int_Int2_d [0])
          \incrHP_mergeCTmain_map'_Int_Int_selected [1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \incrHP_mergeCTmain_map'_Int_Int_select  <= 2'd0;
    else
      \incrHP_mergeCTmain_map'_Int_Int_select  <= (\incrHP_mergeCTmain_map'_Int_Int_r  ? 2'd0 :
                                                   \incrHP_mergeCTmain_map'_Int_Int_selected );
  always_comb
    if (\incrHP_mergeCTmain_map'_Int_Int_selected [0])
      \incrHP_mergeCTmain_map'_Int_Int_d  = goFor_5_d;
    else if (\incrHP_mergeCTmain_map'_Int_Int_selected [1])
      \incrHP_mergeCTmain_map'_Int_Int_d  = \incrHP_CTmain_map'_Int_Int2_d ;
    else \incrHP_mergeCTmain_map'_Int_Int_d  = 1'd0;
  assign {\incrHP_CTmain_map'_Int_Int2_r ,
          goFor_5_r} = (\incrHP_mergeCTmain_map'_Int_Int_r  ? \incrHP_mergeCTmain_map'_Int_Int_selected  :
                        2'd0);
  
  /* fork (Ty Go) : (incrHP_mergeCTmain_map'_Int_Int_buf,Go) > [(incrHP_CTmain_map'_Int_Int1,Go),
                                                           (incrHP_CTmain_map'_Int_Int2,Go)] */
  logic [1:0] \incrHP_mergeCTmain_map'_Int_Int_buf_emitted ;
  logic [1:0] \incrHP_mergeCTmain_map'_Int_Int_buf_done ;
  assign \incrHP_CTmain_map'_Int_Int1_d  = (\incrHP_mergeCTmain_map'_Int_Int_buf_d [0] && (! \incrHP_mergeCTmain_map'_Int_Int_buf_emitted [0]));
  assign \incrHP_CTmain_map'_Int_Int2_d  = (\incrHP_mergeCTmain_map'_Int_Int_buf_d [0] && (! \incrHP_mergeCTmain_map'_Int_Int_buf_emitted [1]));
  assign \incrHP_mergeCTmain_map'_Int_Int_buf_done  = (\incrHP_mergeCTmain_map'_Int_Int_buf_emitted  | ({\incrHP_CTmain_map'_Int_Int2_d [0],
                                                                                                         \incrHP_CTmain_map'_Int_Int1_d [0]} & {\incrHP_CTmain_map'_Int_Int2_r ,
                                                                                                                                                \incrHP_CTmain_map'_Int_Int1_r }));
  assign \incrHP_mergeCTmain_map'_Int_Int_buf_r  = (& \incrHP_mergeCTmain_map'_Int_Int_buf_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \incrHP_mergeCTmain_map'_Int_Int_buf_emitted  <= 2'd0;
    else
      \incrHP_mergeCTmain_map'_Int_Int_buf_emitted  <= (\incrHP_mergeCTmain_map'_Int_Int_buf_r  ? 2'd0 :
                                                        \incrHP_mergeCTmain_map'_Int_Int_buf_done );
  
  /* op_add (Ty Word16#) : (incrHP_CTmain_map'_Int_Int,Word16#) (forkHP1_CTmain_map'_Int_Int,Word16#) > (addHP_CTmain_map'_Int_Int,Word16#) */
  assign \addHP_CTmain_map'_Int_Int_d  = {(\incrHP_CTmain_map'_Int_Int_d [16:1] + \forkHP1_CTmain_map'_Int_Int_d [16:1]),
                                          (\incrHP_CTmain_map'_Int_Int_d [0] && \forkHP1_CTmain_map'_Int_Int_d [0])};
  assign {\incrHP_CTmain_map'_Int_Int_r ,
          \forkHP1_CTmain_map'_Int_Int_r } = {2 {(\addHP_CTmain_map'_Int_Int_r  && \addHP_CTmain_map'_Int_Int_d [0])}};
  
  /* merge (Ty Word16#) : [(initHP_CTmain_map'_Int_Int,Word16#),
                      (addHP_CTmain_map'_Int_Int,Word16#)] > (mergeHP_CTmain_map'_Int_Int,Word16#) */
  logic [1:0] \mergeHP_CTmain_map'_Int_Int_selected ;
  logic [1:0] \mergeHP_CTmain_map'_Int_Int_select ;
  always_comb
    begin
      \mergeHP_CTmain_map'_Int_Int_selected  = 2'd0;
      if ((| \mergeHP_CTmain_map'_Int_Int_select ))
        \mergeHP_CTmain_map'_Int_Int_selected  = \mergeHP_CTmain_map'_Int_Int_select ;
      else
        if (\initHP_CTmain_map'_Int_Int_d [0])
          \mergeHP_CTmain_map'_Int_Int_selected [0] = 1'd1;
        else if (\addHP_CTmain_map'_Int_Int_d [0])
          \mergeHP_CTmain_map'_Int_Int_selected [1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \mergeHP_CTmain_map'_Int_Int_select  <= 2'd0;
    else
      \mergeHP_CTmain_map'_Int_Int_select  <= (\mergeHP_CTmain_map'_Int_Int_r  ? 2'd0 :
                                               \mergeHP_CTmain_map'_Int_Int_selected );
  always_comb
    if (\mergeHP_CTmain_map'_Int_Int_selected [0])
      \mergeHP_CTmain_map'_Int_Int_d  = \initHP_CTmain_map'_Int_Int_d ;
    else if (\mergeHP_CTmain_map'_Int_Int_selected [1])
      \mergeHP_CTmain_map'_Int_Int_d  = \addHP_CTmain_map'_Int_Int_d ;
    else \mergeHP_CTmain_map'_Int_Int_d  = {16'd0, 1'd0};
  assign {\addHP_CTmain_map'_Int_Int_r ,
          \initHP_CTmain_map'_Int_Int_r } = (\mergeHP_CTmain_map'_Int_Int_r  ? \mergeHP_CTmain_map'_Int_Int_selected  :
                                             2'd0);
  
  /* buf (Ty Go) : (incrHP_mergeCTmain_map'_Int_Int,Go) > (incrHP_mergeCTmain_map'_Int_Int_buf,Go) */
  Go_t \incrHP_mergeCTmain_map'_Int_Int_bufchan_d ;
  logic \incrHP_mergeCTmain_map'_Int_Int_bufchan_r ;
  assign \incrHP_mergeCTmain_map'_Int_Int_r  = ((! \incrHP_mergeCTmain_map'_Int_Int_bufchan_d [0]) || \incrHP_mergeCTmain_map'_Int_Int_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \incrHP_mergeCTmain_map'_Int_Int_bufchan_d  <= 1'd0;
    else
      if (\incrHP_mergeCTmain_map'_Int_Int_r )
        \incrHP_mergeCTmain_map'_Int_Int_bufchan_d  <= \incrHP_mergeCTmain_map'_Int_Int_d ;
  Go_t \incrHP_mergeCTmain_map'_Int_Int_bufchan_buf ;
  assign \incrHP_mergeCTmain_map'_Int_Int_bufchan_r  = (! \incrHP_mergeCTmain_map'_Int_Int_bufchan_buf [0]);
  assign \incrHP_mergeCTmain_map'_Int_Int_buf_d  = (\incrHP_mergeCTmain_map'_Int_Int_bufchan_buf [0] ? \incrHP_mergeCTmain_map'_Int_Int_bufchan_buf  :
                                                    \incrHP_mergeCTmain_map'_Int_Int_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \incrHP_mergeCTmain_map'_Int_Int_bufchan_buf  <= 1'd0;
    else
      if ((\incrHP_mergeCTmain_map'_Int_Int_buf_r  && \incrHP_mergeCTmain_map'_Int_Int_bufchan_buf [0]))
        \incrHP_mergeCTmain_map'_Int_Int_bufchan_buf  <= 1'd0;
      else if (((! \incrHP_mergeCTmain_map'_Int_Int_buf_r ) && (! \incrHP_mergeCTmain_map'_Int_Int_bufchan_buf [0])))
        \incrHP_mergeCTmain_map'_Int_Int_bufchan_buf  <= \incrHP_mergeCTmain_map'_Int_Int_bufchan_d ;
  
  /* buf (Ty Word16#) : (mergeHP_CTmain_map'_Int_Int,Word16#) > (mergeHP_CTmain_map'_Int_Int_buf,Word16#) */
  \Word16#_t  \mergeHP_CTmain_map'_Int_Int_bufchan_d ;
  logic \mergeHP_CTmain_map'_Int_Int_bufchan_r ;
  assign \mergeHP_CTmain_map'_Int_Int_r  = ((! \mergeHP_CTmain_map'_Int_Int_bufchan_d [0]) || \mergeHP_CTmain_map'_Int_Int_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \mergeHP_CTmain_map'_Int_Int_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\mergeHP_CTmain_map'_Int_Int_r )
        \mergeHP_CTmain_map'_Int_Int_bufchan_d  <= \mergeHP_CTmain_map'_Int_Int_d ;
  \Word16#_t  \mergeHP_CTmain_map'_Int_Int_bufchan_buf ;
  assign \mergeHP_CTmain_map'_Int_Int_bufchan_r  = (! \mergeHP_CTmain_map'_Int_Int_bufchan_buf [0]);
  assign \mergeHP_CTmain_map'_Int_Int_buf_d  = (\mergeHP_CTmain_map'_Int_Int_bufchan_buf [0] ? \mergeHP_CTmain_map'_Int_Int_bufchan_buf  :
                                                \mergeHP_CTmain_map'_Int_Int_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \mergeHP_CTmain_map'_Int_Int_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((\mergeHP_CTmain_map'_Int_Int_buf_r  && \mergeHP_CTmain_map'_Int_Int_bufchan_buf [0]))
        \mergeHP_CTmain_map'_Int_Int_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! \mergeHP_CTmain_map'_Int_Int_buf_r ) && (! \mergeHP_CTmain_map'_Int_Int_bufchan_buf [0])))
        \mergeHP_CTmain_map'_Int_Int_bufchan_buf  <= \mergeHP_CTmain_map'_Int_Int_bufchan_d ;
  
  /* fork (Ty Word16#) : (mergeHP_CTmain_map'_Int_Int_buf,Word16#) > [(forkHP1_CTmain_map'_Int_Int,Word16#),
                                                                 (forkHP1_CTmain_map'_Int_In2,Word16#),
                                                                 (forkHP1_CTmain_map'_Int_In3,Word16#)] */
  logic [2:0] \mergeHP_CTmain_map'_Int_Int_buf_emitted ;
  logic [2:0] \mergeHP_CTmain_map'_Int_Int_buf_done ;
  assign \forkHP1_CTmain_map'_Int_Int_d  = {\mergeHP_CTmain_map'_Int_Int_buf_d [16:1],
                                            (\mergeHP_CTmain_map'_Int_Int_buf_d [0] && (! \mergeHP_CTmain_map'_Int_Int_buf_emitted [0]))};
  assign \forkHP1_CTmain_map'_Int_In2_d  = {\mergeHP_CTmain_map'_Int_Int_buf_d [16:1],
                                            (\mergeHP_CTmain_map'_Int_Int_buf_d [0] && (! \mergeHP_CTmain_map'_Int_Int_buf_emitted [1]))};
  assign \forkHP1_CTmain_map'_Int_In3_d  = {\mergeHP_CTmain_map'_Int_Int_buf_d [16:1],
                                            (\mergeHP_CTmain_map'_Int_Int_buf_d [0] && (! \mergeHP_CTmain_map'_Int_Int_buf_emitted [2]))};
  assign \mergeHP_CTmain_map'_Int_Int_buf_done  = (\mergeHP_CTmain_map'_Int_Int_buf_emitted  | ({\forkHP1_CTmain_map'_Int_In3_d [0],
                                                                                                 \forkHP1_CTmain_map'_Int_In2_d [0],
                                                                                                 \forkHP1_CTmain_map'_Int_Int_d [0]} & {\forkHP1_CTmain_map'_Int_In3_r ,
                                                                                                                                        \forkHP1_CTmain_map'_Int_In2_r ,
                                                                                                                                        \forkHP1_CTmain_map'_Int_Int_r }));
  assign \mergeHP_CTmain_map'_Int_Int_buf_r  = (& \mergeHP_CTmain_map'_Int_Int_buf_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \mergeHP_CTmain_map'_Int_Int_buf_emitted  <= 3'd0;
    else
      \mergeHP_CTmain_map'_Int_Int_buf_emitted  <= (\mergeHP_CTmain_map'_Int_Int_buf_r  ? 3'd0 :
                                                    \mergeHP_CTmain_map'_Int_Int_buf_done );
  
  /* mergectrl (Ty C2,
           Ty MemIn_CTmain_map'_Int_Int) : [(dconReadIn_CTmain_map'_Int_Int,MemIn_CTmain_map'_Int_Int),
                                            (dconWriteIn_CTmain_map'_Int_Int,MemIn_CTmain_map'_Int_Int)] > (memMergeChoice_CTmain_map'_Int_Int,C2) (memMergeIn_CTmain_map'_Int_Int,MemIn_CTmain_map'_Int_Int) */
  logic [1:0] \dconReadIn_CTmain_map'_Int_Int_select_d ;
  assign \dconReadIn_CTmain_map'_Int_Int_select_d  = ((| \dconReadIn_CTmain_map'_Int_Int_select_q ) ? \dconReadIn_CTmain_map'_Int_Int_select_q  :
                                                      (\dconReadIn_CTmain_map'_Int_Int_d [0] ? 2'd1 :
                                                       (\dconWriteIn_CTmain_map'_Int_Int_d [0] ? 2'd2 :
                                                        2'd0)));
  logic [1:0] \dconReadIn_CTmain_map'_Int_Int_select_q ;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \dconReadIn_CTmain_map'_Int_Int_select_q  <= 2'd0;
    else
      \dconReadIn_CTmain_map'_Int_Int_select_q  <= (\dconReadIn_CTmain_map'_Int_Int_done  ? 2'd0 :
                                                    \dconReadIn_CTmain_map'_Int_Int_select_d );
  logic [1:0] \dconReadIn_CTmain_map'_Int_Int_emit_q ;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \dconReadIn_CTmain_map'_Int_Int_emit_q  <= 2'd0;
    else
      \dconReadIn_CTmain_map'_Int_Int_emit_q  <= (\dconReadIn_CTmain_map'_Int_Int_done  ? 2'd0 :
                                                  \dconReadIn_CTmain_map'_Int_Int_emit_d );
  logic [1:0] \dconReadIn_CTmain_map'_Int_Int_emit_d ;
  assign \dconReadIn_CTmain_map'_Int_Int_emit_d  = (\dconReadIn_CTmain_map'_Int_Int_emit_q  | ({\memMergeChoice_CTmain_map'_Int_Int_d [0],
                                                                                                \memMergeIn_CTmain_map'_Int_Int_d [0]} & {\memMergeChoice_CTmain_map'_Int_Int_r ,
                                                                                                                                          \memMergeIn_CTmain_map'_Int_Int_r }));
  logic \dconReadIn_CTmain_map'_Int_Int_done ;
  assign \dconReadIn_CTmain_map'_Int_Int_done  = (& \dconReadIn_CTmain_map'_Int_Int_emit_d );
  assign {\dconWriteIn_CTmain_map'_Int_Int_r ,
          \dconReadIn_CTmain_map'_Int_Int_r } = (\dconReadIn_CTmain_map'_Int_Int_done  ? \dconReadIn_CTmain_map'_Int_Int_select_d  :
                                                 2'd0);
  assign \memMergeIn_CTmain_map'_Int_Int_d  = ((\dconReadIn_CTmain_map'_Int_Int_select_d [0] && (! \dconReadIn_CTmain_map'_Int_Int_emit_q [0])) ? \dconReadIn_CTmain_map'_Int_Int_d  :
                                               ((\dconReadIn_CTmain_map'_Int_Int_select_d [1] && (! \dconReadIn_CTmain_map'_Int_Int_emit_q [0])) ? \dconWriteIn_CTmain_map'_Int_Int_d  :
                                                {84'd0, 1'd0}));
  assign \memMergeChoice_CTmain_map'_Int_Int_d  = ((\dconReadIn_CTmain_map'_Int_Int_select_d [0] && (! \dconReadIn_CTmain_map'_Int_Int_emit_q [1])) ? C1_2_dc(1'd1) :
                                                   ((\dconReadIn_CTmain_map'_Int_Int_select_d [1] && (! \dconReadIn_CTmain_map'_Int_Int_emit_q [1])) ? C2_2_dc(1'd1) :
                                                    {1'd0, 1'd0}));
  
  /* bram (Ty MemIn_CTmain_map'_Int_Int,
      Ty MemOut_CTmain_map'_Int_Int) : (memMergeIn_CTmain_map'_Int_Int_dbuf,MemIn_CTmain_map'_Int_Int) > (memOut_CTmain_map'_Int_Int,MemOut_CTmain_map'_Int_Int) */
  logic [66:0] \memMergeIn_CTmain_map'_Int_Int_dbuf_mem [65535:0];
  logic [15:0] \memMergeIn_CTmain_map'_Int_Int_dbuf_address ;
  logic [66:0] \memMergeIn_CTmain_map'_Int_Int_dbuf_din ;
  logic [66:0] \memOut_CTmain_map'_Int_Int_q ;
  logic \memOut_CTmain_map'_Int_Int_valid ;
  logic \memMergeIn_CTmain_map'_Int_Int_dbuf_we ;
  logic \memOut_CTmain_map'_Int_Int_we ;
  assign \memMergeIn_CTmain_map'_Int_Int_dbuf_din  = \memMergeIn_CTmain_map'_Int_Int_dbuf_d [84:18];
  assign \memMergeIn_CTmain_map'_Int_Int_dbuf_address  = \memMergeIn_CTmain_map'_Int_Int_dbuf_d [17:2];
  assign \memMergeIn_CTmain_map'_Int_Int_dbuf_we  = (\memMergeIn_CTmain_map'_Int_Int_dbuf_d [1:1] && \memMergeIn_CTmain_map'_Int_Int_dbuf_d [0]);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        \memOut_CTmain_map'_Int_Int_we  <= 1'd0;
        \memOut_CTmain_map'_Int_Int_valid  <= 1'd0;
      end
    else
      begin
        \memOut_CTmain_map'_Int_Int_we  <= \memMergeIn_CTmain_map'_Int_Int_dbuf_we ;
        \memOut_CTmain_map'_Int_Int_valid  <= \memMergeIn_CTmain_map'_Int_Int_dbuf_d [0];
        if (\memMergeIn_CTmain_map'_Int_Int_dbuf_we )
          begin
            \memMergeIn_CTmain_map'_Int_Int_dbuf_mem [\memMergeIn_CTmain_map'_Int_Int_dbuf_address ] <= \memMergeIn_CTmain_map'_Int_Int_dbuf_din ;
            \memOut_CTmain_map'_Int_Int_q  <= \memMergeIn_CTmain_map'_Int_Int_dbuf_din ;
          end
        else
          \memOut_CTmain_map'_Int_Int_q  <= \memMergeIn_CTmain_map'_Int_Int_dbuf_mem [\memMergeIn_CTmain_map'_Int_Int_dbuf_address ];
      end
  assign \memOut_CTmain_map'_Int_Int_d  = {\memOut_CTmain_map'_Int_Int_q ,
                                           \memOut_CTmain_map'_Int_Int_we ,
                                           \memOut_CTmain_map'_Int_Int_valid };
  assign \memMergeIn_CTmain_map'_Int_Int_dbuf_r  = ((! \memOut_CTmain_map'_Int_Int_valid ) || \memOut_CTmain_map'_Int_Int_r );
  
  /* demux (Ty C2,
       Ty MemOut_CTmain_map'_Int_Int) : (memMergeChoice_CTmain_map'_Int_Int,C2) (memOut_CTmain_map'_Int_Int_dbuf,MemOut_CTmain_map'_Int_Int) > [(memReadOut_CTmain_map'_Int_Int,MemOut_CTmain_map'_Int_Int),
                                                                                                                                                (memWriteOut_CTmain_map'_Int_Int,MemOut_CTmain_map'_Int_Int)] */
  logic [1:0] \memOut_CTmain_map'_Int_Int_dbuf_onehotd ;
  always_comb
    if ((\memMergeChoice_CTmain_map'_Int_Int_d [0] && \memOut_CTmain_map'_Int_Int_dbuf_d [0]))
      unique case (\memMergeChoice_CTmain_map'_Int_Int_d [1:1])
        1'd0: \memOut_CTmain_map'_Int_Int_dbuf_onehotd  = 2'd1;
        1'd1: \memOut_CTmain_map'_Int_Int_dbuf_onehotd  = 2'd2;
        default: \memOut_CTmain_map'_Int_Int_dbuf_onehotd  = 2'd0;
      endcase
    else \memOut_CTmain_map'_Int_Int_dbuf_onehotd  = 2'd0;
  assign \memReadOut_CTmain_map'_Int_Int_d  = {\memOut_CTmain_map'_Int_Int_dbuf_d [68:1],
                                               \memOut_CTmain_map'_Int_Int_dbuf_onehotd [0]};
  assign \memWriteOut_CTmain_map'_Int_Int_d  = {\memOut_CTmain_map'_Int_Int_dbuf_d [68:1],
                                                \memOut_CTmain_map'_Int_Int_dbuf_onehotd [1]};
  assign \memOut_CTmain_map'_Int_Int_dbuf_r  = (| (\memOut_CTmain_map'_Int_Int_dbuf_onehotd  & {\memWriteOut_CTmain_map'_Int_Int_r ,
                                                                                                \memReadOut_CTmain_map'_Int_Int_r }));
  assign \memMergeChoice_CTmain_map'_Int_Int_r  = \memOut_CTmain_map'_Int_Int_dbuf_r ;
  
  /* dbuf (Ty MemIn_CTmain_map'_Int_Int) : (memMergeIn_CTmain_map'_Int_Int_rbuf,MemIn_CTmain_map'_Int_Int) > (memMergeIn_CTmain_map'_Int_Int_dbuf,MemIn_CTmain_map'_Int_Int) */
  assign \memMergeIn_CTmain_map'_Int_Int_rbuf_r  = ((! \memMergeIn_CTmain_map'_Int_Int_dbuf_d [0]) || \memMergeIn_CTmain_map'_Int_Int_dbuf_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \memMergeIn_CTmain_map'_Int_Int_dbuf_d  <= {84'd0, 1'd0};
    else
      if (\memMergeIn_CTmain_map'_Int_Int_rbuf_r )
        \memMergeIn_CTmain_map'_Int_Int_dbuf_d  <= \memMergeIn_CTmain_map'_Int_Int_rbuf_d ;
  
  /* rbuf (Ty MemIn_CTmain_map'_Int_Int) : (memMergeIn_CTmain_map'_Int_Int,MemIn_CTmain_map'_Int_Int) > (memMergeIn_CTmain_map'_Int_Int_rbuf,MemIn_CTmain_map'_Int_Int) */
  \MemIn_CTmain_map'_Int_Int_t  \memMergeIn_CTmain_map'_Int_Int_buf ;
  assign \memMergeIn_CTmain_map'_Int_Int_r  = (! \memMergeIn_CTmain_map'_Int_Int_buf [0]);
  assign \memMergeIn_CTmain_map'_Int_Int_rbuf_d  = (\memMergeIn_CTmain_map'_Int_Int_buf [0] ? \memMergeIn_CTmain_map'_Int_Int_buf  :
                                                    \memMergeIn_CTmain_map'_Int_Int_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \memMergeIn_CTmain_map'_Int_Int_buf  <= {84'd0, 1'd0};
    else
      if ((\memMergeIn_CTmain_map'_Int_Int_rbuf_r  && \memMergeIn_CTmain_map'_Int_Int_buf [0]))
        \memMergeIn_CTmain_map'_Int_Int_buf  <= {84'd0, 1'd0};
      else if (((! \memMergeIn_CTmain_map'_Int_Int_rbuf_r ) && (! \memMergeIn_CTmain_map'_Int_Int_buf [0])))
        \memMergeIn_CTmain_map'_Int_Int_buf  <= \memMergeIn_CTmain_map'_Int_Int_d ;
  
  /* dbuf (Ty MemOut_CTmain_map'_Int_Int) : (memOut_CTmain_map'_Int_Int_rbuf,MemOut_CTmain_map'_Int_Int) > (memOut_CTmain_map'_Int_Int_dbuf,MemOut_CTmain_map'_Int_Int) */
  assign \memOut_CTmain_map'_Int_Int_rbuf_r  = ((! \memOut_CTmain_map'_Int_Int_dbuf_d [0]) || \memOut_CTmain_map'_Int_Int_dbuf_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \memOut_CTmain_map'_Int_Int_dbuf_d  <= {68'd0, 1'd0};
    else
      if (\memOut_CTmain_map'_Int_Int_rbuf_r )
        \memOut_CTmain_map'_Int_Int_dbuf_d  <= \memOut_CTmain_map'_Int_Int_rbuf_d ;
  
  /* rbuf (Ty MemOut_CTmain_map'_Int_Int) : (memOut_CTmain_map'_Int_Int,MemOut_CTmain_map'_Int_Int) > (memOut_CTmain_map'_Int_Int_rbuf,MemOut_CTmain_map'_Int_Int) */
  \MemOut_CTmain_map'_Int_Int_t  \memOut_CTmain_map'_Int_Int_buf ;
  assign \memOut_CTmain_map'_Int_Int_r  = (! \memOut_CTmain_map'_Int_Int_buf [0]);
  assign \memOut_CTmain_map'_Int_Int_rbuf_d  = (\memOut_CTmain_map'_Int_Int_buf [0] ? \memOut_CTmain_map'_Int_Int_buf  :
                                                \memOut_CTmain_map'_Int_Int_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \memOut_CTmain_map'_Int_Int_buf  <= {68'd0, 1'd0};
    else
      if ((\memOut_CTmain_map'_Int_Int_rbuf_r  && \memOut_CTmain_map'_Int_Int_buf [0]))
        \memOut_CTmain_map'_Int_Int_buf  <= {68'd0, 1'd0};
      else if (((! \memOut_CTmain_map'_Int_Int_rbuf_r ) && (! \memOut_CTmain_map'_Int_Int_buf [0])))
        \memOut_CTmain_map'_Int_Int_buf  <= \memOut_CTmain_map'_Int_Int_d ;
  
  /* destruct (Ty Pointer_CTmain_map'_Int_Int,
          Dcon Pointer_CTmain_map'_Int_Int) : (scfarg_0_2_1_argbuf,Pointer_CTmain_map'_Int_Int) > [(destructReadIn_CTmain_map'_Int_Int,Word16#)] */
  assign \destructReadIn_CTmain_map'_Int_Int_d  = {scfarg_0_2_1_argbuf_d[16:1],
                                                   scfarg_0_2_1_argbuf_d[0]};
  assign scfarg_0_2_1_argbuf_r = \destructReadIn_CTmain_map'_Int_Int_r ;
  
  /* dcon (Ty MemIn_CTmain_map'_Int_Int,
      Dcon ReadIn_CTmain_map'_Int_Int) : [(destructReadIn_CTmain_map'_Int_Int,Word16#)] > (dconReadIn_CTmain_map'_Int_Int,MemIn_CTmain_map'_Int_Int) */
  assign \dconReadIn_CTmain_map'_Int_Int_d  = \ReadIn_CTmain_map'_Int_Int_dc ((& {\destructReadIn_CTmain_map'_Int_Int_d [0]}), \destructReadIn_CTmain_map'_Int_Int_d );
  assign {\destructReadIn_CTmain_map'_Int_Int_r } = {1 {(\dconReadIn_CTmain_map'_Int_Int_r  && \dconReadIn_CTmain_map'_Int_Int_d [0])}};
  
  /* destruct (Ty MemOut_CTmain_map'_Int_Int,
          Dcon ReadOut_CTmain_map'_Int_Int) : (memReadOut_CTmain_map'_Int_Int,MemOut_CTmain_map'_Int_Int) > [(readPointer_CTmain_map'_Int_Intscfarg_0_2_1_argbuf,CTmain_map'_Int_Int)] */
  assign \readPointer_CTmain_map'_Int_Intscfarg_0_2_1_argbuf_d  = {\memReadOut_CTmain_map'_Int_Int_d [68:2],
                                                                   \memReadOut_CTmain_map'_Int_Int_d [0]};
  assign \memReadOut_CTmain_map'_Int_Int_r  = \readPointer_CTmain_map'_Int_Intscfarg_0_2_1_argbuf_r ;
  
  /* mergectrl (Ty C5,
           Ty CTmain_map'_Int_Int) : [(lizzieLet14_1_argbuf,CTmain_map'_Int_Int),
                                      (lizzieLet23_1_argbuf,CTmain_map'_Int_Int),
                                      (lizzieLet35_1_argbuf,CTmain_map'_Int_Int),
                                      (lizzieLet36_1_argbuf,CTmain_map'_Int_Int),
                                      (lizzieLet37_1_argbuf,CTmain_map'_Int_Int)] > (writeMerge_choice_CTmain_map'_Int_Int,C5) (writeMerge_data_CTmain_map'_Int_Int,CTmain_map'_Int_Int) */
  logic [4:0] lizzieLet14_1_argbuf_select_d;
  assign lizzieLet14_1_argbuf_select_d = ((| lizzieLet14_1_argbuf_select_q) ? lizzieLet14_1_argbuf_select_q :
                                          (lizzieLet14_1_argbuf_d[0] ? 5'd1 :
                                           (lizzieLet23_1_argbuf_d[0] ? 5'd2 :
                                            (lizzieLet35_1_argbuf_d[0] ? 5'd4 :
                                             (lizzieLet36_1_argbuf_d[0] ? 5'd8 :
                                              (lizzieLet37_1_argbuf_d[0] ? 5'd16 :
                                               5'd0))))));
  logic [4:0] lizzieLet14_1_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet14_1_argbuf_select_q <= 5'd0;
    else
      lizzieLet14_1_argbuf_select_q <= (lizzieLet14_1_argbuf_done ? 5'd0 :
                                        lizzieLet14_1_argbuf_select_d);
  logic [1:0] lizzieLet14_1_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet14_1_argbuf_emit_q <= 2'd0;
    else
      lizzieLet14_1_argbuf_emit_q <= (lizzieLet14_1_argbuf_done ? 2'd0 :
                                      lizzieLet14_1_argbuf_emit_d);
  logic [1:0] lizzieLet14_1_argbuf_emit_d;
  assign lizzieLet14_1_argbuf_emit_d = (lizzieLet14_1_argbuf_emit_q | ({\writeMerge_choice_CTmain_map'_Int_Int_d [0],
                                                                        \writeMerge_data_CTmain_map'_Int_Int_d [0]} & {\writeMerge_choice_CTmain_map'_Int_Int_r ,
                                                                                                                       \writeMerge_data_CTmain_map'_Int_Int_r }));
  logic lizzieLet14_1_argbuf_done;
  assign lizzieLet14_1_argbuf_done = (& lizzieLet14_1_argbuf_emit_d);
  assign {lizzieLet37_1_argbuf_r,
          lizzieLet36_1_argbuf_r,
          lizzieLet35_1_argbuf_r,
          lizzieLet23_1_argbuf_r,
          lizzieLet14_1_argbuf_r} = (lizzieLet14_1_argbuf_done ? lizzieLet14_1_argbuf_select_d :
                                     5'd0);
  assign \writeMerge_data_CTmain_map'_Int_Int_d  = ((lizzieLet14_1_argbuf_select_d[0] && (! lizzieLet14_1_argbuf_emit_q[0])) ? lizzieLet14_1_argbuf_d :
                                                    ((lizzieLet14_1_argbuf_select_d[1] && (! lizzieLet14_1_argbuf_emit_q[0])) ? lizzieLet23_1_argbuf_d :
                                                     ((lizzieLet14_1_argbuf_select_d[2] && (! lizzieLet14_1_argbuf_emit_q[0])) ? lizzieLet35_1_argbuf_d :
                                                      ((lizzieLet14_1_argbuf_select_d[3] && (! lizzieLet14_1_argbuf_emit_q[0])) ? lizzieLet36_1_argbuf_d :
                                                       ((lizzieLet14_1_argbuf_select_d[4] && (! lizzieLet14_1_argbuf_emit_q[0])) ? lizzieLet37_1_argbuf_d :
                                                        {67'd0, 1'd0})))));
  assign \writeMerge_choice_CTmain_map'_Int_Int_d  = ((lizzieLet14_1_argbuf_select_d[0] && (! lizzieLet14_1_argbuf_emit_q[1])) ? C1_5_dc(1'd1) :
                                                      ((lizzieLet14_1_argbuf_select_d[1] && (! lizzieLet14_1_argbuf_emit_q[1])) ? C2_5_dc(1'd1) :
                                                       ((lizzieLet14_1_argbuf_select_d[2] && (! lizzieLet14_1_argbuf_emit_q[1])) ? C3_5_dc(1'd1) :
                                                        ((lizzieLet14_1_argbuf_select_d[3] && (! lizzieLet14_1_argbuf_emit_q[1])) ? C4_5_dc(1'd1) :
                                                         ((lizzieLet14_1_argbuf_select_d[4] && (! lizzieLet14_1_argbuf_emit_q[1])) ? C5_5_dc(1'd1) :
                                                          {3'd0, 1'd0})))));
  
  /* demux (Ty C5,
       Ty Pointer_CTmain_map'_Int_Int) : (writeMerge_choice_CTmain_map'_Int_Int,C5) (demuxWriteResult_CTmain_map'_Int_Int,Pointer_CTmain_map'_Int_Int) > [(writeCTmain_map'_Int_IntlizzieLet14_1_argbuf,Pointer_CTmain_map'_Int_Int),
                                                                                                                                                          (writeCTmain_map'_Int_IntlizzieLet23_1_argbuf,Pointer_CTmain_map'_Int_Int),
                                                                                                                                                          (writeCTmain_map'_Int_IntlizzieLet35_1_argbuf,Pointer_CTmain_map'_Int_Int),
                                                                                                                                                          (writeCTmain_map'_Int_IntlizzieLet36_1_argbuf,Pointer_CTmain_map'_Int_Int),
                                                                                                                                                          (writeCTmain_map'_Int_IntlizzieLet37_1_argbuf,Pointer_CTmain_map'_Int_Int)] */
  logic [4:0] \demuxWriteResult_CTmain_map'_Int_Int_onehotd ;
  always_comb
    if ((\writeMerge_choice_CTmain_map'_Int_Int_d [0] && \demuxWriteResult_CTmain_map'_Int_Int_d [0]))
      unique case (\writeMerge_choice_CTmain_map'_Int_Int_d [3:1])
        3'd0: \demuxWriteResult_CTmain_map'_Int_Int_onehotd  = 5'd1;
        3'd1: \demuxWriteResult_CTmain_map'_Int_Int_onehotd  = 5'd2;
        3'd2: \demuxWriteResult_CTmain_map'_Int_Int_onehotd  = 5'd4;
        3'd3: \demuxWriteResult_CTmain_map'_Int_Int_onehotd  = 5'd8;
        3'd4: \demuxWriteResult_CTmain_map'_Int_Int_onehotd  = 5'd16;
        default: \demuxWriteResult_CTmain_map'_Int_Int_onehotd  = 5'd0;
      endcase
    else \demuxWriteResult_CTmain_map'_Int_Int_onehotd  = 5'd0;
  assign \writeCTmain_map'_Int_IntlizzieLet14_1_argbuf_d  = {\demuxWriteResult_CTmain_map'_Int_Int_d [16:1],
                                                             \demuxWriteResult_CTmain_map'_Int_Int_onehotd [0]};
  assign \writeCTmain_map'_Int_IntlizzieLet23_1_argbuf_d  = {\demuxWriteResult_CTmain_map'_Int_Int_d [16:1],
                                                             \demuxWriteResult_CTmain_map'_Int_Int_onehotd [1]};
  assign \writeCTmain_map'_Int_IntlizzieLet35_1_argbuf_d  = {\demuxWriteResult_CTmain_map'_Int_Int_d [16:1],
                                                             \demuxWriteResult_CTmain_map'_Int_Int_onehotd [2]};
  assign \writeCTmain_map'_Int_IntlizzieLet36_1_argbuf_d  = {\demuxWriteResult_CTmain_map'_Int_Int_d [16:1],
                                                             \demuxWriteResult_CTmain_map'_Int_Int_onehotd [3]};
  assign \writeCTmain_map'_Int_IntlizzieLet37_1_argbuf_d  = {\demuxWriteResult_CTmain_map'_Int_Int_d [16:1],
                                                             \demuxWriteResult_CTmain_map'_Int_Int_onehotd [4]};
  assign \demuxWriteResult_CTmain_map'_Int_Int_r  = (| (\demuxWriteResult_CTmain_map'_Int_Int_onehotd  & {\writeCTmain_map'_Int_IntlizzieLet37_1_argbuf_r ,
                                                                                                          \writeCTmain_map'_Int_IntlizzieLet36_1_argbuf_r ,
                                                                                                          \writeCTmain_map'_Int_IntlizzieLet35_1_argbuf_r ,
                                                                                                          \writeCTmain_map'_Int_IntlizzieLet23_1_argbuf_r ,
                                                                                                          \writeCTmain_map'_Int_IntlizzieLet14_1_argbuf_r }));
  assign \writeMerge_choice_CTmain_map'_Int_Int_r  = \demuxWriteResult_CTmain_map'_Int_Int_r ;
  
  /* dcon (Ty MemIn_CTmain_map'_Int_Int,
      Dcon WriteIn_CTmain_map'_Int_Int) : [(forkHP1_CTmain_map'_Int_In2,Word16#),
                                           (writeMerge_data_CTmain_map'_Int_Int,CTmain_map'_Int_Int)] > (dconWriteIn_CTmain_map'_Int_Int,MemIn_CTmain_map'_Int_Int) */
  assign \dconWriteIn_CTmain_map'_Int_Int_d  = \WriteIn_CTmain_map'_Int_Int_dc ((& {\forkHP1_CTmain_map'_Int_In2_d [0],
                                                                                    \writeMerge_data_CTmain_map'_Int_Int_d [0]}), \forkHP1_CTmain_map'_Int_In2_d , \writeMerge_data_CTmain_map'_Int_Int_d );
  assign {\forkHP1_CTmain_map'_Int_In2_r ,
          \writeMerge_data_CTmain_map'_Int_Int_r } = {2 {(\dconWriteIn_CTmain_map'_Int_Int_r  && \dconWriteIn_CTmain_map'_Int_Int_d [0])}};
  
  /* dcon (Ty Pointer_CTmain_map'_Int_Int,
      Dcon Pointer_CTmain_map'_Int_Int) : [(forkHP1_CTmain_map'_Int_In3,Word16#)] > (dconPtr_CTmain_map'_Int_Int,Pointer_CTmain_map'_Int_Int) */
  assign \dconPtr_CTmain_map'_Int_Int_d  = \Pointer_CTmain_map'_Int_Int_dc ((& {\forkHP1_CTmain_map'_Int_In3_d [0]}), \forkHP1_CTmain_map'_Int_In3_d );
  assign {\forkHP1_CTmain_map'_Int_In3_r } = {1 {(\dconPtr_CTmain_map'_Int_Int_r  && \dconPtr_CTmain_map'_Int_Int_d [0])}};
  
  /* demux (Ty MemOut_CTmain_map'_Int_Int,
       Ty Pointer_CTmain_map'_Int_Int) : (memWriteOut_CTmain_map'_Int_Int,MemOut_CTmain_map'_Int_Int) (dconPtr_CTmain_map'_Int_Int,Pointer_CTmain_map'_Int_Int) > [(_37,Pointer_CTmain_map'_Int_Int),
                                                                                                                                                                   (demuxWriteResult_CTmain_map'_Int_Int,Pointer_CTmain_map'_Int_Int)] */
  logic [1:0] \dconPtr_CTmain_map'_Int_Int_onehotd ;
  always_comb
    if ((\memWriteOut_CTmain_map'_Int_Int_d [0] && \dconPtr_CTmain_map'_Int_Int_d [0]))
      unique case (\memWriteOut_CTmain_map'_Int_Int_d [1:1])
        1'd0: \dconPtr_CTmain_map'_Int_Int_onehotd  = 2'd1;
        1'd1: \dconPtr_CTmain_map'_Int_Int_onehotd  = 2'd2;
        default: \dconPtr_CTmain_map'_Int_Int_onehotd  = 2'd0;
      endcase
    else \dconPtr_CTmain_map'_Int_Int_onehotd  = 2'd0;
  assign _37_d = {\dconPtr_CTmain_map'_Int_Int_d [16:1],
                  \dconPtr_CTmain_map'_Int_Int_onehotd [0]};
  assign \demuxWriteResult_CTmain_map'_Int_Int_d  = {\dconPtr_CTmain_map'_Int_Int_d [16:1],
                                                     \dconPtr_CTmain_map'_Int_Int_onehotd [1]};
  assign \dconPtr_CTmain_map'_Int_Int_r  = (| (\dconPtr_CTmain_map'_Int_Int_onehotd  & {\demuxWriteResult_CTmain_map'_Int_Int_r ,
                                                                                        _37_r}));
  assign \memWriteOut_CTmain_map'_Int_Int_r  = \dconPtr_CTmain_map'_Int_Int_r ;
  
  /* const (Ty Word16#,
       Lit 0) : (goFor_6,Go) > (initHP_CTmap''_map''_Int_Int_Int,Word16#) */
  assign \initHP_CTmap''_map''_Int_Int_Int_d  = {16'd0,
                                                 goFor_6_d[0]};
  assign goFor_6_r = \initHP_CTmap''_map''_Int_Int_Int_r ;
  
  /* const (Ty Word16#,
       Lit 1) : (incrHP_CTmap''_map''_Int_Int_Int1,Go) > (incrHP_CTmap''_map''_Int_Int_Int,Word16#) */
  assign \incrHP_CTmap''_map''_Int_Int_Int_d  = {16'd1,
                                                 \incrHP_CTmap''_map''_Int_Int_Int1_d [0]};
  assign \incrHP_CTmap''_map''_Int_Int_Int1_r  = \incrHP_CTmap''_map''_Int_Int_Int_r ;
  
  /* merge (Ty Go) : [(goFor_7,Go),
                 (incrHP_CTmap''_map''_Int_Int_Int2,Go)] > (incrHP_mergeCTmap''_map''_Int_Int_Int,Go) */
  logic [1:0] \incrHP_mergeCTmap''_map''_Int_Int_Int_selected ;
  logic [1:0] \incrHP_mergeCTmap''_map''_Int_Int_Int_select ;
  always_comb
    begin
      \incrHP_mergeCTmap''_map''_Int_Int_Int_selected  = 2'd0;
      if ((| \incrHP_mergeCTmap''_map''_Int_Int_Int_select ))
        \incrHP_mergeCTmap''_map''_Int_Int_Int_selected  = \incrHP_mergeCTmap''_map''_Int_Int_Int_select ;
      else
        if (goFor_7_d[0])
          \incrHP_mergeCTmap''_map''_Int_Int_Int_selected [0] = 1'd1;
        else if (\incrHP_CTmap''_map''_Int_Int_Int2_d [0])
          \incrHP_mergeCTmap''_map''_Int_Int_Int_selected [1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \incrHP_mergeCTmap''_map''_Int_Int_Int_select  <= 2'd0;
    else
      \incrHP_mergeCTmap''_map''_Int_Int_Int_select  <= (\incrHP_mergeCTmap''_map''_Int_Int_Int_r  ? 2'd0 :
                                                         \incrHP_mergeCTmap''_map''_Int_Int_Int_selected );
  always_comb
    if (\incrHP_mergeCTmap''_map''_Int_Int_Int_selected [0])
      \incrHP_mergeCTmap''_map''_Int_Int_Int_d  = goFor_7_d;
    else if (\incrHP_mergeCTmap''_map''_Int_Int_Int_selected [1])
      \incrHP_mergeCTmap''_map''_Int_Int_Int_d  = \incrHP_CTmap''_map''_Int_Int_Int2_d ;
    else \incrHP_mergeCTmap''_map''_Int_Int_Int_d  = 1'd0;
  assign {\incrHP_CTmap''_map''_Int_Int_Int2_r ,
          goFor_7_r} = (\incrHP_mergeCTmap''_map''_Int_Int_Int_r  ? \incrHP_mergeCTmap''_map''_Int_Int_Int_selected  :
                        2'd0);
  
  /* fork (Ty Go) : (incrHP_mergeCTmap''_map''_Int_Int_Int_buf,Go) > [(incrHP_CTmap''_map''_Int_Int_Int1,Go),
                                                                 (incrHP_CTmap''_map''_Int_Int_Int2,Go)] */
  logic [1:0] \incrHP_mergeCTmap''_map''_Int_Int_Int_buf_emitted ;
  logic [1:0] \incrHP_mergeCTmap''_map''_Int_Int_Int_buf_done ;
  assign \incrHP_CTmap''_map''_Int_Int_Int1_d  = (\incrHP_mergeCTmap''_map''_Int_Int_Int_buf_d [0] && (! \incrHP_mergeCTmap''_map''_Int_Int_Int_buf_emitted [0]));
  assign \incrHP_CTmap''_map''_Int_Int_Int2_d  = (\incrHP_mergeCTmap''_map''_Int_Int_Int_buf_d [0] && (! \incrHP_mergeCTmap''_map''_Int_Int_Int_buf_emitted [1]));
  assign \incrHP_mergeCTmap''_map''_Int_Int_Int_buf_done  = (\incrHP_mergeCTmap''_map''_Int_Int_Int_buf_emitted  | ({\incrHP_CTmap''_map''_Int_Int_Int2_d [0],
                                                                                                                     \incrHP_CTmap''_map''_Int_Int_Int1_d [0]} & {\incrHP_CTmap''_map''_Int_Int_Int2_r ,
                                                                                                                                                                  \incrHP_CTmap''_map''_Int_Int_Int1_r }));
  assign \incrHP_mergeCTmap''_map''_Int_Int_Int_buf_r  = (& \incrHP_mergeCTmap''_map''_Int_Int_Int_buf_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \incrHP_mergeCTmap''_map''_Int_Int_Int_buf_emitted  <= 2'd0;
    else
      \incrHP_mergeCTmap''_map''_Int_Int_Int_buf_emitted  <= (\incrHP_mergeCTmap''_map''_Int_Int_Int_buf_r  ? 2'd0 :
                                                              \incrHP_mergeCTmap''_map''_Int_Int_Int_buf_done );
  
  /* op_add (Ty Word16#) : (incrHP_CTmap''_map''_Int_Int_Int,Word16#) (forkHP1_CTmap''_map''_Int_Int_Int,Word16#) > (addHP_CTmap''_map''_Int_Int_Int,Word16#) */
  assign \addHP_CTmap''_map''_Int_Int_Int_d  = {(\incrHP_CTmap''_map''_Int_Int_Int_d [16:1] + \forkHP1_CTmap''_map''_Int_Int_Int_d [16:1]),
                                                (\incrHP_CTmap''_map''_Int_Int_Int_d [0] && \forkHP1_CTmap''_map''_Int_Int_Int_d [0])};
  assign {\incrHP_CTmap''_map''_Int_Int_Int_r ,
          \forkHP1_CTmap''_map''_Int_Int_Int_r } = {2 {(\addHP_CTmap''_map''_Int_Int_Int_r  && \addHP_CTmap''_map''_Int_Int_Int_d [0])}};
  
  /* merge (Ty Word16#) : [(initHP_CTmap''_map''_Int_Int_Int,Word16#),
                      (addHP_CTmap''_map''_Int_Int_Int,Word16#)] > (mergeHP_CTmap''_map''_Int_Int_Int,Word16#) */
  logic [1:0] \mergeHP_CTmap''_map''_Int_Int_Int_selected ;
  logic [1:0] \mergeHP_CTmap''_map''_Int_Int_Int_select ;
  always_comb
    begin
      \mergeHP_CTmap''_map''_Int_Int_Int_selected  = 2'd0;
      if ((| \mergeHP_CTmap''_map''_Int_Int_Int_select ))
        \mergeHP_CTmap''_map''_Int_Int_Int_selected  = \mergeHP_CTmap''_map''_Int_Int_Int_select ;
      else
        if (\initHP_CTmap''_map''_Int_Int_Int_d [0])
          \mergeHP_CTmap''_map''_Int_Int_Int_selected [0] = 1'd1;
        else if (\addHP_CTmap''_map''_Int_Int_Int_d [0])
          \mergeHP_CTmap''_map''_Int_Int_Int_selected [1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \mergeHP_CTmap''_map''_Int_Int_Int_select  <= 2'd0;
    else
      \mergeHP_CTmap''_map''_Int_Int_Int_select  <= (\mergeHP_CTmap''_map''_Int_Int_Int_r  ? 2'd0 :
                                                     \mergeHP_CTmap''_map''_Int_Int_Int_selected );
  always_comb
    if (\mergeHP_CTmap''_map''_Int_Int_Int_selected [0])
      \mergeHP_CTmap''_map''_Int_Int_Int_d  = \initHP_CTmap''_map''_Int_Int_Int_d ;
    else if (\mergeHP_CTmap''_map''_Int_Int_Int_selected [1])
      \mergeHP_CTmap''_map''_Int_Int_Int_d  = \addHP_CTmap''_map''_Int_Int_Int_d ;
    else \mergeHP_CTmap''_map''_Int_Int_Int_d  = {16'd0, 1'd0};
  assign {\addHP_CTmap''_map''_Int_Int_Int_r ,
          \initHP_CTmap''_map''_Int_Int_Int_r } = (\mergeHP_CTmap''_map''_Int_Int_Int_r  ? \mergeHP_CTmap''_map''_Int_Int_Int_selected  :
                                                   2'd0);
  
  /* buf (Ty Go) : (incrHP_mergeCTmap''_map''_Int_Int_Int,Go) > (incrHP_mergeCTmap''_map''_Int_Int_Int_buf,Go) */
  Go_t \incrHP_mergeCTmap''_map''_Int_Int_Int_bufchan_d ;
  logic \incrHP_mergeCTmap''_map''_Int_Int_Int_bufchan_r ;
  assign \incrHP_mergeCTmap''_map''_Int_Int_Int_r  = ((! \incrHP_mergeCTmap''_map''_Int_Int_Int_bufchan_d [0]) || \incrHP_mergeCTmap''_map''_Int_Int_Int_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \incrHP_mergeCTmap''_map''_Int_Int_Int_bufchan_d  <= 1'd0;
    else
      if (\incrHP_mergeCTmap''_map''_Int_Int_Int_r )
        \incrHP_mergeCTmap''_map''_Int_Int_Int_bufchan_d  <= \incrHP_mergeCTmap''_map''_Int_Int_Int_d ;
  Go_t \incrHP_mergeCTmap''_map''_Int_Int_Int_bufchan_buf ;
  assign \incrHP_mergeCTmap''_map''_Int_Int_Int_bufchan_r  = (! \incrHP_mergeCTmap''_map''_Int_Int_Int_bufchan_buf [0]);
  assign \incrHP_mergeCTmap''_map''_Int_Int_Int_buf_d  = (\incrHP_mergeCTmap''_map''_Int_Int_Int_bufchan_buf [0] ? \incrHP_mergeCTmap''_map''_Int_Int_Int_bufchan_buf  :
                                                          \incrHP_mergeCTmap''_map''_Int_Int_Int_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \incrHP_mergeCTmap''_map''_Int_Int_Int_bufchan_buf  <= 1'd0;
    else
      if ((\incrHP_mergeCTmap''_map''_Int_Int_Int_buf_r  && \incrHP_mergeCTmap''_map''_Int_Int_Int_bufchan_buf [0]))
        \incrHP_mergeCTmap''_map''_Int_Int_Int_bufchan_buf  <= 1'd0;
      else if (((! \incrHP_mergeCTmap''_map''_Int_Int_Int_buf_r ) && (! \incrHP_mergeCTmap''_map''_Int_Int_Int_bufchan_buf [0])))
        \incrHP_mergeCTmap''_map''_Int_Int_Int_bufchan_buf  <= \incrHP_mergeCTmap''_map''_Int_Int_Int_bufchan_d ;
  
  /* buf (Ty Word16#) : (mergeHP_CTmap''_map''_Int_Int_Int,Word16#) > (mergeHP_CTmap''_map''_Int_Int_Int_buf,Word16#) */
  \Word16#_t  \mergeHP_CTmap''_map''_Int_Int_Int_bufchan_d ;
  logic \mergeHP_CTmap''_map''_Int_Int_Int_bufchan_r ;
  assign \mergeHP_CTmap''_map''_Int_Int_Int_r  = ((! \mergeHP_CTmap''_map''_Int_Int_Int_bufchan_d [0]) || \mergeHP_CTmap''_map''_Int_Int_Int_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \mergeHP_CTmap''_map''_Int_Int_Int_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\mergeHP_CTmap''_map''_Int_Int_Int_r )
        \mergeHP_CTmap''_map''_Int_Int_Int_bufchan_d  <= \mergeHP_CTmap''_map''_Int_Int_Int_d ;
  \Word16#_t  \mergeHP_CTmap''_map''_Int_Int_Int_bufchan_buf ;
  assign \mergeHP_CTmap''_map''_Int_Int_Int_bufchan_r  = (! \mergeHP_CTmap''_map''_Int_Int_Int_bufchan_buf [0]);
  assign \mergeHP_CTmap''_map''_Int_Int_Int_buf_d  = (\mergeHP_CTmap''_map''_Int_Int_Int_bufchan_buf [0] ? \mergeHP_CTmap''_map''_Int_Int_Int_bufchan_buf  :
                                                      \mergeHP_CTmap''_map''_Int_Int_Int_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \mergeHP_CTmap''_map''_Int_Int_Int_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((\mergeHP_CTmap''_map''_Int_Int_Int_buf_r  && \mergeHP_CTmap''_map''_Int_Int_Int_bufchan_buf [0]))
        \mergeHP_CTmap''_map''_Int_Int_Int_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! \mergeHP_CTmap''_map''_Int_Int_Int_buf_r ) && (! \mergeHP_CTmap''_map''_Int_Int_Int_bufchan_buf [0])))
        \mergeHP_CTmap''_map''_Int_Int_Int_bufchan_buf  <= \mergeHP_CTmap''_map''_Int_Int_Int_bufchan_d ;
  
  /* fork (Ty Word16#) : (mergeHP_CTmap''_map''_Int_Int_Int_buf,Word16#) > [(forkHP1_CTmap''_map''_Int_Int_Int,Word16#),
                                                                       (forkHP1_CTmap''_map''_Int_Int_In2,Word16#),
                                                                       (forkHP1_CTmap''_map''_Int_Int_In3,Word16#)] */
  logic [2:0] \mergeHP_CTmap''_map''_Int_Int_Int_buf_emitted ;
  logic [2:0] \mergeHP_CTmap''_map''_Int_Int_Int_buf_done ;
  assign \forkHP1_CTmap''_map''_Int_Int_Int_d  = {\mergeHP_CTmap''_map''_Int_Int_Int_buf_d [16:1],
                                                  (\mergeHP_CTmap''_map''_Int_Int_Int_buf_d [0] && (! \mergeHP_CTmap''_map''_Int_Int_Int_buf_emitted [0]))};
  assign \forkHP1_CTmap''_map''_Int_Int_In2_d  = {\mergeHP_CTmap''_map''_Int_Int_Int_buf_d [16:1],
                                                  (\mergeHP_CTmap''_map''_Int_Int_Int_buf_d [0] && (! \mergeHP_CTmap''_map''_Int_Int_Int_buf_emitted [1]))};
  assign \forkHP1_CTmap''_map''_Int_Int_In3_d  = {\mergeHP_CTmap''_map''_Int_Int_Int_buf_d [16:1],
                                                  (\mergeHP_CTmap''_map''_Int_Int_Int_buf_d [0] && (! \mergeHP_CTmap''_map''_Int_Int_Int_buf_emitted [2]))};
  assign \mergeHP_CTmap''_map''_Int_Int_Int_buf_done  = (\mergeHP_CTmap''_map''_Int_Int_Int_buf_emitted  | ({\forkHP1_CTmap''_map''_Int_Int_In3_d [0],
                                                                                                             \forkHP1_CTmap''_map''_Int_Int_In2_d [0],
                                                                                                             \forkHP1_CTmap''_map''_Int_Int_Int_d [0]} & {\forkHP1_CTmap''_map''_Int_Int_In3_r ,
                                                                                                                                                          \forkHP1_CTmap''_map''_Int_Int_In2_r ,
                                                                                                                                                          \forkHP1_CTmap''_map''_Int_Int_Int_r }));
  assign \mergeHP_CTmap''_map''_Int_Int_Int_buf_r  = (& \mergeHP_CTmap''_map''_Int_Int_Int_buf_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \mergeHP_CTmap''_map''_Int_Int_Int_buf_emitted  <= 3'd0;
    else
      \mergeHP_CTmap''_map''_Int_Int_Int_buf_emitted  <= (\mergeHP_CTmap''_map''_Int_Int_Int_buf_r  ? 3'd0 :
                                                          \mergeHP_CTmap''_map''_Int_Int_Int_buf_done );
  
  /* mergectrl (Ty C2,
           Ty MemIn_CTmap''_map''_Int_Int_Int) : [(dconReadIn_CTmap''_map''_Int_Int_Int,MemIn_CTmap''_map''_Int_Int_Int),
                                                  (dconWriteIn_CTmap''_map''_Int_Int_Int,MemIn_CTmap''_map''_Int_Int_Int)] > (memMergeChoice_CTmap''_map''_Int_Int_Int,C2) (memMergeIn_CTmap''_map''_Int_Int_Int,MemIn_CTmap''_map''_Int_Int_Int) */
  logic [1:0] \dconReadIn_CTmap''_map''_Int_Int_Int_select_d ;
  assign \dconReadIn_CTmap''_map''_Int_Int_Int_select_d  = ((| \dconReadIn_CTmap''_map''_Int_Int_Int_select_q ) ? \dconReadIn_CTmap''_map''_Int_Int_Int_select_q  :
                                                            (\dconReadIn_CTmap''_map''_Int_Int_Int_d [0] ? 2'd1 :
                                                             (\dconWriteIn_CTmap''_map''_Int_Int_Int_d [0] ? 2'd2 :
                                                              2'd0)));
  logic [1:0] \dconReadIn_CTmap''_map''_Int_Int_Int_select_q ;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \dconReadIn_CTmap''_map''_Int_Int_Int_select_q  <= 2'd0;
    else
      \dconReadIn_CTmap''_map''_Int_Int_Int_select_q  <= (\dconReadIn_CTmap''_map''_Int_Int_Int_done  ? 2'd0 :
                                                          \dconReadIn_CTmap''_map''_Int_Int_Int_select_d );
  logic [1:0] \dconReadIn_CTmap''_map''_Int_Int_Int_emit_q ;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \dconReadIn_CTmap''_map''_Int_Int_Int_emit_q  <= 2'd0;
    else
      \dconReadIn_CTmap''_map''_Int_Int_Int_emit_q  <= (\dconReadIn_CTmap''_map''_Int_Int_Int_done  ? 2'd0 :
                                                        \dconReadIn_CTmap''_map''_Int_Int_Int_emit_d );
  logic [1:0] \dconReadIn_CTmap''_map''_Int_Int_Int_emit_d ;
  assign \dconReadIn_CTmap''_map''_Int_Int_Int_emit_d  = (\dconReadIn_CTmap''_map''_Int_Int_Int_emit_q  | ({\memMergeChoice_CTmap''_map''_Int_Int_Int_d [0],
                                                                                                            \memMergeIn_CTmap''_map''_Int_Int_Int_d [0]} & {\memMergeChoice_CTmap''_map''_Int_Int_Int_r ,
                                                                                                                                                            \memMergeIn_CTmap''_map''_Int_Int_Int_r }));
  logic \dconReadIn_CTmap''_map''_Int_Int_Int_done ;
  assign \dconReadIn_CTmap''_map''_Int_Int_Int_done  = (& \dconReadIn_CTmap''_map''_Int_Int_Int_emit_d );
  assign {\dconWriteIn_CTmap''_map''_Int_Int_Int_r ,
          \dconReadIn_CTmap''_map''_Int_Int_Int_r } = (\dconReadIn_CTmap''_map''_Int_Int_Int_done  ? \dconReadIn_CTmap''_map''_Int_Int_Int_select_d  :
                                                       2'd0);
  assign \memMergeIn_CTmap''_map''_Int_Int_Int_d  = ((\dconReadIn_CTmap''_map''_Int_Int_Int_select_d [0] && (! \dconReadIn_CTmap''_map''_Int_Int_Int_emit_q [0])) ? \dconReadIn_CTmap''_map''_Int_Int_Int_d  :
                                                     ((\dconReadIn_CTmap''_map''_Int_Int_Int_select_d [1] && (! \dconReadIn_CTmap''_map''_Int_Int_Int_emit_q [0])) ? \dconWriteIn_CTmap''_map''_Int_Int_Int_d  :
                                                      {116'd0, 1'd0}));
  assign \memMergeChoice_CTmap''_map''_Int_Int_Int_d  = ((\dconReadIn_CTmap''_map''_Int_Int_Int_select_d [0] && (! \dconReadIn_CTmap''_map''_Int_Int_Int_emit_q [1])) ? C1_2_dc(1'd1) :
                                                         ((\dconReadIn_CTmap''_map''_Int_Int_Int_select_d [1] && (! \dconReadIn_CTmap''_map''_Int_Int_Int_emit_q [1])) ? C2_2_dc(1'd1) :
                                                          {1'd0, 1'd0}));
  
  /* bram (Ty MemIn_CTmap''_map''_Int_Int_Int,
      Ty MemOut_CTmap''_map''_Int_Int_Int) : (memMergeIn_CTmap''_map''_Int_Int_Int_dbuf,MemIn_CTmap''_map''_Int_Int_Int) > (memOut_CTmap''_map''_Int_Int_Int,MemOut_CTmap''_map''_Int_Int_Int) */
  logic [98:0] \memMergeIn_CTmap''_map''_Int_Int_Int_dbuf_mem [65535:0];
  logic [15:0] \memMergeIn_CTmap''_map''_Int_Int_Int_dbuf_address ;
  logic [98:0] \memMergeIn_CTmap''_map''_Int_Int_Int_dbuf_din ;
  logic [98:0] \memOut_CTmap''_map''_Int_Int_Int_q ;
  logic \memOut_CTmap''_map''_Int_Int_Int_valid ;
  logic \memMergeIn_CTmap''_map''_Int_Int_Int_dbuf_we ;
  logic \memOut_CTmap''_map''_Int_Int_Int_we ;
  assign \memMergeIn_CTmap''_map''_Int_Int_Int_dbuf_din  = \memMergeIn_CTmap''_map''_Int_Int_Int_dbuf_d [116:18];
  assign \memMergeIn_CTmap''_map''_Int_Int_Int_dbuf_address  = \memMergeIn_CTmap''_map''_Int_Int_Int_dbuf_d [17:2];
  assign \memMergeIn_CTmap''_map''_Int_Int_Int_dbuf_we  = (\memMergeIn_CTmap''_map''_Int_Int_Int_dbuf_d [1:1] && \memMergeIn_CTmap''_map''_Int_Int_Int_dbuf_d [0]);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        \memOut_CTmap''_map''_Int_Int_Int_we  <= 1'd0;
        \memOut_CTmap''_map''_Int_Int_Int_valid  <= 1'd0;
      end
    else
      begin
        \memOut_CTmap''_map''_Int_Int_Int_we  <= \memMergeIn_CTmap''_map''_Int_Int_Int_dbuf_we ;
        \memOut_CTmap''_map''_Int_Int_Int_valid  <= \memMergeIn_CTmap''_map''_Int_Int_Int_dbuf_d [0];
        if (\memMergeIn_CTmap''_map''_Int_Int_Int_dbuf_we )
          begin
            \memMergeIn_CTmap''_map''_Int_Int_Int_dbuf_mem [\memMergeIn_CTmap''_map''_Int_Int_Int_dbuf_address ] <= \memMergeIn_CTmap''_map''_Int_Int_Int_dbuf_din ;
            \memOut_CTmap''_map''_Int_Int_Int_q  <= \memMergeIn_CTmap''_map''_Int_Int_Int_dbuf_din ;
          end
        else
          \memOut_CTmap''_map''_Int_Int_Int_q  <= \memMergeIn_CTmap''_map''_Int_Int_Int_dbuf_mem [\memMergeIn_CTmap''_map''_Int_Int_Int_dbuf_address ];
      end
  assign \memOut_CTmap''_map''_Int_Int_Int_d  = {\memOut_CTmap''_map''_Int_Int_Int_q ,
                                                 \memOut_CTmap''_map''_Int_Int_Int_we ,
                                                 \memOut_CTmap''_map''_Int_Int_Int_valid };
  assign \memMergeIn_CTmap''_map''_Int_Int_Int_dbuf_r  = ((! \memOut_CTmap''_map''_Int_Int_Int_valid ) || \memOut_CTmap''_map''_Int_Int_Int_r );
  
  /* demux (Ty C2,
       Ty MemOut_CTmap''_map''_Int_Int_Int) : (memMergeChoice_CTmap''_map''_Int_Int_Int,C2) (memOut_CTmap''_map''_Int_Int_Int_dbuf,MemOut_CTmap''_map''_Int_Int_Int) > [(memReadOut_CTmap''_map''_Int_Int_Int,MemOut_CTmap''_map''_Int_Int_Int),
                                                                                                                                                                        (memWriteOut_CTmap''_map''_Int_Int_Int,MemOut_CTmap''_map''_Int_Int_Int)] */
  logic [1:0] \memOut_CTmap''_map''_Int_Int_Int_dbuf_onehotd ;
  always_comb
    if ((\memMergeChoice_CTmap''_map''_Int_Int_Int_d [0] && \memOut_CTmap''_map''_Int_Int_Int_dbuf_d [0]))
      unique case (\memMergeChoice_CTmap''_map''_Int_Int_Int_d [1:1])
        1'd0: \memOut_CTmap''_map''_Int_Int_Int_dbuf_onehotd  = 2'd1;
        1'd1: \memOut_CTmap''_map''_Int_Int_Int_dbuf_onehotd  = 2'd2;
        default: \memOut_CTmap''_map''_Int_Int_Int_dbuf_onehotd  = 2'd0;
      endcase
    else \memOut_CTmap''_map''_Int_Int_Int_dbuf_onehotd  = 2'd0;
  assign \memReadOut_CTmap''_map''_Int_Int_Int_d  = {\memOut_CTmap''_map''_Int_Int_Int_dbuf_d [100:1],
                                                     \memOut_CTmap''_map''_Int_Int_Int_dbuf_onehotd [0]};
  assign \memWriteOut_CTmap''_map''_Int_Int_Int_d  = {\memOut_CTmap''_map''_Int_Int_Int_dbuf_d [100:1],
                                                      \memOut_CTmap''_map''_Int_Int_Int_dbuf_onehotd [1]};
  assign \memOut_CTmap''_map''_Int_Int_Int_dbuf_r  = (| (\memOut_CTmap''_map''_Int_Int_Int_dbuf_onehotd  & {\memWriteOut_CTmap''_map''_Int_Int_Int_r ,
                                                                                                            \memReadOut_CTmap''_map''_Int_Int_Int_r }));
  assign \memMergeChoice_CTmap''_map''_Int_Int_Int_r  = \memOut_CTmap''_map''_Int_Int_Int_dbuf_r ;
  
  /* dbuf (Ty MemIn_CTmap''_map''_Int_Int_Int) : (memMergeIn_CTmap''_map''_Int_Int_Int_rbuf,MemIn_CTmap''_map''_Int_Int_Int) > (memMergeIn_CTmap''_map''_Int_Int_Int_dbuf,MemIn_CTmap''_map''_Int_Int_Int) */
  assign \memMergeIn_CTmap''_map''_Int_Int_Int_rbuf_r  = ((! \memMergeIn_CTmap''_map''_Int_Int_Int_dbuf_d [0]) || \memMergeIn_CTmap''_map''_Int_Int_Int_dbuf_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \memMergeIn_CTmap''_map''_Int_Int_Int_dbuf_d  <= {116'd0, 1'd0};
    else
      if (\memMergeIn_CTmap''_map''_Int_Int_Int_rbuf_r )
        \memMergeIn_CTmap''_map''_Int_Int_Int_dbuf_d  <= \memMergeIn_CTmap''_map''_Int_Int_Int_rbuf_d ;
  
  /* rbuf (Ty MemIn_CTmap''_map''_Int_Int_Int) : (memMergeIn_CTmap''_map''_Int_Int_Int,MemIn_CTmap''_map''_Int_Int_Int) > (memMergeIn_CTmap''_map''_Int_Int_Int_rbuf,MemIn_CTmap''_map''_Int_Int_Int) */
  \MemIn_CTmap''_map''_Int_Int_Int_t  \memMergeIn_CTmap''_map''_Int_Int_Int_buf ;
  assign \memMergeIn_CTmap''_map''_Int_Int_Int_r  = (! \memMergeIn_CTmap''_map''_Int_Int_Int_buf [0]);
  assign \memMergeIn_CTmap''_map''_Int_Int_Int_rbuf_d  = (\memMergeIn_CTmap''_map''_Int_Int_Int_buf [0] ? \memMergeIn_CTmap''_map''_Int_Int_Int_buf  :
                                                          \memMergeIn_CTmap''_map''_Int_Int_Int_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \memMergeIn_CTmap''_map''_Int_Int_Int_buf  <= {116'd0, 1'd0};
    else
      if ((\memMergeIn_CTmap''_map''_Int_Int_Int_rbuf_r  && \memMergeIn_CTmap''_map''_Int_Int_Int_buf [0]))
        \memMergeIn_CTmap''_map''_Int_Int_Int_buf  <= {116'd0, 1'd0};
      else if (((! \memMergeIn_CTmap''_map''_Int_Int_Int_rbuf_r ) && (! \memMergeIn_CTmap''_map''_Int_Int_Int_buf [0])))
        \memMergeIn_CTmap''_map''_Int_Int_Int_buf  <= \memMergeIn_CTmap''_map''_Int_Int_Int_d ;
  
  /* dbuf (Ty MemOut_CTmap''_map''_Int_Int_Int) : (memOut_CTmap''_map''_Int_Int_Int_rbuf,MemOut_CTmap''_map''_Int_Int_Int) > (memOut_CTmap''_map''_Int_Int_Int_dbuf,MemOut_CTmap''_map''_Int_Int_Int) */
  assign \memOut_CTmap''_map''_Int_Int_Int_rbuf_r  = ((! \memOut_CTmap''_map''_Int_Int_Int_dbuf_d [0]) || \memOut_CTmap''_map''_Int_Int_Int_dbuf_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \memOut_CTmap''_map''_Int_Int_Int_dbuf_d  <= {100'd0, 1'd0};
    else
      if (\memOut_CTmap''_map''_Int_Int_Int_rbuf_r )
        \memOut_CTmap''_map''_Int_Int_Int_dbuf_d  <= \memOut_CTmap''_map''_Int_Int_Int_rbuf_d ;
  
  /* rbuf (Ty MemOut_CTmap''_map''_Int_Int_Int) : (memOut_CTmap''_map''_Int_Int_Int,MemOut_CTmap''_map''_Int_Int_Int) > (memOut_CTmap''_map''_Int_Int_Int_rbuf,MemOut_CTmap''_map''_Int_Int_Int) */
  \MemOut_CTmap''_map''_Int_Int_Int_t  \memOut_CTmap''_map''_Int_Int_Int_buf ;
  assign \memOut_CTmap''_map''_Int_Int_Int_r  = (! \memOut_CTmap''_map''_Int_Int_Int_buf [0]);
  assign \memOut_CTmap''_map''_Int_Int_Int_rbuf_d  = (\memOut_CTmap''_map''_Int_Int_Int_buf [0] ? \memOut_CTmap''_map''_Int_Int_Int_buf  :
                                                      \memOut_CTmap''_map''_Int_Int_Int_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \memOut_CTmap''_map''_Int_Int_Int_buf  <= {100'd0, 1'd0};
    else
      if ((\memOut_CTmap''_map''_Int_Int_Int_rbuf_r  && \memOut_CTmap''_map''_Int_Int_Int_buf [0]))
        \memOut_CTmap''_map''_Int_Int_Int_buf  <= {100'd0, 1'd0};
      else if (((! \memOut_CTmap''_map''_Int_Int_Int_rbuf_r ) && (! \memOut_CTmap''_map''_Int_Int_Int_buf [0])))
        \memOut_CTmap''_map''_Int_Int_Int_buf  <= \memOut_CTmap''_map''_Int_Int_Int_d ;
  
  /* destruct (Ty Pointer_CTmap''_map''_Int_Int_Int,
          Dcon Pointer_CTmap''_map''_Int_Int_Int) : (scfarg_0_3_1_argbuf,Pointer_CTmap''_map''_Int_Int_Int) > [(destructReadIn_CTmap''_map''_Int_Int_Int,Word16#)] */
  assign \destructReadIn_CTmap''_map''_Int_Int_Int_d  = {scfarg_0_3_1_argbuf_d[16:1],
                                                         scfarg_0_3_1_argbuf_d[0]};
  assign scfarg_0_3_1_argbuf_r = \destructReadIn_CTmap''_map''_Int_Int_Int_r ;
  
  /* dcon (Ty MemIn_CTmap''_map''_Int_Int_Int,
      Dcon ReadIn_CTmap''_map''_Int_Int_Int) : [(destructReadIn_CTmap''_map''_Int_Int_Int,Word16#)] > (dconReadIn_CTmap''_map''_Int_Int_Int,MemIn_CTmap''_map''_Int_Int_Int) */
  assign \dconReadIn_CTmap''_map''_Int_Int_Int_d  = \ReadIn_CTmap''_map''_Int_Int_Int_dc ((& {\destructReadIn_CTmap''_map''_Int_Int_Int_d [0]}), \destructReadIn_CTmap''_map''_Int_Int_Int_d );
  assign {\destructReadIn_CTmap''_map''_Int_Int_Int_r } = {1 {(\dconReadIn_CTmap''_map''_Int_Int_Int_r  && \dconReadIn_CTmap''_map''_Int_Int_Int_d [0])}};
  
  /* destruct (Ty MemOut_CTmap''_map''_Int_Int_Int,
          Dcon ReadOut_CTmap''_map''_Int_Int_Int) : (memReadOut_CTmap''_map''_Int_Int_Int,MemOut_CTmap''_map''_Int_Int_Int) > [(readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf,CTmap''_map''_Int_Int_Int)] */
  assign \readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf_d  = {\memReadOut_CTmap''_map''_Int_Int_Int_d [100:2],
                                                                         \memReadOut_CTmap''_map''_Int_Int_Int_d [0]};
  assign \memReadOut_CTmap''_map''_Int_Int_Int_r  = \readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf_r ;
  
  /* mergectrl (Ty C5,
           Ty CTmap''_map''_Int_Int_Int) : [(lizzieLet20_1_argbuf,CTmap''_map''_Int_Int_Int),
                                            (lizzieLet24_1_argbuf,CTmap''_map''_Int_Int_Int),
                                            (lizzieLet40_1_argbuf,CTmap''_map''_Int_Int_Int),
                                            (lizzieLet41_1_argbuf,CTmap''_map''_Int_Int_Int),
                                            (lizzieLet42_1_argbuf,CTmap''_map''_Int_Int_Int)] > (writeMerge_choice_CTmap''_map''_Int_Int_Int,C5) (writeMerge_data_CTmap''_map''_Int_Int_Int,CTmap''_map''_Int_Int_Int) */
  logic [4:0] lizzieLet20_1_argbuf_select_d;
  assign lizzieLet20_1_argbuf_select_d = ((| lizzieLet20_1_argbuf_select_q) ? lizzieLet20_1_argbuf_select_q :
                                          (lizzieLet20_1_argbuf_d[0] ? 5'd1 :
                                           (lizzieLet24_1_argbuf_d[0] ? 5'd2 :
                                            (lizzieLet40_1_argbuf_d[0] ? 5'd4 :
                                             (lizzieLet41_1_argbuf_d[0] ? 5'd8 :
                                              (lizzieLet42_1_argbuf_d[0] ? 5'd16 :
                                               5'd0))))));
  logic [4:0] lizzieLet20_1_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet20_1_argbuf_select_q <= 5'd0;
    else
      lizzieLet20_1_argbuf_select_q <= (lizzieLet20_1_argbuf_done ? 5'd0 :
                                        lizzieLet20_1_argbuf_select_d);
  logic [1:0] lizzieLet20_1_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet20_1_argbuf_emit_q <= 2'd0;
    else
      lizzieLet20_1_argbuf_emit_q <= (lizzieLet20_1_argbuf_done ? 2'd0 :
                                      lizzieLet20_1_argbuf_emit_d);
  logic [1:0] lizzieLet20_1_argbuf_emit_d;
  assign lizzieLet20_1_argbuf_emit_d = (lizzieLet20_1_argbuf_emit_q | ({\writeMerge_choice_CTmap''_map''_Int_Int_Int_d [0],
                                                                        \writeMerge_data_CTmap''_map''_Int_Int_Int_d [0]} & {\writeMerge_choice_CTmap''_map''_Int_Int_Int_r ,
                                                                                                                             \writeMerge_data_CTmap''_map''_Int_Int_Int_r }));
  logic lizzieLet20_1_argbuf_done;
  assign lizzieLet20_1_argbuf_done = (& lizzieLet20_1_argbuf_emit_d);
  assign {lizzieLet42_1_argbuf_r,
          lizzieLet41_1_argbuf_r,
          lizzieLet40_1_argbuf_r,
          lizzieLet24_1_argbuf_r,
          lizzieLet20_1_argbuf_r} = (lizzieLet20_1_argbuf_done ? lizzieLet20_1_argbuf_select_d :
                                     5'd0);
  assign \writeMerge_data_CTmap''_map''_Int_Int_Int_d  = ((lizzieLet20_1_argbuf_select_d[0] && (! lizzieLet20_1_argbuf_emit_q[0])) ? lizzieLet20_1_argbuf_d :
                                                          ((lizzieLet20_1_argbuf_select_d[1] && (! lizzieLet20_1_argbuf_emit_q[0])) ? lizzieLet24_1_argbuf_d :
                                                           ((lizzieLet20_1_argbuf_select_d[2] && (! lizzieLet20_1_argbuf_emit_q[0])) ? lizzieLet40_1_argbuf_d :
                                                            ((lizzieLet20_1_argbuf_select_d[3] && (! lizzieLet20_1_argbuf_emit_q[0])) ? lizzieLet41_1_argbuf_d :
                                                             ((lizzieLet20_1_argbuf_select_d[4] && (! lizzieLet20_1_argbuf_emit_q[0])) ? lizzieLet42_1_argbuf_d :
                                                              {99'd0, 1'd0})))));
  assign \writeMerge_choice_CTmap''_map''_Int_Int_Int_d  = ((lizzieLet20_1_argbuf_select_d[0] && (! lizzieLet20_1_argbuf_emit_q[1])) ? C1_5_dc(1'd1) :
                                                            ((lizzieLet20_1_argbuf_select_d[1] && (! lizzieLet20_1_argbuf_emit_q[1])) ? C2_5_dc(1'd1) :
                                                             ((lizzieLet20_1_argbuf_select_d[2] && (! lizzieLet20_1_argbuf_emit_q[1])) ? C3_5_dc(1'd1) :
                                                              ((lizzieLet20_1_argbuf_select_d[3] && (! lizzieLet20_1_argbuf_emit_q[1])) ? C4_5_dc(1'd1) :
                                                               ((lizzieLet20_1_argbuf_select_d[4] && (! lizzieLet20_1_argbuf_emit_q[1])) ? C5_5_dc(1'd1) :
                                                                {3'd0, 1'd0})))));
  
  /* demux (Ty C5,
       Ty Pointer_CTmap''_map''_Int_Int_Int) : (writeMerge_choice_CTmap''_map''_Int_Int_Int,C5) (demuxWriteResult_CTmap''_map''_Int_Int_Int,Pointer_CTmap''_map''_Int_Int_Int) > [(writeCTmap''_map''_Int_Int_IntlizzieLet20_1_argbuf,Pointer_CTmap''_map''_Int_Int_Int),
                                                                                                                                                                                  (writeCTmap''_map''_Int_Int_IntlizzieLet24_1_argbuf,Pointer_CTmap''_map''_Int_Int_Int),
                                                                                                                                                                                  (writeCTmap''_map''_Int_Int_IntlizzieLet40_1_argbuf,Pointer_CTmap''_map''_Int_Int_Int),
                                                                                                                                                                                  (writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf,Pointer_CTmap''_map''_Int_Int_Int),
                                                                                                                                                                                  (writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf,Pointer_CTmap''_map''_Int_Int_Int)] */
  logic [4:0] \demuxWriteResult_CTmap''_map''_Int_Int_Int_onehotd ;
  always_comb
    if ((\writeMerge_choice_CTmap''_map''_Int_Int_Int_d [0] && \demuxWriteResult_CTmap''_map''_Int_Int_Int_d [0]))
      unique case (\writeMerge_choice_CTmap''_map''_Int_Int_Int_d [3:1])
        3'd0: \demuxWriteResult_CTmap''_map''_Int_Int_Int_onehotd  = 5'd1;
        3'd1: \demuxWriteResult_CTmap''_map''_Int_Int_Int_onehotd  = 5'd2;
        3'd2: \demuxWriteResult_CTmap''_map''_Int_Int_Int_onehotd  = 5'd4;
        3'd3: \demuxWriteResult_CTmap''_map''_Int_Int_Int_onehotd  = 5'd8;
        3'd4: \demuxWriteResult_CTmap''_map''_Int_Int_Int_onehotd  = 5'd16;
        default:
          \demuxWriteResult_CTmap''_map''_Int_Int_Int_onehotd  = 5'd0;
      endcase
    else \demuxWriteResult_CTmap''_map''_Int_Int_Int_onehotd  = 5'd0;
  assign \writeCTmap''_map''_Int_Int_IntlizzieLet20_1_argbuf_d  = {\demuxWriteResult_CTmap''_map''_Int_Int_Int_d [16:1],
                                                                   \demuxWriteResult_CTmap''_map''_Int_Int_Int_onehotd [0]};
  assign \writeCTmap''_map''_Int_Int_IntlizzieLet24_1_argbuf_d  = {\demuxWriteResult_CTmap''_map''_Int_Int_Int_d [16:1],
                                                                   \demuxWriteResult_CTmap''_map''_Int_Int_Int_onehotd [1]};
  assign \writeCTmap''_map''_Int_Int_IntlizzieLet40_1_argbuf_d  = {\demuxWriteResult_CTmap''_map''_Int_Int_Int_d [16:1],
                                                                   \demuxWriteResult_CTmap''_map''_Int_Int_Int_onehotd [2]};
  assign \writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf_d  = {\demuxWriteResult_CTmap''_map''_Int_Int_Int_d [16:1],
                                                                   \demuxWriteResult_CTmap''_map''_Int_Int_Int_onehotd [3]};
  assign \writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf_d  = {\demuxWriteResult_CTmap''_map''_Int_Int_Int_d [16:1],
                                                                   \demuxWriteResult_CTmap''_map''_Int_Int_Int_onehotd [4]};
  assign \demuxWriteResult_CTmap''_map''_Int_Int_Int_r  = (| (\demuxWriteResult_CTmap''_map''_Int_Int_Int_onehotd  & {\writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf_r ,
                                                                                                                      \writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf_r ,
                                                                                                                      \writeCTmap''_map''_Int_Int_IntlizzieLet40_1_argbuf_r ,
                                                                                                                      \writeCTmap''_map''_Int_Int_IntlizzieLet24_1_argbuf_r ,
                                                                                                                      \writeCTmap''_map''_Int_Int_IntlizzieLet20_1_argbuf_r }));
  assign \writeMerge_choice_CTmap''_map''_Int_Int_Int_r  = \demuxWriteResult_CTmap''_map''_Int_Int_Int_r ;
  
  /* dcon (Ty MemIn_CTmap''_map''_Int_Int_Int,
      Dcon WriteIn_CTmap''_map''_Int_Int_Int) : [(forkHP1_CTmap''_map''_Int_Int_In2,Word16#),
                                                 (writeMerge_data_CTmap''_map''_Int_Int_Int,CTmap''_map''_Int_Int_Int)] > (dconWriteIn_CTmap''_map''_Int_Int_Int,MemIn_CTmap''_map''_Int_Int_Int) */
  assign \dconWriteIn_CTmap''_map''_Int_Int_Int_d  = \WriteIn_CTmap''_map''_Int_Int_Int_dc ((& {\forkHP1_CTmap''_map''_Int_Int_In2_d [0],
                                                                                                \writeMerge_data_CTmap''_map''_Int_Int_Int_d [0]}), \forkHP1_CTmap''_map''_Int_Int_In2_d , \writeMerge_data_CTmap''_map''_Int_Int_Int_d );
  assign {\forkHP1_CTmap''_map''_Int_Int_In2_r ,
          \writeMerge_data_CTmap''_map''_Int_Int_Int_r } = {2 {(\dconWriteIn_CTmap''_map''_Int_Int_Int_r  && \dconWriteIn_CTmap''_map''_Int_Int_Int_d [0])}};
  
  /* dcon (Ty Pointer_CTmap''_map''_Int_Int_Int,
      Dcon Pointer_CTmap''_map''_Int_Int_Int) : [(forkHP1_CTmap''_map''_Int_Int_In3,Word16#)] > (dconPtr_CTmap''_map''_Int_Int_Int,Pointer_CTmap''_map''_Int_Int_Int) */
  assign \dconPtr_CTmap''_map''_Int_Int_Int_d  = \Pointer_CTmap''_map''_Int_Int_Int_dc ((& {\forkHP1_CTmap''_map''_Int_Int_In3_d [0]}), \forkHP1_CTmap''_map''_Int_Int_In3_d );
  assign {\forkHP1_CTmap''_map''_Int_Int_In3_r } = {1 {(\dconPtr_CTmap''_map''_Int_Int_Int_r  && \dconPtr_CTmap''_map''_Int_Int_Int_d [0])}};
  
  /* demux (Ty MemOut_CTmap''_map''_Int_Int_Int,
       Ty Pointer_CTmap''_map''_Int_Int_Int) : (memWriteOut_CTmap''_map''_Int_Int_Int,MemOut_CTmap''_map''_Int_Int_Int) (dconPtr_CTmap''_map''_Int_Int_Int,Pointer_CTmap''_map''_Int_Int_Int) > [(_36,Pointer_CTmap''_map''_Int_Int_Int),
                                                                                                                                                                                                 (demuxWriteResult_CTmap''_map''_Int_Int_Int,Pointer_CTmap''_map''_Int_Int_Int)] */
  logic [1:0] \dconPtr_CTmap''_map''_Int_Int_Int_onehotd ;
  always_comb
    if ((\memWriteOut_CTmap''_map''_Int_Int_Int_d [0] && \dconPtr_CTmap''_map''_Int_Int_Int_d [0]))
      unique case (\memWriteOut_CTmap''_map''_Int_Int_Int_d [1:1])
        1'd0: \dconPtr_CTmap''_map''_Int_Int_Int_onehotd  = 2'd1;
        1'd1: \dconPtr_CTmap''_map''_Int_Int_Int_onehotd  = 2'd2;
        default: \dconPtr_CTmap''_map''_Int_Int_Int_onehotd  = 2'd0;
      endcase
    else \dconPtr_CTmap''_map''_Int_Int_Int_onehotd  = 2'd0;
  assign _36_d = {\dconPtr_CTmap''_map''_Int_Int_Int_d [16:1],
                  \dconPtr_CTmap''_map''_Int_Int_Int_onehotd [0]};
  assign \demuxWriteResult_CTmap''_map''_Int_Int_Int_d  = {\dconPtr_CTmap''_map''_Int_Int_Int_d [16:1],
                                                           \dconPtr_CTmap''_map''_Int_Int_Int_onehotd [1]};
  assign \dconPtr_CTmap''_map''_Int_Int_Int_r  = (| (\dconPtr_CTmap''_map''_Int_Int_Int_onehotd  & {\demuxWriteResult_CTmap''_map''_Int_Int_Int_r ,
                                                                                                    _36_r}));
  assign \memWriteOut_CTmap''_map''_Int_Int_Int_r  = \dconPtr_CTmap''_map''_Int_Int_Int_r ;
  
  /* const (Ty Word16#,
       Lit 0) : (goFor_8,Go) > (initHP_CTkron_kron_Int_Int_Int,Word16#) */
  assign initHP_CTkron_kron_Int_Int_Int_d = {16'd0, goFor_8_d[0]};
  assign goFor_8_r = initHP_CTkron_kron_Int_Int_Int_r;
  
  /* const (Ty Word16#,
       Lit 1) : (incrHP_CTkron_kron_Int_Int_Int1,Go) > (incrHP_CTkron_kron_Int_Int_Int,Word16#) */
  assign incrHP_CTkron_kron_Int_Int_Int_d = {16'd1,
                                             incrHP_CTkron_kron_Int_Int_Int1_d[0]};
  assign incrHP_CTkron_kron_Int_Int_Int1_r = incrHP_CTkron_kron_Int_Int_Int_r;
  
  /* merge (Ty Go) : [(goFor_9,Go),
                 (incrHP_CTkron_kron_Int_Int_Int2,Go)] > (incrHP_mergeCTkron_kron_Int_Int_Int,Go) */
  logic [1:0] incrHP_mergeCTkron_kron_Int_Int_Int_selected;
  logic [1:0] incrHP_mergeCTkron_kron_Int_Int_Int_select;
  always_comb
    begin
      incrHP_mergeCTkron_kron_Int_Int_Int_selected = 2'd0;
      if ((| incrHP_mergeCTkron_kron_Int_Int_Int_select))
        incrHP_mergeCTkron_kron_Int_Int_Int_selected = incrHP_mergeCTkron_kron_Int_Int_Int_select;
      else
        if (goFor_9_d[0])
          incrHP_mergeCTkron_kron_Int_Int_Int_selected[0] = 1'd1;
        else if (incrHP_CTkron_kron_Int_Int_Int2_d[0])
          incrHP_mergeCTkron_kron_Int_Int_Int_selected[1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      incrHP_mergeCTkron_kron_Int_Int_Int_select <= 2'd0;
    else
      incrHP_mergeCTkron_kron_Int_Int_Int_select <= (incrHP_mergeCTkron_kron_Int_Int_Int_r ? 2'd0 :
                                                     incrHP_mergeCTkron_kron_Int_Int_Int_selected);
  always_comb
    if (incrHP_mergeCTkron_kron_Int_Int_Int_selected[0])
      incrHP_mergeCTkron_kron_Int_Int_Int_d = goFor_9_d;
    else if (incrHP_mergeCTkron_kron_Int_Int_Int_selected[1])
      incrHP_mergeCTkron_kron_Int_Int_Int_d = incrHP_CTkron_kron_Int_Int_Int2_d;
    else incrHP_mergeCTkron_kron_Int_Int_Int_d = 1'd0;
  assign {incrHP_CTkron_kron_Int_Int_Int2_r,
          goFor_9_r} = (incrHP_mergeCTkron_kron_Int_Int_Int_r ? incrHP_mergeCTkron_kron_Int_Int_Int_selected :
                        2'd0);
  
  /* fork (Ty Go) : (incrHP_mergeCTkron_kron_Int_Int_Int_buf,Go) > [(incrHP_CTkron_kron_Int_Int_Int1,Go),
                                                               (incrHP_CTkron_kron_Int_Int_Int2,Go)] */
  logic [1:0] incrHP_mergeCTkron_kron_Int_Int_Int_buf_emitted;
  logic [1:0] incrHP_mergeCTkron_kron_Int_Int_Int_buf_done;
  assign incrHP_CTkron_kron_Int_Int_Int1_d = (incrHP_mergeCTkron_kron_Int_Int_Int_buf_d[0] && (! incrHP_mergeCTkron_kron_Int_Int_Int_buf_emitted[0]));
  assign incrHP_CTkron_kron_Int_Int_Int2_d = (incrHP_mergeCTkron_kron_Int_Int_Int_buf_d[0] && (! incrHP_mergeCTkron_kron_Int_Int_Int_buf_emitted[1]));
  assign incrHP_mergeCTkron_kron_Int_Int_Int_buf_done = (incrHP_mergeCTkron_kron_Int_Int_Int_buf_emitted | ({incrHP_CTkron_kron_Int_Int_Int2_d[0],
                                                                                                             incrHP_CTkron_kron_Int_Int_Int1_d[0]} & {incrHP_CTkron_kron_Int_Int_Int2_r,
                                                                                                                                                      incrHP_CTkron_kron_Int_Int_Int1_r}));
  assign incrHP_mergeCTkron_kron_Int_Int_Int_buf_r = (& incrHP_mergeCTkron_kron_Int_Int_Int_buf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      incrHP_mergeCTkron_kron_Int_Int_Int_buf_emitted <= 2'd0;
    else
      incrHP_mergeCTkron_kron_Int_Int_Int_buf_emitted <= (incrHP_mergeCTkron_kron_Int_Int_Int_buf_r ? 2'd0 :
                                                          incrHP_mergeCTkron_kron_Int_Int_Int_buf_done);
  
  /* op_add (Ty Word16#) : (incrHP_CTkron_kron_Int_Int_Int,Word16#) (forkHP1_CTkron_kron_Int_Int_Int,Word16#) > (addHP_CTkron_kron_Int_Int_Int,Word16#) */
  assign addHP_CTkron_kron_Int_Int_Int_d = {(incrHP_CTkron_kron_Int_Int_Int_d[16:1] + forkHP1_CTkron_kron_Int_Int_Int_d[16:1]),
                                            (incrHP_CTkron_kron_Int_Int_Int_d[0] && forkHP1_CTkron_kron_Int_Int_Int_d[0])};
  assign {incrHP_CTkron_kron_Int_Int_Int_r,
          forkHP1_CTkron_kron_Int_Int_Int_r} = {2 {(addHP_CTkron_kron_Int_Int_Int_r && addHP_CTkron_kron_Int_Int_Int_d[0])}};
  
  /* merge (Ty Word16#) : [(initHP_CTkron_kron_Int_Int_Int,Word16#),
                      (addHP_CTkron_kron_Int_Int_Int,Word16#)] > (mergeHP_CTkron_kron_Int_Int_Int,Word16#) */
  logic [1:0] mergeHP_CTkron_kron_Int_Int_Int_selected;
  logic [1:0] mergeHP_CTkron_kron_Int_Int_Int_select;
  always_comb
    begin
      mergeHP_CTkron_kron_Int_Int_Int_selected = 2'd0;
      if ((| mergeHP_CTkron_kron_Int_Int_Int_select))
        mergeHP_CTkron_kron_Int_Int_Int_selected = mergeHP_CTkron_kron_Int_Int_Int_select;
      else
        if (initHP_CTkron_kron_Int_Int_Int_d[0])
          mergeHP_CTkron_kron_Int_Int_Int_selected[0] = 1'd1;
        else if (addHP_CTkron_kron_Int_Int_Int_d[0])
          mergeHP_CTkron_kron_Int_Int_Int_selected[1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      mergeHP_CTkron_kron_Int_Int_Int_select <= 2'd0;
    else
      mergeHP_CTkron_kron_Int_Int_Int_select <= (mergeHP_CTkron_kron_Int_Int_Int_r ? 2'd0 :
                                                 mergeHP_CTkron_kron_Int_Int_Int_selected);
  always_comb
    if (mergeHP_CTkron_kron_Int_Int_Int_selected[0])
      mergeHP_CTkron_kron_Int_Int_Int_d = initHP_CTkron_kron_Int_Int_Int_d;
    else if (mergeHP_CTkron_kron_Int_Int_Int_selected[1])
      mergeHP_CTkron_kron_Int_Int_Int_d = addHP_CTkron_kron_Int_Int_Int_d;
    else mergeHP_CTkron_kron_Int_Int_Int_d = {16'd0, 1'd0};
  assign {addHP_CTkron_kron_Int_Int_Int_r,
          initHP_CTkron_kron_Int_Int_Int_r} = (mergeHP_CTkron_kron_Int_Int_Int_r ? mergeHP_CTkron_kron_Int_Int_Int_selected :
                                               2'd0);
  
  /* buf (Ty Go) : (incrHP_mergeCTkron_kron_Int_Int_Int,Go) > (incrHP_mergeCTkron_kron_Int_Int_Int_buf,Go) */
  Go_t incrHP_mergeCTkron_kron_Int_Int_Int_bufchan_d;
  logic incrHP_mergeCTkron_kron_Int_Int_Int_bufchan_r;
  assign incrHP_mergeCTkron_kron_Int_Int_Int_r = ((! incrHP_mergeCTkron_kron_Int_Int_Int_bufchan_d[0]) || incrHP_mergeCTkron_kron_Int_Int_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      incrHP_mergeCTkron_kron_Int_Int_Int_bufchan_d <= 1'd0;
    else
      if (incrHP_mergeCTkron_kron_Int_Int_Int_r)
        incrHP_mergeCTkron_kron_Int_Int_Int_bufchan_d <= incrHP_mergeCTkron_kron_Int_Int_Int_d;
  Go_t incrHP_mergeCTkron_kron_Int_Int_Int_bufchan_buf;
  assign incrHP_mergeCTkron_kron_Int_Int_Int_bufchan_r = (! incrHP_mergeCTkron_kron_Int_Int_Int_bufchan_buf[0]);
  assign incrHP_mergeCTkron_kron_Int_Int_Int_buf_d = (incrHP_mergeCTkron_kron_Int_Int_Int_bufchan_buf[0] ? incrHP_mergeCTkron_kron_Int_Int_Int_bufchan_buf :
                                                      incrHP_mergeCTkron_kron_Int_Int_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      incrHP_mergeCTkron_kron_Int_Int_Int_bufchan_buf <= 1'd0;
    else
      if ((incrHP_mergeCTkron_kron_Int_Int_Int_buf_r && incrHP_mergeCTkron_kron_Int_Int_Int_bufchan_buf[0]))
        incrHP_mergeCTkron_kron_Int_Int_Int_bufchan_buf <= 1'd0;
      else if (((! incrHP_mergeCTkron_kron_Int_Int_Int_buf_r) && (! incrHP_mergeCTkron_kron_Int_Int_Int_bufchan_buf[0])))
        incrHP_mergeCTkron_kron_Int_Int_Int_bufchan_buf <= incrHP_mergeCTkron_kron_Int_Int_Int_bufchan_d;
  
  /* buf (Ty Word16#) : (mergeHP_CTkron_kron_Int_Int_Int,Word16#) > (mergeHP_CTkron_kron_Int_Int_Int_buf,Word16#) */
  \Word16#_t  mergeHP_CTkron_kron_Int_Int_Int_bufchan_d;
  logic mergeHP_CTkron_kron_Int_Int_Int_bufchan_r;
  assign mergeHP_CTkron_kron_Int_Int_Int_r = ((! mergeHP_CTkron_kron_Int_Int_Int_bufchan_d[0]) || mergeHP_CTkron_kron_Int_Int_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      mergeHP_CTkron_kron_Int_Int_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (mergeHP_CTkron_kron_Int_Int_Int_r)
        mergeHP_CTkron_kron_Int_Int_Int_bufchan_d <= mergeHP_CTkron_kron_Int_Int_Int_d;
  \Word16#_t  mergeHP_CTkron_kron_Int_Int_Int_bufchan_buf;
  assign mergeHP_CTkron_kron_Int_Int_Int_bufchan_r = (! mergeHP_CTkron_kron_Int_Int_Int_bufchan_buf[0]);
  assign mergeHP_CTkron_kron_Int_Int_Int_buf_d = (mergeHP_CTkron_kron_Int_Int_Int_bufchan_buf[0] ? mergeHP_CTkron_kron_Int_Int_Int_bufchan_buf :
                                                  mergeHP_CTkron_kron_Int_Int_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      mergeHP_CTkron_kron_Int_Int_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((mergeHP_CTkron_kron_Int_Int_Int_buf_r && mergeHP_CTkron_kron_Int_Int_Int_bufchan_buf[0]))
        mergeHP_CTkron_kron_Int_Int_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! mergeHP_CTkron_kron_Int_Int_Int_buf_r) && (! mergeHP_CTkron_kron_Int_Int_Int_bufchan_buf[0])))
        mergeHP_CTkron_kron_Int_Int_Int_bufchan_buf <= mergeHP_CTkron_kron_Int_Int_Int_bufchan_d;
  
  /* fork (Ty Word16#) : (mergeHP_CTkron_kron_Int_Int_Int_buf,Word16#) > [(forkHP1_CTkron_kron_Int_Int_Int,Word16#),
                                                                     (forkHP1_CTkron_kron_Int_Int_In2,Word16#),
                                                                     (forkHP1_CTkron_kron_Int_Int_In3,Word16#)] */
  logic [2:0] mergeHP_CTkron_kron_Int_Int_Int_buf_emitted;
  logic [2:0] mergeHP_CTkron_kron_Int_Int_Int_buf_done;
  assign forkHP1_CTkron_kron_Int_Int_Int_d = {mergeHP_CTkron_kron_Int_Int_Int_buf_d[16:1],
                                              (mergeHP_CTkron_kron_Int_Int_Int_buf_d[0] && (! mergeHP_CTkron_kron_Int_Int_Int_buf_emitted[0]))};
  assign forkHP1_CTkron_kron_Int_Int_In2_d = {mergeHP_CTkron_kron_Int_Int_Int_buf_d[16:1],
                                              (mergeHP_CTkron_kron_Int_Int_Int_buf_d[0] && (! mergeHP_CTkron_kron_Int_Int_Int_buf_emitted[1]))};
  assign forkHP1_CTkron_kron_Int_Int_In3_d = {mergeHP_CTkron_kron_Int_Int_Int_buf_d[16:1],
                                              (mergeHP_CTkron_kron_Int_Int_Int_buf_d[0] && (! mergeHP_CTkron_kron_Int_Int_Int_buf_emitted[2]))};
  assign mergeHP_CTkron_kron_Int_Int_Int_buf_done = (mergeHP_CTkron_kron_Int_Int_Int_buf_emitted | ({forkHP1_CTkron_kron_Int_Int_In3_d[0],
                                                                                                     forkHP1_CTkron_kron_Int_Int_In2_d[0],
                                                                                                     forkHP1_CTkron_kron_Int_Int_Int_d[0]} & {forkHP1_CTkron_kron_Int_Int_In3_r,
                                                                                                                                              forkHP1_CTkron_kron_Int_Int_In2_r,
                                                                                                                                              forkHP1_CTkron_kron_Int_Int_Int_r}));
  assign mergeHP_CTkron_kron_Int_Int_Int_buf_r = (& mergeHP_CTkron_kron_Int_Int_Int_buf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      mergeHP_CTkron_kron_Int_Int_Int_buf_emitted <= 3'd0;
    else
      mergeHP_CTkron_kron_Int_Int_Int_buf_emitted <= (mergeHP_CTkron_kron_Int_Int_Int_buf_r ? 3'd0 :
                                                      mergeHP_CTkron_kron_Int_Int_Int_buf_done);
  
  /* mergectrl (Ty C2,
           Ty MemIn_CTkron_kron_Int_Int_Int) : [(dconReadIn_CTkron_kron_Int_Int_Int,MemIn_CTkron_kron_Int_Int_Int),
                                                (dconWriteIn_CTkron_kron_Int_Int_Int,MemIn_CTkron_kron_Int_Int_Int)] > (memMergeChoice_CTkron_kron_Int_Int_Int,C2) (memMergeIn_CTkron_kron_Int_Int_Int,MemIn_CTkron_kron_Int_Int_Int) */
  logic [1:0] dconReadIn_CTkron_kron_Int_Int_Int_select_d;
  assign dconReadIn_CTkron_kron_Int_Int_Int_select_d = ((| dconReadIn_CTkron_kron_Int_Int_Int_select_q) ? dconReadIn_CTkron_kron_Int_Int_Int_select_q :
                                                        (dconReadIn_CTkron_kron_Int_Int_Int_d[0] ? 2'd1 :
                                                         (dconWriteIn_CTkron_kron_Int_Int_Int_d[0] ? 2'd2 :
                                                          2'd0)));
  logic [1:0] dconReadIn_CTkron_kron_Int_Int_Int_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      dconReadIn_CTkron_kron_Int_Int_Int_select_q <= 2'd0;
    else
      dconReadIn_CTkron_kron_Int_Int_Int_select_q <= (dconReadIn_CTkron_kron_Int_Int_Int_done ? 2'd0 :
                                                      dconReadIn_CTkron_kron_Int_Int_Int_select_d);
  logic [1:0] dconReadIn_CTkron_kron_Int_Int_Int_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      dconReadIn_CTkron_kron_Int_Int_Int_emit_q <= 2'd0;
    else
      dconReadIn_CTkron_kron_Int_Int_Int_emit_q <= (dconReadIn_CTkron_kron_Int_Int_Int_done ? 2'd0 :
                                                    dconReadIn_CTkron_kron_Int_Int_Int_emit_d);
  logic [1:0] dconReadIn_CTkron_kron_Int_Int_Int_emit_d;
  assign dconReadIn_CTkron_kron_Int_Int_Int_emit_d = (dconReadIn_CTkron_kron_Int_Int_Int_emit_q | ({memMergeChoice_CTkron_kron_Int_Int_Int_d[0],
                                                                                                    memMergeIn_CTkron_kron_Int_Int_Int_d[0]} & {memMergeChoice_CTkron_kron_Int_Int_Int_r,
                                                                                                                                                memMergeIn_CTkron_kron_Int_Int_Int_r}));
  logic dconReadIn_CTkron_kron_Int_Int_Int_done;
  assign dconReadIn_CTkron_kron_Int_Int_Int_done = (& dconReadIn_CTkron_kron_Int_Int_Int_emit_d);
  assign {dconWriteIn_CTkron_kron_Int_Int_Int_r,
          dconReadIn_CTkron_kron_Int_Int_Int_r} = (dconReadIn_CTkron_kron_Int_Int_Int_done ? dconReadIn_CTkron_kron_Int_Int_Int_select_d :
                                                   2'd0);
  assign memMergeIn_CTkron_kron_Int_Int_Int_d = ((dconReadIn_CTkron_kron_Int_Int_Int_select_d[0] && (! dconReadIn_CTkron_kron_Int_Int_Int_emit_q[0])) ? dconReadIn_CTkron_kron_Int_Int_Int_d :
                                                 ((dconReadIn_CTkron_kron_Int_Int_Int_select_d[1] && (! dconReadIn_CTkron_kron_Int_Int_Int_emit_q[0])) ? dconWriteIn_CTkron_kron_Int_Int_Int_d :
                                                  {100'd0, 1'd0}));
  assign memMergeChoice_CTkron_kron_Int_Int_Int_d = ((dconReadIn_CTkron_kron_Int_Int_Int_select_d[0] && (! dconReadIn_CTkron_kron_Int_Int_Int_emit_q[1])) ? C1_2_dc(1'd1) :
                                                     ((dconReadIn_CTkron_kron_Int_Int_Int_select_d[1] && (! dconReadIn_CTkron_kron_Int_Int_Int_emit_q[1])) ? C2_2_dc(1'd1) :
                                                      {1'd0, 1'd0}));
  
  /* bram (Ty MemIn_CTkron_kron_Int_Int_Int,
      Ty MemOut_CTkron_kron_Int_Int_Int) : (memMergeIn_CTkron_kron_Int_Int_Int_dbuf,MemIn_CTkron_kron_Int_Int_Int) > (memOut_CTkron_kron_Int_Int_Int,MemOut_CTkron_kron_Int_Int_Int) */
  logic [82:0] memMergeIn_CTkron_kron_Int_Int_Int_dbuf_mem[65535:0];
  logic [15:0] memMergeIn_CTkron_kron_Int_Int_Int_dbuf_address;
  logic [82:0] memMergeIn_CTkron_kron_Int_Int_Int_dbuf_din;
  logic [82:0] memOut_CTkron_kron_Int_Int_Int_q;
  logic memOut_CTkron_kron_Int_Int_Int_valid;
  logic memMergeIn_CTkron_kron_Int_Int_Int_dbuf_we;
  logic memOut_CTkron_kron_Int_Int_Int_we;
  assign memMergeIn_CTkron_kron_Int_Int_Int_dbuf_din = memMergeIn_CTkron_kron_Int_Int_Int_dbuf_d[100:18];
  assign memMergeIn_CTkron_kron_Int_Int_Int_dbuf_address = memMergeIn_CTkron_kron_Int_Int_Int_dbuf_d[17:2];
  assign memMergeIn_CTkron_kron_Int_Int_Int_dbuf_we = (memMergeIn_CTkron_kron_Int_Int_Int_dbuf_d[1:1] && memMergeIn_CTkron_kron_Int_Int_Int_dbuf_d[0]);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        memOut_CTkron_kron_Int_Int_Int_we <= 1'd0;
        memOut_CTkron_kron_Int_Int_Int_valid <= 1'd0;
      end
    else
      begin
        memOut_CTkron_kron_Int_Int_Int_we <= memMergeIn_CTkron_kron_Int_Int_Int_dbuf_we;
        memOut_CTkron_kron_Int_Int_Int_valid <= memMergeIn_CTkron_kron_Int_Int_Int_dbuf_d[0];
        if (memMergeIn_CTkron_kron_Int_Int_Int_dbuf_we)
          begin
            memMergeIn_CTkron_kron_Int_Int_Int_dbuf_mem[memMergeIn_CTkron_kron_Int_Int_Int_dbuf_address] <= memMergeIn_CTkron_kron_Int_Int_Int_dbuf_din;
            memOut_CTkron_kron_Int_Int_Int_q <= memMergeIn_CTkron_kron_Int_Int_Int_dbuf_din;
          end
        else
          memOut_CTkron_kron_Int_Int_Int_q <= memMergeIn_CTkron_kron_Int_Int_Int_dbuf_mem[memMergeIn_CTkron_kron_Int_Int_Int_dbuf_address];
      end
  assign memOut_CTkron_kron_Int_Int_Int_d = {memOut_CTkron_kron_Int_Int_Int_q,
                                             memOut_CTkron_kron_Int_Int_Int_we,
                                             memOut_CTkron_kron_Int_Int_Int_valid};
  assign memMergeIn_CTkron_kron_Int_Int_Int_dbuf_r = ((! memOut_CTkron_kron_Int_Int_Int_valid) || memOut_CTkron_kron_Int_Int_Int_r);
  
  /* demux (Ty C2,
       Ty MemOut_CTkron_kron_Int_Int_Int) : (memMergeChoice_CTkron_kron_Int_Int_Int,C2) (memOut_CTkron_kron_Int_Int_Int_dbuf,MemOut_CTkron_kron_Int_Int_Int) > [(memReadOut_CTkron_kron_Int_Int_Int,MemOut_CTkron_kron_Int_Int_Int),
                                                                                                                                                                (memWriteOut_CTkron_kron_Int_Int_Int,MemOut_CTkron_kron_Int_Int_Int)] */
  logic [1:0] memOut_CTkron_kron_Int_Int_Int_dbuf_onehotd;
  always_comb
    if ((memMergeChoice_CTkron_kron_Int_Int_Int_d[0] && memOut_CTkron_kron_Int_Int_Int_dbuf_d[0]))
      unique case (memMergeChoice_CTkron_kron_Int_Int_Int_d[1:1])
        1'd0: memOut_CTkron_kron_Int_Int_Int_dbuf_onehotd = 2'd1;
        1'd1: memOut_CTkron_kron_Int_Int_Int_dbuf_onehotd = 2'd2;
        default: memOut_CTkron_kron_Int_Int_Int_dbuf_onehotd = 2'd0;
      endcase
    else memOut_CTkron_kron_Int_Int_Int_dbuf_onehotd = 2'd0;
  assign memReadOut_CTkron_kron_Int_Int_Int_d = {memOut_CTkron_kron_Int_Int_Int_dbuf_d[84:1],
                                                 memOut_CTkron_kron_Int_Int_Int_dbuf_onehotd[0]};
  assign memWriteOut_CTkron_kron_Int_Int_Int_d = {memOut_CTkron_kron_Int_Int_Int_dbuf_d[84:1],
                                                  memOut_CTkron_kron_Int_Int_Int_dbuf_onehotd[1]};
  assign memOut_CTkron_kron_Int_Int_Int_dbuf_r = (| (memOut_CTkron_kron_Int_Int_Int_dbuf_onehotd & {memWriteOut_CTkron_kron_Int_Int_Int_r,
                                                                                                    memReadOut_CTkron_kron_Int_Int_Int_r}));
  assign memMergeChoice_CTkron_kron_Int_Int_Int_r = memOut_CTkron_kron_Int_Int_Int_dbuf_r;
  
  /* dbuf (Ty MemIn_CTkron_kron_Int_Int_Int) : (memMergeIn_CTkron_kron_Int_Int_Int_rbuf,MemIn_CTkron_kron_Int_Int_Int) > (memMergeIn_CTkron_kron_Int_Int_Int_dbuf,MemIn_CTkron_kron_Int_Int_Int) */
  assign memMergeIn_CTkron_kron_Int_Int_Int_rbuf_r = ((! memMergeIn_CTkron_kron_Int_Int_Int_dbuf_d[0]) || memMergeIn_CTkron_kron_Int_Int_Int_dbuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      memMergeIn_CTkron_kron_Int_Int_Int_dbuf_d <= {100'd0, 1'd0};
    else
      if (memMergeIn_CTkron_kron_Int_Int_Int_rbuf_r)
        memMergeIn_CTkron_kron_Int_Int_Int_dbuf_d <= memMergeIn_CTkron_kron_Int_Int_Int_rbuf_d;
  
  /* rbuf (Ty MemIn_CTkron_kron_Int_Int_Int) : (memMergeIn_CTkron_kron_Int_Int_Int,MemIn_CTkron_kron_Int_Int_Int) > (memMergeIn_CTkron_kron_Int_Int_Int_rbuf,MemIn_CTkron_kron_Int_Int_Int) */
  MemIn_CTkron_kron_Int_Int_Int_t memMergeIn_CTkron_kron_Int_Int_Int_buf;
  assign memMergeIn_CTkron_kron_Int_Int_Int_r = (! memMergeIn_CTkron_kron_Int_Int_Int_buf[0]);
  assign memMergeIn_CTkron_kron_Int_Int_Int_rbuf_d = (memMergeIn_CTkron_kron_Int_Int_Int_buf[0] ? memMergeIn_CTkron_kron_Int_Int_Int_buf :
                                                      memMergeIn_CTkron_kron_Int_Int_Int_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      memMergeIn_CTkron_kron_Int_Int_Int_buf <= {100'd0, 1'd0};
    else
      if ((memMergeIn_CTkron_kron_Int_Int_Int_rbuf_r && memMergeIn_CTkron_kron_Int_Int_Int_buf[0]))
        memMergeIn_CTkron_kron_Int_Int_Int_buf <= {100'd0, 1'd0};
      else if (((! memMergeIn_CTkron_kron_Int_Int_Int_rbuf_r) && (! memMergeIn_CTkron_kron_Int_Int_Int_buf[0])))
        memMergeIn_CTkron_kron_Int_Int_Int_buf <= memMergeIn_CTkron_kron_Int_Int_Int_d;
  
  /* dbuf (Ty MemOut_CTkron_kron_Int_Int_Int) : (memOut_CTkron_kron_Int_Int_Int_rbuf,MemOut_CTkron_kron_Int_Int_Int) > (memOut_CTkron_kron_Int_Int_Int_dbuf,MemOut_CTkron_kron_Int_Int_Int) */
  assign memOut_CTkron_kron_Int_Int_Int_rbuf_r = ((! memOut_CTkron_kron_Int_Int_Int_dbuf_d[0]) || memOut_CTkron_kron_Int_Int_Int_dbuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      memOut_CTkron_kron_Int_Int_Int_dbuf_d <= {84'd0, 1'd0};
    else
      if (memOut_CTkron_kron_Int_Int_Int_rbuf_r)
        memOut_CTkron_kron_Int_Int_Int_dbuf_d <= memOut_CTkron_kron_Int_Int_Int_rbuf_d;
  
  /* rbuf (Ty MemOut_CTkron_kron_Int_Int_Int) : (memOut_CTkron_kron_Int_Int_Int,MemOut_CTkron_kron_Int_Int_Int) > (memOut_CTkron_kron_Int_Int_Int_rbuf,MemOut_CTkron_kron_Int_Int_Int) */
  MemOut_CTkron_kron_Int_Int_Int_t memOut_CTkron_kron_Int_Int_Int_buf;
  assign memOut_CTkron_kron_Int_Int_Int_r = (! memOut_CTkron_kron_Int_Int_Int_buf[0]);
  assign memOut_CTkron_kron_Int_Int_Int_rbuf_d = (memOut_CTkron_kron_Int_Int_Int_buf[0] ? memOut_CTkron_kron_Int_Int_Int_buf :
                                                  memOut_CTkron_kron_Int_Int_Int_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      memOut_CTkron_kron_Int_Int_Int_buf <= {84'd0, 1'd0};
    else
      if ((memOut_CTkron_kron_Int_Int_Int_rbuf_r && memOut_CTkron_kron_Int_Int_Int_buf[0]))
        memOut_CTkron_kron_Int_Int_Int_buf <= {84'd0, 1'd0};
      else if (((! memOut_CTkron_kron_Int_Int_Int_rbuf_r) && (! memOut_CTkron_kron_Int_Int_Int_buf[0])))
        memOut_CTkron_kron_Int_Int_Int_buf <= memOut_CTkron_kron_Int_Int_Int_d;
  
  /* destruct (Ty Pointer_CTkron_kron_Int_Int_Int,
          Dcon Pointer_CTkron_kron_Int_Int_Int) : (scfarg_0_1_1_argbuf,Pointer_CTkron_kron_Int_Int_Int) > [(destructReadIn_CTkron_kron_Int_Int_Int,Word16#)] */
  assign destructReadIn_CTkron_kron_Int_Int_Int_d = {scfarg_0_1_1_argbuf_d[16:1],
                                                     scfarg_0_1_1_argbuf_d[0]};
  assign scfarg_0_1_1_argbuf_r = destructReadIn_CTkron_kron_Int_Int_Int_r;
  
  /* dcon (Ty MemIn_CTkron_kron_Int_Int_Int,
      Dcon ReadIn_CTkron_kron_Int_Int_Int) : [(destructReadIn_CTkron_kron_Int_Int_Int,Word16#)] > (dconReadIn_CTkron_kron_Int_Int_Int,MemIn_CTkron_kron_Int_Int_Int) */
  assign dconReadIn_CTkron_kron_Int_Int_Int_d = ReadIn_CTkron_kron_Int_Int_Int_dc((& {destructReadIn_CTkron_kron_Int_Int_Int_d[0]}), destructReadIn_CTkron_kron_Int_Int_Int_d);
  assign {destructReadIn_CTkron_kron_Int_Int_Int_r} = {1 {(dconReadIn_CTkron_kron_Int_Int_Int_r && dconReadIn_CTkron_kron_Int_Int_Int_d[0])}};
  
  /* destruct (Ty MemOut_CTkron_kron_Int_Int_Int,
          Dcon ReadOut_CTkron_kron_Int_Int_Int) : (memReadOut_CTkron_kron_Int_Int_Int,MemOut_CTkron_kron_Int_Int_Int) > [(readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf,CTkron_kron_Int_Int_Int)] */
  assign readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf_d = {memReadOut_CTkron_kron_Int_Int_Int_d[84:2],
                                                                     memReadOut_CTkron_kron_Int_Int_Int_d[0]};
  assign memReadOut_CTkron_kron_Int_Int_Int_r = readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf_r;
  
  /* mergectrl (Ty C5,
           Ty CTkron_kron_Int_Int_Int) : [(lizzieLet22_1_argbuf,CTkron_kron_Int_Int_Int),
                                          (lizzieLet30_1_argbuf,CTkron_kron_Int_Int_Int),
                                          (lizzieLet31_1_argbuf,CTkron_kron_Int_Int_Int),
                                          (lizzieLet32_1_argbuf,CTkron_kron_Int_Int_Int),
                                          (lizzieLet8_1_argbuf,CTkron_kron_Int_Int_Int)] > (writeMerge_choice_CTkron_kron_Int_Int_Int,C5) (writeMerge_data_CTkron_kron_Int_Int_Int,CTkron_kron_Int_Int_Int) */
  logic [4:0] lizzieLet22_1_argbuf_select_d;
  assign lizzieLet22_1_argbuf_select_d = ((| lizzieLet22_1_argbuf_select_q) ? lizzieLet22_1_argbuf_select_q :
                                          (lizzieLet22_1_argbuf_d[0] ? 5'd1 :
                                           (lizzieLet30_1_argbuf_d[0] ? 5'd2 :
                                            (lizzieLet31_1_argbuf_d[0] ? 5'd4 :
                                             (lizzieLet32_1_argbuf_d[0] ? 5'd8 :
                                              (lizzieLet8_1_argbuf_d[0] ? 5'd16 :
                                               5'd0))))));
  logic [4:0] lizzieLet22_1_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet22_1_argbuf_select_q <= 5'd0;
    else
      lizzieLet22_1_argbuf_select_q <= (lizzieLet22_1_argbuf_done ? 5'd0 :
                                        lizzieLet22_1_argbuf_select_d);
  logic [1:0] lizzieLet22_1_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet22_1_argbuf_emit_q <= 2'd0;
    else
      lizzieLet22_1_argbuf_emit_q <= (lizzieLet22_1_argbuf_done ? 2'd0 :
                                      lizzieLet22_1_argbuf_emit_d);
  logic [1:0] lizzieLet22_1_argbuf_emit_d;
  assign lizzieLet22_1_argbuf_emit_d = (lizzieLet22_1_argbuf_emit_q | ({writeMerge_choice_CTkron_kron_Int_Int_Int_d[0],
                                                                        writeMerge_data_CTkron_kron_Int_Int_Int_d[0]} & {writeMerge_choice_CTkron_kron_Int_Int_Int_r,
                                                                                                                         writeMerge_data_CTkron_kron_Int_Int_Int_r}));
  logic lizzieLet22_1_argbuf_done;
  assign lizzieLet22_1_argbuf_done = (& lizzieLet22_1_argbuf_emit_d);
  assign {lizzieLet8_1_argbuf_r,
          lizzieLet32_1_argbuf_r,
          lizzieLet31_1_argbuf_r,
          lizzieLet30_1_argbuf_r,
          lizzieLet22_1_argbuf_r} = (lizzieLet22_1_argbuf_done ? lizzieLet22_1_argbuf_select_d :
                                     5'd0);
  assign writeMerge_data_CTkron_kron_Int_Int_Int_d = ((lizzieLet22_1_argbuf_select_d[0] && (! lizzieLet22_1_argbuf_emit_q[0])) ? lizzieLet22_1_argbuf_d :
                                                      ((lizzieLet22_1_argbuf_select_d[1] && (! lizzieLet22_1_argbuf_emit_q[0])) ? lizzieLet30_1_argbuf_d :
                                                       ((lizzieLet22_1_argbuf_select_d[2] && (! lizzieLet22_1_argbuf_emit_q[0])) ? lizzieLet31_1_argbuf_d :
                                                        ((lizzieLet22_1_argbuf_select_d[3] && (! lizzieLet22_1_argbuf_emit_q[0])) ? lizzieLet32_1_argbuf_d :
                                                         ((lizzieLet22_1_argbuf_select_d[4] && (! lizzieLet22_1_argbuf_emit_q[0])) ? lizzieLet8_1_argbuf_d :
                                                          {83'd0, 1'd0})))));
  assign writeMerge_choice_CTkron_kron_Int_Int_Int_d = ((lizzieLet22_1_argbuf_select_d[0] && (! lizzieLet22_1_argbuf_emit_q[1])) ? C1_5_dc(1'd1) :
                                                        ((lizzieLet22_1_argbuf_select_d[1] && (! lizzieLet22_1_argbuf_emit_q[1])) ? C2_5_dc(1'd1) :
                                                         ((lizzieLet22_1_argbuf_select_d[2] && (! lizzieLet22_1_argbuf_emit_q[1])) ? C3_5_dc(1'd1) :
                                                          ((lizzieLet22_1_argbuf_select_d[3] && (! lizzieLet22_1_argbuf_emit_q[1])) ? C4_5_dc(1'd1) :
                                                           ((lizzieLet22_1_argbuf_select_d[4] && (! lizzieLet22_1_argbuf_emit_q[1])) ? C5_5_dc(1'd1) :
                                                            {3'd0, 1'd0})))));
  
  /* demux (Ty C5,
       Ty Pointer_CTkron_kron_Int_Int_Int) : (writeMerge_choice_CTkron_kron_Int_Int_Int,C5) (demuxWriteResult_CTkron_kron_Int_Int_Int,Pointer_CTkron_kron_Int_Int_Int) > [(writeCTkron_kron_Int_Int_IntlizzieLet22_1_argbuf,Pointer_CTkron_kron_Int_Int_Int),
                                                                                                                                                                          (writeCTkron_kron_Int_Int_IntlizzieLet30_1_argbuf,Pointer_CTkron_kron_Int_Int_Int),
                                                                                                                                                                          (writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf,Pointer_CTkron_kron_Int_Int_Int),
                                                                                                                                                                          (writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf,Pointer_CTkron_kron_Int_Int_Int),
                                                                                                                                                                          (writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf,Pointer_CTkron_kron_Int_Int_Int)] */
  logic [4:0] demuxWriteResult_CTkron_kron_Int_Int_Int_onehotd;
  always_comb
    if ((writeMerge_choice_CTkron_kron_Int_Int_Int_d[0] && demuxWriteResult_CTkron_kron_Int_Int_Int_d[0]))
      unique case (writeMerge_choice_CTkron_kron_Int_Int_Int_d[3:1])
        3'd0: demuxWriteResult_CTkron_kron_Int_Int_Int_onehotd = 5'd1;
        3'd1: demuxWriteResult_CTkron_kron_Int_Int_Int_onehotd = 5'd2;
        3'd2: demuxWriteResult_CTkron_kron_Int_Int_Int_onehotd = 5'd4;
        3'd3: demuxWriteResult_CTkron_kron_Int_Int_Int_onehotd = 5'd8;
        3'd4: demuxWriteResult_CTkron_kron_Int_Int_Int_onehotd = 5'd16;
        default: demuxWriteResult_CTkron_kron_Int_Int_Int_onehotd = 5'd0;
      endcase
    else demuxWriteResult_CTkron_kron_Int_Int_Int_onehotd = 5'd0;
  assign writeCTkron_kron_Int_Int_IntlizzieLet22_1_argbuf_d = {demuxWriteResult_CTkron_kron_Int_Int_Int_d[16:1],
                                                               demuxWriteResult_CTkron_kron_Int_Int_Int_onehotd[0]};
  assign writeCTkron_kron_Int_Int_IntlizzieLet30_1_argbuf_d = {demuxWriteResult_CTkron_kron_Int_Int_Int_d[16:1],
                                                               demuxWriteResult_CTkron_kron_Int_Int_Int_onehotd[1]};
  assign writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf_d = {demuxWriteResult_CTkron_kron_Int_Int_Int_d[16:1],
                                                               demuxWriteResult_CTkron_kron_Int_Int_Int_onehotd[2]};
  assign writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf_d = {demuxWriteResult_CTkron_kron_Int_Int_Int_d[16:1],
                                                               demuxWriteResult_CTkron_kron_Int_Int_Int_onehotd[3]};
  assign writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf_d = {demuxWriteResult_CTkron_kron_Int_Int_Int_d[16:1],
                                                              demuxWriteResult_CTkron_kron_Int_Int_Int_onehotd[4]};
  assign demuxWriteResult_CTkron_kron_Int_Int_Int_r = (| (demuxWriteResult_CTkron_kron_Int_Int_Int_onehotd & {writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf_r,
                                                                                                              writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf_r,
                                                                                                              writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf_r,
                                                                                                              writeCTkron_kron_Int_Int_IntlizzieLet30_1_argbuf_r,
                                                                                                              writeCTkron_kron_Int_Int_IntlizzieLet22_1_argbuf_r}));
  assign writeMerge_choice_CTkron_kron_Int_Int_Int_r = demuxWriteResult_CTkron_kron_Int_Int_Int_r;
  
  /* dcon (Ty MemIn_CTkron_kron_Int_Int_Int,
      Dcon WriteIn_CTkron_kron_Int_Int_Int) : [(forkHP1_CTkron_kron_Int_Int_In2,Word16#),
                                               (writeMerge_data_CTkron_kron_Int_Int_Int,CTkron_kron_Int_Int_Int)] > (dconWriteIn_CTkron_kron_Int_Int_Int,MemIn_CTkron_kron_Int_Int_Int) */
  assign dconWriteIn_CTkron_kron_Int_Int_Int_d = WriteIn_CTkron_kron_Int_Int_Int_dc((& {forkHP1_CTkron_kron_Int_Int_In2_d[0],
                                                                                        writeMerge_data_CTkron_kron_Int_Int_Int_d[0]}), forkHP1_CTkron_kron_Int_Int_In2_d, writeMerge_data_CTkron_kron_Int_Int_Int_d);
  assign {forkHP1_CTkron_kron_Int_Int_In2_r,
          writeMerge_data_CTkron_kron_Int_Int_Int_r} = {2 {(dconWriteIn_CTkron_kron_Int_Int_Int_r && dconWriteIn_CTkron_kron_Int_Int_Int_d[0])}};
  
  /* dcon (Ty Pointer_CTkron_kron_Int_Int_Int,
      Dcon Pointer_CTkron_kron_Int_Int_Int) : [(forkHP1_CTkron_kron_Int_Int_In3,Word16#)] > (dconPtr_CTkron_kron_Int_Int_Int,Pointer_CTkron_kron_Int_Int_Int) */
  assign dconPtr_CTkron_kron_Int_Int_Int_d = Pointer_CTkron_kron_Int_Int_Int_dc((& {forkHP1_CTkron_kron_Int_Int_In3_d[0]}), forkHP1_CTkron_kron_Int_Int_In3_d);
  assign {forkHP1_CTkron_kron_Int_Int_In3_r} = {1 {(dconPtr_CTkron_kron_Int_Int_Int_r && dconPtr_CTkron_kron_Int_Int_Int_d[0])}};
  
  /* demux (Ty MemOut_CTkron_kron_Int_Int_Int,
       Ty Pointer_CTkron_kron_Int_Int_Int) : (memWriteOut_CTkron_kron_Int_Int_Int,MemOut_CTkron_kron_Int_Int_Int) (dconPtr_CTkron_kron_Int_Int_Int,Pointer_CTkron_kron_Int_Int_Int) > [(_35,Pointer_CTkron_kron_Int_Int_Int),
                                                                                                                                                                                       (demuxWriteResult_CTkron_kron_Int_Int_Int,Pointer_CTkron_kron_Int_Int_Int)] */
  logic [1:0] dconPtr_CTkron_kron_Int_Int_Int_onehotd;
  always_comb
    if ((memWriteOut_CTkron_kron_Int_Int_Int_d[0] && dconPtr_CTkron_kron_Int_Int_Int_d[0]))
      unique case (memWriteOut_CTkron_kron_Int_Int_Int_d[1:1])
        1'd0: dconPtr_CTkron_kron_Int_Int_Int_onehotd = 2'd1;
        1'd1: dconPtr_CTkron_kron_Int_Int_Int_onehotd = 2'd2;
        default: dconPtr_CTkron_kron_Int_Int_Int_onehotd = 2'd0;
      endcase
    else dconPtr_CTkron_kron_Int_Int_Int_onehotd = 2'd0;
  assign _35_d = {dconPtr_CTkron_kron_Int_Int_Int_d[16:1],
                  dconPtr_CTkron_kron_Int_Int_Int_onehotd[0]};
  assign demuxWriteResult_CTkron_kron_Int_Int_Int_d = {dconPtr_CTkron_kron_Int_Int_Int_d[16:1],
                                                       dconPtr_CTkron_kron_Int_Int_Int_onehotd[1]};
  assign dconPtr_CTkron_kron_Int_Int_Int_r = (| (dconPtr_CTkron_kron_Int_Int_Int_onehotd & {demuxWriteResult_CTkron_kron_Int_Int_Int_r,
                                                                                            _35_r}));
  assign memWriteOut_CTkron_kron_Int_Int_Int_r = dconPtr_CTkron_kron_Int_Int_Int_r;
  
  /* buf (Ty Go) : (goFork,Go) > (go_1_argbuf,Go) */
  Go_t goFork_bufchan_d;
  logic goFork_bufchan_r;
  assign goFork_r = ((! goFork_bufchan_d[0]) || goFork_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) goFork_bufchan_d <= 1'd0;
    else if (goFork_r) goFork_bufchan_d <= goFork_d;
  Go_t goFork_bufchan_buf;
  assign goFork_bufchan_r = (! goFork_bufchan_buf[0]);
  assign go_1_argbuf_d = (goFork_bufchan_buf[0] ? goFork_bufchan_buf :
                          goFork_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) goFork_bufchan_buf <= 1'd0;
    else
      if ((go_1_argbuf_r && goFork_bufchan_buf[0]))
        goFork_bufchan_buf <= 1'd0;
      else if (((! go_1_argbuf_r) && (! goFork_bufchan_buf[0])))
        goFork_bufchan_buf <= goFork_bufchan_d;
  
  /* source (Ty Go) : > (sourceGo,Go) */
  
  /* source (Ty Pointer_QTree_Int) : > (w1svB_1_1,Pointer_QTree_Int) */
  
  /* source (Ty Pointer_QTree_Int) : > (wsvA_1_0,Pointer_QTree_Int) */
  
  /* destruct (Ty TupGo___Pointer_QTree_Int___Pointer_QTree_Int,
          Dcon TupGo___Pointer_QTree_Int___Pointer_QTree_Int) : ($wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Int_1,TupGo___Pointer_QTree_Int___Pointer_QTree_Int) > [($wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intgo_7,Go),
                                                                                                                                                                         ($wmainTupGo___Pointer_QTree_Int___Pointer_QTree_IntwsvA,Pointer_QTree_Int),
                                                                                                                                                                         ($wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intw1svB,Pointer_QTree_Int)] */
  logic [2:0] \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Int_1_emitted ;
  logic [2:0] \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Int_1_done ;
  assign \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intgo_7_d  = (\$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Int_1_d [0] && (! \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Int_1_emitted [0]));
  assign \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_IntwsvA_d  = {\$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Int_1_d [16:1],
                                                                        (\$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Int_1_d [0] && (! \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Int_1_emitted [1]))};
  assign \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intw1svB_d  = {\$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Int_1_d [32:17],
                                                                         (\$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Int_1_d [0] && (! \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Int_1_emitted [2]))};
  assign \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Int_1_done  = (\$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Int_1_emitted  | ({\$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intw1svB_d [0],
                                                                                                                                             \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_IntwsvA_d [0],
                                                                                                                                             \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intgo_7_d [0]} & {\$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intw1svB_r ,
                                                                                                                                                                                                                \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_IntwsvA_r ,
                                                                                                                                                                                                                \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intgo_7_r }));
  assign \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Int_1_r  = (& \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Int_1_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Int_1_emitted  <= 3'd0;
    else
      \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Int_1_emitted  <= (\$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Int_1_r  ? 3'd0 :
                                                                          \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Int_1_done );
  
  /* fork (Ty Go) : ($wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intgo_7,Go) > [(go_7_1,Go),
                                                                               (go_7_2,Go),
                                                                               (go_7_3,Go),
                                                                               (go_7_4,Go),
                                                                               (go_7_5,Go),
                                                                               (go_7_6,Go),
                                                                               (go_7_7,Go)] */
  logic [6:0] \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intgo_7_emitted ;
  logic [6:0] \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intgo_7_done ;
  assign go_7_1_d = (\$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intgo_7_d [0] && (! \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intgo_7_emitted [0]));
  assign go_7_2_d = (\$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intgo_7_d [0] && (! \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intgo_7_emitted [1]));
  assign go_7_3_d = (\$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intgo_7_d [0] && (! \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intgo_7_emitted [2]));
  assign go_7_4_d = (\$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intgo_7_d [0] && (! \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intgo_7_emitted [3]));
  assign go_7_5_d = (\$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intgo_7_d [0] && (! \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intgo_7_emitted [4]));
  assign go_7_6_d = (\$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intgo_7_d [0] && (! \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intgo_7_emitted [5]));
  assign go_7_7_d = (\$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intgo_7_d [0] && (! \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intgo_7_emitted [6]));
  assign \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intgo_7_done  = (\$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intgo_7_emitted  | ({go_7_7_d[0],
                                                                                                                                                 go_7_6_d[0],
                                                                                                                                                 go_7_5_d[0],
                                                                                                                                                 go_7_4_d[0],
                                                                                                                                                 go_7_3_d[0],
                                                                                                                                                 go_7_2_d[0],
                                                                                                                                                 go_7_1_d[0]} & {go_7_7_r,
                                                                                                                                                                 go_7_6_r,
                                                                                                                                                                 go_7_5_r,
                                                                                                                                                                 go_7_4_r,
                                                                                                                                                                 go_7_3_r,
                                                                                                                                                                 go_7_2_r,
                                                                                                                                                                 go_7_1_r}));
  assign \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intgo_7_r  = (& \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intgo_7_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intgo_7_emitted  <= 7'd0;
    else
      \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intgo_7_emitted  <= (\$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intgo_7_r  ? 7'd0 :
                                                                            \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intgo_7_done );
  
  /* buf (Ty Pointer_QTree_Int) : ($wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intw1svB,Pointer_QTree_Int) > (w1svB_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intw1svB_bufchan_d ;
  logic \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intw1svB_bufchan_r ;
  assign \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intw1svB_r  = ((! \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intw1svB_bufchan_d [0]) || \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intw1svB_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intw1svB_bufchan_d  <= {16'd0,
                                                                               1'd0};
    else
      if (\$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intw1svB_r )
        \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intw1svB_bufchan_d  <= \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intw1svB_d ;
  Pointer_QTree_Int_t \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intw1svB_bufchan_buf ;
  assign \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intw1svB_bufchan_r  = (! \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intw1svB_bufchan_buf [0]);
  assign w1svB_1_argbuf_d = (\$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intw1svB_bufchan_buf [0] ? \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intw1svB_bufchan_buf  :
                             \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intw1svB_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intw1svB_bufchan_buf  <= {16'd0,
                                                                                 1'd0};
    else
      if ((w1svB_1_argbuf_r && \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intw1svB_bufchan_buf [0]))
        \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intw1svB_bufchan_buf  <= {16'd0,
                                                                                   1'd0};
      else if (((! w1svB_1_argbuf_r) && (! \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intw1svB_bufchan_buf [0])))
        \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intw1svB_bufchan_buf  <= \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intw1svB_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Int) : ($wmainTupGo___Pointer_QTree_Int___Pointer_QTree_IntwsvA,Pointer_QTree_Int) > (wsvA_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_IntwsvA_bufchan_d ;
  logic \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_IntwsvA_bufchan_r ;
  assign \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_IntwsvA_r  = ((! \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_IntwsvA_bufchan_d [0]) || \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_IntwsvA_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_IntwsvA_bufchan_d  <= {16'd0,
                                                                              1'd0};
    else
      if (\$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_IntwsvA_r )
        \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_IntwsvA_bufchan_d  <= \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_IntwsvA_d ;
  Pointer_QTree_Int_t \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_IntwsvA_bufchan_buf ;
  assign \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_IntwsvA_bufchan_r  = (! \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_IntwsvA_bufchan_buf [0]);
  assign wsvA_1_argbuf_d = (\$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_IntwsvA_bufchan_buf [0] ? \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_IntwsvA_bufchan_buf  :
                            \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_IntwsvA_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_IntwsvA_bufchan_buf  <= {16'd0,
                                                                                1'd0};
    else
      if ((wsvA_1_argbuf_r && \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_IntwsvA_bufchan_buf [0]))
        \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_IntwsvA_bufchan_buf  <= {16'd0,
                                                                                  1'd0};
      else if (((! wsvA_1_argbuf_r) && (! \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_IntwsvA_bufchan_buf [0])))
        \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_IntwsvA_bufchan_buf  <= \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_IntwsvA_bufchan_d ;
  
  /* dcon (Ty Int,Dcon I#) : [($wmain_resbuf,Int#)] > (es_0_1I#,Int) */
  assign \es_0_1I#_d  = \I#_dc ((& {\$wmain_resbuf_d [0]}), \$wmain_resbuf_d );
  assign {\$wmain_resbuf_r } = {1 {(\es_0_1I#_r  && \es_0_1I#_d [0])}};
  
  /* destruct (Ty TupGo___Pointer_QTree_Int,
          Dcon TupGo___Pointer_QTree_Int) : ($wnnz_IntTupGo___Pointer_QTree_Int_1,TupGo___Pointer_QTree_Int) > [($wnnz_IntTupGo___Pointer_QTree_Intgo_8,Go),
                                                                                                                ($wnnz_IntTupGo___Pointer_QTree_Intwsvt,Pointer_QTree_Int)] */
  logic [1:0] \$wnnz_IntTupGo___Pointer_QTree_Int_1_emitted ;
  logic [1:0] \$wnnz_IntTupGo___Pointer_QTree_Int_1_done ;
  assign \$wnnz_IntTupGo___Pointer_QTree_Intgo_8_d  = (\$wnnz_IntTupGo___Pointer_QTree_Int_1_d [0] && (! \$wnnz_IntTupGo___Pointer_QTree_Int_1_emitted [0]));
  assign \$wnnz_IntTupGo___Pointer_QTree_Intwsvt_d  = {\$wnnz_IntTupGo___Pointer_QTree_Int_1_d [16:1],
                                                       (\$wnnz_IntTupGo___Pointer_QTree_Int_1_d [0] && (! \$wnnz_IntTupGo___Pointer_QTree_Int_1_emitted [1]))};
  assign \$wnnz_IntTupGo___Pointer_QTree_Int_1_done  = (\$wnnz_IntTupGo___Pointer_QTree_Int_1_emitted  | ({\$wnnz_IntTupGo___Pointer_QTree_Intwsvt_d [0],
                                                                                                           \$wnnz_IntTupGo___Pointer_QTree_Intgo_8_d [0]} & {\$wnnz_IntTupGo___Pointer_QTree_Intwsvt_r ,
                                                                                                                                                             \$wnnz_IntTupGo___Pointer_QTree_Intgo_8_r }));
  assign \$wnnz_IntTupGo___Pointer_QTree_Int_1_r  = (& \$wnnz_IntTupGo___Pointer_QTree_Int_1_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \$wnnz_IntTupGo___Pointer_QTree_Int_1_emitted  <= 2'd0;
    else
      \$wnnz_IntTupGo___Pointer_QTree_Int_1_emitted  <= (\$wnnz_IntTupGo___Pointer_QTree_Int_1_r  ? 2'd0 :
                                                         \$wnnz_IntTupGo___Pointer_QTree_Int_1_done );
  
  /* fork (Ty Go) : ($wnnz_IntTupGo___Pointer_QTree_Intgo_8,Go) > [(go_8_1,Go),
                                                              (go_8_2,Go)] */
  logic [1:0] \$wnnz_IntTupGo___Pointer_QTree_Intgo_8_emitted ;
  logic [1:0] \$wnnz_IntTupGo___Pointer_QTree_Intgo_8_done ;
  assign go_8_1_d = (\$wnnz_IntTupGo___Pointer_QTree_Intgo_8_d [0] && (! \$wnnz_IntTupGo___Pointer_QTree_Intgo_8_emitted [0]));
  assign go_8_2_d = (\$wnnz_IntTupGo___Pointer_QTree_Intgo_8_d [0] && (! \$wnnz_IntTupGo___Pointer_QTree_Intgo_8_emitted [1]));
  assign \$wnnz_IntTupGo___Pointer_QTree_Intgo_8_done  = (\$wnnz_IntTupGo___Pointer_QTree_Intgo_8_emitted  | ({go_8_2_d[0],
                                                                                                               go_8_1_d[0]} & {go_8_2_r,
                                                                                                                               go_8_1_r}));
  assign \$wnnz_IntTupGo___Pointer_QTree_Intgo_8_r  = (& \$wnnz_IntTupGo___Pointer_QTree_Intgo_8_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \$wnnz_IntTupGo___Pointer_QTree_Intgo_8_emitted  <= 2'd0;
    else
      \$wnnz_IntTupGo___Pointer_QTree_Intgo_8_emitted  <= (\$wnnz_IntTupGo___Pointer_QTree_Intgo_8_r  ? 2'd0 :
                                                           \$wnnz_IntTupGo___Pointer_QTree_Intgo_8_done );
  
  /* buf (Ty Pointer_QTree_Int) : ($wnnz_IntTupGo___Pointer_QTree_Intwsvt,Pointer_QTree_Int) > (wsvt_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t \$wnnz_IntTupGo___Pointer_QTree_Intwsvt_bufchan_d ;
  logic \$wnnz_IntTupGo___Pointer_QTree_Intwsvt_bufchan_r ;
  assign \$wnnz_IntTupGo___Pointer_QTree_Intwsvt_r  = ((! \$wnnz_IntTupGo___Pointer_QTree_Intwsvt_bufchan_d [0]) || \$wnnz_IntTupGo___Pointer_QTree_Intwsvt_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \$wnnz_IntTupGo___Pointer_QTree_Intwsvt_bufchan_d  <= {16'd0,
                                                             1'd0};
    else
      if (\$wnnz_IntTupGo___Pointer_QTree_Intwsvt_r )
        \$wnnz_IntTupGo___Pointer_QTree_Intwsvt_bufchan_d  <= \$wnnz_IntTupGo___Pointer_QTree_Intwsvt_d ;
  Pointer_QTree_Int_t \$wnnz_IntTupGo___Pointer_QTree_Intwsvt_bufchan_buf ;
  assign \$wnnz_IntTupGo___Pointer_QTree_Intwsvt_bufchan_r  = (! \$wnnz_IntTupGo___Pointer_QTree_Intwsvt_bufchan_buf [0]);
  assign wsvt_1_argbuf_d = (\$wnnz_IntTupGo___Pointer_QTree_Intwsvt_bufchan_buf [0] ? \$wnnz_IntTupGo___Pointer_QTree_Intwsvt_bufchan_buf  :
                            \$wnnz_IntTupGo___Pointer_QTree_Intwsvt_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \$wnnz_IntTupGo___Pointer_QTree_Intwsvt_bufchan_buf  <= {16'd0,
                                                               1'd0};
    else
      if ((wsvt_1_argbuf_r && \$wnnz_IntTupGo___Pointer_QTree_Intwsvt_bufchan_buf [0]))
        \$wnnz_IntTupGo___Pointer_QTree_Intwsvt_bufchan_buf  <= {16'd0,
                                                                 1'd0};
      else if (((! wsvt_1_argbuf_r) && (! \$wnnz_IntTupGo___Pointer_QTree_Intwsvt_bufchan_buf [0])))
        \$wnnz_IntTupGo___Pointer_QTree_Intwsvt_bufchan_buf  <= \$wnnz_IntTupGo___Pointer_QTree_Intwsvt_bufchan_d ;
  
  /* buf (Ty Int#) : ($wnnz_Int_resbuf,Int#) > ($wmain_resbuf,Int#) */
  \Int#_t  \$wnnz_Int_resbuf_bufchan_d ;
  logic \$wnnz_Int_resbuf_bufchan_r ;
  assign \$wnnz_Int_resbuf_r  = ((! \$wnnz_Int_resbuf_bufchan_d [0]) || \$wnnz_Int_resbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \$wnnz_Int_resbuf_bufchan_d  <= {32'd0, 1'd0};
    else
      if (\$wnnz_Int_resbuf_r )
        \$wnnz_Int_resbuf_bufchan_d  <= \$wnnz_Int_resbuf_d ;
  \Int#_t  \$wnnz_Int_resbuf_bufchan_buf ;
  assign \$wnnz_Int_resbuf_bufchan_r  = (! \$wnnz_Int_resbuf_bufchan_buf [0]);
  assign \$wmain_resbuf_d  = (\$wnnz_Int_resbuf_bufchan_buf [0] ? \$wnnz_Int_resbuf_bufchan_buf  :
                              \$wnnz_Int_resbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \$wnnz_Int_resbuf_bufchan_buf  <= {32'd0, 1'd0};
    else
      if ((\$wmain_resbuf_r  && \$wnnz_Int_resbuf_bufchan_buf [0]))
        \$wnnz_Int_resbuf_bufchan_buf  <= {32'd0, 1'd0};
      else if (((! \$wmain_resbuf_r ) && (! \$wnnz_Int_resbuf_bufchan_buf [0])))
        \$wnnz_Int_resbuf_bufchan_buf  <= \$wnnz_Int_resbuf_bufchan_d ;
  
  /* mergectrl (Ty C2,
           Ty TupGo___MyDTInt_Bool___Int) : [(applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1,TupGo___MyDTInt_Bool___Int),
                                             (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int2,TupGo___MyDTInt_Bool___Int)] > (applyfnInt_Bool_5_choice,C2) (applyfnInt_Bool_5_data,TupGo___MyDTInt_Bool___Int) */
  logic [1:0] applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_select_d;
  assign applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_select_d = ((| applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_select_q) ? applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_select_q :
                                                                   (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_d[0] ? 2'd1 :
                                                                    (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int2_d[0] ? 2'd2 :
                                                                     2'd0)));
  logic [1:0] applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_select_q <= 2'd0;
    else
      applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_select_q <= (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_done ? 2'd0 :
                                                                 applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_select_d);
  logic [1:0] applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_emit_q <= 2'd0;
    else
      applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_emit_q <= (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_done ? 2'd0 :
                                                               applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_emit_d);
  logic [1:0] applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_emit_d;
  assign applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_emit_d = (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_emit_q | ({applyfnInt_Bool_5_choice_d[0],
                                                                                                                          applyfnInt_Bool_5_data_d[0]} & {applyfnInt_Bool_5_choice_r,
                                                                                                                                                          applyfnInt_Bool_5_data_r}));
  logic applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_done;
  assign applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_done = (& applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_emit_d);
  assign {applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int2_r,
          applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_r} = (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_done ? applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_select_d :
                                                              2'd0);
  assign applyfnInt_Bool_5_data_d = ((applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_select_d[0] && (! applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_emit_q[0])) ? applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_d :
                                     ((applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_select_d[1] && (! applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_emit_q[0])) ? applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int2_d :
                                      {32'd0, 1'd0}));
  assign applyfnInt_Bool_5_choice_d = ((applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_select_d[0] && (! applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_emit_q[1])) ? C1_2_dc(1'd1) :
                                       ((applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_select_d[1] && (! applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_emit_q[1])) ? C2_2_dc(1'd1) :
                                        {1'd0, 1'd0}));
  
  /* fork (Ty MyDTInt_Bool) : (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0,MyDTInt_Bool) > [(arg0_1,MyDTInt_Bool),
                                                                                           (arg0_2,MyDTInt_Bool),
                                                                                           (arg0_3,MyDTInt_Bool)] */
  logic [2:0] applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_emitted;
  logic [2:0] applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_done;
  assign arg0_1_d = (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_d[0] && (! applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_emitted[0]));
  assign arg0_2_d = (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_d[0] && (! applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_emitted[1]));
  assign arg0_3_d = (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_d[0] && (! applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_emitted[2]));
  assign applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_done = (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_emitted | ({arg0_3_d[0],
                                                                                                                             arg0_2_d[0],
                                                                                                                             arg0_1_d[0]} & {arg0_3_r,
                                                                                                                                             arg0_2_r,
                                                                                                                                             arg0_1_r}));
  assign applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_r = (& applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_emitted <= 3'd0;
    else
      applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_emitted <= (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_r ? 3'd0 :
                                                                  applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_done);
  
  /* buf (Ty MyBool) : (applyfnInt_Bool_5_1,MyBool) > (applyfnInt_Bool_5_resbuf,MyBool) */
  MyBool_t applyfnInt_Bool_5_1_bufchan_d;
  logic applyfnInt_Bool_5_1_bufchan_r;
  assign applyfnInt_Bool_5_1_r = ((! applyfnInt_Bool_5_1_bufchan_d[0]) || applyfnInt_Bool_5_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) applyfnInt_Bool_5_1_bufchan_d <= {1'd0, 1'd0};
    else
      if (applyfnInt_Bool_5_1_r)
        applyfnInt_Bool_5_1_bufchan_d <= applyfnInt_Bool_5_1_d;
  MyBool_t applyfnInt_Bool_5_1_bufchan_buf;
  assign applyfnInt_Bool_5_1_bufchan_r = (! applyfnInt_Bool_5_1_bufchan_buf[0]);
  assign applyfnInt_Bool_5_resbuf_d = (applyfnInt_Bool_5_1_bufchan_buf[0] ? applyfnInt_Bool_5_1_bufchan_buf :
                                       applyfnInt_Bool_5_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Bool_5_1_bufchan_buf <= {1'd0, 1'd0};
    else
      if ((applyfnInt_Bool_5_resbuf_r && applyfnInt_Bool_5_1_bufchan_buf[0]))
        applyfnInt_Bool_5_1_bufchan_buf <= {1'd0, 1'd0};
      else if (((! applyfnInt_Bool_5_resbuf_r) && (! applyfnInt_Bool_5_1_bufchan_buf[0])))
        applyfnInt_Bool_5_1_bufchan_buf <= applyfnInt_Bool_5_1_bufchan_d;
  
  /* buf (Ty MyBool) : (applyfnInt_Bool_5_2,MyBool) > (applyfnInt_Bool_5_2_argbuf,MyBool) */
  MyBool_t applyfnInt_Bool_5_2_bufchan_d;
  logic applyfnInt_Bool_5_2_bufchan_r;
  assign applyfnInt_Bool_5_2_r = ((! applyfnInt_Bool_5_2_bufchan_d[0]) || applyfnInt_Bool_5_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) applyfnInt_Bool_5_2_bufchan_d <= {1'd0, 1'd0};
    else
      if (applyfnInt_Bool_5_2_r)
        applyfnInt_Bool_5_2_bufchan_d <= applyfnInt_Bool_5_2_d;
  MyBool_t applyfnInt_Bool_5_2_bufchan_buf;
  assign applyfnInt_Bool_5_2_bufchan_r = (! applyfnInt_Bool_5_2_bufchan_buf[0]);
  assign applyfnInt_Bool_5_2_argbuf_d = (applyfnInt_Bool_5_2_bufchan_buf[0] ? applyfnInt_Bool_5_2_bufchan_buf :
                                         applyfnInt_Bool_5_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Bool_5_2_bufchan_buf <= {1'd0, 1'd0};
    else
      if ((applyfnInt_Bool_5_2_argbuf_r && applyfnInt_Bool_5_2_bufchan_buf[0]))
        applyfnInt_Bool_5_2_bufchan_buf <= {1'd0, 1'd0};
      else if (((! applyfnInt_Bool_5_2_argbuf_r) && (! applyfnInt_Bool_5_2_bufchan_buf[0])))
        applyfnInt_Bool_5_2_bufchan_buf <= applyfnInt_Bool_5_2_bufchan_d;
  
  /* fork (Ty MyBool) : (applyfnInt_Bool_5_2_argbuf,MyBool) > [(es_0_4_1,MyBool),
                                                          (es_0_4_2,MyBool),
                                                          (es_0_4_3,MyBool)] */
  logic [2:0] applyfnInt_Bool_5_2_argbuf_emitted;
  logic [2:0] applyfnInt_Bool_5_2_argbuf_done;
  assign es_0_4_1_d = {applyfnInt_Bool_5_2_argbuf_d[1:1],
                       (applyfnInt_Bool_5_2_argbuf_d[0] && (! applyfnInt_Bool_5_2_argbuf_emitted[0]))};
  assign es_0_4_2_d = {applyfnInt_Bool_5_2_argbuf_d[1:1],
                       (applyfnInt_Bool_5_2_argbuf_d[0] && (! applyfnInt_Bool_5_2_argbuf_emitted[1]))};
  assign es_0_4_3_d = {applyfnInt_Bool_5_2_argbuf_d[1:1],
                       (applyfnInt_Bool_5_2_argbuf_d[0] && (! applyfnInt_Bool_5_2_argbuf_emitted[2]))};
  assign applyfnInt_Bool_5_2_argbuf_done = (applyfnInt_Bool_5_2_argbuf_emitted | ({es_0_4_3_d[0],
                                                                                   es_0_4_2_d[0],
                                                                                   es_0_4_1_d[0]} & {es_0_4_3_r,
                                                                                                     es_0_4_2_r,
                                                                                                     es_0_4_1_r}));
  assign applyfnInt_Bool_5_2_argbuf_r = (& applyfnInt_Bool_5_2_argbuf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) applyfnInt_Bool_5_2_argbuf_emitted <= 3'd0;
    else
      applyfnInt_Bool_5_2_argbuf_emitted <= (applyfnInt_Bool_5_2_argbuf_r ? 3'd0 :
                                             applyfnInt_Bool_5_2_argbuf_done);
  
  /* demux (Ty C2,
       Ty MyBool) : (applyfnInt_Bool_5_choice,C2) (lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux,MyBool) > [(applyfnInt_Bool_5_1,MyBool),
                                                                                                                                 (applyfnInt_Bool_5_2,MyBool)] */
  logic [1:0] lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_onehotd;
  always_comb
    if ((applyfnInt_Bool_5_choice_d[0] && lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_d[0]))
      unique case (applyfnInt_Bool_5_choice_d[1:1])
        1'd0:
          lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_onehotd = 2'd1;
        1'd1:
          lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_onehotd = 2'd2;
        default:
          lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_onehotd = 2'd0;
      endcase
    else
      lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_onehotd = 2'd0;
  assign applyfnInt_Bool_5_1_d = {lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_d[1:1],
                                  lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_onehotd[0]};
  assign applyfnInt_Bool_5_2_d = {lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_d[1:1],
                                  lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_onehotd[1]};
  assign lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_r = (| (lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_onehotd & {applyfnInt_Bool_5_2_r,
                                                                                                                                                                  applyfnInt_Bool_5_1_r}));
  assign applyfnInt_Bool_5_choice_r = lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_r;
  
  /* destruct (Ty TupGo___MyDTInt_Bool___Int,
          Dcon TupGo___MyDTInt_Bool___Int) : (applyfnInt_Bool_5_data,TupGo___MyDTInt_Bool___Int) > [(applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intgo_9,Go),
                                                                                                    (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0,MyDTInt_Bool),
                                                                                                    (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg1,Int)] */
  logic [2:0] applyfnInt_Bool_5_data_emitted;
  logic [2:0] applyfnInt_Bool_5_data_done;
  assign applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intgo_9_d = (applyfnInt_Bool_5_data_d[0] && (! applyfnInt_Bool_5_data_emitted[0]));
  assign applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_d = (applyfnInt_Bool_5_data_d[0] && (! applyfnInt_Bool_5_data_emitted[1]));
  assign applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg1_d = {applyfnInt_Bool_5_data_d[32:1],
                                                              (applyfnInt_Bool_5_data_d[0] && (! applyfnInt_Bool_5_data_emitted[2]))};
  assign applyfnInt_Bool_5_data_done = (applyfnInt_Bool_5_data_emitted | ({applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg1_d[0],
                                                                           applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_d[0],
                                                                           applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intgo_9_d[0]} & {applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg1_r,
                                                                                                                                    applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_r,
                                                                                                                                    applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intgo_9_r}));
  assign applyfnInt_Bool_5_data_r = (& applyfnInt_Bool_5_data_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) applyfnInt_Bool_5_data_emitted <= 3'd0;
    else
      applyfnInt_Bool_5_data_emitted <= (applyfnInt_Bool_5_data_r ? 3'd0 :
                                         applyfnInt_Bool_5_data_done);
  
  /* fork (Ty MyBool) : (applyfnInt_Bool_5_resbuf,MyBool) > [(es_0_5_1,MyBool),
                                                        (es_0_5_2,MyBool),
                                                        (es_0_5_3,MyBool)] */
  logic [2:0] applyfnInt_Bool_5_resbuf_emitted;
  logic [2:0] applyfnInt_Bool_5_resbuf_done;
  assign es_0_5_1_d = {applyfnInt_Bool_5_resbuf_d[1:1],
                       (applyfnInt_Bool_5_resbuf_d[0] && (! applyfnInt_Bool_5_resbuf_emitted[0]))};
  assign es_0_5_2_d = {applyfnInt_Bool_5_resbuf_d[1:1],
                       (applyfnInt_Bool_5_resbuf_d[0] && (! applyfnInt_Bool_5_resbuf_emitted[1]))};
  assign es_0_5_3_d = {applyfnInt_Bool_5_resbuf_d[1:1],
                       (applyfnInt_Bool_5_resbuf_d[0] && (! applyfnInt_Bool_5_resbuf_emitted[2]))};
  assign applyfnInt_Bool_5_resbuf_done = (applyfnInt_Bool_5_resbuf_emitted | ({es_0_5_3_d[0],
                                                                               es_0_5_2_d[0],
                                                                               es_0_5_1_d[0]} & {es_0_5_3_r,
                                                                                                 es_0_5_2_r,
                                                                                                 es_0_5_1_r}));
  assign applyfnInt_Bool_5_resbuf_r = (& applyfnInt_Bool_5_resbuf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) applyfnInt_Bool_5_resbuf_emitted <= 3'd0;
    else
      applyfnInt_Bool_5_resbuf_emitted <= (applyfnInt_Bool_5_resbuf_r ? 3'd0 :
                                           applyfnInt_Bool_5_resbuf_done);
  
  /* destruct (Ty TupGo___MyDTInt_Int___Int,
          Dcon TupGo___MyDTInt_Int___Int) : (applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1,TupGo___MyDTInt_Int___Int) > [(applyfnInt_Int_5TupGo___MyDTInt_Int___Intgo_10,Go),
                                                                                                                       (applyfnInt_Int_5TupGo___MyDTInt_Int___Intarg0_2,MyDTInt_Int),
                                                                                                                       (applyfnInt_Int_5TupGo___MyDTInt_Int___Intarg1_1,Int)] */
  logic [2:0] applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_emitted;
  logic [2:0] applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_done;
  assign applyfnInt_Int_5TupGo___MyDTInt_Int___Intgo_10_d = (applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_d[0] && (! applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_emitted[0]));
  assign applyfnInt_Int_5TupGo___MyDTInt_Int___Intarg0_2_d = (applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_d[0] && (! applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_emitted[1]));
  assign applyfnInt_Int_5TupGo___MyDTInt_Int___Intarg1_1_d = {applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_d[32:1],
                                                              (applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_d[0] && (! applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_emitted[2]))};
  assign applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_done = (applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_emitted | ({applyfnInt_Int_5TupGo___MyDTInt_Int___Intarg1_1_d[0],
                                                                                                                     applyfnInt_Int_5TupGo___MyDTInt_Int___Intarg0_2_d[0],
                                                                                                                     applyfnInt_Int_5TupGo___MyDTInt_Int___Intgo_10_d[0]} & {applyfnInt_Int_5TupGo___MyDTInt_Int___Intarg1_1_r,
                                                                                                                                                                             applyfnInt_Int_5TupGo___MyDTInt_Int___Intarg0_2_r,
                                                                                                                                                                             applyfnInt_Int_5TupGo___MyDTInt_Int___Intgo_10_r}));
  assign applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_r = (& applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_emitted <= 3'd0;
    else
      applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_emitted <= (applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_r ? 3'd0 :
                                                              applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_done);
  
  /* fork (Ty MyDTInt_Int) : (applyfnInt_Int_5TupGo___MyDTInt_Int___Intarg0_2,MyDTInt_Int) > [(arg0_2_1,MyDTInt_Int),
                                                                                         (arg0_2_2,MyDTInt_Int),
                                                                                         (arg0_2_3,MyDTInt_Int)] */
  logic [2:0] applyfnInt_Int_5TupGo___MyDTInt_Int___Intarg0_2_emitted;
  logic [2:0] applyfnInt_Int_5TupGo___MyDTInt_Int___Intarg0_2_done;
  assign arg0_2_1_d = (applyfnInt_Int_5TupGo___MyDTInt_Int___Intarg0_2_d[0] && (! applyfnInt_Int_5TupGo___MyDTInt_Int___Intarg0_2_emitted[0]));
  assign arg0_2_2_d = (applyfnInt_Int_5TupGo___MyDTInt_Int___Intarg0_2_d[0] && (! applyfnInt_Int_5TupGo___MyDTInt_Int___Intarg0_2_emitted[1]));
  assign arg0_2_3_d = (applyfnInt_Int_5TupGo___MyDTInt_Int___Intarg0_2_d[0] && (! applyfnInt_Int_5TupGo___MyDTInt_Int___Intarg0_2_emitted[2]));
  assign applyfnInt_Int_5TupGo___MyDTInt_Int___Intarg0_2_done = (applyfnInt_Int_5TupGo___MyDTInt_Int___Intarg0_2_emitted | ({arg0_2_3_d[0],
                                                                                                                             arg0_2_2_d[0],
                                                                                                                             arg0_2_1_d[0]} & {arg0_2_3_r,
                                                                                                                                               arg0_2_2_r,
                                                                                                                                               arg0_2_1_r}));
  assign applyfnInt_Int_5TupGo___MyDTInt_Int___Intarg0_2_r = (& applyfnInt_Int_5TupGo___MyDTInt_Int___Intarg0_2_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_5TupGo___MyDTInt_Int___Intarg0_2_emitted <= 3'd0;
    else
      applyfnInt_Int_5TupGo___MyDTInt_Int___Intarg0_2_emitted <= (applyfnInt_Int_5TupGo___MyDTInt_Int___Intarg0_2_r ? 3'd0 :
                                                                  applyfnInt_Int_5TupGo___MyDTInt_Int___Intarg0_2_done);
  
  /* fork (Ty Int) : (applyfnInt_Int_5_resbuf,Int) > [(xacr_1,Int),
                                                 (xacr_2,Int)] */
  logic [1:0] applyfnInt_Int_5_resbuf_emitted;
  logic [1:0] applyfnInt_Int_5_resbuf_done;
  assign xacr_1_d = {applyfnInt_Int_5_resbuf_d[32:1],
                     (applyfnInt_Int_5_resbuf_d[0] && (! applyfnInt_Int_5_resbuf_emitted[0]))};
  assign xacr_2_d = {applyfnInt_Int_5_resbuf_d[32:1],
                     (applyfnInt_Int_5_resbuf_d[0] && (! applyfnInt_Int_5_resbuf_emitted[1]))};
  assign applyfnInt_Int_5_resbuf_done = (applyfnInt_Int_5_resbuf_emitted | ({xacr_2_d[0],
                                                                             xacr_1_d[0]} & {xacr_2_r,
                                                                                             xacr_1_r}));
  assign applyfnInt_Int_5_resbuf_r = (& applyfnInt_Int_5_resbuf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) applyfnInt_Int_5_resbuf_emitted <= 2'd0;
    else
      applyfnInt_Int_5_resbuf_emitted <= (applyfnInt_Int_5_resbuf_r ? 2'd0 :
                                          applyfnInt_Int_5_resbuf_done);
  
  /* destruct (Ty TupMyDTInt_Int_Int___Int___Int,
          Dcon TupMyDTInt_Int_Int___Int___Int) : (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1,TupMyDTInt_Int_Int___Int___Int) > [(applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_4,MyDTInt_Int_Int),
                                                                                                                                          (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg2,Int),
                                                                                                                                          (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg1_2,Int)] */
  logic [2:0] applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_emitted;
  logic [2:0] applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_done;
  assign applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_4_d = (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_d[0] && (! applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_emitted[0]));
  assign applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg2_d = {applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_d[32:1],
                                                                     (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_d[0] && (! applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_emitted[1]))};
  assign applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg1_2_d = {applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_d[64:33],
                                                                       (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_d[0] && (! applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_emitted[2]))};
  assign applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_done = (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_emitted | ({applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg1_2_d[0],
                                                                                                                                       applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg2_d[0],
                                                                                                                                       applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_4_d[0]} & {applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg1_2_r,
                                                                                                                                                                                                         applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg2_r,
                                                                                                                                                                                                         applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_4_r}));
  assign applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_r = (& applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_emitted <= 3'd0;
    else
      applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_emitted <= (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_r ? 3'd0 :
                                                                       applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_done);
  
  /* fork (Ty MyDTInt_Int_Int) : (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_4,MyDTInt_Int_Int) > [(arg0_4_1,MyDTInt_Int_Int),
                                                                                                          (arg0_4_2,MyDTInt_Int_Int),
                                                                                                          (arg0_4_3,MyDTInt_Int_Int)] */
  logic [2:0] applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_4_emitted;
  logic [2:0] applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_4_done;
  assign arg0_4_1_d = (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_4_d[0] && (! applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_4_emitted[0]));
  assign arg0_4_2_d = (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_4_d[0] && (! applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_4_emitted[1]));
  assign arg0_4_3_d = (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_4_d[0] && (! applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_4_emitted[2]));
  assign applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_4_done = (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_4_emitted | ({arg0_4_3_d[0],
                                                                                                                                               arg0_4_2_d[0],
                                                                                                                                               arg0_4_1_d[0]} & {arg0_4_3_r,
                                                                                                                                                                 arg0_4_2_r,
                                                                                                                                                                 arg0_4_1_r}));
  assign applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_4_r = (& applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_4_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_4_emitted <= 3'd0;
    else
      applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_4_emitted <= (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_4_r ? 3'd0 :
                                                                           applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_4_done);
  
  /* fork (Ty Int) : (applyfnInt_Int_Int_5_resbuf,Int) > [(xacr_1_1,Int),
                                                     (xacr_1_2,Int)] */
  logic [1:0] applyfnInt_Int_Int_5_resbuf_emitted;
  logic [1:0] applyfnInt_Int_Int_5_resbuf_done;
  assign xacr_1_1_d = {applyfnInt_Int_Int_5_resbuf_d[32:1],
                       (applyfnInt_Int_Int_5_resbuf_d[0] && (! applyfnInt_Int_Int_5_resbuf_emitted[0]))};
  assign xacr_1_2_d = {applyfnInt_Int_Int_5_resbuf_d[32:1],
                       (applyfnInt_Int_Int_5_resbuf_d[0] && (! applyfnInt_Int_Int_5_resbuf_emitted[1]))};
  assign applyfnInt_Int_Int_5_resbuf_done = (applyfnInt_Int_Int_5_resbuf_emitted | ({xacr_1_2_d[0],
                                                                                     xacr_1_1_d[0]} & {xacr_1_2_r,
                                                                                                       xacr_1_1_r}));
  assign applyfnInt_Int_Int_5_resbuf_r = (& applyfnInt_Int_Int_5_resbuf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) applyfnInt_Int_Int_5_resbuf_emitted <= 2'd0;
    else
      applyfnInt_Int_Int_5_resbuf_emitted <= (applyfnInt_Int_Int_5_resbuf_r ? 2'd0 :
                                              applyfnInt_Int_Int_5_resbuf_done);
  
  /* demux (Ty MyDTInt_Bool,
       Ty Int) : (arg0_1,MyDTInt_Bool) (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg1,Int) > [(arg0_1Dcon_eqZero,Int)] */
  assign arg0_1Dcon_eqZero_d = {applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg1_d[32:1],
                                (arg0_1_d[0] && applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg1_d[0])};
  assign applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg1_r = (arg0_1Dcon_eqZero_r && (arg0_1_d[0] && applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg1_d[0]));
  assign arg0_1_r = (arg0_1Dcon_eqZero_r && (arg0_1_d[0] && applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg1_d[0]));
  
  /* fork (Ty Int) : (arg0_1Dcon_eqZero,Int) > [(arg0_1Dcon_eqZero_1,Int),
                                           (arg0_1Dcon_eqZero_2,Int),
                                           (arg0_1Dcon_eqZero_3,Int),
                                           (arg0_1Dcon_eqZero_4,Int)] */
  logic [3:0] arg0_1Dcon_eqZero_emitted;
  logic [3:0] arg0_1Dcon_eqZero_done;
  assign arg0_1Dcon_eqZero_1_d = {arg0_1Dcon_eqZero_d[32:1],
                                  (arg0_1Dcon_eqZero_d[0] && (! arg0_1Dcon_eqZero_emitted[0]))};
  assign arg0_1Dcon_eqZero_2_d = {arg0_1Dcon_eqZero_d[32:1],
                                  (arg0_1Dcon_eqZero_d[0] && (! arg0_1Dcon_eqZero_emitted[1]))};
  assign arg0_1Dcon_eqZero_3_d = {arg0_1Dcon_eqZero_d[32:1],
                                  (arg0_1Dcon_eqZero_d[0] && (! arg0_1Dcon_eqZero_emitted[2]))};
  assign arg0_1Dcon_eqZero_4_d = {arg0_1Dcon_eqZero_d[32:1],
                                  (arg0_1Dcon_eqZero_d[0] && (! arg0_1Dcon_eqZero_emitted[3]))};
  assign arg0_1Dcon_eqZero_done = (arg0_1Dcon_eqZero_emitted | ({arg0_1Dcon_eqZero_4_d[0],
                                                                 arg0_1Dcon_eqZero_3_d[0],
                                                                 arg0_1Dcon_eqZero_2_d[0],
                                                                 arg0_1Dcon_eqZero_1_d[0]} & {arg0_1Dcon_eqZero_4_r,
                                                                                              arg0_1Dcon_eqZero_3_r,
                                                                                              arg0_1Dcon_eqZero_2_r,
                                                                                              arg0_1Dcon_eqZero_1_r}));
  assign arg0_1Dcon_eqZero_r = (& arg0_1Dcon_eqZero_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) arg0_1Dcon_eqZero_emitted <= 4'd0;
    else
      arg0_1Dcon_eqZero_emitted <= (arg0_1Dcon_eqZero_r ? 4'd0 :
                                    arg0_1Dcon_eqZero_done);
  
  /* destruct (Ty Int,
          Dcon I#) : (arg0_1Dcon_eqZero_1I#,Int) > [(x1aqk_destruct,Int#)] */
  assign x1aqk_destruct_d = {\arg0_1Dcon_eqZero_1I#_d [32:1],
                             \arg0_1Dcon_eqZero_1I#_d [0]};
  assign \arg0_1Dcon_eqZero_1I#_r  = x1aqk_destruct_r;
  
  /* demux (Ty Int,
       Ty Int) : (arg0_1Dcon_eqZero_2,Int) (arg0_1Dcon_eqZero_1,Int) > [(arg0_1Dcon_eqZero_1I#,Int)] */
  assign \arg0_1Dcon_eqZero_1I#_d  = {arg0_1Dcon_eqZero_1_d[32:1],
                                      (arg0_1Dcon_eqZero_2_d[0] && arg0_1Dcon_eqZero_1_d[0])};
  assign arg0_1Dcon_eqZero_1_r = (\arg0_1Dcon_eqZero_1I#_r  && (arg0_1Dcon_eqZero_2_d[0] && arg0_1Dcon_eqZero_1_d[0]));
  assign arg0_1Dcon_eqZero_2_r = (\arg0_1Dcon_eqZero_1I#_r  && (arg0_1Dcon_eqZero_2_d[0] && arg0_1Dcon_eqZero_1_d[0]));
  
  /* demux (Ty Int,
       Ty Go) : (arg0_1Dcon_eqZero_3,Int) (arg0_2Dcon_eqZero,Go) > [(arg0_1Dcon_eqZero_3I#,Go)] */
  assign \arg0_1Dcon_eqZero_3I#_d  = (arg0_1Dcon_eqZero_3_d[0] && arg0_2Dcon_eqZero_d[0]);
  assign arg0_2Dcon_eqZero_r = (\arg0_1Dcon_eqZero_3I#_r  && (arg0_1Dcon_eqZero_3_d[0] && arg0_2Dcon_eqZero_d[0]));
  assign arg0_1Dcon_eqZero_3_r = (\arg0_1Dcon_eqZero_3I#_r  && (arg0_1Dcon_eqZero_3_d[0] && arg0_2Dcon_eqZero_d[0]));
  
  /* fork (Ty Go) : (arg0_1Dcon_eqZero_3I#,Go) > [(arg0_1Dcon_eqZero_3I#_1,Go),
                                             (arg0_1Dcon_eqZero_3I#_2,Go),
                                             (arg0_1Dcon_eqZero_3I#_3,Go)] */
  logic [2:0] \arg0_1Dcon_eqZero_3I#_emitted ;
  logic [2:0] \arg0_1Dcon_eqZero_3I#_done ;
  assign \arg0_1Dcon_eqZero_3I#_1_d  = (\arg0_1Dcon_eqZero_3I#_d [0] && (! \arg0_1Dcon_eqZero_3I#_emitted [0]));
  assign \arg0_1Dcon_eqZero_3I#_2_d  = (\arg0_1Dcon_eqZero_3I#_d [0] && (! \arg0_1Dcon_eqZero_3I#_emitted [1]));
  assign \arg0_1Dcon_eqZero_3I#_3_d  = (\arg0_1Dcon_eqZero_3I#_d [0] && (! \arg0_1Dcon_eqZero_3I#_emitted [2]));
  assign \arg0_1Dcon_eqZero_3I#_done  = (\arg0_1Dcon_eqZero_3I#_emitted  | ({\arg0_1Dcon_eqZero_3I#_3_d [0],
                                                                             \arg0_1Dcon_eqZero_3I#_2_d [0],
                                                                             \arg0_1Dcon_eqZero_3I#_1_d [0]} & {\arg0_1Dcon_eqZero_3I#_3_r ,
                                                                                                                \arg0_1Dcon_eqZero_3I#_2_r ,
                                                                                                                \arg0_1Dcon_eqZero_3I#_1_r }));
  assign \arg0_1Dcon_eqZero_3I#_r  = (& \arg0_1Dcon_eqZero_3I#_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \arg0_1Dcon_eqZero_3I#_emitted  <= 3'd0;
    else
      \arg0_1Dcon_eqZero_3I#_emitted  <= (\arg0_1Dcon_eqZero_3I#_r  ? 3'd0 :
                                          \arg0_1Dcon_eqZero_3I#_done );
  
  /* buf (Ty Go) : (arg0_1Dcon_eqZero_3I#_1,Go) > (arg0_1Dcon_eqZero_3I#_1_argbuf,Go) */
  Go_t \arg0_1Dcon_eqZero_3I#_1_bufchan_d ;
  logic \arg0_1Dcon_eqZero_3I#_1_bufchan_r ;
  assign \arg0_1Dcon_eqZero_3I#_1_r  = ((! \arg0_1Dcon_eqZero_3I#_1_bufchan_d [0]) || \arg0_1Dcon_eqZero_3I#_1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \arg0_1Dcon_eqZero_3I#_1_bufchan_d  <= 1'd0;
    else
      if (\arg0_1Dcon_eqZero_3I#_1_r )
        \arg0_1Dcon_eqZero_3I#_1_bufchan_d  <= \arg0_1Dcon_eqZero_3I#_1_d ;
  Go_t \arg0_1Dcon_eqZero_3I#_1_bufchan_buf ;
  assign \arg0_1Dcon_eqZero_3I#_1_bufchan_r  = (! \arg0_1Dcon_eqZero_3I#_1_bufchan_buf [0]);
  assign \arg0_1Dcon_eqZero_3I#_1_argbuf_d  = (\arg0_1Dcon_eqZero_3I#_1_bufchan_buf [0] ? \arg0_1Dcon_eqZero_3I#_1_bufchan_buf  :
                                               \arg0_1Dcon_eqZero_3I#_1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \arg0_1Dcon_eqZero_3I#_1_bufchan_buf  <= 1'd0;
    else
      if ((\arg0_1Dcon_eqZero_3I#_1_argbuf_r  && \arg0_1Dcon_eqZero_3I#_1_bufchan_buf [0]))
        \arg0_1Dcon_eqZero_3I#_1_bufchan_buf  <= 1'd0;
      else if (((! \arg0_1Dcon_eqZero_3I#_1_argbuf_r ) && (! \arg0_1Dcon_eqZero_3I#_1_bufchan_buf [0])))
        \arg0_1Dcon_eqZero_3I#_1_bufchan_buf  <= \arg0_1Dcon_eqZero_3I#_1_bufchan_d ;
  
  /* const (Ty Int#,
       Lit 0) : (arg0_1Dcon_eqZero_3I#_1_argbuf,Go) > (arg0_1Dcon_eqZero_3I#_1_argbuf_0,Int#) */
  assign \arg0_1Dcon_eqZero_3I#_1_argbuf_0_d  = {32'd0,
                                                 \arg0_1Dcon_eqZero_3I#_1_argbuf_d [0]};
  assign \arg0_1Dcon_eqZero_3I#_1_argbuf_r  = \arg0_1Dcon_eqZero_3I#_1_argbuf_0_r ;
  
  /* op_eq (Ty Int#) : (arg0_1Dcon_eqZero_3I#_1_argbuf_0,Int#) (x1aqk_destruct,Int#) > (lizzieLet1_1wild1X1h_1_Eq,Bool) */
  assign lizzieLet1_1wild1X1h_1_Eq_d = {(\arg0_1Dcon_eqZero_3I#_1_argbuf_0_d [32:1] == x1aqk_destruct_d[32:1]),
                                        (\arg0_1Dcon_eqZero_3I#_1_argbuf_0_d [0] && x1aqk_destruct_d[0])};
  assign {\arg0_1Dcon_eqZero_3I#_1_argbuf_0_r ,
          x1aqk_destruct_r} = {2 {(lizzieLet1_1wild1X1h_1_Eq_r && lizzieLet1_1wild1X1h_1_Eq_d[0])}};
  
  /* buf (Ty Go) : (arg0_1Dcon_eqZero_3I#_2,Go) > (arg0_1Dcon_eqZero_3I#_2_argbuf,Go) */
  Go_t \arg0_1Dcon_eqZero_3I#_2_bufchan_d ;
  logic \arg0_1Dcon_eqZero_3I#_2_bufchan_r ;
  assign \arg0_1Dcon_eqZero_3I#_2_r  = ((! \arg0_1Dcon_eqZero_3I#_2_bufchan_d [0]) || \arg0_1Dcon_eqZero_3I#_2_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \arg0_1Dcon_eqZero_3I#_2_bufchan_d  <= 1'd0;
    else
      if (\arg0_1Dcon_eqZero_3I#_2_r )
        \arg0_1Dcon_eqZero_3I#_2_bufchan_d  <= \arg0_1Dcon_eqZero_3I#_2_d ;
  Go_t \arg0_1Dcon_eqZero_3I#_2_bufchan_buf ;
  assign \arg0_1Dcon_eqZero_3I#_2_bufchan_r  = (! \arg0_1Dcon_eqZero_3I#_2_bufchan_buf [0]);
  assign \arg0_1Dcon_eqZero_3I#_2_argbuf_d  = (\arg0_1Dcon_eqZero_3I#_2_bufchan_buf [0] ? \arg0_1Dcon_eqZero_3I#_2_bufchan_buf  :
                                               \arg0_1Dcon_eqZero_3I#_2_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \arg0_1Dcon_eqZero_3I#_2_bufchan_buf  <= 1'd0;
    else
      if ((\arg0_1Dcon_eqZero_3I#_2_argbuf_r  && \arg0_1Dcon_eqZero_3I#_2_bufchan_buf [0]))
        \arg0_1Dcon_eqZero_3I#_2_bufchan_buf  <= 1'd0;
      else if (((! \arg0_1Dcon_eqZero_3I#_2_argbuf_r ) && (! \arg0_1Dcon_eqZero_3I#_2_bufchan_buf [0])))
        \arg0_1Dcon_eqZero_3I#_2_bufchan_buf  <= \arg0_1Dcon_eqZero_3I#_2_bufchan_d ;
  
  /* dcon (Ty TupGo___Bool,
      Dcon TupGo___Bool) : [(arg0_1Dcon_eqZero_3I#_2_argbuf,Go),
                            (lizzieLet2_1_argbuf,Bool)] > (boolConvert_1TupGo___Bool_1,TupGo___Bool) */
  assign boolConvert_1TupGo___Bool_1_d = TupGo___Bool_dc((& {\arg0_1Dcon_eqZero_3I#_2_argbuf_d [0],
                                                             lizzieLet2_1_argbuf_d[0]}), \arg0_1Dcon_eqZero_3I#_2_argbuf_d , lizzieLet2_1_argbuf_d);
  assign {\arg0_1Dcon_eqZero_3I#_2_argbuf_r ,
          lizzieLet2_1_argbuf_r} = {2 {(boolConvert_1TupGo___Bool_1_r && boolConvert_1TupGo___Bool_1_d[0])}};
  
  /* mux (Ty Int,
     Ty MyBool) : (arg0_1Dcon_eqZero_4,Int) [(lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux,MyBool)] > (lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux,MyBool) */
  assign lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_d = {lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_d[1:1],
                                                                             (arg0_1Dcon_eqZero_4_d[0] && lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_d[0])};
  assign lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_r = (lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_r && (arg0_1Dcon_eqZero_4_d[0] && lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_d[0]));
  assign arg0_1Dcon_eqZero_4_r = (lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_r && (arg0_1Dcon_eqZero_4_d[0] && lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_d[0]));
  
  /* demux (Ty MyDTInt_Bool,
       Ty Go) : (arg0_2,MyDTInt_Bool) (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intgo_9,Go) > [(arg0_2Dcon_eqZero,Go)] */
  assign arg0_2Dcon_eqZero_d = (arg0_2_d[0] && applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intgo_9_d[0]);
  assign applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intgo_9_r = (arg0_2Dcon_eqZero_r && (arg0_2_d[0] && applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intgo_9_d[0]));
  assign arg0_2_r = (arg0_2Dcon_eqZero_r && (arg0_2_d[0] && applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intgo_9_d[0]));
  
  /* demux (Ty MyDTInt_Int,
       Ty Int) : (arg0_2_1,MyDTInt_Int) (applyfnInt_Int_5TupGo___MyDTInt_Int___Intarg1_1,Int) > [(arg0_2_1Dcon_main1,Int)] */
  assign arg0_2_1Dcon_main1_d = {applyfnInt_Int_5TupGo___MyDTInt_Int___Intarg1_1_d[32:1],
                                 (arg0_2_1_d[0] && applyfnInt_Int_5TupGo___MyDTInt_Int___Intarg1_1_d[0])};
  assign applyfnInt_Int_5TupGo___MyDTInt_Int___Intarg1_1_r = (arg0_2_1Dcon_main1_r && (arg0_2_1_d[0] && applyfnInt_Int_5TupGo___MyDTInt_Int___Intarg1_1_d[0]));
  assign arg0_2_1_r = (arg0_2_1Dcon_main1_r && (arg0_2_1_d[0] && applyfnInt_Int_5TupGo___MyDTInt_Int___Intarg1_1_d[0]));
  
  /* fork (Ty Int) : (arg0_2_1Dcon_main1,Int) > [(arg0_2_1Dcon_main1_1,Int),
                                            (arg0_2_1Dcon_main1_2,Int),
                                            (arg0_2_1Dcon_main1_3,Int),
                                            (arg0_2_1Dcon_main1_4,Int)] */
  logic [3:0] arg0_2_1Dcon_main1_emitted;
  logic [3:0] arg0_2_1Dcon_main1_done;
  assign arg0_2_1Dcon_main1_1_d = {arg0_2_1Dcon_main1_d[32:1],
                                   (arg0_2_1Dcon_main1_d[0] && (! arg0_2_1Dcon_main1_emitted[0]))};
  assign arg0_2_1Dcon_main1_2_d = {arg0_2_1Dcon_main1_d[32:1],
                                   (arg0_2_1Dcon_main1_d[0] && (! arg0_2_1Dcon_main1_emitted[1]))};
  assign arg0_2_1Dcon_main1_3_d = {arg0_2_1Dcon_main1_d[32:1],
                                   (arg0_2_1Dcon_main1_d[0] && (! arg0_2_1Dcon_main1_emitted[2]))};
  assign arg0_2_1Dcon_main1_4_d = {arg0_2_1Dcon_main1_d[32:1],
                                   (arg0_2_1Dcon_main1_d[0] && (! arg0_2_1Dcon_main1_emitted[3]))};
  assign arg0_2_1Dcon_main1_done = (arg0_2_1Dcon_main1_emitted | ({arg0_2_1Dcon_main1_4_d[0],
                                                                   arg0_2_1Dcon_main1_3_d[0],
                                                                   arg0_2_1Dcon_main1_2_d[0],
                                                                   arg0_2_1Dcon_main1_1_d[0]} & {arg0_2_1Dcon_main1_4_r,
                                                                                                 arg0_2_1Dcon_main1_3_r,
                                                                                                 arg0_2_1Dcon_main1_2_r,
                                                                                                 arg0_2_1Dcon_main1_1_r}));
  assign arg0_2_1Dcon_main1_r = (& arg0_2_1Dcon_main1_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) arg0_2_1Dcon_main1_emitted <= 4'd0;
    else
      arg0_2_1Dcon_main1_emitted <= (arg0_2_1Dcon_main1_r ? 4'd0 :
                                     arg0_2_1Dcon_main1_done);
  
  /* destruct (Ty Int,
          Dcon I#) : (arg0_2_1Dcon_main1_1I#,Int) > [(xaqa_destruct,Int#)] */
  assign xaqa_destruct_d = {\arg0_2_1Dcon_main1_1I#_d [32:1],
                            \arg0_2_1Dcon_main1_1I#_d [0]};
  assign \arg0_2_1Dcon_main1_1I#_r  = xaqa_destruct_r;
  
  /* demux (Ty Int,
       Ty Int) : (arg0_2_1Dcon_main1_2,Int) (arg0_2_1Dcon_main1_1,Int) > [(arg0_2_1Dcon_main1_1I#,Int)] */
  assign \arg0_2_1Dcon_main1_1I#_d  = {arg0_2_1Dcon_main1_1_d[32:1],
                                       (arg0_2_1Dcon_main1_2_d[0] && arg0_2_1Dcon_main1_1_d[0])};
  assign arg0_2_1Dcon_main1_1_r = (\arg0_2_1Dcon_main1_1I#_r  && (arg0_2_1Dcon_main1_2_d[0] && arg0_2_1Dcon_main1_1_d[0]));
  assign arg0_2_1Dcon_main1_2_r = (\arg0_2_1Dcon_main1_1I#_r  && (arg0_2_1Dcon_main1_2_d[0] && arg0_2_1Dcon_main1_1_d[0]));
  
  /* demux (Ty Int,
       Ty Go) : (arg0_2_1Dcon_main1_3,Int) (arg0_2_2Dcon_main1,Go) > [(arg0_2_1Dcon_main1_3I#,Go)] */
  assign \arg0_2_1Dcon_main1_3I#_d  = (arg0_2_1Dcon_main1_3_d[0] && arg0_2_2Dcon_main1_d[0]);
  assign arg0_2_2Dcon_main1_r = (\arg0_2_1Dcon_main1_3I#_r  && (arg0_2_1Dcon_main1_3_d[0] && arg0_2_2Dcon_main1_d[0]));
  assign arg0_2_1Dcon_main1_3_r = (\arg0_2_1Dcon_main1_3I#_r  && (arg0_2_1Dcon_main1_3_d[0] && arg0_2_2Dcon_main1_d[0]));
  
  /* buf (Ty Go) : (arg0_2_1Dcon_main1_3I#,Go) > (arg0_2_1Dcon_main1_3I#_1_argbuf,Go) */
  Go_t \arg0_2_1Dcon_main1_3I#_bufchan_d ;
  logic \arg0_2_1Dcon_main1_3I#_bufchan_r ;
  assign \arg0_2_1Dcon_main1_3I#_r  = ((! \arg0_2_1Dcon_main1_3I#_bufchan_d [0]) || \arg0_2_1Dcon_main1_3I#_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \arg0_2_1Dcon_main1_3I#_bufchan_d  <= 1'd0;
    else
      if (\arg0_2_1Dcon_main1_3I#_r )
        \arg0_2_1Dcon_main1_3I#_bufchan_d  <= \arg0_2_1Dcon_main1_3I#_d ;
  Go_t \arg0_2_1Dcon_main1_3I#_bufchan_buf ;
  assign \arg0_2_1Dcon_main1_3I#_bufchan_r  = (! \arg0_2_1Dcon_main1_3I#_bufchan_buf [0]);
  assign \arg0_2_1Dcon_main1_3I#_1_argbuf_d  = (\arg0_2_1Dcon_main1_3I#_bufchan_buf [0] ? \arg0_2_1Dcon_main1_3I#_bufchan_buf  :
                                                \arg0_2_1Dcon_main1_3I#_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \arg0_2_1Dcon_main1_3I#_bufchan_buf  <= 1'd0;
    else
      if ((\arg0_2_1Dcon_main1_3I#_1_argbuf_r  && \arg0_2_1Dcon_main1_3I#_bufchan_buf [0]))
        \arg0_2_1Dcon_main1_3I#_bufchan_buf  <= 1'd0;
      else if (((! \arg0_2_1Dcon_main1_3I#_1_argbuf_r ) && (! \arg0_2_1Dcon_main1_3I#_bufchan_buf [0])))
        \arg0_2_1Dcon_main1_3I#_bufchan_buf  <= \arg0_2_1Dcon_main1_3I#_bufchan_d ;
  
  /* const (Ty Int#,
       Lit 2) : (arg0_2_1Dcon_main1_3I#_1_argbuf,Go) > (arg0_2_1Dcon_main1_3I#_1_argbuf_2,Int#) */
  assign \arg0_2_1Dcon_main1_3I#_1_argbuf_2_d  = {32'd2,
                                                  \arg0_2_1Dcon_main1_3I#_1_argbuf_d [0]};
  assign \arg0_2_1Dcon_main1_3I#_1_argbuf_r  = \arg0_2_1Dcon_main1_3I#_1_argbuf_2_r ;
  
  /* mux (Ty Int,
     Ty Int) : (arg0_2_1Dcon_main1_4,Int) [(es_0_2_1I#,Int)] > (es_0_2_1I#_mux,Int) */
  assign \es_0_2_1I#_mux_d  = {\es_0_2_1I#_d [32:1],
                               (arg0_2_1Dcon_main1_4_d[0] && \es_0_2_1I#_d [0])};
  assign \es_0_2_1I#_r  = (\es_0_2_1I#_mux_r  && (arg0_2_1Dcon_main1_4_d[0] && \es_0_2_1I#_d [0]));
  assign arg0_2_1Dcon_main1_4_r = (\es_0_2_1I#_mux_r  && (arg0_2_1Dcon_main1_4_d[0] && \es_0_2_1I#_d [0]));
  
  /* demux (Ty MyDTInt_Int,
       Ty Go) : (arg0_2_2,MyDTInt_Int) (applyfnInt_Int_5TupGo___MyDTInt_Int___Intgo_10,Go) > [(arg0_2_2Dcon_main1,Go)] */
  assign arg0_2_2Dcon_main1_d = (arg0_2_2_d[0] && applyfnInt_Int_5TupGo___MyDTInt_Int___Intgo_10_d[0]);
  assign applyfnInt_Int_5TupGo___MyDTInt_Int___Intgo_10_r = (arg0_2_2Dcon_main1_r && (arg0_2_2_d[0] && applyfnInt_Int_5TupGo___MyDTInt_Int___Intgo_10_d[0]));
  assign arg0_2_2_r = (arg0_2_2Dcon_main1_r && (arg0_2_2_d[0] && applyfnInt_Int_5TupGo___MyDTInt_Int___Intgo_10_d[0]));
  
  /* mux (Ty MyDTInt_Int,
     Ty Int) : (arg0_2_3,MyDTInt_Int) [(es_0_2_1I#_mux,Int)] > (es_0_2_1I#_mux_mux,Int) */
  assign \es_0_2_1I#_mux_mux_d  = {\es_0_2_1I#_mux_d [32:1],
                                   (arg0_2_3_d[0] && \es_0_2_1I#_mux_d [0])};
  assign \es_0_2_1I#_mux_r  = (\es_0_2_1I#_mux_mux_r  && (arg0_2_3_d[0] && \es_0_2_1I#_mux_d [0]));
  assign arg0_2_3_r = (\es_0_2_1I#_mux_mux_r  && (arg0_2_3_d[0] && \es_0_2_1I#_mux_d [0]));
  
  /* mux (Ty MyDTInt_Bool,
     Ty MyBool) : (arg0_3,MyDTInt_Bool) [(lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux,MyBool)] > (lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux,MyBool) */
  assign lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_d = {lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_d[1:1],
                                                                                 (arg0_3_d[0] && lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_d[0])};
  assign lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_r = (lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_r && (arg0_3_d[0] && lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_d[0]));
  assign arg0_3_r = (lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_r && (arg0_3_d[0] && lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_d[0]));
  
  /* demux (Ty MyDTInt_Int_Int,
       Ty Int) : (arg0_4_1,MyDTInt_Int_Int) (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg1_2,Int) > [(arg0_4_1Dcon_$fNumInt_$c*,Int)] */
  assign \arg0_4_1Dcon_$fNumInt_$ctimes_d  = {applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg1_2_d[32:1],
                                              (arg0_4_1_d[0] && applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg1_2_d[0])};
  assign applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg1_2_r = (\arg0_4_1Dcon_$fNumInt_$ctimes_r  && (arg0_4_1_d[0] && applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg1_2_d[0]));
  assign arg0_4_1_r = (\arg0_4_1Dcon_$fNumInt_$ctimes_r  && (arg0_4_1_d[0] && applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg1_2_d[0]));
  
  /* demux (Ty MyDTInt_Int_Int,
       Ty Int) : (arg0_4_2,MyDTInt_Int_Int) (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg2,Int) > [(arg0_4_2Dcon_$fNumInt_$c*,Int)] */
  assign \arg0_4_2Dcon_$fNumInt_$ctimes_d  = {applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg2_d[32:1],
                                              (arg0_4_2_d[0] && applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg2_d[0])};
  assign applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg2_r = (\arg0_4_2Dcon_$fNumInt_$ctimes_r  && (arg0_4_2_d[0] && applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg2_d[0]));
  assign arg0_4_2_r = (\arg0_4_2Dcon_$fNumInt_$ctimes_r  && (arg0_4_2_d[0] && applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg2_d[0]));
  
  /* fork (Ty Int) : (arg0_4_2Dcon_$fNumInt_$c*,Int) > [(arg0_4_2Dcon_$fNumInt_$c*_1,Int),
                                                   (arg0_4_2Dcon_$fNumInt_$c*_2,Int),
                                                   (arg0_4_2Dcon_$fNumInt_$c*_3,Int),
                                                   (arg0_4_2Dcon_$fNumInt_$c*_4,Int)] */
  logic [3:0] \arg0_4_2Dcon_$fNumInt_$ctimes_emitted ;
  logic [3:0] \arg0_4_2Dcon_$fNumInt_$ctimes_done ;
  assign \arg0_4_2Dcon_$fNumInt_$ctimes_1_d  = {\arg0_4_2Dcon_$fNumInt_$ctimes_d [32:1],
                                                (\arg0_4_2Dcon_$fNumInt_$ctimes_d [0] && (! \arg0_4_2Dcon_$fNumInt_$ctimes_emitted [0]))};
  assign \arg0_4_2Dcon_$fNumInt_$ctimes_2_d  = {\arg0_4_2Dcon_$fNumInt_$ctimes_d [32:1],
                                                (\arg0_4_2Dcon_$fNumInt_$ctimes_d [0] && (! \arg0_4_2Dcon_$fNumInt_$ctimes_emitted [1]))};
  assign \arg0_4_2Dcon_$fNumInt_$ctimes_3_d  = {\arg0_4_2Dcon_$fNumInt_$ctimes_d [32:1],
                                                (\arg0_4_2Dcon_$fNumInt_$ctimes_d [0] && (! \arg0_4_2Dcon_$fNumInt_$ctimes_emitted [2]))};
  assign \arg0_4_2Dcon_$fNumInt_$ctimes_4_d  = {\arg0_4_2Dcon_$fNumInt_$ctimes_d [32:1],
                                                (\arg0_4_2Dcon_$fNumInt_$ctimes_d [0] && (! \arg0_4_2Dcon_$fNumInt_$ctimes_emitted [3]))};
  assign \arg0_4_2Dcon_$fNumInt_$ctimes_done  = (\arg0_4_2Dcon_$fNumInt_$ctimes_emitted  | ({\arg0_4_2Dcon_$fNumInt_$ctimes_4_d [0],
                                                                                             \arg0_4_2Dcon_$fNumInt_$ctimes_3_d [0],
                                                                                             \arg0_4_2Dcon_$fNumInt_$ctimes_2_d [0],
                                                                                             \arg0_4_2Dcon_$fNumInt_$ctimes_1_d [0]} & {\arg0_4_2Dcon_$fNumInt_$ctimes_4_r ,
                                                                                                                                        \arg0_4_2Dcon_$fNumInt_$ctimes_3_r ,
                                                                                                                                        \arg0_4_2Dcon_$fNumInt_$ctimes_2_r ,
                                                                                                                                        \arg0_4_2Dcon_$fNumInt_$ctimes_1_r }));
  assign \arg0_4_2Dcon_$fNumInt_$ctimes_r  = (& \arg0_4_2Dcon_$fNumInt_$ctimes_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \arg0_4_2Dcon_$fNumInt_$ctimes_emitted  <= 4'd0;
    else
      \arg0_4_2Dcon_$fNumInt_$ctimes_emitted  <= (\arg0_4_2Dcon_$fNumInt_$ctimes_r  ? 4'd0 :
                                                  \arg0_4_2Dcon_$fNumInt_$ctimes_done );
  
  /* destruct (Ty Int,
          Dcon I#) : (arg0_4_2Dcon_$fNumInt_$c*_1I#,Int) > [(xa1m0_destruct,Int#)] */
  assign xa1m0_destruct_d = {\arg0_4_2Dcon_$fNumInt_$ctimes_1I#_d [32:1],
                             \arg0_4_2Dcon_$fNumInt_$ctimes_1I#_d [0]};
  assign \arg0_4_2Dcon_$fNumInt_$ctimes_1I#_r  = xa1m0_destruct_r;
  
  /* demux (Ty Int,
       Ty Int) : (arg0_4_2Dcon_$fNumInt_$c*_2,Int) (arg0_4_2Dcon_$fNumInt_$c*_1,Int) > [(arg0_4_2Dcon_$fNumInt_$c*_1I#,Int)] */
  assign \arg0_4_2Dcon_$fNumInt_$ctimes_1I#_d  = {\arg0_4_2Dcon_$fNumInt_$ctimes_1_d [32:1],
                                                  (\arg0_4_2Dcon_$fNumInt_$ctimes_2_d [0] && \arg0_4_2Dcon_$fNumInt_$ctimes_1_d [0])};
  assign \arg0_4_2Dcon_$fNumInt_$ctimes_1_r  = (\arg0_4_2Dcon_$fNumInt_$ctimes_1I#_r  && (\arg0_4_2Dcon_$fNumInt_$ctimes_2_d [0] && \arg0_4_2Dcon_$fNumInt_$ctimes_1_d [0]));
  assign \arg0_4_2Dcon_$fNumInt_$ctimes_2_r  = (\arg0_4_2Dcon_$fNumInt_$ctimes_1I#_r  && (\arg0_4_2Dcon_$fNumInt_$ctimes_2_d [0] && \arg0_4_2Dcon_$fNumInt_$ctimes_1_d [0]));
  
  /* demux (Ty Int,
       Ty Int) : (arg0_4_2Dcon_$fNumInt_$c*_3,Int) (arg0_4_1Dcon_$fNumInt_$c*,Int) > [(arg0_4_2Dcon_$fNumInt_$c*_3I#,Int)] */
  assign \arg0_4_2Dcon_$fNumInt_$ctimes_3I#_d  = {\arg0_4_1Dcon_$fNumInt_$ctimes_d [32:1],
                                                  (\arg0_4_2Dcon_$fNumInt_$ctimes_3_d [0] && \arg0_4_1Dcon_$fNumInt_$ctimes_d [0])};
  assign \arg0_4_1Dcon_$fNumInt_$ctimes_r  = (\arg0_4_2Dcon_$fNumInt_$ctimes_3I#_r  && (\arg0_4_2Dcon_$fNumInt_$ctimes_3_d [0] && \arg0_4_1Dcon_$fNumInt_$ctimes_d [0]));
  assign \arg0_4_2Dcon_$fNumInt_$ctimes_3_r  = (\arg0_4_2Dcon_$fNumInt_$ctimes_3I#_r  && (\arg0_4_2Dcon_$fNumInt_$ctimes_3_d [0] && \arg0_4_1Dcon_$fNumInt_$ctimes_d [0]));
  
  /* fork (Ty Int) : (arg0_4_2Dcon_$fNumInt_$c*_3I#,Int) > [(arg0_4_2Dcon_$fNumInt_$c*_3I#_1,Int),
                                                       (arg0_4_2Dcon_$fNumInt_$c*_3I#_2,Int),
                                                       (arg0_4_2Dcon_$fNumInt_$c*_3I#_3,Int),
                                                       (arg0_4_2Dcon_$fNumInt_$c*_3I#_4,Int)] */
  logic [3:0] \arg0_4_2Dcon_$fNumInt_$ctimes_3I#_emitted ;
  logic [3:0] \arg0_4_2Dcon_$fNumInt_$ctimes_3I#_done ;
  assign \arg0_4_2Dcon_$fNumInt_$ctimes_3I#_1_d  = {\arg0_4_2Dcon_$fNumInt_$ctimes_3I#_d [32:1],
                                                    (\arg0_4_2Dcon_$fNumInt_$ctimes_3I#_d [0] && (! \arg0_4_2Dcon_$fNumInt_$ctimes_3I#_emitted [0]))};
  assign \arg0_4_2Dcon_$fNumInt_$ctimes_3I#_2_d  = {\arg0_4_2Dcon_$fNumInt_$ctimes_3I#_d [32:1],
                                                    (\arg0_4_2Dcon_$fNumInt_$ctimes_3I#_d [0] && (! \arg0_4_2Dcon_$fNumInt_$ctimes_3I#_emitted [1]))};
  assign \arg0_4_2Dcon_$fNumInt_$ctimes_3I#_3_d  = {\arg0_4_2Dcon_$fNumInt_$ctimes_3I#_d [32:1],
                                                    (\arg0_4_2Dcon_$fNumInt_$ctimes_3I#_d [0] && (! \arg0_4_2Dcon_$fNumInt_$ctimes_3I#_emitted [2]))};
  assign \arg0_4_2Dcon_$fNumInt_$ctimes_3I#_4_d  = {\arg0_4_2Dcon_$fNumInt_$ctimes_3I#_d [32:1],
                                                    (\arg0_4_2Dcon_$fNumInt_$ctimes_3I#_d [0] && (! \arg0_4_2Dcon_$fNumInt_$ctimes_3I#_emitted [3]))};
  assign \arg0_4_2Dcon_$fNumInt_$ctimes_3I#_done  = (\arg0_4_2Dcon_$fNumInt_$ctimes_3I#_emitted  | ({\arg0_4_2Dcon_$fNumInt_$ctimes_3I#_4_d [0],
                                                                                                     \arg0_4_2Dcon_$fNumInt_$ctimes_3I#_3_d [0],
                                                                                                     \arg0_4_2Dcon_$fNumInt_$ctimes_3I#_2_d [0],
                                                                                                     \arg0_4_2Dcon_$fNumInt_$ctimes_3I#_1_d [0]} & {\arg0_4_2Dcon_$fNumInt_$ctimes_3I#_4_r ,
                                                                                                                                                    \arg0_4_2Dcon_$fNumInt_$ctimes_3I#_3_r ,
                                                                                                                                                    \arg0_4_2Dcon_$fNumInt_$ctimes_3I#_2_r ,
                                                                                                                                                    \arg0_4_2Dcon_$fNumInt_$ctimes_3I#_1_r }));
  assign \arg0_4_2Dcon_$fNumInt_$ctimes_3I#_r  = (& \arg0_4_2Dcon_$fNumInt_$ctimes_3I#_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \arg0_4_2Dcon_$fNumInt_$ctimes_3I#_emitted  <= 4'd0;
    else
      \arg0_4_2Dcon_$fNumInt_$ctimes_3I#_emitted  <= (\arg0_4_2Dcon_$fNumInt_$ctimes_3I#_r  ? 4'd0 :
                                                      \arg0_4_2Dcon_$fNumInt_$ctimes_3I#_done );
  
  /* destruct (Ty Int,
          Dcon I#) : (arg0_4_2Dcon_$fNumInt_$c*_3I#_1I#,Int) > [(ya1m1_destruct,Int#)] */
  assign ya1m1_destruct_d = {\arg0_4_2Dcon_$fNumInt_$ctimes_3I#_1I#_d [32:1],
                             \arg0_4_2Dcon_$fNumInt_$ctimes_3I#_1I#_d [0]};
  assign \arg0_4_2Dcon_$fNumInt_$ctimes_3I#_1I#_r  = ya1m1_destruct_r;
  
  /* demux (Ty Int,
       Ty Int) : (arg0_4_2Dcon_$fNumInt_$c*_3I#_2,Int) (arg0_4_2Dcon_$fNumInt_$c*_3I#_1,Int) > [(arg0_4_2Dcon_$fNumInt_$c*_3I#_1I#,Int)] */
  assign \arg0_4_2Dcon_$fNumInt_$ctimes_3I#_1I#_d  = {\arg0_4_2Dcon_$fNumInt_$ctimes_3I#_1_d [32:1],
                                                      (\arg0_4_2Dcon_$fNumInt_$ctimes_3I#_2_d [0] && \arg0_4_2Dcon_$fNumInt_$ctimes_3I#_1_d [0])};
  assign \arg0_4_2Dcon_$fNumInt_$ctimes_3I#_1_r  = (\arg0_4_2Dcon_$fNumInt_$ctimes_3I#_1I#_r  && (\arg0_4_2Dcon_$fNumInt_$ctimes_3I#_2_d [0] && \arg0_4_2Dcon_$fNumInt_$ctimes_3I#_1_d [0]));
  assign \arg0_4_2Dcon_$fNumInt_$ctimes_3I#_2_r  = (\arg0_4_2Dcon_$fNumInt_$ctimes_3I#_1I#_r  && (\arg0_4_2Dcon_$fNumInt_$ctimes_3I#_2_d [0] && \arg0_4_2Dcon_$fNumInt_$ctimes_3I#_1_d [0]));
  
  /* demux (Ty Int,
       Ty Int#) : (arg0_4_2Dcon_$fNumInt_$c*_3I#_3,Int) (xa1m0_destruct,Int#) > [(arg0_4_2Dcon_$fNumInt_$c*_3I#_3I#,Int#)] */
  assign \arg0_4_2Dcon_$fNumInt_$ctimes_3I#_3I#_d  = {xa1m0_destruct_d[32:1],
                                                      (\arg0_4_2Dcon_$fNumInt_$ctimes_3I#_3_d [0] && xa1m0_destruct_d[0])};
  assign xa1m0_destruct_r = (\arg0_4_2Dcon_$fNumInt_$ctimes_3I#_3I#_r  && (\arg0_4_2Dcon_$fNumInt_$ctimes_3I#_3_d [0] && xa1m0_destruct_d[0]));
  assign \arg0_4_2Dcon_$fNumInt_$ctimes_3I#_3_r  = (\arg0_4_2Dcon_$fNumInt_$ctimes_3I#_3I#_r  && (\arg0_4_2Dcon_$fNumInt_$ctimes_3I#_3_d [0] && xa1m0_destruct_d[0]));
  
  /* op_mul (Ty Int#) : (arg0_4_2Dcon_$fNumInt_$c*_3I#_3I#,Int#) (ya1m1_destruct,Int#) > (arg0_4_2Dcon_$fNumInt_$c*_3I#_3I#_1ya1m1_1_Mul32,Int#) */
  assign \arg0_4_2Dcon_$fNumInt_$ctimes_3I#_3I#_1ya1m1_1_Mul32_d  = {(\arg0_4_2Dcon_$fNumInt_$ctimes_3I#_3I#_d [32:1] * ya1m1_destruct_d[32:1]),
                                                                     (\arg0_4_2Dcon_$fNumInt_$ctimes_3I#_3I#_d [0] && ya1m1_destruct_d[0])};
  assign {\arg0_4_2Dcon_$fNumInt_$ctimes_3I#_3I#_r ,
          ya1m1_destruct_r} = {2 {(\arg0_4_2Dcon_$fNumInt_$ctimes_3I#_3I#_1ya1m1_1_Mul32_r  && \arg0_4_2Dcon_$fNumInt_$ctimes_3I#_3I#_1ya1m1_1_Mul32_d [0])}};
  
  /* dcon (Ty Int,
      Dcon I#) : [(arg0_4_2Dcon_$fNumInt_$c*_3I#_3I#_1ya1m1_1_Mul32,Int#)] > (es_0_3_1I#,Int) */
  assign \es_0_3_1I#_d  = \I#_dc ((& {\arg0_4_2Dcon_$fNumInt_$ctimes_3I#_3I#_1ya1m1_1_Mul32_d [0]}), \arg0_4_2Dcon_$fNumInt_$ctimes_3I#_3I#_1ya1m1_1_Mul32_d );
  assign {\arg0_4_2Dcon_$fNumInt_$ctimes_3I#_3I#_1ya1m1_1_Mul32_r } = {1 {(\es_0_3_1I#_r  && \es_0_3_1I#_d [0])}};
  
  /* mux (Ty Int,
     Ty Int) : (arg0_4_2Dcon_$fNumInt_$c*_3I#_4,Int) [(es_0_3_1I#,Int)] > (es_0_3_1I#_mux,Int) */
  assign \es_0_3_1I#_mux_d  = {\es_0_3_1I#_d [32:1],
                               (\arg0_4_2Dcon_$fNumInt_$ctimes_3I#_4_d [0] && \es_0_3_1I#_d [0])};
  assign \es_0_3_1I#_r  = (\es_0_3_1I#_mux_r  && (\arg0_4_2Dcon_$fNumInt_$ctimes_3I#_4_d [0] && \es_0_3_1I#_d [0]));
  assign \arg0_4_2Dcon_$fNumInt_$ctimes_3I#_4_r  = (\es_0_3_1I#_mux_r  && (\arg0_4_2Dcon_$fNumInt_$ctimes_3I#_4_d [0] && \es_0_3_1I#_d [0]));
  
  /* mux (Ty Int,
     Ty Int) : (arg0_4_2Dcon_$fNumInt_$c*_4,Int) [(es_0_3_1I#_mux,Int)] > (es_0_3_1I#_mux_mux,Int) */
  assign \es_0_3_1I#_mux_mux_d  = {\es_0_3_1I#_mux_d [32:1],
                                   (\arg0_4_2Dcon_$fNumInt_$ctimes_4_d [0] && \es_0_3_1I#_mux_d [0])};
  assign \es_0_3_1I#_mux_r  = (\es_0_3_1I#_mux_mux_r  && (\arg0_4_2Dcon_$fNumInt_$ctimes_4_d [0] && \es_0_3_1I#_mux_d [0]));
  assign \arg0_4_2Dcon_$fNumInt_$ctimes_4_r  = (\es_0_3_1I#_mux_mux_r  && (\arg0_4_2Dcon_$fNumInt_$ctimes_4_d [0] && \es_0_3_1I#_mux_d [0]));
  
  /* mux (Ty MyDTInt_Int_Int,
     Ty Int) : (arg0_4_3,MyDTInt_Int_Int) [(es_0_3_1I#_mux_mux,Int)] > (es_0_3_1I#_mux_mux_mux,Int) */
  assign \es_0_3_1I#_mux_mux_mux_d  = {\es_0_3_1I#_mux_mux_d [32:1],
                                       (arg0_4_3_d[0] && \es_0_3_1I#_mux_mux_d [0])};
  assign \es_0_3_1I#_mux_mux_r  = (\es_0_3_1I#_mux_mux_mux_r  && (arg0_4_3_d[0] && \es_0_3_1I#_mux_mux_d [0]));
  assign arg0_4_3_r = (\es_0_3_1I#_mux_mux_mux_r  && (arg0_4_3_d[0] && \es_0_3_1I#_mux_mux_d [0]));
  
  /* destruct (Ty TupGo___Bool,
          Dcon TupGo___Bool) : (boolConvert_1TupGo___Bool_1,TupGo___Bool) > [(boolConvert_1TupGo___Boolgo_1,Go),
                                                                             (boolConvert_1TupGo___Boolbool,Bool)] */
  logic [1:0] boolConvert_1TupGo___Bool_1_emitted;
  logic [1:0] boolConvert_1TupGo___Bool_1_done;
  assign boolConvert_1TupGo___Boolgo_1_d = (boolConvert_1TupGo___Bool_1_d[0] && (! boolConvert_1TupGo___Bool_1_emitted[0]));
  assign boolConvert_1TupGo___Boolbool_d = {boolConvert_1TupGo___Bool_1_d[1:1],
                                            (boolConvert_1TupGo___Bool_1_d[0] && (! boolConvert_1TupGo___Bool_1_emitted[1]))};
  assign boolConvert_1TupGo___Bool_1_done = (boolConvert_1TupGo___Bool_1_emitted | ({boolConvert_1TupGo___Boolbool_d[0],
                                                                                     boolConvert_1TupGo___Boolgo_1_d[0]} & {boolConvert_1TupGo___Boolbool_r,
                                                                                                                            boolConvert_1TupGo___Boolgo_1_r}));
  assign boolConvert_1TupGo___Bool_1_r = (& boolConvert_1TupGo___Bool_1_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) boolConvert_1TupGo___Bool_1_emitted <= 2'd0;
    else
      boolConvert_1TupGo___Bool_1_emitted <= (boolConvert_1TupGo___Bool_1_r ? 2'd0 :
                                              boolConvert_1TupGo___Bool_1_done);
  
  /* fork (Ty Bool) : (boolConvert_1TupGo___Boolbool,Bool) > [(bool_1,Bool),
                                                         (bool_2,Bool)] */
  logic [1:0] boolConvert_1TupGo___Boolbool_emitted;
  logic [1:0] boolConvert_1TupGo___Boolbool_done;
  assign bool_1_d = {boolConvert_1TupGo___Boolbool_d[1:1],
                     (boolConvert_1TupGo___Boolbool_d[0] && (! boolConvert_1TupGo___Boolbool_emitted[0]))};
  assign bool_2_d = {boolConvert_1TupGo___Boolbool_d[1:1],
                     (boolConvert_1TupGo___Boolbool_d[0] && (! boolConvert_1TupGo___Boolbool_emitted[1]))};
  assign boolConvert_1TupGo___Boolbool_done = (boolConvert_1TupGo___Boolbool_emitted | ({bool_2_d[0],
                                                                                         bool_1_d[0]} & {bool_2_r,
                                                                                                         bool_1_r}));
  assign boolConvert_1TupGo___Boolbool_r = (& boolConvert_1TupGo___Boolbool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) boolConvert_1TupGo___Boolbool_emitted <= 2'd0;
    else
      boolConvert_1TupGo___Boolbool_emitted <= (boolConvert_1TupGo___Boolbool_r ? 2'd0 :
                                                boolConvert_1TupGo___Boolbool_done);
  
  /* fork (Ty MyBool) : (boolConvert_1_resbuf,MyBool) > [(lizzieLet3_1,MyBool),
                                                    (lizzieLet3_2,MyBool)] */
  logic [1:0] boolConvert_1_resbuf_emitted;
  logic [1:0] boolConvert_1_resbuf_done;
  assign lizzieLet3_1_d = {boolConvert_1_resbuf_d[1:1],
                           (boolConvert_1_resbuf_d[0] && (! boolConvert_1_resbuf_emitted[0]))};
  assign lizzieLet3_2_d = {boolConvert_1_resbuf_d[1:1],
                           (boolConvert_1_resbuf_d[0] && (! boolConvert_1_resbuf_emitted[1]))};
  assign boolConvert_1_resbuf_done = (boolConvert_1_resbuf_emitted | ({lizzieLet3_2_d[0],
                                                                       lizzieLet3_1_d[0]} & {lizzieLet3_2_r,
                                                                                             lizzieLet3_1_r}));
  assign boolConvert_1_resbuf_r = (& boolConvert_1_resbuf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) boolConvert_1_resbuf_emitted <= 2'd0;
    else
      boolConvert_1_resbuf_emitted <= (boolConvert_1_resbuf_r ? 2'd0 :
                                       boolConvert_1_resbuf_done);
  
  /* demux (Ty Bool,
       Ty Go) : (bool_1,Bool) (boolConvert_1TupGo___Boolgo_1,Go) > [(bool_1False,Go),
                                                                    (bool_1True,Go)] */
  logic [1:0] boolConvert_1TupGo___Boolgo_1_onehotd;
  always_comb
    if ((bool_1_d[0] && boolConvert_1TupGo___Boolgo_1_d[0]))
      unique case (bool_1_d[1:1])
        1'd0: boolConvert_1TupGo___Boolgo_1_onehotd = 2'd1;
        1'd1: boolConvert_1TupGo___Boolgo_1_onehotd = 2'd2;
        default: boolConvert_1TupGo___Boolgo_1_onehotd = 2'd0;
      endcase
    else boolConvert_1TupGo___Boolgo_1_onehotd = 2'd0;
  assign bool_1False_d = boolConvert_1TupGo___Boolgo_1_onehotd[0];
  assign bool_1True_d = boolConvert_1TupGo___Boolgo_1_onehotd[1];
  assign boolConvert_1TupGo___Boolgo_1_r = (| (boolConvert_1TupGo___Boolgo_1_onehotd & {bool_1True_r,
                                                                                        bool_1False_r}));
  assign bool_1_r = boolConvert_1TupGo___Boolgo_1_r;
  
  /* dcon (Ty MyBool,
      Dcon MyFalse) : [(bool_1False,Go)] > (bool_1False_1MyFalse,MyBool) */
  assign bool_1False_1MyFalse_d = MyFalse_dc((& {bool_1False_d[0]}), bool_1False_d);
  assign {bool_1False_r} = {1 {(bool_1False_1MyFalse_r && bool_1False_1MyFalse_d[0])}};
  
  /* buf (Ty MyBool) : (bool_1False_1MyFalsebool_1True_1MyTrue_mux,MyBool) > (boolConvert_1_resbuf,MyBool) */
  MyBool_t bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_d;
  logic bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_r;
  assign bool_1False_1MyFalsebool_1True_1MyTrue_mux_r = ((! bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_d[0]) || bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_d <= {1'd0,
                                                               1'd0};
    else
      if (bool_1False_1MyFalsebool_1True_1MyTrue_mux_r)
        bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_d <= bool_1False_1MyFalsebool_1True_1MyTrue_mux_d;
  MyBool_t bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_buf;
  assign bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_r = (! bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_buf[0]);
  assign boolConvert_1_resbuf_d = (bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_buf[0] ? bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_buf :
                                   bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_buf <= {1'd0,
                                                                 1'd0};
    else
      if ((boolConvert_1_resbuf_r && bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_buf[0]))
        bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_buf <= {1'd0,
                                                                   1'd0};
      else if (((! boolConvert_1_resbuf_r) && (! bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_buf[0])))
        bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_buf <= bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_d;
  
  /* dcon (Ty MyBool,
      Dcon MyTrue) : [(bool_1True,Go)] > (bool_1True_1MyTrue,MyBool) */
  assign bool_1True_1MyTrue_d = MyTrue_dc((& {bool_1True_d[0]}), bool_1True_d);
  assign {bool_1True_r} = {1 {(bool_1True_1MyTrue_r && bool_1True_1MyTrue_d[0])}};
  
  /* mux (Ty Bool,
     Ty MyBool) : (bool_2,Bool) [(bool_1False_1MyFalse,MyBool),
                                 (bool_1True_1MyTrue,MyBool)] > (bool_1False_1MyFalsebool_1True_1MyTrue_mux,MyBool) */
  logic [1:0] bool_1False_1MyFalsebool_1True_1MyTrue_mux_mux;
  logic [1:0] bool_1False_1MyFalsebool_1True_1MyTrue_mux_onehot;
  always_comb
    unique case (bool_2_d[1:1])
      1'd0:
        {bool_1False_1MyFalsebool_1True_1MyTrue_mux_onehot,
         bool_1False_1MyFalsebool_1True_1MyTrue_mux_mux} = {2'd1,
                                                            bool_1False_1MyFalse_d};
      1'd1:
        {bool_1False_1MyFalsebool_1True_1MyTrue_mux_onehot,
         bool_1False_1MyFalsebool_1True_1MyTrue_mux_mux} = {2'd2,
                                                            bool_1True_1MyTrue_d};
      default:
        {bool_1False_1MyFalsebool_1True_1MyTrue_mux_onehot,
         bool_1False_1MyFalsebool_1True_1MyTrue_mux_mux} = {2'd0,
                                                            {1'd0, 1'd0}};
    endcase
  assign bool_1False_1MyFalsebool_1True_1MyTrue_mux_d = {bool_1False_1MyFalsebool_1True_1MyTrue_mux_mux[1:1],
                                                         (bool_1False_1MyFalsebool_1True_1MyTrue_mux_mux[0] && bool_2_d[0])};
  assign bool_2_r = (bool_1False_1MyFalsebool_1True_1MyTrue_mux_d[0] && bool_1False_1MyFalsebool_1True_1MyTrue_mux_r);
  assign {bool_1True_1MyTrue_r,
          bool_1False_1MyFalse_r} = (bool_2_r ? bool_1False_1MyFalsebool_1True_1MyTrue_mux_onehot :
                                     2'd0);
  
  /* destruct (Ty TupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int,
          Dcon TupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int) : (call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1,TupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int) > [(call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intgo_11,Go),
                                                                                                                                                                                       (call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intwsvt_1,Pointer_QTree_Int),
                                                                                                                                                                                       (call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intsc_0,Pointer_CT$wnnz_Int)] */
  logic [2:0] call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_emitted;
  logic [2:0] call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_done;
  assign call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intgo_11_d = (call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_d[0] && (! call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_emitted[0]));
  assign call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intwsvt_1_d = {call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_d[16:1],
                                                                                  (call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_d[0] && (! call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_emitted[1]))};
  assign call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intsc_0_d = {call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_d[32:17],
                                                                                (call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_d[0] && (! call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_emitted[2]))};
  assign call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_done = (call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_emitted | ({call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intsc_0_d[0],
                                                                                                                                                             call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intwsvt_1_d[0],
                                                                                                                                                             call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intgo_11_d[0]} & {call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intsc_0_r,
                                                                                                                                                                                                                                         call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intwsvt_1_r,
                                                                                                                                                                                                                                         call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intgo_11_r}));
  assign call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_r = (& call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_emitted <= 3'd0;
    else
      call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_emitted <= (call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_r ? 3'd0 :
                                                                                  call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_done);
  
  /* rbuf (Ty Go) : (call_$wnnz_Int_goConst,Go) > (call_$wnnz_Int_initBufi,Go) */
  Go_t call_$wnnz_Int_goConst_buf;
  assign call_$wnnz_Int_goConst_r = (! call_$wnnz_Int_goConst_buf[0]);
  assign call_$wnnz_Int_initBufi_d = (call_$wnnz_Int_goConst_buf[0] ? call_$wnnz_Int_goConst_buf :
                                      call_$wnnz_Int_goConst_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_$wnnz_Int_goConst_buf <= 1'd0;
    else
      if ((call_$wnnz_Int_initBufi_r && call_$wnnz_Int_goConst_buf[0]))
        call_$wnnz_Int_goConst_buf <= 1'd0;
      else if (((! call_$wnnz_Int_initBufi_r) && (! call_$wnnz_Int_goConst_buf[0])))
        call_$wnnz_Int_goConst_buf <= call_$wnnz_Int_goConst_d;
  
  /* mergectrl (Ty C5,Ty Go) : [(call_$wnnz_Int_goMux1,Go),
                           (lizzieLet25_3Lcall_$wnnz_Int3_1_argbuf,Go),
                           (lizzieLet25_3Lcall_$wnnz_Int2_1_argbuf,Go),
                           (lizzieLet25_3Lcall_$wnnz_Int1_1_argbuf,Go),
                           (lizzieLet4_3QNode_Int_1_argbuf,Go)] > (go_11_goMux_choice,C5) (go_11_goMux_data,Go) */
  logic [4:0] call_$wnnz_Int_goMux1_select_d;
  assign call_$wnnz_Int_goMux1_select_d = ((| call_$wnnz_Int_goMux1_select_q) ? call_$wnnz_Int_goMux1_select_q :
                                           (call_$wnnz_Int_goMux1_d[0] ? 5'd1 :
                                            (lizzieLet25_3Lcall_$wnnz_Int3_1_argbuf_d[0] ? 5'd2 :
                                             (lizzieLet25_3Lcall_$wnnz_Int2_1_argbuf_d[0] ? 5'd4 :
                                              (lizzieLet25_3Lcall_$wnnz_Int1_1_argbuf_d[0] ? 5'd8 :
                                               (lizzieLet4_3QNode_Int_1_argbuf_d[0] ? 5'd16 :
                                                5'd0))))));
  logic [4:0] call_$wnnz_Int_goMux1_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_$wnnz_Int_goMux1_select_q <= 5'd0;
    else
      call_$wnnz_Int_goMux1_select_q <= (call_$wnnz_Int_goMux1_done ? 5'd0 :
                                         call_$wnnz_Int_goMux1_select_d);
  logic [1:0] call_$wnnz_Int_goMux1_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_$wnnz_Int_goMux1_emit_q <= 2'd0;
    else
      call_$wnnz_Int_goMux1_emit_q <= (call_$wnnz_Int_goMux1_done ? 2'd0 :
                                       call_$wnnz_Int_goMux1_emit_d);
  logic [1:0] call_$wnnz_Int_goMux1_emit_d;
  assign call_$wnnz_Int_goMux1_emit_d = (call_$wnnz_Int_goMux1_emit_q | ({go_11_goMux_choice_d[0],
                                                                          go_11_goMux_data_d[0]} & {go_11_goMux_choice_r,
                                                                                                    go_11_goMux_data_r}));
  logic call_$wnnz_Int_goMux1_done;
  assign call_$wnnz_Int_goMux1_done = (& call_$wnnz_Int_goMux1_emit_d);
  assign {lizzieLet4_3QNode_Int_1_argbuf_r,
          lizzieLet25_3Lcall_$wnnz_Int1_1_argbuf_r,
          lizzieLet25_3Lcall_$wnnz_Int2_1_argbuf_r,
          lizzieLet25_3Lcall_$wnnz_Int3_1_argbuf_r,
          call_$wnnz_Int_goMux1_r} = (call_$wnnz_Int_goMux1_done ? call_$wnnz_Int_goMux1_select_d :
                                      5'd0);
  assign go_11_goMux_data_d = ((call_$wnnz_Int_goMux1_select_d[0] && (! call_$wnnz_Int_goMux1_emit_q[0])) ? call_$wnnz_Int_goMux1_d :
                               ((call_$wnnz_Int_goMux1_select_d[1] && (! call_$wnnz_Int_goMux1_emit_q[0])) ? lizzieLet25_3Lcall_$wnnz_Int3_1_argbuf_d :
                                ((call_$wnnz_Int_goMux1_select_d[2] && (! call_$wnnz_Int_goMux1_emit_q[0])) ? lizzieLet25_3Lcall_$wnnz_Int2_1_argbuf_d :
                                 ((call_$wnnz_Int_goMux1_select_d[3] && (! call_$wnnz_Int_goMux1_emit_q[0])) ? lizzieLet25_3Lcall_$wnnz_Int1_1_argbuf_d :
                                  ((call_$wnnz_Int_goMux1_select_d[4] && (! call_$wnnz_Int_goMux1_emit_q[0])) ? lizzieLet4_3QNode_Int_1_argbuf_d :
                                   1'd0)))));
  assign go_11_goMux_choice_d = ((call_$wnnz_Int_goMux1_select_d[0] && (! call_$wnnz_Int_goMux1_emit_q[1])) ? C1_5_dc(1'd1) :
                                 ((call_$wnnz_Int_goMux1_select_d[1] && (! call_$wnnz_Int_goMux1_emit_q[1])) ? C2_5_dc(1'd1) :
                                  ((call_$wnnz_Int_goMux1_select_d[2] && (! call_$wnnz_Int_goMux1_emit_q[1])) ? C3_5_dc(1'd1) :
                                   ((call_$wnnz_Int_goMux1_select_d[3] && (! call_$wnnz_Int_goMux1_emit_q[1])) ? C4_5_dc(1'd1) :
                                    ((call_$wnnz_Int_goMux1_select_d[4] && (! call_$wnnz_Int_goMux1_emit_q[1])) ? C5_5_dc(1'd1) :
                                     {3'd0, 1'd0})))));
  
  /* fork (Ty Go) : (call_$wnnz_Int_initBuf,Go) > [(call_$wnnz_Int_unlockFork1,Go),
                                              (call_$wnnz_Int_unlockFork2,Go),
                                              (call_$wnnz_Int_unlockFork3,Go)] */
  logic [2:0] call_$wnnz_Int_initBuf_emitted;
  logic [2:0] call_$wnnz_Int_initBuf_done;
  assign call_$wnnz_Int_unlockFork1_d = (call_$wnnz_Int_initBuf_d[0] && (! call_$wnnz_Int_initBuf_emitted[0]));
  assign call_$wnnz_Int_unlockFork2_d = (call_$wnnz_Int_initBuf_d[0] && (! call_$wnnz_Int_initBuf_emitted[1]));
  assign call_$wnnz_Int_unlockFork3_d = (call_$wnnz_Int_initBuf_d[0] && (! call_$wnnz_Int_initBuf_emitted[2]));
  assign call_$wnnz_Int_initBuf_done = (call_$wnnz_Int_initBuf_emitted | ({call_$wnnz_Int_unlockFork3_d[0],
                                                                           call_$wnnz_Int_unlockFork2_d[0],
                                                                           call_$wnnz_Int_unlockFork1_d[0]} & {call_$wnnz_Int_unlockFork3_r,
                                                                                                               call_$wnnz_Int_unlockFork2_r,
                                                                                                               call_$wnnz_Int_unlockFork1_r}));
  assign call_$wnnz_Int_initBuf_r = (& call_$wnnz_Int_initBuf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_$wnnz_Int_initBuf_emitted <= 3'd0;
    else
      call_$wnnz_Int_initBuf_emitted <= (call_$wnnz_Int_initBuf_r ? 3'd0 :
                                         call_$wnnz_Int_initBuf_done);
  
  /* initbuf (Ty Go,
         Dcon Go) : (call_$wnnz_Int_initBufi,Go) > (call_$wnnz_Int_initBuf,Go) */
  assign call_$wnnz_Int_initBufi_r = ((! call_$wnnz_Int_initBuf_d[0]) || call_$wnnz_Int_initBuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_$wnnz_Int_initBuf_d <= Go_dc(1'd1);
    else
      if (call_$wnnz_Int_initBufi_r)
        call_$wnnz_Int_initBuf_d <= call_$wnnz_Int_initBufi_d;
  
  /* mux (Ty Go,
     Ty Go) : (call_$wnnz_Int_unlockFork1,Go) [(call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intgo_11,Go)] > (call_$wnnz_Int_goMux1,Go) */
  assign call_$wnnz_Int_goMux1_d = (call_$wnnz_Int_unlockFork1_d[0] && call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intgo_11_d[0]);
  assign call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intgo_11_r = (call_$wnnz_Int_goMux1_r && (call_$wnnz_Int_unlockFork1_d[0] && call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intgo_11_d[0]));
  assign call_$wnnz_Int_unlockFork1_r = (call_$wnnz_Int_goMux1_r && (call_$wnnz_Int_unlockFork1_d[0] && call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intgo_11_d[0]));
  
  /* mux (Ty Go,
     Ty Pointer_QTree_Int) : (call_$wnnz_Int_unlockFork2,Go) [(call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intwsvt_1,Pointer_QTree_Int)] > (call_$wnnz_Int_goMux2,Pointer_QTree_Int) */
  assign call_$wnnz_Int_goMux2_d = {call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intwsvt_1_d[16:1],
                                    (call_$wnnz_Int_unlockFork2_d[0] && call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intwsvt_1_d[0])};
  assign call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intwsvt_1_r = (call_$wnnz_Int_goMux2_r && (call_$wnnz_Int_unlockFork2_d[0] && call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intwsvt_1_d[0]));
  assign call_$wnnz_Int_unlockFork2_r = (call_$wnnz_Int_goMux2_r && (call_$wnnz_Int_unlockFork2_d[0] && call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intwsvt_1_d[0]));
  
  /* mux (Ty Go,
     Ty Pointer_CT$wnnz_Int) : (call_$wnnz_Int_unlockFork3,Go) [(call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intsc_0,Pointer_CT$wnnz_Int)] > (call_$wnnz_Int_goMux3,Pointer_CT$wnnz_Int) */
  assign call_$wnnz_Int_goMux3_d = {call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intsc_0_d[16:1],
                                    (call_$wnnz_Int_unlockFork3_d[0] && call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intsc_0_d[0])};
  assign call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intsc_0_r = (call_$wnnz_Int_goMux3_r && (call_$wnnz_Int_unlockFork3_d[0] && call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intsc_0_d[0]));
  assign call_$wnnz_Int_unlockFork3_r = (call_$wnnz_Int_goMux3_r && (call_$wnnz_Int_unlockFork3_d[0] && call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intsc_0_d[0]));
  
  /* destruct (Ty TupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Int,
          Dcon TupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Int) : (call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Int_1,TupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Int) > [(call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Intgo_12,Go),
                                                                                                                                                                                                                                                                                                                                                                                                      (call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_IntisZad2,MyDTInt_Bool),
                                                                                                                                                                                                                                                                                                                                                                                                      (call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Intgad3,MyDTInt_Int_Int),
                                                                                                                                                                                                                                                                                                                                                                                                      (call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Intm1ad4,Pointer_QTree_Int),
                                                                                                                                                                                                                                                                                                                                                                                                      (call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Intm2ad5,Pointer_QTree_Int),
                                                                                                                                                                                                                                                                                                                                                                                                      (call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Intsc_0_1,Pointer_CTkron_kron_Int_Int_Int)] */
  logic [5:0] call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Int_1_emitted;
  logic [5:0] call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Int_1_done;
  assign call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Intgo_12_d = (call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Int_1_d[0] && (! call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Int_1_emitted[0]));
  assign call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_IntisZad2_d = (call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Int_1_d[0] && (! call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Int_1_emitted[1]));
  assign call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Intgad3_d = (call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Int_1_d[0] && (! call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Int_1_emitted[2]));
  assign call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Intm1ad4_d = {call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Int_1_d[16:1],
                                                                                                                                                              (call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Int_1_d[0] && (! call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Int_1_emitted[3]))};
  assign call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Intm2ad5_d = {call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Int_1_d[32:17],
                                                                                                                                                              (call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Int_1_d[0] && (! call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Int_1_emitted[4]))};
  assign call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Intsc_0_1_d = {call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Int_1_d[48:33],
                                                                                                                                                               (call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Int_1_d[0] && (! call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Int_1_emitted[5]))};
  assign call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Int_1_done = (call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Int_1_emitted | ({call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Intsc_0_1_d[0],
                                                                                                                                                                                                                                                                                                                       call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Intm2ad5_d[0],
                                                                                                                                                                                                                                                                                                                       call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Intm1ad4_d[0],
                                                                                                                                                                                                                                                                                                                       call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Intgad3_d[0],
                                                                                                                                                                                                                                                                                                                       call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_IntisZad2_d[0],
                                                                                                                                                                                                                                                                                                                       call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Intgo_12_d[0]} & {call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Intsc_0_1_r,
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Intm2ad5_r,
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Intm1ad4_r,
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Intgad3_r,
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_IntisZad2_r,
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Intgo_12_r}));
  assign call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Int_1_r = (& call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Int_1_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Int_1_emitted <= 6'd0;
    else
      call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Int_1_emitted <= (call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Int_1_r ? 6'd0 :
                                                                                                                                                               call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Int_1_done);
  
  /* rbuf (Ty Go) : (call_kron_kron_Int_Int_Int_goConst,Go) > (call_kron_kron_Int_Int_Int_initBufi,Go) */
  Go_t call_kron_kron_Int_Int_Int_goConst_buf;
  assign call_kron_kron_Int_Int_Int_goConst_r = (! call_kron_kron_Int_Int_Int_goConst_buf[0]);
  assign call_kron_kron_Int_Int_Int_initBufi_d = (call_kron_kron_Int_Int_Int_goConst_buf[0] ? call_kron_kron_Int_Int_Int_goConst_buf :
                                                  call_kron_kron_Int_Int_Int_goConst_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      call_kron_kron_Int_Int_Int_goConst_buf <= 1'd0;
    else
      if ((call_kron_kron_Int_Int_Int_initBufi_r && call_kron_kron_Int_Int_Int_goConst_buf[0]))
        call_kron_kron_Int_Int_Int_goConst_buf <= 1'd0;
      else if (((! call_kron_kron_Int_Int_Int_initBufi_r) && (! call_kron_kron_Int_Int_Int_goConst_buf[0])))
        call_kron_kron_Int_Int_Int_goConst_buf <= call_kron_kron_Int_Int_Int_goConst_d;
  
  /* mergectrl (Ty C5,Ty Go) : [(call_kron_kron_Int_Int_Int_goMux1,Go),
                           (lizzieLet29_3Lcall_kron_kron_Int_Int_Int3_1_argbuf,Go),
                           (lizzieLet29_3Lcall_kron_kron_Int_Int_Int2_1_argbuf,Go),
                           (lizzieLet29_3Lcall_kron_kron_Int_Int_Int1_1_argbuf,Go),
                           (lizzieLet6_4QNode_Int_1_argbuf,Go)] > (go_12_goMux_choice,C5) (go_12_goMux_data,Go) */
  logic [4:0] call_kron_kron_Int_Int_Int_goMux1_select_d;
  assign call_kron_kron_Int_Int_Int_goMux1_select_d = ((| call_kron_kron_Int_Int_Int_goMux1_select_q) ? call_kron_kron_Int_Int_Int_goMux1_select_q :
                                                       (call_kron_kron_Int_Int_Int_goMux1_d[0] ? 5'd1 :
                                                        (lizzieLet29_3Lcall_kron_kron_Int_Int_Int3_1_argbuf_d[0] ? 5'd2 :
                                                         (lizzieLet29_3Lcall_kron_kron_Int_Int_Int2_1_argbuf_d[0] ? 5'd4 :
                                                          (lizzieLet29_3Lcall_kron_kron_Int_Int_Int1_1_argbuf_d[0] ? 5'd8 :
                                                           (lizzieLet6_4QNode_Int_1_argbuf_d[0] ? 5'd16 :
                                                            5'd0))))));
  logic [4:0] call_kron_kron_Int_Int_Int_goMux1_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      call_kron_kron_Int_Int_Int_goMux1_select_q <= 5'd0;
    else
      call_kron_kron_Int_Int_Int_goMux1_select_q <= (call_kron_kron_Int_Int_Int_goMux1_done ? 5'd0 :
                                                     call_kron_kron_Int_Int_Int_goMux1_select_d);
  logic [1:0] call_kron_kron_Int_Int_Int_goMux1_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      call_kron_kron_Int_Int_Int_goMux1_emit_q <= 2'd0;
    else
      call_kron_kron_Int_Int_Int_goMux1_emit_q <= (call_kron_kron_Int_Int_Int_goMux1_done ? 2'd0 :
                                                   call_kron_kron_Int_Int_Int_goMux1_emit_d);
  logic [1:0] call_kron_kron_Int_Int_Int_goMux1_emit_d;
  assign call_kron_kron_Int_Int_Int_goMux1_emit_d = (call_kron_kron_Int_Int_Int_goMux1_emit_q | ({go_12_goMux_choice_d[0],
                                                                                                  go_12_goMux_data_d[0]} & {go_12_goMux_choice_r,
                                                                                                                            go_12_goMux_data_r}));
  logic call_kron_kron_Int_Int_Int_goMux1_done;
  assign call_kron_kron_Int_Int_Int_goMux1_done = (& call_kron_kron_Int_Int_Int_goMux1_emit_d);
  assign {lizzieLet6_4QNode_Int_1_argbuf_r,
          lizzieLet29_3Lcall_kron_kron_Int_Int_Int1_1_argbuf_r,
          lizzieLet29_3Lcall_kron_kron_Int_Int_Int2_1_argbuf_r,
          lizzieLet29_3Lcall_kron_kron_Int_Int_Int3_1_argbuf_r,
          call_kron_kron_Int_Int_Int_goMux1_r} = (call_kron_kron_Int_Int_Int_goMux1_done ? call_kron_kron_Int_Int_Int_goMux1_select_d :
                                                  5'd0);
  assign go_12_goMux_data_d = ((call_kron_kron_Int_Int_Int_goMux1_select_d[0] && (! call_kron_kron_Int_Int_Int_goMux1_emit_q[0])) ? call_kron_kron_Int_Int_Int_goMux1_d :
                               ((call_kron_kron_Int_Int_Int_goMux1_select_d[1] && (! call_kron_kron_Int_Int_Int_goMux1_emit_q[0])) ? lizzieLet29_3Lcall_kron_kron_Int_Int_Int3_1_argbuf_d :
                                ((call_kron_kron_Int_Int_Int_goMux1_select_d[2] && (! call_kron_kron_Int_Int_Int_goMux1_emit_q[0])) ? lizzieLet29_3Lcall_kron_kron_Int_Int_Int2_1_argbuf_d :
                                 ((call_kron_kron_Int_Int_Int_goMux1_select_d[3] && (! call_kron_kron_Int_Int_Int_goMux1_emit_q[0])) ? lizzieLet29_3Lcall_kron_kron_Int_Int_Int1_1_argbuf_d :
                                  ((call_kron_kron_Int_Int_Int_goMux1_select_d[4] && (! call_kron_kron_Int_Int_Int_goMux1_emit_q[0])) ? lizzieLet6_4QNode_Int_1_argbuf_d :
                                   1'd0)))));
  assign go_12_goMux_choice_d = ((call_kron_kron_Int_Int_Int_goMux1_select_d[0] && (! call_kron_kron_Int_Int_Int_goMux1_emit_q[1])) ? C1_5_dc(1'd1) :
                                 ((call_kron_kron_Int_Int_Int_goMux1_select_d[1] && (! call_kron_kron_Int_Int_Int_goMux1_emit_q[1])) ? C2_5_dc(1'd1) :
                                  ((call_kron_kron_Int_Int_Int_goMux1_select_d[2] && (! call_kron_kron_Int_Int_Int_goMux1_emit_q[1])) ? C3_5_dc(1'd1) :
                                   ((call_kron_kron_Int_Int_Int_goMux1_select_d[3] && (! call_kron_kron_Int_Int_Int_goMux1_emit_q[1])) ? C4_5_dc(1'd1) :
                                    ((call_kron_kron_Int_Int_Int_goMux1_select_d[4] && (! call_kron_kron_Int_Int_Int_goMux1_emit_q[1])) ? C5_5_dc(1'd1) :
                                     {3'd0, 1'd0})))));
  
  /* fork (Ty Go) : (call_kron_kron_Int_Int_Int_initBuf,Go) > [(call_kron_kron_Int_Int_Int_unlockFork1,Go),
                                                          (call_kron_kron_Int_Int_Int_unlockFork2,Go),
                                                          (call_kron_kron_Int_Int_Int_unlockFork3,Go),
                                                          (call_kron_kron_Int_Int_Int_unlockFork4,Go),
                                                          (call_kron_kron_Int_Int_Int_unlockFork5,Go),
                                                          (call_kron_kron_Int_Int_Int_unlockFork6,Go)] */
  logic [5:0] call_kron_kron_Int_Int_Int_initBuf_emitted;
  logic [5:0] call_kron_kron_Int_Int_Int_initBuf_done;
  assign call_kron_kron_Int_Int_Int_unlockFork1_d = (call_kron_kron_Int_Int_Int_initBuf_d[0] && (! call_kron_kron_Int_Int_Int_initBuf_emitted[0]));
  assign call_kron_kron_Int_Int_Int_unlockFork2_d = (call_kron_kron_Int_Int_Int_initBuf_d[0] && (! call_kron_kron_Int_Int_Int_initBuf_emitted[1]));
  assign call_kron_kron_Int_Int_Int_unlockFork3_d = (call_kron_kron_Int_Int_Int_initBuf_d[0] && (! call_kron_kron_Int_Int_Int_initBuf_emitted[2]));
  assign call_kron_kron_Int_Int_Int_unlockFork4_d = (call_kron_kron_Int_Int_Int_initBuf_d[0] && (! call_kron_kron_Int_Int_Int_initBuf_emitted[3]));
  assign call_kron_kron_Int_Int_Int_unlockFork5_d = (call_kron_kron_Int_Int_Int_initBuf_d[0] && (! call_kron_kron_Int_Int_Int_initBuf_emitted[4]));
  assign call_kron_kron_Int_Int_Int_unlockFork6_d = (call_kron_kron_Int_Int_Int_initBuf_d[0] && (! call_kron_kron_Int_Int_Int_initBuf_emitted[5]));
  assign call_kron_kron_Int_Int_Int_initBuf_done = (call_kron_kron_Int_Int_Int_initBuf_emitted | ({call_kron_kron_Int_Int_Int_unlockFork6_d[0],
                                                                                                   call_kron_kron_Int_Int_Int_unlockFork5_d[0],
                                                                                                   call_kron_kron_Int_Int_Int_unlockFork4_d[0],
                                                                                                   call_kron_kron_Int_Int_Int_unlockFork3_d[0],
                                                                                                   call_kron_kron_Int_Int_Int_unlockFork2_d[0],
                                                                                                   call_kron_kron_Int_Int_Int_unlockFork1_d[0]} & {call_kron_kron_Int_Int_Int_unlockFork6_r,
                                                                                                                                                   call_kron_kron_Int_Int_Int_unlockFork5_r,
                                                                                                                                                   call_kron_kron_Int_Int_Int_unlockFork4_r,
                                                                                                                                                   call_kron_kron_Int_Int_Int_unlockFork3_r,
                                                                                                                                                   call_kron_kron_Int_Int_Int_unlockFork2_r,
                                                                                                                                                   call_kron_kron_Int_Int_Int_unlockFork1_r}));
  assign call_kron_kron_Int_Int_Int_initBuf_r = (& call_kron_kron_Int_Int_Int_initBuf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      call_kron_kron_Int_Int_Int_initBuf_emitted <= 6'd0;
    else
      call_kron_kron_Int_Int_Int_initBuf_emitted <= (call_kron_kron_Int_Int_Int_initBuf_r ? 6'd0 :
                                                     call_kron_kron_Int_Int_Int_initBuf_done);
  
  /* initbuf (Ty Go,
         Dcon Go) : (call_kron_kron_Int_Int_Int_initBufi,Go) > (call_kron_kron_Int_Int_Int_initBuf,Go) */
  assign call_kron_kron_Int_Int_Int_initBufi_r = ((! call_kron_kron_Int_Int_Int_initBuf_d[0]) || call_kron_kron_Int_Int_Int_initBuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      call_kron_kron_Int_Int_Int_initBuf_d <= Go_dc(1'd1);
    else
      if (call_kron_kron_Int_Int_Int_initBufi_r)
        call_kron_kron_Int_Int_Int_initBuf_d <= call_kron_kron_Int_Int_Int_initBufi_d;
  
  /* mux (Ty Go,
     Ty Go) : (call_kron_kron_Int_Int_Int_unlockFork1,Go) [(call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Intgo_12,Go)] > (call_kron_kron_Int_Int_Int_goMux1,Go) */
  assign call_kron_kron_Int_Int_Int_goMux1_d = (call_kron_kron_Int_Int_Int_unlockFork1_d[0] && call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Intgo_12_d[0]);
  assign call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Intgo_12_r = (call_kron_kron_Int_Int_Int_goMux1_r && (call_kron_kron_Int_Int_Int_unlockFork1_d[0] && call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Intgo_12_d[0]));
  assign call_kron_kron_Int_Int_Int_unlockFork1_r = (call_kron_kron_Int_Int_Int_goMux1_r && (call_kron_kron_Int_Int_Int_unlockFork1_d[0] && call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Intgo_12_d[0]));
  
  /* mux (Ty Go,
     Ty MyDTInt_Bool) : (call_kron_kron_Int_Int_Int_unlockFork2,Go) [(call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_IntisZad2,MyDTInt_Bool)] > (call_kron_kron_Int_Int_Int_goMux2,MyDTInt_Bool) */
  assign call_kron_kron_Int_Int_Int_goMux2_d = (call_kron_kron_Int_Int_Int_unlockFork2_d[0] && call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_IntisZad2_d[0]);
  assign call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_IntisZad2_r = (call_kron_kron_Int_Int_Int_goMux2_r && (call_kron_kron_Int_Int_Int_unlockFork2_d[0] && call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_IntisZad2_d[0]));
  assign call_kron_kron_Int_Int_Int_unlockFork2_r = (call_kron_kron_Int_Int_Int_goMux2_r && (call_kron_kron_Int_Int_Int_unlockFork2_d[0] && call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_IntisZad2_d[0]));
  
  /* mux (Ty Go,
     Ty MyDTInt_Int_Int) : (call_kron_kron_Int_Int_Int_unlockFork3,Go) [(call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Intgad3,MyDTInt_Int_Int)] > (call_kron_kron_Int_Int_Int_goMux3,MyDTInt_Int_Int) */
  assign call_kron_kron_Int_Int_Int_goMux3_d = (call_kron_kron_Int_Int_Int_unlockFork3_d[0] && call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Intgad3_d[0]);
  assign call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Intgad3_r = (call_kron_kron_Int_Int_Int_goMux3_r && (call_kron_kron_Int_Int_Int_unlockFork3_d[0] && call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Intgad3_d[0]));
  assign call_kron_kron_Int_Int_Int_unlockFork3_r = (call_kron_kron_Int_Int_Int_goMux3_r && (call_kron_kron_Int_Int_Int_unlockFork3_d[0] && call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Intgad3_d[0]));
  
  /* mux (Ty Go,
     Ty Pointer_QTree_Int) : (call_kron_kron_Int_Int_Int_unlockFork4,Go) [(call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Intm1ad4,Pointer_QTree_Int)] > (call_kron_kron_Int_Int_Int_goMux4,Pointer_QTree_Int) */
  assign call_kron_kron_Int_Int_Int_goMux4_d = {call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Intm1ad4_d[16:1],
                                                (call_kron_kron_Int_Int_Int_unlockFork4_d[0] && call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Intm1ad4_d[0])};
  assign call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Intm1ad4_r = (call_kron_kron_Int_Int_Int_goMux4_r && (call_kron_kron_Int_Int_Int_unlockFork4_d[0] && call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Intm1ad4_d[0]));
  assign call_kron_kron_Int_Int_Int_unlockFork4_r = (call_kron_kron_Int_Int_Int_goMux4_r && (call_kron_kron_Int_Int_Int_unlockFork4_d[0] && call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Intm1ad4_d[0]));
  
  /* mux (Ty Go,
     Ty Pointer_QTree_Int) : (call_kron_kron_Int_Int_Int_unlockFork5,Go) [(call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Intm2ad5,Pointer_QTree_Int)] > (call_kron_kron_Int_Int_Int_goMux5,Pointer_QTree_Int) */
  assign call_kron_kron_Int_Int_Int_goMux5_d = {call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Intm2ad5_d[16:1],
                                                (call_kron_kron_Int_Int_Int_unlockFork5_d[0] && call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Intm2ad5_d[0])};
  assign call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Intm2ad5_r = (call_kron_kron_Int_Int_Int_goMux5_r && (call_kron_kron_Int_Int_Int_unlockFork5_d[0] && call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Intm2ad5_d[0]));
  assign call_kron_kron_Int_Int_Int_unlockFork5_r = (call_kron_kron_Int_Int_Int_goMux5_r && (call_kron_kron_Int_Int_Int_unlockFork5_d[0] && call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Intm2ad5_d[0]));
  
  /* mux (Ty Go,
     Ty Pointer_CTkron_kron_Int_Int_Int) : (call_kron_kron_Int_Int_Int_unlockFork6,Go) [(call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Intsc_0_1,Pointer_CTkron_kron_Int_Int_Int)] > (call_kron_kron_Int_Int_Int_goMux6,Pointer_CTkron_kron_Int_Int_Int) */
  assign call_kron_kron_Int_Int_Int_goMux6_d = {call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Intsc_0_1_d[16:1],
                                                (call_kron_kron_Int_Int_Int_unlockFork6_d[0] && call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Intsc_0_1_d[0])};
  assign call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Intsc_0_1_r = (call_kron_kron_Int_Int_Int_goMux6_r && (call_kron_kron_Int_Int_Int_unlockFork6_d[0] && call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Intsc_0_1_d[0]));
  assign call_kron_kron_Int_Int_Int_unlockFork6_r = (call_kron_kron_Int_Int_Int_goMux6_r && (call_kron_kron_Int_Int_Int_unlockFork6_d[0] && call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Intsc_0_1_d[0]));
  
  /* destruct (Ty TupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Int,
          Dcon TupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Int) : (call_main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Int_1,TupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Int) > [(call_main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Intgo_13,Go),
                                                                                                                                                                                                                                                                                                              (call_main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int___Pointer_CTmain_map'_Int_IntisZacL,MyDTInt_Bool),
                                                                                                                                                                                                                                                                                                              (call_main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int___Pointer_CTmain_map'_Int_IntgacM,MyDTInt_Int),
                                                                                                                                                                                                                                                                                                              (call_main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int___Pointer_CTmain_map'_Int_IntmacN,Pointer_QTree_Int),
                                                                                                                                                                                                                                                                                                              (call_main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Intsc_0_2,Pointer_CTmain_map'_Int_Int)] */
  logic [4:0] \call_main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Int_1_emitted ;
  logic [4:0] \call_main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Int_1_done ;
  assign \call_main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Intgo_13_d  = (\call_main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Int_1_d [0] && (! \call_main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Int_1_emitted [0]));
  assign \call_main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int___Pointer_CTmain_map'_Int_IntisZacL_d  = (\call_main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Int_1_d [0] && (! \call_main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Int_1_emitted [1]));
  assign \call_main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int___Pointer_CTmain_map'_Int_IntgacM_d  = (\call_main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Int_1_d [0] && (! \call_main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Int_1_emitted [2]));
  assign \call_main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int___Pointer_CTmain_map'_Int_IntmacN_d  = {\call_main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Int_1_d [16:1],
                                                                                                                               (\call_main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Int_1_d [0] && (! \call_main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Int_1_emitted [3]))};
  assign \call_main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Intsc_0_2_d  = {\call_main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Int_1_d [32:17],
                                                                                                                                 (\call_main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Int_1_d [0] && (! \call_main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Int_1_emitted [4]))};
  assign \call_main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Int_1_done  = (\call_main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Int_1_emitted  | ({\call_main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Intsc_0_2_d [0],
                                                                                                                                                                                                                                                           \call_main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int___Pointer_CTmain_map'_Int_IntmacN_d [0],
                                                                                                                                                                                                                                                           \call_main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int___Pointer_CTmain_map'_Int_IntgacM_d [0],
                                                                                                                                                                                                                                                           \call_main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int___Pointer_CTmain_map'_Int_IntisZacL_d [0],
                                                                                                                                                                                                                                                           \call_main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Intgo_13_d [0]} & {\call_main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Intsc_0_2_r ,
                                                                                                                                                                                                                                                                                                                                                                                      \call_main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int___Pointer_CTmain_map'_Int_IntmacN_r ,
                                                                                                                                                                                                                                                                                                                                                                                      \call_main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int___Pointer_CTmain_map'_Int_IntgacM_r ,
                                                                                                                                                                                                                                                                                                                                                                                      \call_main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int___Pointer_CTmain_map'_Int_IntisZacL_r ,
                                                                                                                                                                                                                                                                                                                                                                                      \call_main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Intgo_13_r }));
  assign \call_main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Int_1_r  = (& \call_main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Int_1_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \call_main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Int_1_emitted  <= 5'd0;
    else
      \call_main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Int_1_emitted  <= (\call_main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Int_1_r  ? 5'd0 :
                                                                                                                                 \call_main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Int_1_done );
  
  /* rbuf (Ty Go) : (call_main_map'_Int_Int_goConst,Go) > (call_main_map'_Int_Int_initBufi,Go) */
  Go_t \call_main_map'_Int_Int_goConst_buf ;
  assign \call_main_map'_Int_Int_goConst_r  = (! \call_main_map'_Int_Int_goConst_buf [0]);
  assign \call_main_map'_Int_Int_initBufi_d  = (\call_main_map'_Int_Int_goConst_buf [0] ? \call_main_map'_Int_Int_goConst_buf  :
                                                \call_main_map'_Int_Int_goConst_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \call_main_map'_Int_Int_goConst_buf  <= 1'd0;
    else
      if ((\call_main_map'_Int_Int_initBufi_r  && \call_main_map'_Int_Int_goConst_buf [0]))
        \call_main_map'_Int_Int_goConst_buf  <= 1'd0;
      else if (((! \call_main_map'_Int_Int_initBufi_r ) && (! \call_main_map'_Int_Int_goConst_buf [0])))
        \call_main_map'_Int_Int_goConst_buf  <= \call_main_map'_Int_Int_goConst_d ;
  
  /* mergectrl (Ty C5,Ty Go) : [(call_main_map'_Int_Int_goMux1,Go),
                           (lizzieLet34_3Lcall_main_map'_Int_Int3_1_argbuf,Go),
                           (lizzieLet34_3Lcall_main_map'_Int_Int2_1_argbuf,Go),
                           (lizzieLet34_3Lcall_main_map'_Int_Int1_1_argbuf,Go),
                           (lizzieLet10_4QNode_Int_1_argbuf,Go)] > (go_13_goMux_choice,C5) (go_13_goMux_data,Go) */
  logic [4:0] \call_main_map'_Int_Int_goMux1_select_d ;
  assign \call_main_map'_Int_Int_goMux1_select_d  = ((| \call_main_map'_Int_Int_goMux1_select_q ) ? \call_main_map'_Int_Int_goMux1_select_q  :
                                                     (\call_main_map'_Int_Int_goMux1_d [0] ? 5'd1 :
                                                      (\lizzieLet34_3Lcall_main_map'_Int_Int3_1_argbuf_d [0] ? 5'd2 :
                                                       (\lizzieLet34_3Lcall_main_map'_Int_Int2_1_argbuf_d [0] ? 5'd4 :
                                                        (\lizzieLet34_3Lcall_main_map'_Int_Int1_1_argbuf_d [0] ? 5'd8 :
                                                         (lizzieLet10_4QNode_Int_1_argbuf_d[0] ? 5'd16 :
                                                          5'd0))))));
  logic [4:0] \call_main_map'_Int_Int_goMux1_select_q ;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \call_main_map'_Int_Int_goMux1_select_q  <= 5'd0;
    else
      \call_main_map'_Int_Int_goMux1_select_q  <= (\call_main_map'_Int_Int_goMux1_done  ? 5'd0 :
                                                   \call_main_map'_Int_Int_goMux1_select_d );
  logic [1:0] \call_main_map'_Int_Int_goMux1_emit_q ;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \call_main_map'_Int_Int_goMux1_emit_q  <= 2'd0;
    else
      \call_main_map'_Int_Int_goMux1_emit_q  <= (\call_main_map'_Int_Int_goMux1_done  ? 2'd0 :
                                                 \call_main_map'_Int_Int_goMux1_emit_d );
  logic [1:0] \call_main_map'_Int_Int_goMux1_emit_d ;
  assign \call_main_map'_Int_Int_goMux1_emit_d  = (\call_main_map'_Int_Int_goMux1_emit_q  | ({go_13_goMux_choice_d[0],
                                                                                              go_13_goMux_data_d[0]} & {go_13_goMux_choice_r,
                                                                                                                        go_13_goMux_data_r}));
  logic \call_main_map'_Int_Int_goMux1_done ;
  assign \call_main_map'_Int_Int_goMux1_done  = (& \call_main_map'_Int_Int_goMux1_emit_d );
  assign {lizzieLet10_4QNode_Int_1_argbuf_r,
          \lizzieLet34_3Lcall_main_map'_Int_Int1_1_argbuf_r ,
          \lizzieLet34_3Lcall_main_map'_Int_Int2_1_argbuf_r ,
          \lizzieLet34_3Lcall_main_map'_Int_Int3_1_argbuf_r ,
          \call_main_map'_Int_Int_goMux1_r } = (\call_main_map'_Int_Int_goMux1_done  ? \call_main_map'_Int_Int_goMux1_select_d  :
                                                5'd0);
  assign go_13_goMux_data_d = ((\call_main_map'_Int_Int_goMux1_select_d [0] && (! \call_main_map'_Int_Int_goMux1_emit_q [0])) ? \call_main_map'_Int_Int_goMux1_d  :
                               ((\call_main_map'_Int_Int_goMux1_select_d [1] && (! \call_main_map'_Int_Int_goMux1_emit_q [0])) ? \lizzieLet34_3Lcall_main_map'_Int_Int3_1_argbuf_d  :
                                ((\call_main_map'_Int_Int_goMux1_select_d [2] && (! \call_main_map'_Int_Int_goMux1_emit_q [0])) ? \lizzieLet34_3Lcall_main_map'_Int_Int2_1_argbuf_d  :
                                 ((\call_main_map'_Int_Int_goMux1_select_d [3] && (! \call_main_map'_Int_Int_goMux1_emit_q [0])) ? \lizzieLet34_3Lcall_main_map'_Int_Int1_1_argbuf_d  :
                                  ((\call_main_map'_Int_Int_goMux1_select_d [4] && (! \call_main_map'_Int_Int_goMux1_emit_q [0])) ? lizzieLet10_4QNode_Int_1_argbuf_d :
                                   1'd0)))));
  assign go_13_goMux_choice_d = ((\call_main_map'_Int_Int_goMux1_select_d [0] && (! \call_main_map'_Int_Int_goMux1_emit_q [1])) ? C1_5_dc(1'd1) :
                                 ((\call_main_map'_Int_Int_goMux1_select_d [1] && (! \call_main_map'_Int_Int_goMux1_emit_q [1])) ? C2_5_dc(1'd1) :
                                  ((\call_main_map'_Int_Int_goMux1_select_d [2] && (! \call_main_map'_Int_Int_goMux1_emit_q [1])) ? C3_5_dc(1'd1) :
                                   ((\call_main_map'_Int_Int_goMux1_select_d [3] && (! \call_main_map'_Int_Int_goMux1_emit_q [1])) ? C4_5_dc(1'd1) :
                                    ((\call_main_map'_Int_Int_goMux1_select_d [4] && (! \call_main_map'_Int_Int_goMux1_emit_q [1])) ? C5_5_dc(1'd1) :
                                     {3'd0, 1'd0})))));
  
  /* fork (Ty Go) : (call_main_map'_Int_Int_initBuf,Go) > [(call_main_map'_Int_Int_unlockFork1,Go),
                                                      (call_main_map'_Int_Int_unlockFork2,Go),
                                                      (call_main_map'_Int_Int_unlockFork3,Go),
                                                      (call_main_map'_Int_Int_unlockFork4,Go),
                                                      (call_main_map'_Int_Int_unlockFork5,Go)] */
  logic [4:0] \call_main_map'_Int_Int_initBuf_emitted ;
  logic [4:0] \call_main_map'_Int_Int_initBuf_done ;
  assign \call_main_map'_Int_Int_unlockFork1_d  = (\call_main_map'_Int_Int_initBuf_d [0] && (! \call_main_map'_Int_Int_initBuf_emitted [0]));
  assign \call_main_map'_Int_Int_unlockFork2_d  = (\call_main_map'_Int_Int_initBuf_d [0] && (! \call_main_map'_Int_Int_initBuf_emitted [1]));
  assign \call_main_map'_Int_Int_unlockFork3_d  = (\call_main_map'_Int_Int_initBuf_d [0] && (! \call_main_map'_Int_Int_initBuf_emitted [2]));
  assign \call_main_map'_Int_Int_unlockFork4_d  = (\call_main_map'_Int_Int_initBuf_d [0] && (! \call_main_map'_Int_Int_initBuf_emitted [3]));
  assign \call_main_map'_Int_Int_unlockFork5_d  = (\call_main_map'_Int_Int_initBuf_d [0] && (! \call_main_map'_Int_Int_initBuf_emitted [4]));
  assign \call_main_map'_Int_Int_initBuf_done  = (\call_main_map'_Int_Int_initBuf_emitted  | ({\call_main_map'_Int_Int_unlockFork5_d [0],
                                                                                               \call_main_map'_Int_Int_unlockFork4_d [0],
                                                                                               \call_main_map'_Int_Int_unlockFork3_d [0],
                                                                                               \call_main_map'_Int_Int_unlockFork2_d [0],
                                                                                               \call_main_map'_Int_Int_unlockFork1_d [0]} & {\call_main_map'_Int_Int_unlockFork5_r ,
                                                                                                                                             \call_main_map'_Int_Int_unlockFork4_r ,
                                                                                                                                             \call_main_map'_Int_Int_unlockFork3_r ,
                                                                                                                                             \call_main_map'_Int_Int_unlockFork2_r ,
                                                                                                                                             \call_main_map'_Int_Int_unlockFork1_r }));
  assign \call_main_map'_Int_Int_initBuf_r  = (& \call_main_map'_Int_Int_initBuf_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \call_main_map'_Int_Int_initBuf_emitted  <= 5'd0;
    else
      \call_main_map'_Int_Int_initBuf_emitted  <= (\call_main_map'_Int_Int_initBuf_r  ? 5'd0 :
                                                   \call_main_map'_Int_Int_initBuf_done );
  
  /* initbuf (Ty Go,
         Dcon Go) : (call_main_map'_Int_Int_initBufi,Go) > (call_main_map'_Int_Int_initBuf,Go) */
  assign \call_main_map'_Int_Int_initBufi_r  = ((! \call_main_map'_Int_Int_initBuf_d [0]) || \call_main_map'_Int_Int_initBuf_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \call_main_map'_Int_Int_initBuf_d  <= Go_dc(1'd1);
    else
      if (\call_main_map'_Int_Int_initBufi_r )
        \call_main_map'_Int_Int_initBuf_d  <= \call_main_map'_Int_Int_initBufi_d ;
  
  /* mux (Ty Go,
     Ty Go) : (call_main_map'_Int_Int_unlockFork1,Go) [(call_main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Intgo_13,Go)] > (call_main_map'_Int_Int_goMux1,Go) */
  assign \call_main_map'_Int_Int_goMux1_d  = (\call_main_map'_Int_Int_unlockFork1_d [0] && \call_main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Intgo_13_d [0]);
  assign \call_main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Intgo_13_r  = (\call_main_map'_Int_Int_goMux1_r  && (\call_main_map'_Int_Int_unlockFork1_d [0] && \call_main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Intgo_13_d [0]));
  assign \call_main_map'_Int_Int_unlockFork1_r  = (\call_main_map'_Int_Int_goMux1_r  && (\call_main_map'_Int_Int_unlockFork1_d [0] && \call_main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Intgo_13_d [0]));
  
  /* mux (Ty Go,
     Ty MyDTInt_Bool) : (call_main_map'_Int_Int_unlockFork2,Go) [(call_main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int___Pointer_CTmain_map'_Int_IntisZacL,MyDTInt_Bool)] > (call_main_map'_Int_Int_goMux2,MyDTInt_Bool) */
  assign \call_main_map'_Int_Int_goMux2_d  = (\call_main_map'_Int_Int_unlockFork2_d [0] && \call_main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int___Pointer_CTmain_map'_Int_IntisZacL_d [0]);
  assign \call_main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int___Pointer_CTmain_map'_Int_IntisZacL_r  = (\call_main_map'_Int_Int_goMux2_r  && (\call_main_map'_Int_Int_unlockFork2_d [0] && \call_main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int___Pointer_CTmain_map'_Int_IntisZacL_d [0]));
  assign \call_main_map'_Int_Int_unlockFork2_r  = (\call_main_map'_Int_Int_goMux2_r  && (\call_main_map'_Int_Int_unlockFork2_d [0] && \call_main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int___Pointer_CTmain_map'_Int_IntisZacL_d [0]));
  
  /* mux (Ty Go,
     Ty MyDTInt_Int) : (call_main_map'_Int_Int_unlockFork3,Go) [(call_main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int___Pointer_CTmain_map'_Int_IntgacM,MyDTInt_Int)] > (call_main_map'_Int_Int_goMux3,MyDTInt_Int) */
  assign \call_main_map'_Int_Int_goMux3_d  = (\call_main_map'_Int_Int_unlockFork3_d [0] && \call_main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int___Pointer_CTmain_map'_Int_IntgacM_d [0]);
  assign \call_main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int___Pointer_CTmain_map'_Int_IntgacM_r  = (\call_main_map'_Int_Int_goMux3_r  && (\call_main_map'_Int_Int_unlockFork3_d [0] && \call_main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int___Pointer_CTmain_map'_Int_IntgacM_d [0]));
  assign \call_main_map'_Int_Int_unlockFork3_r  = (\call_main_map'_Int_Int_goMux3_r  && (\call_main_map'_Int_Int_unlockFork3_d [0] && \call_main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int___Pointer_CTmain_map'_Int_IntgacM_d [0]));
  
  /* mux (Ty Go,
     Ty Pointer_QTree_Int) : (call_main_map'_Int_Int_unlockFork4,Go) [(call_main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int___Pointer_CTmain_map'_Int_IntmacN,Pointer_QTree_Int)] > (call_main_map'_Int_Int_goMux4,Pointer_QTree_Int) */
  assign \call_main_map'_Int_Int_goMux4_d  = {\call_main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int___Pointer_CTmain_map'_Int_IntmacN_d [16:1],
                                              (\call_main_map'_Int_Int_unlockFork4_d [0] && \call_main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int___Pointer_CTmain_map'_Int_IntmacN_d [0])};
  assign \call_main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int___Pointer_CTmain_map'_Int_IntmacN_r  = (\call_main_map'_Int_Int_goMux4_r  && (\call_main_map'_Int_Int_unlockFork4_d [0] && \call_main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int___Pointer_CTmain_map'_Int_IntmacN_d [0]));
  assign \call_main_map'_Int_Int_unlockFork4_r  = (\call_main_map'_Int_Int_goMux4_r  && (\call_main_map'_Int_Int_unlockFork4_d [0] && \call_main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int___Pointer_CTmain_map'_Int_IntmacN_d [0]));
  
  /* mux (Ty Go,
     Ty Pointer_CTmain_map'_Int_Int) : (call_main_map'_Int_Int_unlockFork5,Go) [(call_main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Intsc_0_2,Pointer_CTmain_map'_Int_Int)] > (call_main_map'_Int_Int_goMux5,Pointer_CTmain_map'_Int_Int) */
  assign \call_main_map'_Int_Int_goMux5_d  = {\call_main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Intsc_0_2_d [16:1],
                                              (\call_main_map'_Int_Int_unlockFork5_d [0] && \call_main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Intsc_0_2_d [0])};
  assign \call_main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Intsc_0_2_r  = (\call_main_map'_Int_Int_goMux5_r  && (\call_main_map'_Int_Int_unlockFork5_d [0] && \call_main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Intsc_0_2_d [0]));
  assign \call_main_map'_Int_Int_unlockFork5_r  = (\call_main_map'_Int_Int_goMux5_r  && (\call_main_map'_Int_Int_unlockFork5_d [0] && \call_main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Intsc_0_2_d [0]));
  
  /* destruct (Ty TupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Int,
          Dcon TupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Int) : (call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Int_1,TupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Int) > [(call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Intgo_14,Go),
                                                                                                                                                                                                                                                                                                                                                                    (call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_IntisZacT,MyDTInt_Bool),
                                                                                                                                                                                                                                                                                                                                                                    (call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_IntgacU,MyDTInt_Int_Int),
                                                                                                                                                                                                                                                                                                                                                                    (call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Intv'acV,Int),
                                                                                                                                                                                                                                                                                                                                                                    (call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_IntmacW,Pointer_QTree_Int),
                                                                                                                                                                                                                                                                                                                                                                    (call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Intsc_0_3,Pointer_CTmap''_map''_Int_Int_Int)] */
  logic [5:0] \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Int_1_emitted ;
  logic [5:0] \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Int_1_done ;
  assign \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Intgo_14_d  = (\call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Int_1_d [0] && (! \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Int_1_emitted [0]));
  assign \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_IntisZacT_d  = (\call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Int_1_d [0] && (! \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Int_1_emitted [1]));
  assign \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_IntgacU_d  = (\call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Int_1_d [0] && (! \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Int_1_emitted [2]));
  assign \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Intv'acV_d  = {\call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Int_1_d [32:1],
                                                                                                                                                      (\call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Int_1_d [0] && (! \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Int_1_emitted [3]))};
  assign \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_IntmacW_d  = {\call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Int_1_d [48:33],
                                                                                                                                                     (\call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Int_1_d [0] && (! \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Int_1_emitted [4]))};
  assign \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Intsc_0_3_d  = {\call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Int_1_d [64:49],
                                                                                                                                                       (\call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Int_1_d [0] && (! \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Int_1_emitted [5]))};
  assign \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Int_1_done  = (\call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Int_1_emitted  | ({\call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Intsc_0_3_d [0],
                                                                                                                                                                                                                                                                                                       \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_IntmacW_d [0],
                                                                                                                                                                                                                                                                                                       \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Intv'acV_d [0],
                                                                                                                                                                                                                                                                                                       \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_IntgacU_d [0],
                                                                                                                                                                                                                                                                                                       \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_IntisZacT_d [0],
                                                                                                                                                                                                                                                                                                       \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Intgo_14_d [0]} & {\call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Intsc_0_3_r ,
                                                                                                                                                                                                                                                                                                                                                                                                                                                        \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_IntmacW_r ,
                                                                                                                                                                                                                                                                                                                                                                                                                                                        \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Intv'acV_r ,
                                                                                                                                                                                                                                                                                                                                                                                                                                                        \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_IntgacU_r ,
                                                                                                                                                                                                                                                                                                                                                                                                                                                        \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_IntisZacT_r ,
                                                                                                                                                                                                                                                                                                                                                                                                                                                        \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Intgo_14_r }));
  assign \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Int_1_r  = (& \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Int_1_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Int_1_emitted  <= 6'd0;
    else
      \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Int_1_emitted  <= (\call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Int_1_r  ? 6'd0 :
                                                                                                                                                       \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Int_1_done );
  
  /* rbuf (Ty Go) : (call_map''_map''_Int_Int_Int_goConst,Go) > (call_map''_map''_Int_Int_Int_initBufi,Go) */
  Go_t \call_map''_map''_Int_Int_Int_goConst_buf ;
  assign \call_map''_map''_Int_Int_Int_goConst_r  = (! \call_map''_map''_Int_Int_Int_goConst_buf [0]);
  assign \call_map''_map''_Int_Int_Int_initBufi_d  = (\call_map''_map''_Int_Int_Int_goConst_buf [0] ? \call_map''_map''_Int_Int_Int_goConst_buf  :
                                                      \call_map''_map''_Int_Int_Int_goConst_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \call_map''_map''_Int_Int_Int_goConst_buf  <= 1'd0;
    else
      if ((\call_map''_map''_Int_Int_Int_initBufi_r  && \call_map''_map''_Int_Int_Int_goConst_buf [0]))
        \call_map''_map''_Int_Int_Int_goConst_buf  <= 1'd0;
      else if (((! \call_map''_map''_Int_Int_Int_initBufi_r ) && (! \call_map''_map''_Int_Int_Int_goConst_buf [0])))
        \call_map''_map''_Int_Int_Int_goConst_buf  <= \call_map''_map''_Int_Int_Int_goConst_d ;
  
  /* mergectrl (Ty C5,
           Ty Go) : [(call_map''_map''_Int_Int_Int_goMux1,Go),
                     (lizzieLet39_3Lcall_map''_map''_Int_Int_Int3_1_argbuf,Go),
                     (lizzieLet39_3Lcall_map''_map''_Int_Int_Int2_1_argbuf,Go),
                     (lizzieLet39_3Lcall_map''_map''_Int_Int_Int1_1_argbuf,Go),
                     (lizzieLet16_1_4QNode_Int_1_argbuf,Go)] > (go_14_goMux_choice,C5) (go_14_goMux_data,Go) */
  logic [4:0] \call_map''_map''_Int_Int_Int_goMux1_select_d ;
  assign \call_map''_map''_Int_Int_Int_goMux1_select_d  = ((| \call_map''_map''_Int_Int_Int_goMux1_select_q ) ? \call_map''_map''_Int_Int_Int_goMux1_select_q  :
                                                           (\call_map''_map''_Int_Int_Int_goMux1_d [0] ? 5'd1 :
                                                            (\lizzieLet39_3Lcall_map''_map''_Int_Int_Int3_1_argbuf_d [0] ? 5'd2 :
                                                             (\lizzieLet39_3Lcall_map''_map''_Int_Int_Int2_1_argbuf_d [0] ? 5'd4 :
                                                              (\lizzieLet39_3Lcall_map''_map''_Int_Int_Int1_1_argbuf_d [0] ? 5'd8 :
                                                               (lizzieLet16_1_4QNode_Int_1_argbuf_d[0] ? 5'd16 :
                                                                5'd0))))));
  logic [4:0] \call_map''_map''_Int_Int_Int_goMux1_select_q ;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \call_map''_map''_Int_Int_Int_goMux1_select_q  <= 5'd0;
    else
      \call_map''_map''_Int_Int_Int_goMux1_select_q  <= (\call_map''_map''_Int_Int_Int_goMux1_done  ? 5'd0 :
                                                         \call_map''_map''_Int_Int_Int_goMux1_select_d );
  logic [1:0] \call_map''_map''_Int_Int_Int_goMux1_emit_q ;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \call_map''_map''_Int_Int_Int_goMux1_emit_q  <= 2'd0;
    else
      \call_map''_map''_Int_Int_Int_goMux1_emit_q  <= (\call_map''_map''_Int_Int_Int_goMux1_done  ? 2'd0 :
                                                       \call_map''_map''_Int_Int_Int_goMux1_emit_d );
  logic [1:0] \call_map''_map''_Int_Int_Int_goMux1_emit_d ;
  assign \call_map''_map''_Int_Int_Int_goMux1_emit_d  = (\call_map''_map''_Int_Int_Int_goMux1_emit_q  | ({go_14_goMux_choice_d[0],
                                                                                                          go_14_goMux_data_d[0]} & {go_14_goMux_choice_r,
                                                                                                                                    go_14_goMux_data_r}));
  logic \call_map''_map''_Int_Int_Int_goMux1_done ;
  assign \call_map''_map''_Int_Int_Int_goMux1_done  = (& \call_map''_map''_Int_Int_Int_goMux1_emit_d );
  assign {lizzieLet16_1_4QNode_Int_1_argbuf_r,
          \lizzieLet39_3Lcall_map''_map''_Int_Int_Int1_1_argbuf_r ,
          \lizzieLet39_3Lcall_map''_map''_Int_Int_Int2_1_argbuf_r ,
          \lizzieLet39_3Lcall_map''_map''_Int_Int_Int3_1_argbuf_r ,
          \call_map''_map''_Int_Int_Int_goMux1_r } = (\call_map''_map''_Int_Int_Int_goMux1_done  ? \call_map''_map''_Int_Int_Int_goMux1_select_d  :
                                                      5'd0);
  assign go_14_goMux_data_d = ((\call_map''_map''_Int_Int_Int_goMux1_select_d [0] && (! \call_map''_map''_Int_Int_Int_goMux1_emit_q [0])) ? \call_map''_map''_Int_Int_Int_goMux1_d  :
                               ((\call_map''_map''_Int_Int_Int_goMux1_select_d [1] && (! \call_map''_map''_Int_Int_Int_goMux1_emit_q [0])) ? \lizzieLet39_3Lcall_map''_map''_Int_Int_Int3_1_argbuf_d  :
                                ((\call_map''_map''_Int_Int_Int_goMux1_select_d [2] && (! \call_map''_map''_Int_Int_Int_goMux1_emit_q [0])) ? \lizzieLet39_3Lcall_map''_map''_Int_Int_Int2_1_argbuf_d  :
                                 ((\call_map''_map''_Int_Int_Int_goMux1_select_d [3] && (! \call_map''_map''_Int_Int_Int_goMux1_emit_q [0])) ? \lizzieLet39_3Lcall_map''_map''_Int_Int_Int1_1_argbuf_d  :
                                  ((\call_map''_map''_Int_Int_Int_goMux1_select_d [4] && (! \call_map''_map''_Int_Int_Int_goMux1_emit_q [0])) ? lizzieLet16_1_4QNode_Int_1_argbuf_d :
                                   1'd0)))));
  assign go_14_goMux_choice_d = ((\call_map''_map''_Int_Int_Int_goMux1_select_d [0] && (! \call_map''_map''_Int_Int_Int_goMux1_emit_q [1])) ? C1_5_dc(1'd1) :
                                 ((\call_map''_map''_Int_Int_Int_goMux1_select_d [1] && (! \call_map''_map''_Int_Int_Int_goMux1_emit_q [1])) ? C2_5_dc(1'd1) :
                                  ((\call_map''_map''_Int_Int_Int_goMux1_select_d [2] && (! \call_map''_map''_Int_Int_Int_goMux1_emit_q [1])) ? C3_5_dc(1'd1) :
                                   ((\call_map''_map''_Int_Int_Int_goMux1_select_d [3] && (! \call_map''_map''_Int_Int_Int_goMux1_emit_q [1])) ? C4_5_dc(1'd1) :
                                    ((\call_map''_map''_Int_Int_Int_goMux1_select_d [4] && (! \call_map''_map''_Int_Int_Int_goMux1_emit_q [1])) ? C5_5_dc(1'd1) :
                                     {3'd0, 1'd0})))));
  
  /* fork (Ty Go) : (call_map''_map''_Int_Int_Int_initBuf,Go) > [(call_map''_map''_Int_Int_Int_unlockFork1,Go),
                                                            (call_map''_map''_Int_Int_Int_unlockFork2,Go),
                                                            (call_map''_map''_Int_Int_Int_unlockFork3,Go),
                                                            (call_map''_map''_Int_Int_Int_unlockFork4,Go),
                                                            (call_map''_map''_Int_Int_Int_unlockFork5,Go),
                                                            (call_map''_map''_Int_Int_Int_unlockFork6,Go)] */
  logic [5:0] \call_map''_map''_Int_Int_Int_initBuf_emitted ;
  logic [5:0] \call_map''_map''_Int_Int_Int_initBuf_done ;
  assign \call_map''_map''_Int_Int_Int_unlockFork1_d  = (\call_map''_map''_Int_Int_Int_initBuf_d [0] && (! \call_map''_map''_Int_Int_Int_initBuf_emitted [0]));
  assign \call_map''_map''_Int_Int_Int_unlockFork2_d  = (\call_map''_map''_Int_Int_Int_initBuf_d [0] && (! \call_map''_map''_Int_Int_Int_initBuf_emitted [1]));
  assign \call_map''_map''_Int_Int_Int_unlockFork3_d  = (\call_map''_map''_Int_Int_Int_initBuf_d [0] && (! \call_map''_map''_Int_Int_Int_initBuf_emitted [2]));
  assign \call_map''_map''_Int_Int_Int_unlockFork4_d  = (\call_map''_map''_Int_Int_Int_initBuf_d [0] && (! \call_map''_map''_Int_Int_Int_initBuf_emitted [3]));
  assign \call_map''_map''_Int_Int_Int_unlockFork5_d  = (\call_map''_map''_Int_Int_Int_initBuf_d [0] && (! \call_map''_map''_Int_Int_Int_initBuf_emitted [4]));
  assign \call_map''_map''_Int_Int_Int_unlockFork6_d  = (\call_map''_map''_Int_Int_Int_initBuf_d [0] && (! \call_map''_map''_Int_Int_Int_initBuf_emitted [5]));
  assign \call_map''_map''_Int_Int_Int_initBuf_done  = (\call_map''_map''_Int_Int_Int_initBuf_emitted  | ({\call_map''_map''_Int_Int_Int_unlockFork6_d [0],
                                                                                                           \call_map''_map''_Int_Int_Int_unlockFork5_d [0],
                                                                                                           \call_map''_map''_Int_Int_Int_unlockFork4_d [0],
                                                                                                           \call_map''_map''_Int_Int_Int_unlockFork3_d [0],
                                                                                                           \call_map''_map''_Int_Int_Int_unlockFork2_d [0],
                                                                                                           \call_map''_map''_Int_Int_Int_unlockFork1_d [0]} & {\call_map''_map''_Int_Int_Int_unlockFork6_r ,
                                                                                                                                                               \call_map''_map''_Int_Int_Int_unlockFork5_r ,
                                                                                                                                                               \call_map''_map''_Int_Int_Int_unlockFork4_r ,
                                                                                                                                                               \call_map''_map''_Int_Int_Int_unlockFork3_r ,
                                                                                                                                                               \call_map''_map''_Int_Int_Int_unlockFork2_r ,
                                                                                                                                                               \call_map''_map''_Int_Int_Int_unlockFork1_r }));
  assign \call_map''_map''_Int_Int_Int_initBuf_r  = (& \call_map''_map''_Int_Int_Int_initBuf_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \call_map''_map''_Int_Int_Int_initBuf_emitted  <= 6'd0;
    else
      \call_map''_map''_Int_Int_Int_initBuf_emitted  <= (\call_map''_map''_Int_Int_Int_initBuf_r  ? 6'd0 :
                                                         \call_map''_map''_Int_Int_Int_initBuf_done );
  
  /* initbuf (Ty Go,
         Dcon Go) : (call_map''_map''_Int_Int_Int_initBufi,Go) > (call_map''_map''_Int_Int_Int_initBuf,Go) */
  assign \call_map''_map''_Int_Int_Int_initBufi_r  = ((! \call_map''_map''_Int_Int_Int_initBuf_d [0]) || \call_map''_map''_Int_Int_Int_initBuf_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \call_map''_map''_Int_Int_Int_initBuf_d  <= Go_dc(1'd1);
    else
      if (\call_map''_map''_Int_Int_Int_initBufi_r )
        \call_map''_map''_Int_Int_Int_initBuf_d  <= \call_map''_map''_Int_Int_Int_initBufi_d ;
  
  /* mux (Ty Go,
     Ty Go) : (call_map''_map''_Int_Int_Int_unlockFork1,Go) [(call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Intgo_14,Go)] > (call_map''_map''_Int_Int_Int_goMux1,Go) */
  assign \call_map''_map''_Int_Int_Int_goMux1_d  = (\call_map''_map''_Int_Int_Int_unlockFork1_d [0] && \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Intgo_14_d [0]);
  assign \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Intgo_14_r  = (\call_map''_map''_Int_Int_Int_goMux1_r  && (\call_map''_map''_Int_Int_Int_unlockFork1_d [0] && \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Intgo_14_d [0]));
  assign \call_map''_map''_Int_Int_Int_unlockFork1_r  = (\call_map''_map''_Int_Int_Int_goMux1_r  && (\call_map''_map''_Int_Int_Int_unlockFork1_d [0] && \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Intgo_14_d [0]));
  
  /* mux (Ty Go,
     Ty MyDTInt_Bool) : (call_map''_map''_Int_Int_Int_unlockFork2,Go) [(call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_IntisZacT,MyDTInt_Bool)] > (call_map''_map''_Int_Int_Int_goMux2,MyDTInt_Bool) */
  assign \call_map''_map''_Int_Int_Int_goMux2_d  = (\call_map''_map''_Int_Int_Int_unlockFork2_d [0] && \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_IntisZacT_d [0]);
  assign \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_IntisZacT_r  = (\call_map''_map''_Int_Int_Int_goMux2_r  && (\call_map''_map''_Int_Int_Int_unlockFork2_d [0] && \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_IntisZacT_d [0]));
  assign \call_map''_map''_Int_Int_Int_unlockFork2_r  = (\call_map''_map''_Int_Int_Int_goMux2_r  && (\call_map''_map''_Int_Int_Int_unlockFork2_d [0] && \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_IntisZacT_d [0]));
  
  /* mux (Ty Go,
     Ty MyDTInt_Int_Int) : (call_map''_map''_Int_Int_Int_unlockFork3,Go) [(call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_IntgacU,MyDTInt_Int_Int)] > (call_map''_map''_Int_Int_Int_goMux3,MyDTInt_Int_Int) */
  assign \call_map''_map''_Int_Int_Int_goMux3_d  = (\call_map''_map''_Int_Int_Int_unlockFork3_d [0] && \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_IntgacU_d [0]);
  assign \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_IntgacU_r  = (\call_map''_map''_Int_Int_Int_goMux3_r  && (\call_map''_map''_Int_Int_Int_unlockFork3_d [0] && \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_IntgacU_d [0]));
  assign \call_map''_map''_Int_Int_Int_unlockFork3_r  = (\call_map''_map''_Int_Int_Int_goMux3_r  && (\call_map''_map''_Int_Int_Int_unlockFork3_d [0] && \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_IntgacU_d [0]));
  
  /* mux (Ty Go,
     Ty Int) : (call_map''_map''_Int_Int_Int_unlockFork4,Go) [(call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Intv'acV,Int)] > (call_map''_map''_Int_Int_Int_goMux4,Int) */
  assign \call_map''_map''_Int_Int_Int_goMux4_d  = {\call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Intv'acV_d [32:1],
                                                    (\call_map''_map''_Int_Int_Int_unlockFork4_d [0] && \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Intv'acV_d [0])};
  assign \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Intv'acV_r  = (\call_map''_map''_Int_Int_Int_goMux4_r  && (\call_map''_map''_Int_Int_Int_unlockFork4_d [0] && \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Intv'acV_d [0]));
  assign \call_map''_map''_Int_Int_Int_unlockFork4_r  = (\call_map''_map''_Int_Int_Int_goMux4_r  && (\call_map''_map''_Int_Int_Int_unlockFork4_d [0] && \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Intv'acV_d [0]));
  
  /* mux (Ty Go,
     Ty Pointer_QTree_Int) : (call_map''_map''_Int_Int_Int_unlockFork5,Go) [(call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_IntmacW,Pointer_QTree_Int)] > (call_map''_map''_Int_Int_Int_goMux5,Pointer_QTree_Int) */
  assign \call_map''_map''_Int_Int_Int_goMux5_d  = {\call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_IntmacW_d [16:1],
                                                    (\call_map''_map''_Int_Int_Int_unlockFork5_d [0] && \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_IntmacW_d [0])};
  assign \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_IntmacW_r  = (\call_map''_map''_Int_Int_Int_goMux5_r  && (\call_map''_map''_Int_Int_Int_unlockFork5_d [0] && \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_IntmacW_d [0]));
  assign \call_map''_map''_Int_Int_Int_unlockFork5_r  = (\call_map''_map''_Int_Int_Int_goMux5_r  && (\call_map''_map''_Int_Int_Int_unlockFork5_d [0] && \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_IntmacW_d [0]));
  
  /* mux (Ty Go,
     Ty Pointer_CTmap''_map''_Int_Int_Int) : (call_map''_map''_Int_Int_Int_unlockFork6,Go) [(call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Intsc_0_3,Pointer_CTmap''_map''_Int_Int_Int)] > (call_map''_map''_Int_Int_Int_goMux6,Pointer_CTmap''_map''_Int_Int_Int) */
  assign \call_map''_map''_Int_Int_Int_goMux6_d  = {\call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Intsc_0_3_d [16:1],
                                                    (\call_map''_map''_Int_Int_Int_unlockFork6_d [0] && \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Intsc_0_3_d [0])};
  assign \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Intsc_0_3_r  = (\call_map''_map''_Int_Int_Int_goMux6_r  && (\call_map''_map''_Int_Int_Int_unlockFork6_d [0] && \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Intsc_0_3_d [0]));
  assign \call_map''_map''_Int_Int_Int_unlockFork6_r  = (\call_map''_map''_Int_Int_Int_goMux6_r  && (\call_map''_map''_Int_Int_Int_unlockFork6_d [0] && \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Intsc_0_3_d [0]));
  
  /* sink (Ty Int) : (es_0_1I#,Int) > */
  assign {\es_0_1I#_r , \es_0_1I#_dout } = {\es_0_1I#_rout ,
                                            \es_0_1I#_d };
  
  /* buf (Ty Int) : (es_0_2_1I#_mux_mux,Int) > (applyfnInt_Int_5_resbuf,Int) */
  Int_t \es_0_2_1I#_mux_mux_bufchan_d ;
  logic \es_0_2_1I#_mux_mux_bufchan_r ;
  assign \es_0_2_1I#_mux_mux_r  = ((! \es_0_2_1I#_mux_mux_bufchan_d [0]) || \es_0_2_1I#_mux_mux_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \es_0_2_1I#_mux_mux_bufchan_d  <= {32'd0, 1'd0};
    else
      if (\es_0_2_1I#_mux_mux_r )
        \es_0_2_1I#_mux_mux_bufchan_d  <= \es_0_2_1I#_mux_mux_d ;
  Int_t \es_0_2_1I#_mux_mux_bufchan_buf ;
  assign \es_0_2_1I#_mux_mux_bufchan_r  = (! \es_0_2_1I#_mux_mux_bufchan_buf [0]);
  assign applyfnInt_Int_5_resbuf_d = (\es_0_2_1I#_mux_mux_bufchan_buf [0] ? \es_0_2_1I#_mux_mux_bufchan_buf  :
                                      \es_0_2_1I#_mux_mux_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \es_0_2_1I#_mux_mux_bufchan_buf  <= {32'd0, 1'd0};
    else
      if ((applyfnInt_Int_5_resbuf_r && \es_0_2_1I#_mux_mux_bufchan_buf [0]))
        \es_0_2_1I#_mux_mux_bufchan_buf  <= {32'd0, 1'd0};
      else if (((! applyfnInt_Int_5_resbuf_r) && (! \es_0_2_1I#_mux_mux_bufchan_buf [0])))
        \es_0_2_1I#_mux_mux_bufchan_buf  <= \es_0_2_1I#_mux_mux_bufchan_d ;
  
  /* buf (Ty Int) : (es_0_3_1I#_mux_mux_mux,Int) > (applyfnInt_Int_Int_5_resbuf,Int) */
  Int_t \es_0_3_1I#_mux_mux_mux_bufchan_d ;
  logic \es_0_3_1I#_mux_mux_mux_bufchan_r ;
  assign \es_0_3_1I#_mux_mux_mux_r  = ((! \es_0_3_1I#_mux_mux_mux_bufchan_d [0]) || \es_0_3_1I#_mux_mux_mux_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \es_0_3_1I#_mux_mux_mux_bufchan_d  <= {32'd0, 1'd0};
    else
      if (\es_0_3_1I#_mux_mux_mux_r )
        \es_0_3_1I#_mux_mux_mux_bufchan_d  <= \es_0_3_1I#_mux_mux_mux_d ;
  Int_t \es_0_3_1I#_mux_mux_mux_bufchan_buf ;
  assign \es_0_3_1I#_mux_mux_mux_bufchan_r  = (! \es_0_3_1I#_mux_mux_mux_bufchan_buf [0]);
  assign applyfnInt_Int_Int_5_resbuf_d = (\es_0_3_1I#_mux_mux_mux_bufchan_buf [0] ? \es_0_3_1I#_mux_mux_mux_bufchan_buf  :
                                          \es_0_3_1I#_mux_mux_mux_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \es_0_3_1I#_mux_mux_mux_bufchan_buf  <= {32'd0, 1'd0};
    else
      if ((applyfnInt_Int_Int_5_resbuf_r && \es_0_3_1I#_mux_mux_mux_bufchan_buf [0]))
        \es_0_3_1I#_mux_mux_mux_bufchan_buf  <= {32'd0, 1'd0};
      else if (((! applyfnInt_Int_Int_5_resbuf_r) && (! \es_0_3_1I#_mux_mux_mux_bufchan_buf [0])))
        \es_0_3_1I#_mux_mux_mux_bufchan_buf  <= \es_0_3_1I#_mux_mux_mux_bufchan_d ;
  
  /* demux (Ty MyBool,
       Ty Go) : (es_0_4_1,MyBool) (lizzieLet10_4QVal_Int_3,Go) > [(es_0_4_1MyFalse,Go),
                                                                  (es_0_4_1MyTrue,Go)] */
  logic [1:0] lizzieLet10_4QVal_Int_3_onehotd;
  always_comb
    if ((es_0_4_1_d[0] && lizzieLet10_4QVal_Int_3_d[0]))
      unique case (es_0_4_1_d[1:1])
        1'd0: lizzieLet10_4QVal_Int_3_onehotd = 2'd1;
        1'd1: lizzieLet10_4QVal_Int_3_onehotd = 2'd2;
        default: lizzieLet10_4QVal_Int_3_onehotd = 2'd0;
      endcase
    else lizzieLet10_4QVal_Int_3_onehotd = 2'd0;
  assign es_0_4_1MyFalse_d = lizzieLet10_4QVal_Int_3_onehotd[0];
  assign es_0_4_1MyTrue_d = lizzieLet10_4QVal_Int_3_onehotd[1];
  assign lizzieLet10_4QVal_Int_3_r = (| (lizzieLet10_4QVal_Int_3_onehotd & {es_0_4_1MyTrue_r,
                                                                            es_0_4_1MyFalse_r}));
  assign es_0_4_1_r = lizzieLet10_4QVal_Int_3_r;
  
  /* buf (Ty Go) : (es_0_4_1MyFalse,Go) > (es_0_4_1MyFalse_1_argbuf,Go) */
  Go_t es_0_4_1MyFalse_bufchan_d;
  logic es_0_4_1MyFalse_bufchan_r;
  assign es_0_4_1MyFalse_r = ((! es_0_4_1MyFalse_bufchan_d[0]) || es_0_4_1MyFalse_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_0_4_1MyFalse_bufchan_d <= 1'd0;
    else
      if (es_0_4_1MyFalse_r)
        es_0_4_1MyFalse_bufchan_d <= es_0_4_1MyFalse_d;
  Go_t es_0_4_1MyFalse_bufchan_buf;
  assign es_0_4_1MyFalse_bufchan_r = (! es_0_4_1MyFalse_bufchan_buf[0]);
  assign es_0_4_1MyFalse_1_argbuf_d = (es_0_4_1MyFalse_bufchan_buf[0] ? es_0_4_1MyFalse_bufchan_buf :
                                       es_0_4_1MyFalse_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_0_4_1MyFalse_bufchan_buf <= 1'd0;
    else
      if ((es_0_4_1MyFalse_1_argbuf_r && es_0_4_1MyFalse_bufchan_buf[0]))
        es_0_4_1MyFalse_bufchan_buf <= 1'd0;
      else if (((! es_0_4_1MyFalse_1_argbuf_r) && (! es_0_4_1MyFalse_bufchan_buf[0])))
        es_0_4_1MyFalse_bufchan_buf <= es_0_4_1MyFalse_bufchan_d;
  
  /* fork (Ty Go) : (es_0_4_1MyTrue,Go) > [(es_0_4_1MyTrue_1,Go),
                                      (es_0_4_1MyTrue_2,Go)] */
  logic [1:0] es_0_4_1MyTrue_emitted;
  logic [1:0] es_0_4_1MyTrue_done;
  assign es_0_4_1MyTrue_1_d = (es_0_4_1MyTrue_d[0] && (! es_0_4_1MyTrue_emitted[0]));
  assign es_0_4_1MyTrue_2_d = (es_0_4_1MyTrue_d[0] && (! es_0_4_1MyTrue_emitted[1]));
  assign es_0_4_1MyTrue_done = (es_0_4_1MyTrue_emitted | ({es_0_4_1MyTrue_2_d[0],
                                                           es_0_4_1MyTrue_1_d[0]} & {es_0_4_1MyTrue_2_r,
                                                                                     es_0_4_1MyTrue_1_r}));
  assign es_0_4_1MyTrue_r = (& es_0_4_1MyTrue_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_0_4_1MyTrue_emitted <= 2'd0;
    else
      es_0_4_1MyTrue_emitted <= (es_0_4_1MyTrue_r ? 2'd0 :
                                 es_0_4_1MyTrue_done);
  
  /* dcon (Ty QTree_Int,
      Dcon QNone_Int) : [(es_0_4_1MyTrue_1,Go)] > (es_0_4_1MyTrue_1QNone_Int,QTree_Int) */
  assign es_0_4_1MyTrue_1QNone_Int_d = QNone_Int_dc((& {es_0_4_1MyTrue_1_d[0]}), es_0_4_1MyTrue_1_d);
  assign {es_0_4_1MyTrue_1_r} = {1 {(es_0_4_1MyTrue_1QNone_Int_r && es_0_4_1MyTrue_1QNone_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (es_0_4_1MyTrue_1QNone_Int,QTree_Int) > (lizzieLet13_1_1_argbuf,QTree_Int) */
  QTree_Int_t es_0_4_1MyTrue_1QNone_Int_bufchan_d;
  logic es_0_4_1MyTrue_1QNone_Int_bufchan_r;
  assign es_0_4_1MyTrue_1QNone_Int_r = ((! es_0_4_1MyTrue_1QNone_Int_bufchan_d[0]) || es_0_4_1MyTrue_1QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_0_4_1MyTrue_1QNone_Int_bufchan_d <= {66'd0, 1'd0};
    else
      if (es_0_4_1MyTrue_1QNone_Int_r)
        es_0_4_1MyTrue_1QNone_Int_bufchan_d <= es_0_4_1MyTrue_1QNone_Int_d;
  QTree_Int_t es_0_4_1MyTrue_1QNone_Int_bufchan_buf;
  assign es_0_4_1MyTrue_1QNone_Int_bufchan_r = (! es_0_4_1MyTrue_1QNone_Int_bufchan_buf[0]);
  assign lizzieLet13_1_1_argbuf_d = (es_0_4_1MyTrue_1QNone_Int_bufchan_buf[0] ? es_0_4_1MyTrue_1QNone_Int_bufchan_buf :
                                     es_0_4_1MyTrue_1QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_0_4_1MyTrue_1QNone_Int_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((lizzieLet13_1_1_argbuf_r && es_0_4_1MyTrue_1QNone_Int_bufchan_buf[0]))
        es_0_4_1MyTrue_1QNone_Int_bufchan_buf <= {66'd0, 1'd0};
      else if (((! lizzieLet13_1_1_argbuf_r) && (! es_0_4_1MyTrue_1QNone_Int_bufchan_buf[0])))
        es_0_4_1MyTrue_1QNone_Int_bufchan_buf <= es_0_4_1MyTrue_1QNone_Int_bufchan_d;
  
  /* buf (Ty Go) : (es_0_4_1MyTrue_2,Go) > (es_0_4_1MyTrue_2_argbuf,Go) */
  Go_t es_0_4_1MyTrue_2_bufchan_d;
  logic es_0_4_1MyTrue_2_bufchan_r;
  assign es_0_4_1MyTrue_2_r = ((! es_0_4_1MyTrue_2_bufchan_d[0]) || es_0_4_1MyTrue_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_0_4_1MyTrue_2_bufchan_d <= 1'd0;
    else
      if (es_0_4_1MyTrue_2_r)
        es_0_4_1MyTrue_2_bufchan_d <= es_0_4_1MyTrue_2_d;
  Go_t es_0_4_1MyTrue_2_bufchan_buf;
  assign es_0_4_1MyTrue_2_bufchan_r = (! es_0_4_1MyTrue_2_bufchan_buf[0]);
  assign es_0_4_1MyTrue_2_argbuf_d = (es_0_4_1MyTrue_2_bufchan_buf[0] ? es_0_4_1MyTrue_2_bufchan_buf :
                                      es_0_4_1MyTrue_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_0_4_1MyTrue_2_bufchan_buf <= 1'd0;
    else
      if ((es_0_4_1MyTrue_2_argbuf_r && es_0_4_1MyTrue_2_bufchan_buf[0]))
        es_0_4_1MyTrue_2_bufchan_buf <= 1'd0;
      else if (((! es_0_4_1MyTrue_2_argbuf_r) && (! es_0_4_1MyTrue_2_bufchan_buf[0])))
        es_0_4_1MyTrue_2_bufchan_buf <= es_0_4_1MyTrue_2_bufchan_d;
  
  /* demux (Ty MyBool,
       Ty Pointer_CTmain_map'_Int_Int) : (es_0_4_2,MyBool) (lizzieLet10_6QVal_Int,Pointer_CTmain_map'_Int_Int) > [(es_0_4_2MyFalse,Pointer_CTmain_map'_Int_Int),
                                                                                                                  (es_0_4_2MyTrue,Pointer_CTmain_map'_Int_Int)] */
  logic [1:0] lizzieLet10_6QVal_Int_onehotd;
  always_comb
    if ((es_0_4_2_d[0] && lizzieLet10_6QVal_Int_d[0]))
      unique case (es_0_4_2_d[1:1])
        1'd0: lizzieLet10_6QVal_Int_onehotd = 2'd1;
        1'd1: lizzieLet10_6QVal_Int_onehotd = 2'd2;
        default: lizzieLet10_6QVal_Int_onehotd = 2'd0;
      endcase
    else lizzieLet10_6QVal_Int_onehotd = 2'd0;
  assign es_0_4_2MyFalse_d = {lizzieLet10_6QVal_Int_d[16:1],
                              lizzieLet10_6QVal_Int_onehotd[0]};
  assign es_0_4_2MyTrue_d = {lizzieLet10_6QVal_Int_d[16:1],
                             lizzieLet10_6QVal_Int_onehotd[1]};
  assign lizzieLet10_6QVal_Int_r = (| (lizzieLet10_6QVal_Int_onehotd & {es_0_4_2MyTrue_r,
                                                                        es_0_4_2MyFalse_r}));
  assign es_0_4_2_r = lizzieLet10_6QVal_Int_r;
  
  /* buf (Ty Pointer_CTmain_map'_Int_Int) : (es_0_4_2MyFalse,Pointer_CTmain_map'_Int_Int) > (es_0_4_2MyFalse_1_argbuf,Pointer_CTmain_map'_Int_Int) */
  \Pointer_CTmain_map'_Int_Int_t  es_0_4_2MyFalse_bufchan_d;
  logic es_0_4_2MyFalse_bufchan_r;
  assign es_0_4_2MyFalse_r = ((! es_0_4_2MyFalse_bufchan_d[0]) || es_0_4_2MyFalse_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_0_4_2MyFalse_bufchan_d <= {16'd0, 1'd0};
    else
      if (es_0_4_2MyFalse_r)
        es_0_4_2MyFalse_bufchan_d <= es_0_4_2MyFalse_d;
  \Pointer_CTmain_map'_Int_Int_t  es_0_4_2MyFalse_bufchan_buf;
  assign es_0_4_2MyFalse_bufchan_r = (! es_0_4_2MyFalse_bufchan_buf[0]);
  assign es_0_4_2MyFalse_1_argbuf_d = (es_0_4_2MyFalse_bufchan_buf[0] ? es_0_4_2MyFalse_bufchan_buf :
                                       es_0_4_2MyFalse_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_0_4_2MyFalse_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((es_0_4_2MyFalse_1_argbuf_r && es_0_4_2MyFalse_bufchan_buf[0]))
        es_0_4_2MyFalse_bufchan_buf <= {16'd0, 1'd0};
      else if (((! es_0_4_2MyFalse_1_argbuf_r) && (! es_0_4_2MyFalse_bufchan_buf[0])))
        es_0_4_2MyFalse_bufchan_buf <= es_0_4_2MyFalse_bufchan_d;
  
  /* buf (Ty Pointer_CTmain_map'_Int_Int) : (es_0_4_2MyTrue,Pointer_CTmain_map'_Int_Int) > (es_0_4_2MyTrue_1_argbuf,Pointer_CTmain_map'_Int_Int) */
  \Pointer_CTmain_map'_Int_Int_t  es_0_4_2MyTrue_bufchan_d;
  logic es_0_4_2MyTrue_bufchan_r;
  assign es_0_4_2MyTrue_r = ((! es_0_4_2MyTrue_bufchan_d[0]) || es_0_4_2MyTrue_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_0_4_2MyTrue_bufchan_d <= {16'd0, 1'd0};
    else
      if (es_0_4_2MyTrue_r) es_0_4_2MyTrue_bufchan_d <= es_0_4_2MyTrue_d;
  \Pointer_CTmain_map'_Int_Int_t  es_0_4_2MyTrue_bufchan_buf;
  assign es_0_4_2MyTrue_bufchan_r = (! es_0_4_2MyTrue_bufchan_buf[0]);
  assign es_0_4_2MyTrue_1_argbuf_d = (es_0_4_2MyTrue_bufchan_buf[0] ? es_0_4_2MyTrue_bufchan_buf :
                                      es_0_4_2MyTrue_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_0_4_2MyTrue_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((es_0_4_2MyTrue_1_argbuf_r && es_0_4_2MyTrue_bufchan_buf[0]))
        es_0_4_2MyTrue_bufchan_buf <= {16'd0, 1'd0};
      else if (((! es_0_4_2MyTrue_1_argbuf_r) && (! es_0_4_2MyTrue_bufchan_buf[0])))
        es_0_4_2MyTrue_bufchan_buf <= es_0_4_2MyTrue_bufchan_d;
  
  /* demux (Ty MyBool,
       Ty Int) : (es_0_4_3,MyBool) (xacr_2,Int) > [(es_0_4_3MyFalse,Int),
                                                   (_34,Int)] */
  logic [1:0] xacr_2_onehotd;
  always_comb
    if ((es_0_4_3_d[0] && xacr_2_d[0]))
      unique case (es_0_4_3_d[1:1])
        1'd0: xacr_2_onehotd = 2'd1;
        1'd1: xacr_2_onehotd = 2'd2;
        default: xacr_2_onehotd = 2'd0;
      endcase
    else xacr_2_onehotd = 2'd0;
  assign es_0_4_3MyFalse_d = {xacr_2_d[32:1], xacr_2_onehotd[0]};
  assign _34_d = {xacr_2_d[32:1], xacr_2_onehotd[1]};
  assign xacr_2_r = (| (xacr_2_onehotd & {_34_r,
                                          es_0_4_3MyFalse_r}));
  assign es_0_4_3_r = xacr_2_r;
  
  /* dcon (Ty QTree_Int,
      Dcon QVal_Int) : [(es_0_4_3MyFalse,Int)] > (es_0_4_3MyFalse_1QVal_Int,QTree_Int) */
  assign es_0_4_3MyFalse_1QVal_Int_d = QVal_Int_dc((& {es_0_4_3MyFalse_d[0]}), es_0_4_3MyFalse_d);
  assign {es_0_4_3MyFalse_r} = {1 {(es_0_4_3MyFalse_1QVal_Int_r && es_0_4_3MyFalse_1QVal_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (es_0_4_3MyFalse_1QVal_Int,QTree_Int) > (lizzieLet12_1_1_argbuf,QTree_Int) */
  QTree_Int_t es_0_4_3MyFalse_1QVal_Int_bufchan_d;
  logic es_0_4_3MyFalse_1QVal_Int_bufchan_r;
  assign es_0_4_3MyFalse_1QVal_Int_r = ((! es_0_4_3MyFalse_1QVal_Int_bufchan_d[0]) || es_0_4_3MyFalse_1QVal_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_0_4_3MyFalse_1QVal_Int_bufchan_d <= {66'd0, 1'd0};
    else
      if (es_0_4_3MyFalse_1QVal_Int_r)
        es_0_4_3MyFalse_1QVal_Int_bufchan_d <= es_0_4_3MyFalse_1QVal_Int_d;
  QTree_Int_t es_0_4_3MyFalse_1QVal_Int_bufchan_buf;
  assign es_0_4_3MyFalse_1QVal_Int_bufchan_r = (! es_0_4_3MyFalse_1QVal_Int_bufchan_buf[0]);
  assign lizzieLet12_1_1_argbuf_d = (es_0_4_3MyFalse_1QVal_Int_bufchan_buf[0] ? es_0_4_3MyFalse_1QVal_Int_bufchan_buf :
                                     es_0_4_3MyFalse_1QVal_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_0_4_3MyFalse_1QVal_Int_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((lizzieLet12_1_1_argbuf_r && es_0_4_3MyFalse_1QVal_Int_bufchan_buf[0]))
        es_0_4_3MyFalse_1QVal_Int_bufchan_buf <= {66'd0, 1'd0};
      else if (((! lizzieLet12_1_1_argbuf_r) && (! es_0_4_3MyFalse_1QVal_Int_bufchan_buf[0])))
        es_0_4_3MyFalse_1QVal_Int_bufchan_buf <= es_0_4_3MyFalse_1QVal_Int_bufchan_d;
  
  /* demux (Ty MyBool,
       Ty Go) : (es_0_5_1,MyBool) (lizzieLet16_1_4QVal_Int_2,Go) > [(es_0_5_1MyFalse,Go),
                                                                    (es_0_5_1MyTrue,Go)] */
  logic [1:0] lizzieLet16_1_4QVal_Int_2_onehotd;
  always_comb
    if ((es_0_5_1_d[0] && lizzieLet16_1_4QVal_Int_2_d[0]))
      unique case (es_0_5_1_d[1:1])
        1'd0: lizzieLet16_1_4QVal_Int_2_onehotd = 2'd1;
        1'd1: lizzieLet16_1_4QVal_Int_2_onehotd = 2'd2;
        default: lizzieLet16_1_4QVal_Int_2_onehotd = 2'd0;
      endcase
    else lizzieLet16_1_4QVal_Int_2_onehotd = 2'd0;
  assign es_0_5_1MyFalse_d = lizzieLet16_1_4QVal_Int_2_onehotd[0];
  assign es_0_5_1MyTrue_d = lizzieLet16_1_4QVal_Int_2_onehotd[1];
  assign lizzieLet16_1_4QVal_Int_2_r = (| (lizzieLet16_1_4QVal_Int_2_onehotd & {es_0_5_1MyTrue_r,
                                                                                es_0_5_1MyFalse_r}));
  assign es_0_5_1_r = lizzieLet16_1_4QVal_Int_2_r;
  
  /* buf (Ty Go) : (es_0_5_1MyFalse,Go) > (es_0_5_1MyFalse_1_argbuf,Go) */
  Go_t es_0_5_1MyFalse_bufchan_d;
  logic es_0_5_1MyFalse_bufchan_r;
  assign es_0_5_1MyFalse_r = ((! es_0_5_1MyFalse_bufchan_d[0]) || es_0_5_1MyFalse_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_0_5_1MyFalse_bufchan_d <= 1'd0;
    else
      if (es_0_5_1MyFalse_r)
        es_0_5_1MyFalse_bufchan_d <= es_0_5_1MyFalse_d;
  Go_t es_0_5_1MyFalse_bufchan_buf;
  assign es_0_5_1MyFalse_bufchan_r = (! es_0_5_1MyFalse_bufchan_buf[0]);
  assign es_0_5_1MyFalse_1_argbuf_d = (es_0_5_1MyFalse_bufchan_buf[0] ? es_0_5_1MyFalse_bufchan_buf :
                                       es_0_5_1MyFalse_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_0_5_1MyFalse_bufchan_buf <= 1'd0;
    else
      if ((es_0_5_1MyFalse_1_argbuf_r && es_0_5_1MyFalse_bufchan_buf[0]))
        es_0_5_1MyFalse_bufchan_buf <= 1'd0;
      else if (((! es_0_5_1MyFalse_1_argbuf_r) && (! es_0_5_1MyFalse_bufchan_buf[0])))
        es_0_5_1MyFalse_bufchan_buf <= es_0_5_1MyFalse_bufchan_d;
  
  /* fork (Ty Go) : (es_0_5_1MyTrue,Go) > [(es_0_5_1MyTrue_1,Go),
                                      (es_0_5_1MyTrue_2,Go)] */
  logic [1:0] es_0_5_1MyTrue_emitted;
  logic [1:0] es_0_5_1MyTrue_done;
  assign es_0_5_1MyTrue_1_d = (es_0_5_1MyTrue_d[0] && (! es_0_5_1MyTrue_emitted[0]));
  assign es_0_5_1MyTrue_2_d = (es_0_5_1MyTrue_d[0] && (! es_0_5_1MyTrue_emitted[1]));
  assign es_0_5_1MyTrue_done = (es_0_5_1MyTrue_emitted | ({es_0_5_1MyTrue_2_d[0],
                                                           es_0_5_1MyTrue_1_d[0]} & {es_0_5_1MyTrue_2_r,
                                                                                     es_0_5_1MyTrue_1_r}));
  assign es_0_5_1MyTrue_r = (& es_0_5_1MyTrue_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_0_5_1MyTrue_emitted <= 2'd0;
    else
      es_0_5_1MyTrue_emitted <= (es_0_5_1MyTrue_r ? 2'd0 :
                                 es_0_5_1MyTrue_done);
  
  /* dcon (Ty QTree_Int,
      Dcon QNone_Int) : [(es_0_5_1MyTrue_1,Go)] > (es_0_5_1MyTrue_1QNone_Int,QTree_Int) */
  assign es_0_5_1MyTrue_1QNone_Int_d = QNone_Int_dc((& {es_0_5_1MyTrue_1_d[0]}), es_0_5_1MyTrue_1_d);
  assign {es_0_5_1MyTrue_1_r} = {1 {(es_0_5_1MyTrue_1QNone_Int_r && es_0_5_1MyTrue_1QNone_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (es_0_5_1MyTrue_1QNone_Int,QTree_Int) > (lizzieLet19_1_argbuf,QTree_Int) */
  QTree_Int_t es_0_5_1MyTrue_1QNone_Int_bufchan_d;
  logic es_0_5_1MyTrue_1QNone_Int_bufchan_r;
  assign es_0_5_1MyTrue_1QNone_Int_r = ((! es_0_5_1MyTrue_1QNone_Int_bufchan_d[0]) || es_0_5_1MyTrue_1QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_0_5_1MyTrue_1QNone_Int_bufchan_d <= {66'd0, 1'd0};
    else
      if (es_0_5_1MyTrue_1QNone_Int_r)
        es_0_5_1MyTrue_1QNone_Int_bufchan_d <= es_0_5_1MyTrue_1QNone_Int_d;
  QTree_Int_t es_0_5_1MyTrue_1QNone_Int_bufchan_buf;
  assign es_0_5_1MyTrue_1QNone_Int_bufchan_r = (! es_0_5_1MyTrue_1QNone_Int_bufchan_buf[0]);
  assign lizzieLet19_1_argbuf_d = (es_0_5_1MyTrue_1QNone_Int_bufchan_buf[0] ? es_0_5_1MyTrue_1QNone_Int_bufchan_buf :
                                   es_0_5_1MyTrue_1QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_0_5_1MyTrue_1QNone_Int_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((lizzieLet19_1_argbuf_r && es_0_5_1MyTrue_1QNone_Int_bufchan_buf[0]))
        es_0_5_1MyTrue_1QNone_Int_bufchan_buf <= {66'd0, 1'd0};
      else if (((! lizzieLet19_1_argbuf_r) && (! es_0_5_1MyTrue_1QNone_Int_bufchan_buf[0])))
        es_0_5_1MyTrue_1QNone_Int_bufchan_buf <= es_0_5_1MyTrue_1QNone_Int_bufchan_d;
  
  /* buf (Ty Go) : (es_0_5_1MyTrue_2,Go) > (es_0_5_1MyTrue_2_argbuf,Go) */
  Go_t es_0_5_1MyTrue_2_bufchan_d;
  logic es_0_5_1MyTrue_2_bufchan_r;
  assign es_0_5_1MyTrue_2_r = ((! es_0_5_1MyTrue_2_bufchan_d[0]) || es_0_5_1MyTrue_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_0_5_1MyTrue_2_bufchan_d <= 1'd0;
    else
      if (es_0_5_1MyTrue_2_r)
        es_0_5_1MyTrue_2_bufchan_d <= es_0_5_1MyTrue_2_d;
  Go_t es_0_5_1MyTrue_2_bufchan_buf;
  assign es_0_5_1MyTrue_2_bufchan_r = (! es_0_5_1MyTrue_2_bufchan_buf[0]);
  assign es_0_5_1MyTrue_2_argbuf_d = (es_0_5_1MyTrue_2_bufchan_buf[0] ? es_0_5_1MyTrue_2_bufchan_buf :
                                      es_0_5_1MyTrue_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_0_5_1MyTrue_2_bufchan_buf <= 1'd0;
    else
      if ((es_0_5_1MyTrue_2_argbuf_r && es_0_5_1MyTrue_2_bufchan_buf[0]))
        es_0_5_1MyTrue_2_bufchan_buf <= 1'd0;
      else if (((! es_0_5_1MyTrue_2_argbuf_r) && (! es_0_5_1MyTrue_2_bufchan_buf[0])))
        es_0_5_1MyTrue_2_bufchan_buf <= es_0_5_1MyTrue_2_bufchan_d;
  
  /* demux (Ty MyBool,
       Ty Pointer_CTmap''_map''_Int_Int_Int) : (es_0_5_2,MyBool) (lizzieLet16_1_6QVal_Int,Pointer_CTmap''_map''_Int_Int_Int) > [(es_0_5_2MyFalse,Pointer_CTmap''_map''_Int_Int_Int),
                                                                                                                                (es_0_5_2MyTrue,Pointer_CTmap''_map''_Int_Int_Int)] */
  logic [1:0] lizzieLet16_1_6QVal_Int_onehotd;
  always_comb
    if ((es_0_5_2_d[0] && lizzieLet16_1_6QVal_Int_d[0]))
      unique case (es_0_5_2_d[1:1])
        1'd0: lizzieLet16_1_6QVal_Int_onehotd = 2'd1;
        1'd1: lizzieLet16_1_6QVal_Int_onehotd = 2'd2;
        default: lizzieLet16_1_6QVal_Int_onehotd = 2'd0;
      endcase
    else lizzieLet16_1_6QVal_Int_onehotd = 2'd0;
  assign es_0_5_2MyFalse_d = {lizzieLet16_1_6QVal_Int_d[16:1],
                              lizzieLet16_1_6QVal_Int_onehotd[0]};
  assign es_0_5_2MyTrue_d = {lizzieLet16_1_6QVal_Int_d[16:1],
                             lizzieLet16_1_6QVal_Int_onehotd[1]};
  assign lizzieLet16_1_6QVal_Int_r = (| (lizzieLet16_1_6QVal_Int_onehotd & {es_0_5_2MyTrue_r,
                                                                            es_0_5_2MyFalse_r}));
  assign es_0_5_2_r = lizzieLet16_1_6QVal_Int_r;
  
  /* buf (Ty Pointer_CTmap''_map''_Int_Int_Int) : (es_0_5_2MyFalse,Pointer_CTmap''_map''_Int_Int_Int) > (es_0_5_2MyFalse_1_argbuf,Pointer_CTmap''_map''_Int_Int_Int) */
  \Pointer_CTmap''_map''_Int_Int_Int_t  es_0_5_2MyFalse_bufchan_d;
  logic es_0_5_2MyFalse_bufchan_r;
  assign es_0_5_2MyFalse_r = ((! es_0_5_2MyFalse_bufchan_d[0]) || es_0_5_2MyFalse_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_0_5_2MyFalse_bufchan_d <= {16'd0, 1'd0};
    else
      if (es_0_5_2MyFalse_r)
        es_0_5_2MyFalse_bufchan_d <= es_0_5_2MyFalse_d;
  \Pointer_CTmap''_map''_Int_Int_Int_t  es_0_5_2MyFalse_bufchan_buf;
  assign es_0_5_2MyFalse_bufchan_r = (! es_0_5_2MyFalse_bufchan_buf[0]);
  assign es_0_5_2MyFalse_1_argbuf_d = (es_0_5_2MyFalse_bufchan_buf[0] ? es_0_5_2MyFalse_bufchan_buf :
                                       es_0_5_2MyFalse_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_0_5_2MyFalse_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((es_0_5_2MyFalse_1_argbuf_r && es_0_5_2MyFalse_bufchan_buf[0]))
        es_0_5_2MyFalse_bufchan_buf <= {16'd0, 1'd0};
      else if (((! es_0_5_2MyFalse_1_argbuf_r) && (! es_0_5_2MyFalse_bufchan_buf[0])))
        es_0_5_2MyFalse_bufchan_buf <= es_0_5_2MyFalse_bufchan_d;
  
  /* buf (Ty Pointer_CTmap''_map''_Int_Int_Int) : (es_0_5_2MyTrue,Pointer_CTmap''_map''_Int_Int_Int) > (es_0_5_2MyTrue_1_argbuf,Pointer_CTmap''_map''_Int_Int_Int) */
  \Pointer_CTmap''_map''_Int_Int_Int_t  es_0_5_2MyTrue_bufchan_d;
  logic es_0_5_2MyTrue_bufchan_r;
  assign es_0_5_2MyTrue_r = ((! es_0_5_2MyTrue_bufchan_d[0]) || es_0_5_2MyTrue_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_0_5_2MyTrue_bufchan_d <= {16'd0, 1'd0};
    else
      if (es_0_5_2MyTrue_r) es_0_5_2MyTrue_bufchan_d <= es_0_5_2MyTrue_d;
  \Pointer_CTmap''_map''_Int_Int_Int_t  es_0_5_2MyTrue_bufchan_buf;
  assign es_0_5_2MyTrue_bufchan_r = (! es_0_5_2MyTrue_bufchan_buf[0]);
  assign es_0_5_2MyTrue_1_argbuf_d = (es_0_5_2MyTrue_bufchan_buf[0] ? es_0_5_2MyTrue_bufchan_buf :
                                      es_0_5_2MyTrue_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_0_5_2MyTrue_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((es_0_5_2MyTrue_1_argbuf_r && es_0_5_2MyTrue_bufchan_buf[0]))
        es_0_5_2MyTrue_bufchan_buf <= {16'd0, 1'd0};
      else if (((! es_0_5_2MyTrue_1_argbuf_r) && (! es_0_5_2MyTrue_bufchan_buf[0])))
        es_0_5_2MyTrue_bufchan_buf <= es_0_5_2MyTrue_bufchan_d;
  
  /* demux (Ty MyBool,
       Ty Int) : (es_0_5_3,MyBool) (xacr_1_2,Int) > [(es_0_5_3MyFalse,Int),
                                                     (_33,Int)] */
  logic [1:0] xacr_1_2_onehotd;
  always_comb
    if ((es_0_5_3_d[0] && xacr_1_2_d[0]))
      unique case (es_0_5_3_d[1:1])
        1'd0: xacr_1_2_onehotd = 2'd1;
        1'd1: xacr_1_2_onehotd = 2'd2;
        default: xacr_1_2_onehotd = 2'd0;
      endcase
    else xacr_1_2_onehotd = 2'd0;
  assign es_0_5_3MyFalse_d = {xacr_1_2_d[32:1], xacr_1_2_onehotd[0]};
  assign _33_d = {xacr_1_2_d[32:1], xacr_1_2_onehotd[1]};
  assign xacr_1_2_r = (| (xacr_1_2_onehotd & {_33_r,
                                              es_0_5_3MyFalse_r}));
  assign es_0_5_3_r = xacr_1_2_r;
  
  /* dcon (Ty QTree_Int,
      Dcon QVal_Int) : [(es_0_5_3MyFalse,Int)] > (es_0_5_3MyFalse_1QVal_Int,QTree_Int) */
  assign es_0_5_3MyFalse_1QVal_Int_d = QVal_Int_dc((& {es_0_5_3MyFalse_d[0]}), es_0_5_3MyFalse_d);
  assign {es_0_5_3MyFalse_r} = {1 {(es_0_5_3MyFalse_1QVal_Int_r && es_0_5_3MyFalse_1QVal_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (es_0_5_3MyFalse_1QVal_Int,QTree_Int) > (lizzieLet18_1_argbuf,QTree_Int) */
  QTree_Int_t es_0_5_3MyFalse_1QVal_Int_bufchan_d;
  logic es_0_5_3MyFalse_1QVal_Int_bufchan_r;
  assign es_0_5_3MyFalse_1QVal_Int_r = ((! es_0_5_3MyFalse_1QVal_Int_bufchan_d[0]) || es_0_5_3MyFalse_1QVal_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_0_5_3MyFalse_1QVal_Int_bufchan_d <= {66'd0, 1'd0};
    else
      if (es_0_5_3MyFalse_1QVal_Int_r)
        es_0_5_3MyFalse_1QVal_Int_bufchan_d <= es_0_5_3MyFalse_1QVal_Int_d;
  QTree_Int_t es_0_5_3MyFalse_1QVal_Int_bufchan_buf;
  assign es_0_5_3MyFalse_1QVal_Int_bufchan_r = (! es_0_5_3MyFalse_1QVal_Int_bufchan_buf[0]);
  assign lizzieLet18_1_argbuf_d = (es_0_5_3MyFalse_1QVal_Int_bufchan_buf[0] ? es_0_5_3MyFalse_1QVal_Int_bufchan_buf :
                                   es_0_5_3MyFalse_1QVal_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_0_5_3MyFalse_1QVal_Int_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((lizzieLet18_1_argbuf_r && es_0_5_3MyFalse_1QVal_Int_bufchan_buf[0]))
        es_0_5_3MyFalse_1QVal_Int_bufchan_buf <= {66'd0, 1'd0};
      else if (((! lizzieLet18_1_argbuf_r) && (! es_0_5_3MyFalse_1QVal_Int_bufchan_buf[0])))
        es_0_5_3MyFalse_1QVal_Int_bufchan_buf <= es_0_5_3MyFalse_1QVal_Int_bufchan_d;
  
  /* buf (Ty Int#) : (es_4_1_1lizzieLet25_4Lcall_$wnnz_Int0_1_Add32,Int#) > (contRet_0_1_argbuf,Int#) */
  \Int#_t  es_4_1_1lizzieLet25_4Lcall_$wnnz_Int0_1_Add32_bufchan_d;
  logic es_4_1_1lizzieLet25_4Lcall_$wnnz_Int0_1_Add32_bufchan_r;
  assign es_4_1_1lizzieLet25_4Lcall_$wnnz_Int0_1_Add32_r = ((! es_4_1_1lizzieLet25_4Lcall_$wnnz_Int0_1_Add32_bufchan_d[0]) || es_4_1_1lizzieLet25_4Lcall_$wnnz_Int0_1_Add32_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_4_1_1lizzieLet25_4Lcall_$wnnz_Int0_1_Add32_bufchan_d <= {32'd0,
                                                                  1'd0};
    else
      if (es_4_1_1lizzieLet25_4Lcall_$wnnz_Int0_1_Add32_r)
        es_4_1_1lizzieLet25_4Lcall_$wnnz_Int0_1_Add32_bufchan_d <= es_4_1_1lizzieLet25_4Lcall_$wnnz_Int0_1_Add32_d;
  \Int#_t  es_4_1_1lizzieLet25_4Lcall_$wnnz_Int0_1_Add32_bufchan_buf;
  assign es_4_1_1lizzieLet25_4Lcall_$wnnz_Int0_1_Add32_bufchan_r = (! es_4_1_1lizzieLet25_4Lcall_$wnnz_Int0_1_Add32_bufchan_buf[0]);
  assign contRet_0_1_argbuf_d = (es_4_1_1lizzieLet25_4Lcall_$wnnz_Int0_1_Add32_bufchan_buf[0] ? es_4_1_1lizzieLet25_4Lcall_$wnnz_Int0_1_Add32_bufchan_buf :
                                 es_4_1_1lizzieLet25_4Lcall_$wnnz_Int0_1_Add32_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_4_1_1lizzieLet25_4Lcall_$wnnz_Int0_1_Add32_bufchan_buf <= {32'd0,
                                                                    1'd0};
    else
      if ((contRet_0_1_argbuf_r && es_4_1_1lizzieLet25_4Lcall_$wnnz_Int0_1_Add32_bufchan_buf[0]))
        es_4_1_1lizzieLet25_4Lcall_$wnnz_Int0_1_Add32_bufchan_buf <= {32'd0,
                                                                      1'd0};
      else if (((! contRet_0_1_argbuf_r) && (! es_4_1_1lizzieLet25_4Lcall_$wnnz_Int0_1_Add32_bufchan_buf[0])))
        es_4_1_1lizzieLet25_4Lcall_$wnnz_Int0_1_Add32_bufchan_buf <= es_4_1_1lizzieLet25_4Lcall_$wnnz_Int0_1_Add32_bufchan_d;
  
  /* op_add (Ty Int#) : (es_6_1ww2XwL_1_1_Add32,Int#) (lizzieLet25_4Lcall_$wnnz_Int0,Int#) > (es_4_1_1lizzieLet25_4Lcall_$wnnz_Int0_1_Add32,Int#) */
  assign es_4_1_1lizzieLet25_4Lcall_$wnnz_Int0_1_Add32_d = {(es_6_1ww2XwL_1_1_Add32_d[32:1] + lizzieLet25_4Lcall_$wnnz_Int0_d[32:1]),
                                                            (es_6_1ww2XwL_1_1_Add32_d[0] && lizzieLet25_4Lcall_$wnnz_Int0_d[0])};
  assign {es_6_1ww2XwL_1_1_Add32_r,
          lizzieLet25_4Lcall_$wnnz_Int0_r} = {2 {(es_4_1_1lizzieLet25_4Lcall_$wnnz_Int0_1_Add32_r && es_4_1_1lizzieLet25_4Lcall_$wnnz_Int0_1_Add32_d[0])}};
  
  /* buf (Ty MyDTInt_Int) : (gacM_2_2,MyDTInt_Int) > (gacM_2_2_argbuf,MyDTInt_Int) */
  MyDTInt_Int_t gacM_2_2_bufchan_d;
  logic gacM_2_2_bufchan_r;
  assign gacM_2_2_r = ((! gacM_2_2_bufchan_d[0]) || gacM_2_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) gacM_2_2_bufchan_d <= 1'd0;
    else if (gacM_2_2_r) gacM_2_2_bufchan_d <= gacM_2_2_d;
  MyDTInt_Int_t gacM_2_2_bufchan_buf;
  assign gacM_2_2_bufchan_r = (! gacM_2_2_bufchan_buf[0]);
  assign gacM_2_2_argbuf_d = (gacM_2_2_bufchan_buf[0] ? gacM_2_2_bufchan_buf :
                              gacM_2_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) gacM_2_2_bufchan_buf <= 1'd0;
    else
      if ((gacM_2_2_argbuf_r && gacM_2_2_bufchan_buf[0]))
        gacM_2_2_bufchan_buf <= 1'd0;
      else if (((! gacM_2_2_argbuf_r) && (! gacM_2_2_bufchan_buf[0])))
        gacM_2_2_bufchan_buf <= gacM_2_2_bufchan_d;
  
  /* fork (Ty MyDTInt_Int) : (gacM_2_destruct,MyDTInt_Int) > [(gacM_2_1,MyDTInt_Int),
                                                         (gacM_2_2,MyDTInt_Int)] */
  logic [1:0] gacM_2_destruct_emitted;
  logic [1:0] gacM_2_destruct_done;
  assign gacM_2_1_d = (gacM_2_destruct_d[0] && (! gacM_2_destruct_emitted[0]));
  assign gacM_2_2_d = (gacM_2_destruct_d[0] && (! gacM_2_destruct_emitted[1]));
  assign gacM_2_destruct_done = (gacM_2_destruct_emitted | ({gacM_2_2_d[0],
                                                             gacM_2_1_d[0]} & {gacM_2_2_r,
                                                                               gacM_2_1_r}));
  assign gacM_2_destruct_r = (& gacM_2_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) gacM_2_destruct_emitted <= 2'd0;
    else
      gacM_2_destruct_emitted <= (gacM_2_destruct_r ? 2'd0 :
                                  gacM_2_destruct_done);
  
  /* buf (Ty MyDTInt_Int) : (gacM_3_2,MyDTInt_Int) > (gacM_3_2_argbuf,MyDTInt_Int) */
  MyDTInt_Int_t gacM_3_2_bufchan_d;
  logic gacM_3_2_bufchan_r;
  assign gacM_3_2_r = ((! gacM_3_2_bufchan_d[0]) || gacM_3_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) gacM_3_2_bufchan_d <= 1'd0;
    else if (gacM_3_2_r) gacM_3_2_bufchan_d <= gacM_3_2_d;
  MyDTInt_Int_t gacM_3_2_bufchan_buf;
  assign gacM_3_2_bufchan_r = (! gacM_3_2_bufchan_buf[0]);
  assign gacM_3_2_argbuf_d = (gacM_3_2_bufchan_buf[0] ? gacM_3_2_bufchan_buf :
                              gacM_3_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) gacM_3_2_bufchan_buf <= 1'd0;
    else
      if ((gacM_3_2_argbuf_r && gacM_3_2_bufchan_buf[0]))
        gacM_3_2_bufchan_buf <= 1'd0;
      else if (((! gacM_3_2_argbuf_r) && (! gacM_3_2_bufchan_buf[0])))
        gacM_3_2_bufchan_buf <= gacM_3_2_bufchan_d;
  
  /* fork (Ty MyDTInt_Int) : (gacM_3_destruct,MyDTInt_Int) > [(gacM_3_1,MyDTInt_Int),
                                                         (gacM_3_2,MyDTInt_Int)] */
  logic [1:0] gacM_3_destruct_emitted;
  logic [1:0] gacM_3_destruct_done;
  assign gacM_3_1_d = (gacM_3_destruct_d[0] && (! gacM_3_destruct_emitted[0]));
  assign gacM_3_2_d = (gacM_3_destruct_d[0] && (! gacM_3_destruct_emitted[1]));
  assign gacM_3_destruct_done = (gacM_3_destruct_emitted | ({gacM_3_2_d[0],
                                                             gacM_3_1_d[0]} & {gacM_3_2_r,
                                                                               gacM_3_1_r}));
  assign gacM_3_destruct_r = (& gacM_3_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) gacM_3_destruct_emitted <= 2'd0;
    else
      gacM_3_destruct_emitted <= (gacM_3_destruct_r ? 2'd0 :
                                  gacM_3_destruct_done);
  
  /* buf (Ty MyDTInt_Int) : (gacM_4_destruct,MyDTInt_Int) > (gacM_4_1_argbuf,MyDTInt_Int) */
  MyDTInt_Int_t gacM_4_destruct_bufchan_d;
  logic gacM_4_destruct_bufchan_r;
  assign gacM_4_destruct_r = ((! gacM_4_destruct_bufchan_d[0]) || gacM_4_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) gacM_4_destruct_bufchan_d <= 1'd0;
    else
      if (gacM_4_destruct_r)
        gacM_4_destruct_bufchan_d <= gacM_4_destruct_d;
  MyDTInt_Int_t gacM_4_destruct_bufchan_buf;
  assign gacM_4_destruct_bufchan_r = (! gacM_4_destruct_bufchan_buf[0]);
  assign gacM_4_1_argbuf_d = (gacM_4_destruct_bufchan_buf[0] ? gacM_4_destruct_bufchan_buf :
                              gacM_4_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) gacM_4_destruct_bufchan_buf <= 1'd0;
    else
      if ((gacM_4_1_argbuf_r && gacM_4_destruct_bufchan_buf[0]))
        gacM_4_destruct_bufchan_buf <= 1'd0;
      else if (((! gacM_4_1_argbuf_r) && (! gacM_4_destruct_bufchan_buf[0])))
        gacM_4_destruct_bufchan_buf <= gacM_4_destruct_bufchan_d;
  
  /* buf (Ty MyDTInt_Int_Int) : (gacU_2_2,MyDTInt_Int_Int) > (gacU_2_2_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t gacU_2_2_bufchan_d;
  logic gacU_2_2_bufchan_r;
  assign gacU_2_2_r = ((! gacU_2_2_bufchan_d[0]) || gacU_2_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) gacU_2_2_bufchan_d <= 1'd0;
    else if (gacU_2_2_r) gacU_2_2_bufchan_d <= gacU_2_2_d;
  MyDTInt_Int_Int_t gacU_2_2_bufchan_buf;
  assign gacU_2_2_bufchan_r = (! gacU_2_2_bufchan_buf[0]);
  assign gacU_2_2_argbuf_d = (gacU_2_2_bufchan_buf[0] ? gacU_2_2_bufchan_buf :
                              gacU_2_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) gacU_2_2_bufchan_buf <= 1'd0;
    else
      if ((gacU_2_2_argbuf_r && gacU_2_2_bufchan_buf[0]))
        gacU_2_2_bufchan_buf <= 1'd0;
      else if (((! gacU_2_2_argbuf_r) && (! gacU_2_2_bufchan_buf[0])))
        gacU_2_2_bufchan_buf <= gacU_2_2_bufchan_d;
  
  /* fork (Ty MyDTInt_Int_Int) : (gacU_2_destruct,MyDTInt_Int_Int) > [(gacU_2_1,MyDTInt_Int_Int),
                                                                 (gacU_2_2,MyDTInt_Int_Int)] */
  logic [1:0] gacU_2_destruct_emitted;
  logic [1:0] gacU_2_destruct_done;
  assign gacU_2_1_d = (gacU_2_destruct_d[0] && (! gacU_2_destruct_emitted[0]));
  assign gacU_2_2_d = (gacU_2_destruct_d[0] && (! gacU_2_destruct_emitted[1]));
  assign gacU_2_destruct_done = (gacU_2_destruct_emitted | ({gacU_2_2_d[0],
                                                             gacU_2_1_d[0]} & {gacU_2_2_r,
                                                                               gacU_2_1_r}));
  assign gacU_2_destruct_r = (& gacU_2_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) gacU_2_destruct_emitted <= 2'd0;
    else
      gacU_2_destruct_emitted <= (gacU_2_destruct_r ? 2'd0 :
                                  gacU_2_destruct_done);
  
  /* buf (Ty MyDTInt_Int_Int) : (gacU_3_2,MyDTInt_Int_Int) > (gacU_3_2_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t gacU_3_2_bufchan_d;
  logic gacU_3_2_bufchan_r;
  assign gacU_3_2_r = ((! gacU_3_2_bufchan_d[0]) || gacU_3_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) gacU_3_2_bufchan_d <= 1'd0;
    else if (gacU_3_2_r) gacU_3_2_bufchan_d <= gacU_3_2_d;
  MyDTInt_Int_Int_t gacU_3_2_bufchan_buf;
  assign gacU_3_2_bufchan_r = (! gacU_3_2_bufchan_buf[0]);
  assign gacU_3_2_argbuf_d = (gacU_3_2_bufchan_buf[0] ? gacU_3_2_bufchan_buf :
                              gacU_3_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) gacU_3_2_bufchan_buf <= 1'd0;
    else
      if ((gacU_3_2_argbuf_r && gacU_3_2_bufchan_buf[0]))
        gacU_3_2_bufchan_buf <= 1'd0;
      else if (((! gacU_3_2_argbuf_r) && (! gacU_3_2_bufchan_buf[0])))
        gacU_3_2_bufchan_buf <= gacU_3_2_bufchan_d;
  
  /* fork (Ty MyDTInt_Int_Int) : (gacU_3_destruct,MyDTInt_Int_Int) > [(gacU_3_1,MyDTInt_Int_Int),
                                                                 (gacU_3_2,MyDTInt_Int_Int)] */
  logic [1:0] gacU_3_destruct_emitted;
  logic [1:0] gacU_3_destruct_done;
  assign gacU_3_1_d = (gacU_3_destruct_d[0] && (! gacU_3_destruct_emitted[0]));
  assign gacU_3_2_d = (gacU_3_destruct_d[0] && (! gacU_3_destruct_emitted[1]));
  assign gacU_3_destruct_done = (gacU_3_destruct_emitted | ({gacU_3_2_d[0],
                                                             gacU_3_1_d[0]} & {gacU_3_2_r,
                                                                               gacU_3_1_r}));
  assign gacU_3_destruct_r = (& gacU_3_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) gacU_3_destruct_emitted <= 2'd0;
    else
      gacU_3_destruct_emitted <= (gacU_3_destruct_r ? 2'd0 :
                                  gacU_3_destruct_done);
  
  /* buf (Ty MyDTInt_Int_Int) : (gacU_4_destruct,MyDTInt_Int_Int) > (gacU_4_1_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t gacU_4_destruct_bufchan_d;
  logic gacU_4_destruct_bufchan_r;
  assign gacU_4_destruct_r = ((! gacU_4_destruct_bufchan_d[0]) || gacU_4_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) gacU_4_destruct_bufchan_d <= 1'd0;
    else
      if (gacU_4_destruct_r)
        gacU_4_destruct_bufchan_d <= gacU_4_destruct_d;
  MyDTInt_Int_Int_t gacU_4_destruct_bufchan_buf;
  assign gacU_4_destruct_bufchan_r = (! gacU_4_destruct_bufchan_buf[0]);
  assign gacU_4_1_argbuf_d = (gacU_4_destruct_bufchan_buf[0] ? gacU_4_destruct_bufchan_buf :
                              gacU_4_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) gacU_4_destruct_bufchan_buf <= 1'd0;
    else
      if ((gacU_4_1_argbuf_r && gacU_4_destruct_bufchan_buf[0]))
        gacU_4_destruct_bufchan_buf <= 1'd0;
      else if (((! gacU_4_1_argbuf_r) && (! gacU_4_destruct_bufchan_buf[0])))
        gacU_4_destruct_bufchan_buf <= gacU_4_destruct_bufchan_d;
  
  /* buf (Ty MyDTInt_Int_Int) : (gad3_2_2,MyDTInt_Int_Int) > (gad3_2_2_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t gad3_2_2_bufchan_d;
  logic gad3_2_2_bufchan_r;
  assign gad3_2_2_r = ((! gad3_2_2_bufchan_d[0]) || gad3_2_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) gad3_2_2_bufchan_d <= 1'd0;
    else if (gad3_2_2_r) gad3_2_2_bufchan_d <= gad3_2_2_d;
  MyDTInt_Int_Int_t gad3_2_2_bufchan_buf;
  assign gad3_2_2_bufchan_r = (! gad3_2_2_bufchan_buf[0]);
  assign gad3_2_2_argbuf_d = (gad3_2_2_bufchan_buf[0] ? gad3_2_2_bufchan_buf :
                              gad3_2_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) gad3_2_2_bufchan_buf <= 1'd0;
    else
      if ((gad3_2_2_argbuf_r && gad3_2_2_bufchan_buf[0]))
        gad3_2_2_bufchan_buf <= 1'd0;
      else if (((! gad3_2_2_argbuf_r) && (! gad3_2_2_bufchan_buf[0])))
        gad3_2_2_bufchan_buf <= gad3_2_2_bufchan_d;
  
  /* fork (Ty MyDTInt_Int_Int) : (gad3_2_destruct,MyDTInt_Int_Int) > [(gad3_2_1,MyDTInt_Int_Int),
                                                                 (gad3_2_2,MyDTInt_Int_Int)] */
  logic [1:0] gad3_2_destruct_emitted;
  logic [1:0] gad3_2_destruct_done;
  assign gad3_2_1_d = (gad3_2_destruct_d[0] && (! gad3_2_destruct_emitted[0]));
  assign gad3_2_2_d = (gad3_2_destruct_d[0] && (! gad3_2_destruct_emitted[1]));
  assign gad3_2_destruct_done = (gad3_2_destruct_emitted | ({gad3_2_2_d[0],
                                                             gad3_2_1_d[0]} & {gad3_2_2_r,
                                                                               gad3_2_1_r}));
  assign gad3_2_destruct_r = (& gad3_2_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) gad3_2_destruct_emitted <= 2'd0;
    else
      gad3_2_destruct_emitted <= (gad3_2_destruct_r ? 2'd0 :
                                  gad3_2_destruct_done);
  
  /* buf (Ty MyDTInt_Int_Int) : (gad3_3_2,MyDTInt_Int_Int) > (gad3_3_2_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t gad3_3_2_bufchan_d;
  logic gad3_3_2_bufchan_r;
  assign gad3_3_2_r = ((! gad3_3_2_bufchan_d[0]) || gad3_3_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) gad3_3_2_bufchan_d <= 1'd0;
    else if (gad3_3_2_r) gad3_3_2_bufchan_d <= gad3_3_2_d;
  MyDTInt_Int_Int_t gad3_3_2_bufchan_buf;
  assign gad3_3_2_bufchan_r = (! gad3_3_2_bufchan_buf[0]);
  assign gad3_3_2_argbuf_d = (gad3_3_2_bufchan_buf[0] ? gad3_3_2_bufchan_buf :
                              gad3_3_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) gad3_3_2_bufchan_buf <= 1'd0;
    else
      if ((gad3_3_2_argbuf_r && gad3_3_2_bufchan_buf[0]))
        gad3_3_2_bufchan_buf <= 1'd0;
      else if (((! gad3_3_2_argbuf_r) && (! gad3_3_2_bufchan_buf[0])))
        gad3_3_2_bufchan_buf <= gad3_3_2_bufchan_d;
  
  /* fork (Ty MyDTInt_Int_Int) : (gad3_3_destruct,MyDTInt_Int_Int) > [(gad3_3_1,MyDTInt_Int_Int),
                                                                 (gad3_3_2,MyDTInt_Int_Int)] */
  logic [1:0] gad3_3_destruct_emitted;
  logic [1:0] gad3_3_destruct_done;
  assign gad3_3_1_d = (gad3_3_destruct_d[0] && (! gad3_3_destruct_emitted[0]));
  assign gad3_3_2_d = (gad3_3_destruct_d[0] && (! gad3_3_destruct_emitted[1]));
  assign gad3_3_destruct_done = (gad3_3_destruct_emitted | ({gad3_3_2_d[0],
                                                             gad3_3_1_d[0]} & {gad3_3_2_r,
                                                                               gad3_3_1_r}));
  assign gad3_3_destruct_r = (& gad3_3_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) gad3_3_destruct_emitted <= 2'd0;
    else
      gad3_3_destruct_emitted <= (gad3_3_destruct_r ? 2'd0 :
                                  gad3_3_destruct_done);
  
  /* buf (Ty MyDTInt_Int_Int) : (gad3_4_destruct,MyDTInt_Int_Int) > (gad3_4_1_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t gad3_4_destruct_bufchan_d;
  logic gad3_4_destruct_bufchan_r;
  assign gad3_4_destruct_r = ((! gad3_4_destruct_bufchan_d[0]) || gad3_4_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) gad3_4_destruct_bufchan_d <= 1'd0;
    else
      if (gad3_4_destruct_r)
        gad3_4_destruct_bufchan_d <= gad3_4_destruct_d;
  MyDTInt_Int_Int_t gad3_4_destruct_bufchan_buf;
  assign gad3_4_destruct_bufchan_r = (! gad3_4_destruct_bufchan_buf[0]);
  assign gad3_4_1_argbuf_d = (gad3_4_destruct_bufchan_buf[0] ? gad3_4_destruct_bufchan_buf :
                              gad3_4_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) gad3_4_destruct_bufchan_buf <= 1'd0;
    else
      if ((gad3_4_1_argbuf_r && gad3_4_destruct_bufchan_buf[0]))
        gad3_4_destruct_bufchan_buf <= 1'd0;
      else if (((! gad3_4_1_argbuf_r) && (! gad3_4_destruct_bufchan_buf[0])))
        gad3_4_destruct_bufchan_buf <= gad3_4_destruct_bufchan_d;
  
  /* fork (Ty C5) : (go_11_goMux_choice,C5) > [(go_11_goMux_choice_1,C5),
                                          (go_11_goMux_choice_2,C5)] */
  logic [1:0] go_11_goMux_choice_emitted;
  logic [1:0] go_11_goMux_choice_done;
  assign go_11_goMux_choice_1_d = {go_11_goMux_choice_d[3:1],
                                   (go_11_goMux_choice_d[0] && (! go_11_goMux_choice_emitted[0]))};
  assign go_11_goMux_choice_2_d = {go_11_goMux_choice_d[3:1],
                                   (go_11_goMux_choice_d[0] && (! go_11_goMux_choice_emitted[1]))};
  assign go_11_goMux_choice_done = (go_11_goMux_choice_emitted | ({go_11_goMux_choice_2_d[0],
                                                                   go_11_goMux_choice_1_d[0]} & {go_11_goMux_choice_2_r,
                                                                                                 go_11_goMux_choice_1_r}));
  assign go_11_goMux_choice_r = (& go_11_goMux_choice_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_11_goMux_choice_emitted <= 2'd0;
    else
      go_11_goMux_choice_emitted <= (go_11_goMux_choice_r ? 2'd0 :
                                     go_11_goMux_choice_done);
  
  /* mux (Ty C5,
     Ty Pointer_QTree_Int) : (go_11_goMux_choice_1,C5) [(call_$wnnz_Int_goMux2,Pointer_QTree_Int),
                                                        (q2ac1_1_1_argbuf,Pointer_QTree_Int),
                                                        (q3ac2_2_1_argbuf,Pointer_QTree_Int),
                                                        (q4ac3_3_1_argbuf,Pointer_QTree_Int),
                                                        (q1ac0_1_argbuf,Pointer_QTree_Int)] > (wsvt_1_goMux_mux,Pointer_QTree_Int) */
  logic [16:0] wsvt_1_goMux_mux_mux;
  logic [4:0] wsvt_1_goMux_mux_onehot;
  always_comb
    unique case (go_11_goMux_choice_1_d[3:1])
      3'd0:
        {wsvt_1_goMux_mux_onehot, wsvt_1_goMux_mux_mux} = {5'd1,
                                                           call_$wnnz_Int_goMux2_d};
      3'd1:
        {wsvt_1_goMux_mux_onehot, wsvt_1_goMux_mux_mux} = {5'd2,
                                                           q2ac1_1_1_argbuf_d};
      3'd2:
        {wsvt_1_goMux_mux_onehot, wsvt_1_goMux_mux_mux} = {5'd4,
                                                           q3ac2_2_1_argbuf_d};
      3'd3:
        {wsvt_1_goMux_mux_onehot, wsvt_1_goMux_mux_mux} = {5'd8,
                                                           q4ac3_3_1_argbuf_d};
      3'd4:
        {wsvt_1_goMux_mux_onehot, wsvt_1_goMux_mux_mux} = {5'd16,
                                                           q1ac0_1_argbuf_d};
      default:
        {wsvt_1_goMux_mux_onehot, wsvt_1_goMux_mux_mux} = {5'd0,
                                                           {16'd0, 1'd0}};
    endcase
  assign wsvt_1_goMux_mux_d = {wsvt_1_goMux_mux_mux[16:1],
                               (wsvt_1_goMux_mux_mux[0] && go_11_goMux_choice_1_d[0])};
  assign go_11_goMux_choice_1_r = (wsvt_1_goMux_mux_d[0] && wsvt_1_goMux_mux_r);
  assign {q1ac0_1_argbuf_r,
          q4ac3_3_1_argbuf_r,
          q3ac2_2_1_argbuf_r,
          q2ac1_1_1_argbuf_r,
          call_$wnnz_Int_goMux2_r} = (go_11_goMux_choice_1_r ? wsvt_1_goMux_mux_onehot :
                                      5'd0);
  
  /* mux (Ty C5,
     Ty Pointer_CT$wnnz_Int) : (go_11_goMux_choice_2,C5) [(call_$wnnz_Int_goMux3,Pointer_CT$wnnz_Int),
                                                          (sca2_1_argbuf,Pointer_CT$wnnz_Int),
                                                          (sca1_1_argbuf,Pointer_CT$wnnz_Int),
                                                          (sca0_1_argbuf,Pointer_CT$wnnz_Int),
                                                          (sca3_1_argbuf,Pointer_CT$wnnz_Int)] > (sc_0_goMux_mux,Pointer_CT$wnnz_Int) */
  logic [16:0] sc_0_goMux_mux_mux;
  logic [4:0] sc_0_goMux_mux_onehot;
  always_comb
    unique case (go_11_goMux_choice_2_d[3:1])
      3'd0:
        {sc_0_goMux_mux_onehot, sc_0_goMux_mux_mux} = {5'd1,
                                                       call_$wnnz_Int_goMux3_d};
      3'd1:
        {sc_0_goMux_mux_onehot, sc_0_goMux_mux_mux} = {5'd2,
                                                       sca2_1_argbuf_d};
      3'd2:
        {sc_0_goMux_mux_onehot, sc_0_goMux_mux_mux} = {5'd4,
                                                       sca1_1_argbuf_d};
      3'd3:
        {sc_0_goMux_mux_onehot, sc_0_goMux_mux_mux} = {5'd8,
                                                       sca0_1_argbuf_d};
      3'd4:
        {sc_0_goMux_mux_onehot, sc_0_goMux_mux_mux} = {5'd16,
                                                       sca3_1_argbuf_d};
      default:
        {sc_0_goMux_mux_onehot, sc_0_goMux_mux_mux} = {5'd0,
                                                       {16'd0, 1'd0}};
    endcase
  assign sc_0_goMux_mux_d = {sc_0_goMux_mux_mux[16:1],
                             (sc_0_goMux_mux_mux[0] && go_11_goMux_choice_2_d[0])};
  assign go_11_goMux_choice_2_r = (sc_0_goMux_mux_d[0] && sc_0_goMux_mux_r);
  assign {sca3_1_argbuf_r,
          sca0_1_argbuf_r,
          sca1_1_argbuf_r,
          sca2_1_argbuf_r,
          call_$wnnz_Int_goMux3_r} = (go_11_goMux_choice_2_r ? sc_0_goMux_mux_onehot :
                                      5'd0);
  
  /* fork (Ty C5) : (go_12_goMux_choice,C5) > [(go_12_goMux_choice_1,C5),
                                          (go_12_goMux_choice_2,C5),
                                          (go_12_goMux_choice_3,C5),
                                          (go_12_goMux_choice_4,C5),
                                          (go_12_goMux_choice_5,C5)] */
  logic [4:0] go_12_goMux_choice_emitted;
  logic [4:0] go_12_goMux_choice_done;
  assign go_12_goMux_choice_1_d = {go_12_goMux_choice_d[3:1],
                                   (go_12_goMux_choice_d[0] && (! go_12_goMux_choice_emitted[0]))};
  assign go_12_goMux_choice_2_d = {go_12_goMux_choice_d[3:1],
                                   (go_12_goMux_choice_d[0] && (! go_12_goMux_choice_emitted[1]))};
  assign go_12_goMux_choice_3_d = {go_12_goMux_choice_d[3:1],
                                   (go_12_goMux_choice_d[0] && (! go_12_goMux_choice_emitted[2]))};
  assign go_12_goMux_choice_4_d = {go_12_goMux_choice_d[3:1],
                                   (go_12_goMux_choice_d[0] && (! go_12_goMux_choice_emitted[3]))};
  assign go_12_goMux_choice_5_d = {go_12_goMux_choice_d[3:1],
                                   (go_12_goMux_choice_d[0] && (! go_12_goMux_choice_emitted[4]))};
  assign go_12_goMux_choice_done = (go_12_goMux_choice_emitted | ({go_12_goMux_choice_5_d[0],
                                                                   go_12_goMux_choice_4_d[0],
                                                                   go_12_goMux_choice_3_d[0],
                                                                   go_12_goMux_choice_2_d[0],
                                                                   go_12_goMux_choice_1_d[0]} & {go_12_goMux_choice_5_r,
                                                                                                 go_12_goMux_choice_4_r,
                                                                                                 go_12_goMux_choice_3_r,
                                                                                                 go_12_goMux_choice_2_r,
                                                                                                 go_12_goMux_choice_1_r}));
  assign go_12_goMux_choice_r = (& go_12_goMux_choice_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_12_goMux_choice_emitted <= 5'd0;
    else
      go_12_goMux_choice_emitted <= (go_12_goMux_choice_r ? 5'd0 :
                                     go_12_goMux_choice_done);
  
  /* mux (Ty C5,
     Ty MyDTInt_Bool) : (go_12_goMux_choice_1,C5) [(call_kron_kron_Int_Int_Int_goMux2,MyDTInt_Bool),
                                                   (isZad2_2_2_argbuf,MyDTInt_Bool),
                                                   (isZad2_3_2_argbuf,MyDTInt_Bool),
                                                   (isZad2_4_1_argbuf,MyDTInt_Bool),
                                                   (lizzieLet6_5QNode_Int_2_argbuf,MyDTInt_Bool)] > (isZad2_goMux_mux,MyDTInt_Bool) */
  logic [0:0] isZad2_goMux_mux_mux;
  logic [4:0] isZad2_goMux_mux_onehot;
  always_comb
    unique case (go_12_goMux_choice_1_d[3:1])
      3'd0:
        {isZad2_goMux_mux_onehot, isZad2_goMux_mux_mux} = {5'd1,
                                                           call_kron_kron_Int_Int_Int_goMux2_d};
      3'd1:
        {isZad2_goMux_mux_onehot, isZad2_goMux_mux_mux} = {5'd2,
                                                           isZad2_2_2_argbuf_d};
      3'd2:
        {isZad2_goMux_mux_onehot, isZad2_goMux_mux_mux} = {5'd4,
                                                           isZad2_3_2_argbuf_d};
      3'd3:
        {isZad2_goMux_mux_onehot, isZad2_goMux_mux_mux} = {5'd8,
                                                           isZad2_4_1_argbuf_d};
      3'd4:
        {isZad2_goMux_mux_onehot, isZad2_goMux_mux_mux} = {5'd16,
                                                           lizzieLet6_5QNode_Int_2_argbuf_d};
      default:
        {isZad2_goMux_mux_onehot, isZad2_goMux_mux_mux} = {5'd0, 1'd0};
    endcase
  assign isZad2_goMux_mux_d = (isZad2_goMux_mux_mux[0] && go_12_goMux_choice_1_d[0]);
  assign go_12_goMux_choice_1_r = (isZad2_goMux_mux_d[0] && isZad2_goMux_mux_r);
  assign {lizzieLet6_5QNode_Int_2_argbuf_r,
          isZad2_4_1_argbuf_r,
          isZad2_3_2_argbuf_r,
          isZad2_2_2_argbuf_r,
          call_kron_kron_Int_Int_Int_goMux2_r} = (go_12_goMux_choice_1_r ? isZad2_goMux_mux_onehot :
                                                  5'd0);
  
  /* mux (Ty C5,
     Ty MyDTInt_Int_Int) : (go_12_goMux_choice_2,C5) [(call_kron_kron_Int_Int_Int_goMux3,MyDTInt_Int_Int),
                                                      (gad3_2_2_argbuf,MyDTInt_Int_Int),
                                                      (gad3_3_2_argbuf,MyDTInt_Int_Int),
                                                      (gad3_4_1_argbuf,MyDTInt_Int_Int),
                                                      (lizzieLet6_3QNode_Int_2_argbuf,MyDTInt_Int_Int)] > (gad3_goMux_mux,MyDTInt_Int_Int) */
  logic [0:0] gad3_goMux_mux_mux;
  logic [4:0] gad3_goMux_mux_onehot;
  always_comb
    unique case (go_12_goMux_choice_2_d[3:1])
      3'd0:
        {gad3_goMux_mux_onehot, gad3_goMux_mux_mux} = {5'd1,
                                                       call_kron_kron_Int_Int_Int_goMux3_d};
      3'd1:
        {gad3_goMux_mux_onehot, gad3_goMux_mux_mux} = {5'd2,
                                                       gad3_2_2_argbuf_d};
      3'd2:
        {gad3_goMux_mux_onehot, gad3_goMux_mux_mux} = {5'd4,
                                                       gad3_3_2_argbuf_d};
      3'd3:
        {gad3_goMux_mux_onehot, gad3_goMux_mux_mux} = {5'd8,
                                                       gad3_4_1_argbuf_d};
      3'd4:
        {gad3_goMux_mux_onehot, gad3_goMux_mux_mux} = {5'd16,
                                                       lizzieLet6_3QNode_Int_2_argbuf_d};
      default:
        {gad3_goMux_mux_onehot, gad3_goMux_mux_mux} = {5'd0, 1'd0};
    endcase
  assign gad3_goMux_mux_d = (gad3_goMux_mux_mux[0] && go_12_goMux_choice_2_d[0]);
  assign go_12_goMux_choice_2_r = (gad3_goMux_mux_d[0] && gad3_goMux_mux_r);
  assign {lizzieLet6_3QNode_Int_2_argbuf_r,
          gad3_4_1_argbuf_r,
          gad3_3_2_argbuf_r,
          gad3_2_2_argbuf_r,
          call_kron_kron_Int_Int_Int_goMux3_r} = (go_12_goMux_choice_2_r ? gad3_goMux_mux_onehot :
                                                  5'd0);
  
  /* mux (Ty C5,
     Ty Pointer_QTree_Int) : (go_12_goMux_choice_3,C5) [(call_kron_kron_Int_Int_Int_goMux4,Pointer_QTree_Int),
                                                        (q3ad9_1_1_argbuf,Pointer_QTree_Int),
                                                        (q2ad8_2_1_argbuf,Pointer_QTree_Int),
                                                        (q1ad7_3_1_argbuf,Pointer_QTree_Int),
                                                        (q4ada_1_argbuf,Pointer_QTree_Int)] > (m1ad4_goMux_mux,Pointer_QTree_Int) */
  logic [16:0] m1ad4_goMux_mux_mux;
  logic [4:0] m1ad4_goMux_mux_onehot;
  always_comb
    unique case (go_12_goMux_choice_3_d[3:1])
      3'd0:
        {m1ad4_goMux_mux_onehot, m1ad4_goMux_mux_mux} = {5'd1,
                                                         call_kron_kron_Int_Int_Int_goMux4_d};
      3'd1:
        {m1ad4_goMux_mux_onehot, m1ad4_goMux_mux_mux} = {5'd2,
                                                         q3ad9_1_1_argbuf_d};
      3'd2:
        {m1ad4_goMux_mux_onehot, m1ad4_goMux_mux_mux} = {5'd4,
                                                         q2ad8_2_1_argbuf_d};
      3'd3:
        {m1ad4_goMux_mux_onehot, m1ad4_goMux_mux_mux} = {5'd8,
                                                         q1ad7_3_1_argbuf_d};
      3'd4:
        {m1ad4_goMux_mux_onehot, m1ad4_goMux_mux_mux} = {5'd16,
                                                         q4ada_1_argbuf_d};
      default:
        {m1ad4_goMux_mux_onehot, m1ad4_goMux_mux_mux} = {5'd0,
                                                         {16'd0, 1'd0}};
    endcase
  assign m1ad4_goMux_mux_d = {m1ad4_goMux_mux_mux[16:1],
                              (m1ad4_goMux_mux_mux[0] && go_12_goMux_choice_3_d[0])};
  assign go_12_goMux_choice_3_r = (m1ad4_goMux_mux_d[0] && m1ad4_goMux_mux_r);
  assign {q4ada_1_argbuf_r,
          q1ad7_3_1_argbuf_r,
          q2ad8_2_1_argbuf_r,
          q3ad9_1_1_argbuf_r,
          call_kron_kron_Int_Int_Int_goMux4_r} = (go_12_goMux_choice_3_r ? m1ad4_goMux_mux_onehot :
                                                  5'd0);
  
  /* mux (Ty C5,
     Ty Pointer_QTree_Int) : (go_12_goMux_choice_4,C5) [(call_kron_kron_Int_Int_Int_goMux5,Pointer_QTree_Int),
                                                        (m2ad5_2_2_argbuf,Pointer_QTree_Int),
                                                        (m2ad5_3_2_argbuf,Pointer_QTree_Int),
                                                        (m2ad5_4_1_argbuf,Pointer_QTree_Int),
                                                        (lizzieLet6_6QNode_Int_2_argbuf,Pointer_QTree_Int)] > (m2ad5_goMux_mux,Pointer_QTree_Int) */
  logic [16:0] m2ad5_goMux_mux_mux;
  logic [4:0] m2ad5_goMux_mux_onehot;
  always_comb
    unique case (go_12_goMux_choice_4_d[3:1])
      3'd0:
        {m2ad5_goMux_mux_onehot, m2ad5_goMux_mux_mux} = {5'd1,
                                                         call_kron_kron_Int_Int_Int_goMux5_d};
      3'd1:
        {m2ad5_goMux_mux_onehot, m2ad5_goMux_mux_mux} = {5'd2,
                                                         m2ad5_2_2_argbuf_d};
      3'd2:
        {m2ad5_goMux_mux_onehot, m2ad5_goMux_mux_mux} = {5'd4,
                                                         m2ad5_3_2_argbuf_d};
      3'd3:
        {m2ad5_goMux_mux_onehot, m2ad5_goMux_mux_mux} = {5'd8,
                                                         m2ad5_4_1_argbuf_d};
      3'd4:
        {m2ad5_goMux_mux_onehot, m2ad5_goMux_mux_mux} = {5'd16,
                                                         lizzieLet6_6QNode_Int_2_argbuf_d};
      default:
        {m2ad5_goMux_mux_onehot, m2ad5_goMux_mux_mux} = {5'd0,
                                                         {16'd0, 1'd0}};
    endcase
  assign m2ad5_goMux_mux_d = {m2ad5_goMux_mux_mux[16:1],
                              (m2ad5_goMux_mux_mux[0] && go_12_goMux_choice_4_d[0])};
  assign go_12_goMux_choice_4_r = (m2ad5_goMux_mux_d[0] && m2ad5_goMux_mux_r);
  assign {lizzieLet6_6QNode_Int_2_argbuf_r,
          m2ad5_4_1_argbuf_r,
          m2ad5_3_2_argbuf_r,
          m2ad5_2_2_argbuf_r,
          call_kron_kron_Int_Int_Int_goMux5_r} = (go_12_goMux_choice_4_r ? m2ad5_goMux_mux_onehot :
                                                  5'd0);
  
  /* mux (Ty C5,
     Ty Pointer_CTkron_kron_Int_Int_Int) : (go_12_goMux_choice_5,C5) [(call_kron_kron_Int_Int_Int_goMux6,Pointer_CTkron_kron_Int_Int_Int),
                                                                      (sca2_1_1_argbuf,Pointer_CTkron_kron_Int_Int_Int),
                                                                      (sca1_1_1_argbuf,Pointer_CTkron_kron_Int_Int_Int),
                                                                      (sca0_1_1_argbuf,Pointer_CTkron_kron_Int_Int_Int),
                                                                      (sca3_1_1_argbuf,Pointer_CTkron_kron_Int_Int_Int)] > (sc_0_1_goMux_mux,Pointer_CTkron_kron_Int_Int_Int) */
  logic [16:0] sc_0_1_goMux_mux_mux;
  logic [4:0] sc_0_1_goMux_mux_onehot;
  always_comb
    unique case (go_12_goMux_choice_5_d[3:1])
      3'd0:
        {sc_0_1_goMux_mux_onehot, sc_0_1_goMux_mux_mux} = {5'd1,
                                                           call_kron_kron_Int_Int_Int_goMux6_d};
      3'd1:
        {sc_0_1_goMux_mux_onehot, sc_0_1_goMux_mux_mux} = {5'd2,
                                                           sca2_1_1_argbuf_d};
      3'd2:
        {sc_0_1_goMux_mux_onehot, sc_0_1_goMux_mux_mux} = {5'd4,
                                                           sca1_1_1_argbuf_d};
      3'd3:
        {sc_0_1_goMux_mux_onehot, sc_0_1_goMux_mux_mux} = {5'd8,
                                                           sca0_1_1_argbuf_d};
      3'd4:
        {sc_0_1_goMux_mux_onehot, sc_0_1_goMux_mux_mux} = {5'd16,
                                                           sca3_1_1_argbuf_d};
      default:
        {sc_0_1_goMux_mux_onehot, sc_0_1_goMux_mux_mux} = {5'd0,
                                                           {16'd0, 1'd0}};
    endcase
  assign sc_0_1_goMux_mux_d = {sc_0_1_goMux_mux_mux[16:1],
                               (sc_0_1_goMux_mux_mux[0] && go_12_goMux_choice_5_d[0])};
  assign go_12_goMux_choice_5_r = (sc_0_1_goMux_mux_d[0] && sc_0_1_goMux_mux_r);
  assign {sca3_1_1_argbuf_r,
          sca0_1_1_argbuf_r,
          sca1_1_1_argbuf_r,
          sca2_1_1_argbuf_r,
          call_kron_kron_Int_Int_Int_goMux6_r} = (go_12_goMux_choice_5_r ? sc_0_1_goMux_mux_onehot :
                                                  5'd0);
  
  /* fork (Ty C5) : (go_13_goMux_choice,C5) > [(go_13_goMux_choice_1,C5),
                                          (go_13_goMux_choice_2,C5),
                                          (go_13_goMux_choice_3,C5),
                                          (go_13_goMux_choice_4,C5)] */
  logic [3:0] go_13_goMux_choice_emitted;
  logic [3:0] go_13_goMux_choice_done;
  assign go_13_goMux_choice_1_d = {go_13_goMux_choice_d[3:1],
                                   (go_13_goMux_choice_d[0] && (! go_13_goMux_choice_emitted[0]))};
  assign go_13_goMux_choice_2_d = {go_13_goMux_choice_d[3:1],
                                   (go_13_goMux_choice_d[0] && (! go_13_goMux_choice_emitted[1]))};
  assign go_13_goMux_choice_3_d = {go_13_goMux_choice_d[3:1],
                                   (go_13_goMux_choice_d[0] && (! go_13_goMux_choice_emitted[2]))};
  assign go_13_goMux_choice_4_d = {go_13_goMux_choice_d[3:1],
                                   (go_13_goMux_choice_d[0] && (! go_13_goMux_choice_emitted[3]))};
  assign go_13_goMux_choice_done = (go_13_goMux_choice_emitted | ({go_13_goMux_choice_4_d[0],
                                                                   go_13_goMux_choice_3_d[0],
                                                                   go_13_goMux_choice_2_d[0],
                                                                   go_13_goMux_choice_1_d[0]} & {go_13_goMux_choice_4_r,
                                                                                                 go_13_goMux_choice_3_r,
                                                                                                 go_13_goMux_choice_2_r,
                                                                                                 go_13_goMux_choice_1_r}));
  assign go_13_goMux_choice_r = (& go_13_goMux_choice_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_13_goMux_choice_emitted <= 4'd0;
    else
      go_13_goMux_choice_emitted <= (go_13_goMux_choice_r ? 4'd0 :
                                     go_13_goMux_choice_done);
  
  /* mux (Ty C5,
     Ty MyDTInt_Bool) : (go_13_goMux_choice_1,C5) [(call_main_map'_Int_Int_goMux2,MyDTInt_Bool),
                                                   (isZacL_2_2_argbuf,MyDTInt_Bool),
                                                   (isZacL_3_2_argbuf,MyDTInt_Bool),
                                                   (isZacL_4_1_argbuf,MyDTInt_Bool),
                                                   (lizzieLet10_5QNode_Int_2_argbuf,MyDTInt_Bool)] > (isZacL_goMux_mux,MyDTInt_Bool) */
  logic [0:0] isZacL_goMux_mux_mux;
  logic [4:0] isZacL_goMux_mux_onehot;
  always_comb
    unique case (go_13_goMux_choice_1_d[3:1])
      3'd0:
        {isZacL_goMux_mux_onehot, isZacL_goMux_mux_mux} = {5'd1,
                                                           \call_main_map'_Int_Int_goMux2_d };
      3'd1:
        {isZacL_goMux_mux_onehot, isZacL_goMux_mux_mux} = {5'd2,
                                                           isZacL_2_2_argbuf_d};
      3'd2:
        {isZacL_goMux_mux_onehot, isZacL_goMux_mux_mux} = {5'd4,
                                                           isZacL_3_2_argbuf_d};
      3'd3:
        {isZacL_goMux_mux_onehot, isZacL_goMux_mux_mux} = {5'd8,
                                                           isZacL_4_1_argbuf_d};
      3'd4:
        {isZacL_goMux_mux_onehot, isZacL_goMux_mux_mux} = {5'd16,
                                                           lizzieLet10_5QNode_Int_2_argbuf_d};
      default:
        {isZacL_goMux_mux_onehot, isZacL_goMux_mux_mux} = {5'd0, 1'd0};
    endcase
  assign isZacL_goMux_mux_d = (isZacL_goMux_mux_mux[0] && go_13_goMux_choice_1_d[0]);
  assign go_13_goMux_choice_1_r = (isZacL_goMux_mux_d[0] && isZacL_goMux_mux_r);
  assign {lizzieLet10_5QNode_Int_2_argbuf_r,
          isZacL_4_1_argbuf_r,
          isZacL_3_2_argbuf_r,
          isZacL_2_2_argbuf_r,
          \call_main_map'_Int_Int_goMux2_r } = (go_13_goMux_choice_1_r ? isZacL_goMux_mux_onehot :
                                                5'd0);
  
  /* mux (Ty C5,
     Ty MyDTInt_Int) : (go_13_goMux_choice_2,C5) [(call_main_map'_Int_Int_goMux3,MyDTInt_Int),
                                                  (gacM_2_2_argbuf,MyDTInt_Int),
                                                  (gacM_3_2_argbuf,MyDTInt_Int),
                                                  (gacM_4_1_argbuf,MyDTInt_Int),
                                                  (lizzieLet10_3QNode_Int_2_argbuf,MyDTInt_Int)] > (gacM_goMux_mux,MyDTInt_Int) */
  logic [0:0] gacM_goMux_mux_mux;
  logic [4:0] gacM_goMux_mux_onehot;
  always_comb
    unique case (go_13_goMux_choice_2_d[3:1])
      3'd0:
        {gacM_goMux_mux_onehot, gacM_goMux_mux_mux} = {5'd1,
                                                       \call_main_map'_Int_Int_goMux3_d };
      3'd1:
        {gacM_goMux_mux_onehot, gacM_goMux_mux_mux} = {5'd2,
                                                       gacM_2_2_argbuf_d};
      3'd2:
        {gacM_goMux_mux_onehot, gacM_goMux_mux_mux} = {5'd4,
                                                       gacM_3_2_argbuf_d};
      3'd3:
        {gacM_goMux_mux_onehot, gacM_goMux_mux_mux} = {5'd8,
                                                       gacM_4_1_argbuf_d};
      3'd4:
        {gacM_goMux_mux_onehot, gacM_goMux_mux_mux} = {5'd16,
                                                       lizzieLet10_3QNode_Int_2_argbuf_d};
      default:
        {gacM_goMux_mux_onehot, gacM_goMux_mux_mux} = {5'd0, 1'd0};
    endcase
  assign gacM_goMux_mux_d = (gacM_goMux_mux_mux[0] && go_13_goMux_choice_2_d[0]);
  assign go_13_goMux_choice_2_r = (gacM_goMux_mux_d[0] && gacM_goMux_mux_r);
  assign {lizzieLet10_3QNode_Int_2_argbuf_r,
          gacM_4_1_argbuf_r,
          gacM_3_2_argbuf_r,
          gacM_2_2_argbuf_r,
          \call_main_map'_Int_Int_goMux3_r } = (go_13_goMux_choice_2_r ? gacM_goMux_mux_onehot :
                                                5'd0);
  
  /* mux (Ty C5,
     Ty Pointer_QTree_Int) : (go_13_goMux_choice_3,C5) [(call_main_map'_Int_Int_goMux4,Pointer_QTree_Int),
                                                        (q3acR_1_1_argbuf,Pointer_QTree_Int),
                                                        (q2acQ_2_1_argbuf,Pointer_QTree_Int),
                                                        (q1acP_3_1_argbuf,Pointer_QTree_Int),
                                                        (q4acS_1_argbuf,Pointer_QTree_Int)] > (macN_goMux_mux,Pointer_QTree_Int) */
  logic [16:0] macN_goMux_mux_mux;
  logic [4:0] macN_goMux_mux_onehot;
  always_comb
    unique case (go_13_goMux_choice_3_d[3:1])
      3'd0:
        {macN_goMux_mux_onehot, macN_goMux_mux_mux} = {5'd1,
                                                       \call_main_map'_Int_Int_goMux4_d };
      3'd1:
        {macN_goMux_mux_onehot, macN_goMux_mux_mux} = {5'd2,
                                                       q3acR_1_1_argbuf_d};
      3'd2:
        {macN_goMux_mux_onehot, macN_goMux_mux_mux} = {5'd4,
                                                       q2acQ_2_1_argbuf_d};
      3'd3:
        {macN_goMux_mux_onehot, macN_goMux_mux_mux} = {5'd8,
                                                       q1acP_3_1_argbuf_d};
      3'd4:
        {macN_goMux_mux_onehot, macN_goMux_mux_mux} = {5'd16,
                                                       q4acS_1_argbuf_d};
      default:
        {macN_goMux_mux_onehot, macN_goMux_mux_mux} = {5'd0,
                                                       {16'd0, 1'd0}};
    endcase
  assign macN_goMux_mux_d = {macN_goMux_mux_mux[16:1],
                             (macN_goMux_mux_mux[0] && go_13_goMux_choice_3_d[0])};
  assign go_13_goMux_choice_3_r = (macN_goMux_mux_d[0] && macN_goMux_mux_r);
  assign {q4acS_1_argbuf_r,
          q1acP_3_1_argbuf_r,
          q2acQ_2_1_argbuf_r,
          q3acR_1_1_argbuf_r,
          \call_main_map'_Int_Int_goMux4_r } = (go_13_goMux_choice_3_r ? macN_goMux_mux_onehot :
                                                5'd0);
  
  /* mux (Ty C5,
     Ty Pointer_CTmain_map'_Int_Int) : (go_13_goMux_choice_4,C5) [(call_main_map'_Int_Int_goMux5,Pointer_CTmain_map'_Int_Int),
                                                                  (sca2_2_1_argbuf,Pointer_CTmain_map'_Int_Int),
                                                                  (sca1_2_1_argbuf,Pointer_CTmain_map'_Int_Int),
                                                                  (sca0_2_1_argbuf,Pointer_CTmain_map'_Int_Int),
                                                                  (sca3_2_1_argbuf,Pointer_CTmain_map'_Int_Int)] > (sc_0_2_goMux_mux,Pointer_CTmain_map'_Int_Int) */
  logic [16:0] sc_0_2_goMux_mux_mux;
  logic [4:0] sc_0_2_goMux_mux_onehot;
  always_comb
    unique case (go_13_goMux_choice_4_d[3:1])
      3'd0:
        {sc_0_2_goMux_mux_onehot, sc_0_2_goMux_mux_mux} = {5'd1,
                                                           \call_main_map'_Int_Int_goMux5_d };
      3'd1:
        {sc_0_2_goMux_mux_onehot, sc_0_2_goMux_mux_mux} = {5'd2,
                                                           sca2_2_1_argbuf_d};
      3'd2:
        {sc_0_2_goMux_mux_onehot, sc_0_2_goMux_mux_mux} = {5'd4,
                                                           sca1_2_1_argbuf_d};
      3'd3:
        {sc_0_2_goMux_mux_onehot, sc_0_2_goMux_mux_mux} = {5'd8,
                                                           sca0_2_1_argbuf_d};
      3'd4:
        {sc_0_2_goMux_mux_onehot, sc_0_2_goMux_mux_mux} = {5'd16,
                                                           sca3_2_1_argbuf_d};
      default:
        {sc_0_2_goMux_mux_onehot, sc_0_2_goMux_mux_mux} = {5'd0,
                                                           {16'd0, 1'd0}};
    endcase
  assign sc_0_2_goMux_mux_d = {sc_0_2_goMux_mux_mux[16:1],
                               (sc_0_2_goMux_mux_mux[0] && go_13_goMux_choice_4_d[0])};
  assign go_13_goMux_choice_4_r = (sc_0_2_goMux_mux_d[0] && sc_0_2_goMux_mux_r);
  assign {sca3_2_1_argbuf_r,
          sca0_2_1_argbuf_r,
          sca1_2_1_argbuf_r,
          sca2_2_1_argbuf_r,
          \call_main_map'_Int_Int_goMux5_r } = (go_13_goMux_choice_4_r ? sc_0_2_goMux_mux_onehot :
                                                5'd0);
  
  /* fork (Ty C5) : (go_14_goMux_choice,C5) > [(go_14_goMux_choice_1,C5),
                                          (go_14_goMux_choice_2,C5),
                                          (go_14_goMux_choice_3,C5),
                                          (go_14_goMux_choice_4,C5),
                                          (go_14_goMux_choice_5,C5)] */
  logic [4:0] go_14_goMux_choice_emitted;
  logic [4:0] go_14_goMux_choice_done;
  assign go_14_goMux_choice_1_d = {go_14_goMux_choice_d[3:1],
                                   (go_14_goMux_choice_d[0] && (! go_14_goMux_choice_emitted[0]))};
  assign go_14_goMux_choice_2_d = {go_14_goMux_choice_d[3:1],
                                   (go_14_goMux_choice_d[0] && (! go_14_goMux_choice_emitted[1]))};
  assign go_14_goMux_choice_3_d = {go_14_goMux_choice_d[3:1],
                                   (go_14_goMux_choice_d[0] && (! go_14_goMux_choice_emitted[2]))};
  assign go_14_goMux_choice_4_d = {go_14_goMux_choice_d[3:1],
                                   (go_14_goMux_choice_d[0] && (! go_14_goMux_choice_emitted[3]))};
  assign go_14_goMux_choice_5_d = {go_14_goMux_choice_d[3:1],
                                   (go_14_goMux_choice_d[0] && (! go_14_goMux_choice_emitted[4]))};
  assign go_14_goMux_choice_done = (go_14_goMux_choice_emitted | ({go_14_goMux_choice_5_d[0],
                                                                   go_14_goMux_choice_4_d[0],
                                                                   go_14_goMux_choice_3_d[0],
                                                                   go_14_goMux_choice_2_d[0],
                                                                   go_14_goMux_choice_1_d[0]} & {go_14_goMux_choice_5_r,
                                                                                                 go_14_goMux_choice_4_r,
                                                                                                 go_14_goMux_choice_3_r,
                                                                                                 go_14_goMux_choice_2_r,
                                                                                                 go_14_goMux_choice_1_r}));
  assign go_14_goMux_choice_r = (& go_14_goMux_choice_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_14_goMux_choice_emitted <= 5'd0;
    else
      go_14_goMux_choice_emitted <= (go_14_goMux_choice_r ? 5'd0 :
                                     go_14_goMux_choice_done);
  
  /* mux (Ty C5,
     Ty MyDTInt_Bool) : (go_14_goMux_choice_1,C5) [(call_map''_map''_Int_Int_Int_goMux2,MyDTInt_Bool),
                                                   (isZacT_2_2_argbuf,MyDTInt_Bool),
                                                   (isZacT_3_2_argbuf,MyDTInt_Bool),
                                                   (isZacT_4_1_argbuf,MyDTInt_Bool),
                                                   (lizzieLet16_1_5QNode_Int_2_argbuf,MyDTInt_Bool)] > (isZacT_goMux_mux,MyDTInt_Bool) */
  logic [0:0] isZacT_goMux_mux_mux;
  logic [4:0] isZacT_goMux_mux_onehot;
  always_comb
    unique case (go_14_goMux_choice_1_d[3:1])
      3'd0:
        {isZacT_goMux_mux_onehot, isZacT_goMux_mux_mux} = {5'd1,
                                                           \call_map''_map''_Int_Int_Int_goMux2_d };
      3'd1:
        {isZacT_goMux_mux_onehot, isZacT_goMux_mux_mux} = {5'd2,
                                                           isZacT_2_2_argbuf_d};
      3'd2:
        {isZacT_goMux_mux_onehot, isZacT_goMux_mux_mux} = {5'd4,
                                                           isZacT_3_2_argbuf_d};
      3'd3:
        {isZacT_goMux_mux_onehot, isZacT_goMux_mux_mux} = {5'd8,
                                                           isZacT_4_1_argbuf_d};
      3'd4:
        {isZacT_goMux_mux_onehot, isZacT_goMux_mux_mux} = {5'd16,
                                                           lizzieLet16_1_5QNode_Int_2_argbuf_d};
      default:
        {isZacT_goMux_mux_onehot, isZacT_goMux_mux_mux} = {5'd0, 1'd0};
    endcase
  assign isZacT_goMux_mux_d = (isZacT_goMux_mux_mux[0] && go_14_goMux_choice_1_d[0]);
  assign go_14_goMux_choice_1_r = (isZacT_goMux_mux_d[0] && isZacT_goMux_mux_r);
  assign {lizzieLet16_1_5QNode_Int_2_argbuf_r,
          isZacT_4_1_argbuf_r,
          isZacT_3_2_argbuf_r,
          isZacT_2_2_argbuf_r,
          \call_map''_map''_Int_Int_Int_goMux2_r } = (go_14_goMux_choice_1_r ? isZacT_goMux_mux_onehot :
                                                      5'd0);
  
  /* mux (Ty C5,
     Ty MyDTInt_Int_Int) : (go_14_goMux_choice_2,C5) [(call_map''_map''_Int_Int_Int_goMux3,MyDTInt_Int_Int),
                                                      (gacU_2_2_argbuf,MyDTInt_Int_Int),
                                                      (gacU_3_2_argbuf,MyDTInt_Int_Int),
                                                      (gacU_4_1_argbuf,MyDTInt_Int_Int),
                                                      (lizzieLet16_1_3QNode_Int_2_argbuf,MyDTInt_Int_Int)] > (gacU_goMux_mux,MyDTInt_Int_Int) */
  logic [0:0] gacU_goMux_mux_mux;
  logic [4:0] gacU_goMux_mux_onehot;
  always_comb
    unique case (go_14_goMux_choice_2_d[3:1])
      3'd0:
        {gacU_goMux_mux_onehot, gacU_goMux_mux_mux} = {5'd1,
                                                       \call_map''_map''_Int_Int_Int_goMux3_d };
      3'd1:
        {gacU_goMux_mux_onehot, gacU_goMux_mux_mux} = {5'd2,
                                                       gacU_2_2_argbuf_d};
      3'd2:
        {gacU_goMux_mux_onehot, gacU_goMux_mux_mux} = {5'd4,
                                                       gacU_3_2_argbuf_d};
      3'd3:
        {gacU_goMux_mux_onehot, gacU_goMux_mux_mux} = {5'd8,
                                                       gacU_4_1_argbuf_d};
      3'd4:
        {gacU_goMux_mux_onehot, gacU_goMux_mux_mux} = {5'd16,
                                                       lizzieLet16_1_3QNode_Int_2_argbuf_d};
      default:
        {gacU_goMux_mux_onehot, gacU_goMux_mux_mux} = {5'd0, 1'd0};
    endcase
  assign gacU_goMux_mux_d = (gacU_goMux_mux_mux[0] && go_14_goMux_choice_2_d[0]);
  assign go_14_goMux_choice_2_r = (gacU_goMux_mux_d[0] && gacU_goMux_mux_r);
  assign {lizzieLet16_1_3QNode_Int_2_argbuf_r,
          gacU_4_1_argbuf_r,
          gacU_3_2_argbuf_r,
          gacU_2_2_argbuf_r,
          \call_map''_map''_Int_Int_Int_goMux3_r } = (go_14_goMux_choice_2_r ? gacU_goMux_mux_onehot :
                                                      5'd0);
  
  /* mux (Ty C5,
     Ty Int) : (go_14_goMux_choice_3,C5) [(call_map''_map''_Int_Int_Int_goMux4,Int),
                                          (v'acV_2_2_argbuf,Int),
                                          (v'acV_3_2_argbuf,Int),
                                          (v'acV_4_1_argbuf,Int),
                                          (lizzieLet16_1_7QNode_Int_2_argbuf,Int)] > (v'acV_goMux_mux,Int) */
  logic [32:0] \v'acV_goMux_mux_mux ;
  logic [4:0] \v'acV_goMux_mux_onehot ;
  always_comb
    unique case (go_14_goMux_choice_3_d[3:1])
      3'd0:
        {\v'acV_goMux_mux_onehot , \v'acV_goMux_mux_mux } = {5'd1,
                                                             \call_map''_map''_Int_Int_Int_goMux4_d };
      3'd1:
        {\v'acV_goMux_mux_onehot , \v'acV_goMux_mux_mux } = {5'd2,
                                                             \v'acV_2_2_argbuf_d };
      3'd2:
        {\v'acV_goMux_mux_onehot , \v'acV_goMux_mux_mux } = {5'd4,
                                                             \v'acV_3_2_argbuf_d };
      3'd3:
        {\v'acV_goMux_mux_onehot , \v'acV_goMux_mux_mux } = {5'd8,
                                                             \v'acV_4_1_argbuf_d };
      3'd4:
        {\v'acV_goMux_mux_onehot , \v'acV_goMux_mux_mux } = {5'd16,
                                                             lizzieLet16_1_7QNode_Int_2_argbuf_d};
      default:
        {\v'acV_goMux_mux_onehot , \v'acV_goMux_mux_mux } = {5'd0,
                                                             {32'd0, 1'd0}};
    endcase
  assign \v'acV_goMux_mux_d  = {\v'acV_goMux_mux_mux [32:1],
                                (\v'acV_goMux_mux_mux [0] && go_14_goMux_choice_3_d[0])};
  assign go_14_goMux_choice_3_r = (\v'acV_goMux_mux_d [0] && \v'acV_goMux_mux_r );
  assign {lizzieLet16_1_7QNode_Int_2_argbuf_r,
          \v'acV_4_1_argbuf_r ,
          \v'acV_3_2_argbuf_r ,
          \v'acV_2_2_argbuf_r ,
          \call_map''_map''_Int_Int_Int_goMux4_r } = (go_14_goMux_choice_3_r ? \v'acV_goMux_mux_onehot  :
                                                      5'd0);
  
  /* mux (Ty C5,
     Ty Pointer_QTree_Int) : (go_14_goMux_choice_4,C5) [(call_map''_map''_Int_Int_Int_goMux5,Pointer_QTree_Int),
                                                        (q3ad0_1_1_argbuf,Pointer_QTree_Int),
                                                        (q2acZ_2_1_argbuf,Pointer_QTree_Int),
                                                        (q1acY_3_1_argbuf,Pointer_QTree_Int),
                                                        (q4ad1_1_argbuf,Pointer_QTree_Int)] > (macW_goMux_mux,Pointer_QTree_Int) */
  logic [16:0] macW_goMux_mux_mux;
  logic [4:0] macW_goMux_mux_onehot;
  always_comb
    unique case (go_14_goMux_choice_4_d[3:1])
      3'd0:
        {macW_goMux_mux_onehot, macW_goMux_mux_mux} = {5'd1,
                                                       \call_map''_map''_Int_Int_Int_goMux5_d };
      3'd1:
        {macW_goMux_mux_onehot, macW_goMux_mux_mux} = {5'd2,
                                                       q3ad0_1_1_argbuf_d};
      3'd2:
        {macW_goMux_mux_onehot, macW_goMux_mux_mux} = {5'd4,
                                                       q2acZ_2_1_argbuf_d};
      3'd3:
        {macW_goMux_mux_onehot, macW_goMux_mux_mux} = {5'd8,
                                                       q1acY_3_1_argbuf_d};
      3'd4:
        {macW_goMux_mux_onehot, macW_goMux_mux_mux} = {5'd16,
                                                       q4ad1_1_argbuf_d};
      default:
        {macW_goMux_mux_onehot, macW_goMux_mux_mux} = {5'd0,
                                                       {16'd0, 1'd0}};
    endcase
  assign macW_goMux_mux_d = {macW_goMux_mux_mux[16:1],
                             (macW_goMux_mux_mux[0] && go_14_goMux_choice_4_d[0])};
  assign go_14_goMux_choice_4_r = (macW_goMux_mux_d[0] && macW_goMux_mux_r);
  assign {q4ad1_1_argbuf_r,
          q1acY_3_1_argbuf_r,
          q2acZ_2_1_argbuf_r,
          q3ad0_1_1_argbuf_r,
          \call_map''_map''_Int_Int_Int_goMux5_r } = (go_14_goMux_choice_4_r ? macW_goMux_mux_onehot :
                                                      5'd0);
  
  /* mux (Ty C5,
     Ty Pointer_CTmap''_map''_Int_Int_Int) : (go_14_goMux_choice_5,C5) [(call_map''_map''_Int_Int_Int_goMux6,Pointer_CTmap''_map''_Int_Int_Int),
                                                                        (sca2_3_1_argbuf,Pointer_CTmap''_map''_Int_Int_Int),
                                                                        (sca1_3_1_argbuf,Pointer_CTmap''_map''_Int_Int_Int),
                                                                        (sca0_3_1_argbuf,Pointer_CTmap''_map''_Int_Int_Int),
                                                                        (sca3_3_1_argbuf,Pointer_CTmap''_map''_Int_Int_Int)] > (sc_0_3_goMux_mux,Pointer_CTmap''_map''_Int_Int_Int) */
  logic [16:0] sc_0_3_goMux_mux_mux;
  logic [4:0] sc_0_3_goMux_mux_onehot;
  always_comb
    unique case (go_14_goMux_choice_5_d[3:1])
      3'd0:
        {sc_0_3_goMux_mux_onehot, sc_0_3_goMux_mux_mux} = {5'd1,
                                                           \call_map''_map''_Int_Int_Int_goMux6_d };
      3'd1:
        {sc_0_3_goMux_mux_onehot, sc_0_3_goMux_mux_mux} = {5'd2,
                                                           sca2_3_1_argbuf_d};
      3'd2:
        {sc_0_3_goMux_mux_onehot, sc_0_3_goMux_mux_mux} = {5'd4,
                                                           sca1_3_1_argbuf_d};
      3'd3:
        {sc_0_3_goMux_mux_onehot, sc_0_3_goMux_mux_mux} = {5'd8,
                                                           sca0_3_1_argbuf_d};
      3'd4:
        {sc_0_3_goMux_mux_onehot, sc_0_3_goMux_mux_mux} = {5'd16,
                                                           sca3_3_1_argbuf_d};
      default:
        {sc_0_3_goMux_mux_onehot, sc_0_3_goMux_mux_mux} = {5'd0,
                                                           {16'd0, 1'd0}};
    endcase
  assign sc_0_3_goMux_mux_d = {sc_0_3_goMux_mux_mux[16:1],
                               (sc_0_3_goMux_mux_mux[0] && go_14_goMux_choice_5_d[0])};
  assign go_14_goMux_choice_5_r = (sc_0_3_goMux_mux_d[0] && sc_0_3_goMux_mux_r);
  assign {sca3_3_1_argbuf_r,
          sca0_3_1_argbuf_r,
          sca1_3_1_argbuf_r,
          sca2_3_1_argbuf_r,
          \call_map''_map''_Int_Int_Int_goMux6_r } = (go_14_goMux_choice_5_r ? sc_0_3_goMux_mux_onehot :
                                                      5'd0);
  
  /* dcon (Ty CTkron_kron_Int_Int_Int,
      Dcon Lkron_kron_Int_Int_Intsbos) : [(go_15_1,Go)] > (go_15_1Lkron_kron_Int_Int_Intsbos,CTkron_kron_Int_Int_Int) */
  assign go_15_1Lkron_kron_Int_Int_Intsbos_d = Lkron_kron_Int_Int_Intsbos_dc((& {go_15_1_d[0]}), go_15_1_d);
  assign {go_15_1_r} = {1 {(go_15_1Lkron_kron_Int_Int_Intsbos_r && go_15_1Lkron_kron_Int_Int_Intsbos_d[0])}};
  
  /* buf (Ty CTkron_kron_Int_Int_Int) : (go_15_1Lkron_kron_Int_Int_Intsbos,CTkron_kron_Int_Int_Int) > (lizzieLet22_1_argbuf,CTkron_kron_Int_Int_Int) */
  CTkron_kron_Int_Int_Int_t go_15_1Lkron_kron_Int_Int_Intsbos_bufchan_d;
  logic go_15_1Lkron_kron_Int_Int_Intsbos_bufchan_r;
  assign go_15_1Lkron_kron_Int_Int_Intsbos_r = ((! go_15_1Lkron_kron_Int_Int_Intsbos_bufchan_d[0]) || go_15_1Lkron_kron_Int_Int_Intsbos_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      go_15_1Lkron_kron_Int_Int_Intsbos_bufchan_d <= {83'd0, 1'd0};
    else
      if (go_15_1Lkron_kron_Int_Int_Intsbos_r)
        go_15_1Lkron_kron_Int_Int_Intsbos_bufchan_d <= go_15_1Lkron_kron_Int_Int_Intsbos_d;
  CTkron_kron_Int_Int_Int_t go_15_1Lkron_kron_Int_Int_Intsbos_bufchan_buf;
  assign go_15_1Lkron_kron_Int_Int_Intsbos_bufchan_r = (! go_15_1Lkron_kron_Int_Int_Intsbos_bufchan_buf[0]);
  assign lizzieLet22_1_argbuf_d = (go_15_1Lkron_kron_Int_Int_Intsbos_bufchan_buf[0] ? go_15_1Lkron_kron_Int_Int_Intsbos_bufchan_buf :
                                   go_15_1Lkron_kron_Int_Int_Intsbos_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      go_15_1Lkron_kron_Int_Int_Intsbos_bufchan_buf <= {83'd0, 1'd0};
    else
      if ((lizzieLet22_1_argbuf_r && go_15_1Lkron_kron_Int_Int_Intsbos_bufchan_buf[0]))
        go_15_1Lkron_kron_Int_Int_Intsbos_bufchan_buf <= {83'd0, 1'd0};
      else if (((! lizzieLet22_1_argbuf_r) && (! go_15_1Lkron_kron_Int_Int_Intsbos_bufchan_buf[0])))
        go_15_1Lkron_kron_Int_Int_Intsbos_bufchan_buf <= go_15_1Lkron_kron_Int_Int_Intsbos_bufchan_d;
  
  /* buf (Ty Go) : (go_15_2,Go) > (go_15_2_argbuf,Go) */
  Go_t go_15_2_bufchan_d;
  logic go_15_2_bufchan_r;
  assign go_15_2_r = ((! go_15_2_bufchan_d[0]) || go_15_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_15_2_bufchan_d <= 1'd0;
    else if (go_15_2_r) go_15_2_bufchan_d <= go_15_2_d;
  Go_t go_15_2_bufchan_buf;
  assign go_15_2_bufchan_r = (! go_15_2_bufchan_buf[0]);
  assign go_15_2_argbuf_d = (go_15_2_bufchan_buf[0] ? go_15_2_bufchan_buf :
                             go_15_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_15_2_bufchan_buf <= 1'd0;
    else
      if ((go_15_2_argbuf_r && go_15_2_bufchan_buf[0]))
        go_15_2_bufchan_buf <= 1'd0;
      else if (((! go_15_2_argbuf_r) && (! go_15_2_bufchan_buf[0])))
        go_15_2_bufchan_buf <= go_15_2_bufchan_d;
  
  /* dcon (Ty TupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Int,
      Dcon TupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Int) : [(go_15_2_argbuf,Go),
                                                                                                                                (isZad2_1_1_argbuf,MyDTInt_Bool),
                                                                                                                                (gad3_1_1_argbuf,MyDTInt_Int_Int),
                                                                                                                                (m1ad4_1_1_argbuf,Pointer_QTree_Int),
                                                                                                                                (m2ad5_1_1_argbuf,Pointer_QTree_Int),
                                                                                                                                (lizzieLet14_1_1_argbuf,Pointer_CTkron_kron_Int_Int_Int)] > (call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Int_1,TupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Int) */
  assign call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Int_1_d = TupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Int_dc((& {go_15_2_argbuf_d[0],
                                                                                                                                                                                                                                                                                  isZad2_1_1_argbuf_d[0],
                                                                                                                                                                                                                                                                                  gad3_1_1_argbuf_d[0],
                                                                                                                                                                                                                                                                                  m1ad4_1_1_argbuf_d[0],
                                                                                                                                                                                                                                                                                  m2ad5_1_1_argbuf_d[0],
                                                                                                                                                                                                                                                                                  lizzieLet14_1_1_argbuf_d[0]}), go_15_2_argbuf_d, isZad2_1_1_argbuf_d, gad3_1_1_argbuf_d, m1ad4_1_1_argbuf_d, m2ad5_1_1_argbuf_d, lizzieLet14_1_1_argbuf_d);
  assign {go_15_2_argbuf_r,
          isZad2_1_1_argbuf_r,
          gad3_1_1_argbuf_r,
          m1ad4_1_1_argbuf_r,
          m2ad5_1_1_argbuf_r,
          lizzieLet14_1_1_argbuf_r} = {6 {(call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Int_1_r && call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Int_1_d[0])}};
  
  /* dcon (Ty CTmain_map'_Int_Int,
      Dcon Lmain_map'_Int_Intsbos) : [(go_16_1,Go)] > (go_16_1Lmain_map'_Int_Intsbos,CTmain_map'_Int_Int) */
  assign \go_16_1Lmain_map'_Int_Intsbos_d  = \Lmain_map'_Int_Intsbos_dc ((& {go_16_1_d[0]}), go_16_1_d);
  assign {go_16_1_r} = {1 {(\go_16_1Lmain_map'_Int_Intsbos_r  && \go_16_1Lmain_map'_Int_Intsbos_d [0])}};
  
  /* buf (Ty CTmain_map'_Int_Int) : (go_16_1Lmain_map'_Int_Intsbos,CTmain_map'_Int_Int) > (lizzieLet23_1_argbuf,CTmain_map'_Int_Int) */
  \CTmain_map'_Int_Int_t  \go_16_1Lmain_map'_Int_Intsbos_bufchan_d ;
  logic \go_16_1Lmain_map'_Int_Intsbos_bufchan_r ;
  assign \go_16_1Lmain_map'_Int_Intsbos_r  = ((! \go_16_1Lmain_map'_Int_Intsbos_bufchan_d [0]) || \go_16_1Lmain_map'_Int_Intsbos_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \go_16_1Lmain_map'_Int_Intsbos_bufchan_d  <= {67'd0, 1'd0};
    else
      if (\go_16_1Lmain_map'_Int_Intsbos_r )
        \go_16_1Lmain_map'_Int_Intsbos_bufchan_d  <= \go_16_1Lmain_map'_Int_Intsbos_d ;
  \CTmain_map'_Int_Int_t  \go_16_1Lmain_map'_Int_Intsbos_bufchan_buf ;
  assign \go_16_1Lmain_map'_Int_Intsbos_bufchan_r  = (! \go_16_1Lmain_map'_Int_Intsbos_bufchan_buf [0]);
  assign lizzieLet23_1_argbuf_d = (\go_16_1Lmain_map'_Int_Intsbos_bufchan_buf [0] ? \go_16_1Lmain_map'_Int_Intsbos_bufchan_buf  :
                                   \go_16_1Lmain_map'_Int_Intsbos_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \go_16_1Lmain_map'_Int_Intsbos_bufchan_buf  <= {67'd0, 1'd0};
    else
      if ((lizzieLet23_1_argbuf_r && \go_16_1Lmain_map'_Int_Intsbos_bufchan_buf [0]))
        \go_16_1Lmain_map'_Int_Intsbos_bufchan_buf  <= {67'd0, 1'd0};
      else if (((! lizzieLet23_1_argbuf_r) && (! \go_16_1Lmain_map'_Int_Intsbos_bufchan_buf [0])))
        \go_16_1Lmain_map'_Int_Intsbos_bufchan_buf  <= \go_16_1Lmain_map'_Int_Intsbos_bufchan_d ;
  
  /* buf (Ty Go) : (go_16_2,Go) > (go_16_2_argbuf,Go) */
  Go_t go_16_2_bufchan_d;
  logic go_16_2_bufchan_r;
  assign go_16_2_r = ((! go_16_2_bufchan_d[0]) || go_16_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_16_2_bufchan_d <= 1'd0;
    else if (go_16_2_r) go_16_2_bufchan_d <= go_16_2_d;
  Go_t go_16_2_bufchan_buf;
  assign go_16_2_bufchan_r = (! go_16_2_bufchan_buf[0]);
  assign go_16_2_argbuf_d = (go_16_2_bufchan_buf[0] ? go_16_2_bufchan_buf :
                             go_16_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_16_2_bufchan_buf <= 1'd0;
    else
      if ((go_16_2_argbuf_r && go_16_2_bufchan_buf[0]))
        go_16_2_bufchan_buf <= 1'd0;
      else if (((! go_16_2_argbuf_r) && (! go_16_2_bufchan_buf[0])))
        go_16_2_bufchan_buf <= go_16_2_bufchan_d;
  
  /* dcon (Ty TupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Int,
      Dcon TupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Int) : [(go_16_2_argbuf,Go),
                                                                                                    (isZacL_1_1_argbuf,MyDTInt_Bool),
                                                                                                    (gacM_1_1_argbuf,MyDTInt_Int),
                                                                                                    (macN_1_1_argbuf,Pointer_QTree_Int),
                                                                                                    (lizzieLet5_1_1_argbuf,Pointer_CTmain_map'_Int_Int)] > (call_main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Int_1,TupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Int) */
  assign \call_main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Int_1_d  = \TupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Int_dc ((& {go_16_2_argbuf_d[0],
                                                                                                                                                                                                                          isZacL_1_1_argbuf_d[0],
                                                                                                                                                                                                                          gacM_1_1_argbuf_d[0],
                                                                                                                                                                                                                          macN_1_1_argbuf_d[0],
                                                                                                                                                                                                                          lizzieLet5_1_1_argbuf_d[0]}), go_16_2_argbuf_d, isZacL_1_1_argbuf_d, gacM_1_1_argbuf_d, macN_1_1_argbuf_d, lizzieLet5_1_1_argbuf_d);
  assign {go_16_2_argbuf_r,
          isZacL_1_1_argbuf_r,
          gacM_1_1_argbuf_r,
          macN_1_1_argbuf_r,
          lizzieLet5_1_1_argbuf_r} = {5 {(\call_main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Int_1_r  && \call_main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Int_1_d [0])}};
  
  /* dcon (Ty CTmap''_map''_Int_Int_Int,
      Dcon Lmap''_map''_Int_Int_Intsbos) : [(go_17_1,Go)] > (go_17_1Lmap''_map''_Int_Int_Intsbos,CTmap''_map''_Int_Int_Int) */
  assign \go_17_1Lmap''_map''_Int_Int_Intsbos_d  = \Lmap''_map''_Int_Int_Intsbos_dc ((& {go_17_1_d[0]}), go_17_1_d);
  assign {go_17_1_r} = {1 {(\go_17_1Lmap''_map''_Int_Int_Intsbos_r  && \go_17_1Lmap''_map''_Int_Int_Intsbos_d [0])}};
  
  /* buf (Ty CTmap''_map''_Int_Int_Int) : (go_17_1Lmap''_map''_Int_Int_Intsbos,CTmap''_map''_Int_Int_Int) > (lizzieLet24_1_argbuf,CTmap''_map''_Int_Int_Int) */
  \CTmap''_map''_Int_Int_Int_t  \go_17_1Lmap''_map''_Int_Int_Intsbos_bufchan_d ;
  logic \go_17_1Lmap''_map''_Int_Int_Intsbos_bufchan_r ;
  assign \go_17_1Lmap''_map''_Int_Int_Intsbos_r  = ((! \go_17_1Lmap''_map''_Int_Int_Intsbos_bufchan_d [0]) || \go_17_1Lmap''_map''_Int_Int_Intsbos_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \go_17_1Lmap''_map''_Int_Int_Intsbos_bufchan_d  <= {99'd0, 1'd0};
    else
      if (\go_17_1Lmap''_map''_Int_Int_Intsbos_r )
        \go_17_1Lmap''_map''_Int_Int_Intsbos_bufchan_d  <= \go_17_1Lmap''_map''_Int_Int_Intsbos_d ;
  \CTmap''_map''_Int_Int_Int_t  \go_17_1Lmap''_map''_Int_Int_Intsbos_bufchan_buf ;
  assign \go_17_1Lmap''_map''_Int_Int_Intsbos_bufchan_r  = (! \go_17_1Lmap''_map''_Int_Int_Intsbos_bufchan_buf [0]);
  assign lizzieLet24_1_argbuf_d = (\go_17_1Lmap''_map''_Int_Int_Intsbos_bufchan_buf [0] ? \go_17_1Lmap''_map''_Int_Int_Intsbos_bufchan_buf  :
                                   \go_17_1Lmap''_map''_Int_Int_Intsbos_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \go_17_1Lmap''_map''_Int_Int_Intsbos_bufchan_buf  <= {99'd0, 1'd0};
    else
      if ((lizzieLet24_1_argbuf_r && \go_17_1Lmap''_map''_Int_Int_Intsbos_bufchan_buf [0]))
        \go_17_1Lmap''_map''_Int_Int_Intsbos_bufchan_buf  <= {99'd0, 1'd0};
      else if (((! lizzieLet24_1_argbuf_r) && (! \go_17_1Lmap''_map''_Int_Int_Intsbos_bufchan_buf [0])))
        \go_17_1Lmap''_map''_Int_Int_Intsbos_bufchan_buf  <= \go_17_1Lmap''_map''_Int_Int_Intsbos_bufchan_d ;
  
  /* buf (Ty Go) : (go_17_2,Go) > (go_17_2_argbuf,Go) */
  Go_t go_17_2_bufchan_d;
  logic go_17_2_bufchan_r;
  assign go_17_2_r = ((! go_17_2_bufchan_d[0]) || go_17_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_17_2_bufchan_d <= 1'd0;
    else if (go_17_2_r) go_17_2_bufchan_d <= go_17_2_d;
  Go_t go_17_2_bufchan_buf;
  assign go_17_2_bufchan_r = (! go_17_2_bufchan_buf[0]);
  assign go_17_2_argbuf_d = (go_17_2_bufchan_buf[0] ? go_17_2_bufchan_buf :
                             go_17_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_17_2_bufchan_buf <= 1'd0;
    else
      if ((go_17_2_argbuf_r && go_17_2_bufchan_buf[0]))
        go_17_2_bufchan_buf <= 1'd0;
      else if (((! go_17_2_argbuf_r) && (! go_17_2_bufchan_buf[0])))
        go_17_2_bufchan_buf <= go_17_2_bufchan_d;
  
  /* dcon (Ty TupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Int,
      Dcon TupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Int) : [(go_17_2_argbuf,Go),
                                                                                                                    (isZacT_1_1_argbuf,MyDTInt_Bool),
                                                                                                                    (gacU_1_1_argbuf,MyDTInt_Int_Int),
                                                                                                                    (v'acV_1_1_argbuf,Int),
                                                                                                                    (macW_1_1_argbuf,Pointer_QTree_Int),
                                                                                                                    (lizzieLet10_1_1_argbuf,Pointer_CTmap''_map''_Int_Int_Int)] > (call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Int_1,TupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Int) */
  assign \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Int_1_d  = \TupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Int_dc ((& {go_17_2_argbuf_d[0],
                                                                                                                                                                                                                                                                isZacT_1_1_argbuf_d[0],
                                                                                                                                                                                                                                                                gacU_1_1_argbuf_d[0],
                                                                                                                                                                                                                                                                \v'acV_1_1_argbuf_d [0],
                                                                                                                                                                                                                                                                macW_1_1_argbuf_d[0],
                                                                                                                                                                                                                                                                lizzieLet10_1_1_argbuf_d[0]}), go_17_2_argbuf_d, isZacT_1_1_argbuf_d, gacU_1_1_argbuf_d, \v'acV_1_1_argbuf_d , macW_1_1_argbuf_d, lizzieLet10_1_1_argbuf_d);
  assign {go_17_2_argbuf_r,
          isZacT_1_1_argbuf_r,
          gacU_1_1_argbuf_r,
          \v'acV_1_1_argbuf_r ,
          macW_1_1_argbuf_r,
          lizzieLet10_1_1_argbuf_r} = {6 {(\call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Int_1_r  && \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Int_1_d [0])}};
  
  /* fork (Ty C4) : (go_18_goMux_choice,C4) > [(go_18_goMux_choice_1,C4),
                                          (go_18_goMux_choice_2,C4)] */
  logic [1:0] go_18_goMux_choice_emitted;
  logic [1:0] go_18_goMux_choice_done;
  assign go_18_goMux_choice_1_d = {go_18_goMux_choice_d[2:1],
                                   (go_18_goMux_choice_d[0] && (! go_18_goMux_choice_emitted[0]))};
  assign go_18_goMux_choice_2_d = {go_18_goMux_choice_d[2:1],
                                   (go_18_goMux_choice_d[0] && (! go_18_goMux_choice_emitted[1]))};
  assign go_18_goMux_choice_done = (go_18_goMux_choice_emitted | ({go_18_goMux_choice_2_d[0],
                                                                   go_18_goMux_choice_1_d[0]} & {go_18_goMux_choice_2_r,
                                                                                                 go_18_goMux_choice_1_r}));
  assign go_18_goMux_choice_r = (& go_18_goMux_choice_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_18_goMux_choice_emitted <= 2'd0;
    else
      go_18_goMux_choice_emitted <= (go_18_goMux_choice_r ? 2'd0 :
                                     go_18_goMux_choice_done);
  
  /* mux (Ty C4,
     Ty Int#) : (go_18_goMux_choice_1,C4) [(lizzieLet15_1_argbuf,Int#),
                                           (contRet_0_1_argbuf,Int#),
                                           (lizzieLet16_1_argbuf,Int#),
                                           (lizzieLet15_1_1_argbuf,Int#)] > (srtarg_0_goMux_mux,Int#) */
  logic [32:0] srtarg_0_goMux_mux_mux;
  logic [3:0] srtarg_0_goMux_mux_onehot;
  always_comb
    unique case (go_18_goMux_choice_1_d[2:1])
      2'd0:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {4'd1,
                                                               lizzieLet15_1_argbuf_d};
      2'd1:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {4'd2,
                                                               contRet_0_1_argbuf_d};
      2'd2:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {4'd4,
                                                               lizzieLet16_1_argbuf_d};
      2'd3:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {4'd8,
                                                               lizzieLet15_1_1_argbuf_d};
      default:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {4'd0,
                                                               {32'd0, 1'd0}};
    endcase
  assign srtarg_0_goMux_mux_d = {srtarg_0_goMux_mux_mux[32:1],
                                 (srtarg_0_goMux_mux_mux[0] && go_18_goMux_choice_1_d[0])};
  assign go_18_goMux_choice_1_r = (srtarg_0_goMux_mux_d[0] && srtarg_0_goMux_mux_r);
  assign {lizzieLet15_1_1_argbuf_r,
          lizzieLet16_1_argbuf_r,
          contRet_0_1_argbuf_r,
          lizzieLet15_1_argbuf_r} = (go_18_goMux_choice_1_r ? srtarg_0_goMux_mux_onehot :
                                     4'd0);
  
  /* mux (Ty C4,
     Ty Pointer_CT$wnnz_Int) : (go_18_goMux_choice_2,C4) [(lizzieLet4_4QNone_Int_1_argbuf,Pointer_CT$wnnz_Int),
                                                          (sc_0_7_1_argbuf,Pointer_CT$wnnz_Int),
                                                          (lizzieLet4_4QVal_Int_1_argbuf,Pointer_CT$wnnz_Int),
                                                          (lizzieLet4_4QError_Int_1_argbuf,Pointer_CT$wnnz_Int)] > (scfarg_0_goMux_mux,Pointer_CT$wnnz_Int) */
  logic [16:0] scfarg_0_goMux_mux_mux;
  logic [3:0] scfarg_0_goMux_mux_onehot;
  always_comb
    unique case (go_18_goMux_choice_2_d[2:1])
      2'd0:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {4'd1,
                                                               lizzieLet4_4QNone_Int_1_argbuf_d};
      2'd1:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {4'd2,
                                                               sc_0_7_1_argbuf_d};
      2'd2:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {4'd4,
                                                               lizzieLet4_4QVal_Int_1_argbuf_d};
      2'd3:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {4'd8,
                                                               lizzieLet4_4QError_Int_1_argbuf_d};
      default:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {4'd0,
                                                               {16'd0, 1'd0}};
    endcase
  assign scfarg_0_goMux_mux_d = {scfarg_0_goMux_mux_mux[16:1],
                                 (scfarg_0_goMux_mux_mux[0] && go_18_goMux_choice_2_d[0])};
  assign go_18_goMux_choice_2_r = (scfarg_0_goMux_mux_d[0] && scfarg_0_goMux_mux_r);
  assign {lizzieLet4_4QError_Int_1_argbuf_r,
          lizzieLet4_4QVal_Int_1_argbuf_r,
          sc_0_7_1_argbuf_r,
          lizzieLet4_4QNone_Int_1_argbuf_r} = (go_18_goMux_choice_2_r ? scfarg_0_goMux_mux_onehot :
                                               4'd0);
  
  /* fork (Ty C4) : (go_19_goMux_choice,C4) > [(go_19_goMux_choice_1,C4),
                                          (go_19_goMux_choice_2,C4)] */
  logic [1:0] go_19_goMux_choice_emitted;
  logic [1:0] go_19_goMux_choice_done;
  assign go_19_goMux_choice_1_d = {go_19_goMux_choice_d[2:1],
                                   (go_19_goMux_choice_d[0] && (! go_19_goMux_choice_emitted[0]))};
  assign go_19_goMux_choice_2_d = {go_19_goMux_choice_d[2:1],
                                   (go_19_goMux_choice_d[0] && (! go_19_goMux_choice_emitted[1]))};
  assign go_19_goMux_choice_done = (go_19_goMux_choice_emitted | ({go_19_goMux_choice_2_d[0],
                                                                   go_19_goMux_choice_1_d[0]} & {go_19_goMux_choice_2_r,
                                                                                                 go_19_goMux_choice_1_r}));
  assign go_19_goMux_choice_r = (& go_19_goMux_choice_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_19_goMux_choice_emitted <= 2'd0;
    else
      go_19_goMux_choice_emitted <= (go_19_goMux_choice_r ? 2'd0 :
                                     go_19_goMux_choice_done);
  
  /* mux (Ty C4,
     Ty Pointer_QTree_Int) : (go_19_goMux_choice_1,C4) [(lizzieLet11_1_argbuf,Pointer_QTree_Int),
                                                        (contRet_0_1_1_argbuf,Pointer_QTree_Int),
                                                        (lizzieLet12_1_argbuf,Pointer_QTree_Int),
                                                        (lizzieLet13_1_argbuf,Pointer_QTree_Int)] > (srtarg_0_1_goMux_mux,Pointer_QTree_Int) */
  logic [16:0] srtarg_0_1_goMux_mux_mux;
  logic [3:0] srtarg_0_1_goMux_mux_onehot;
  always_comb
    unique case (go_19_goMux_choice_1_d[2:1])
      2'd0:
        {srtarg_0_1_goMux_mux_onehot, srtarg_0_1_goMux_mux_mux} = {4'd1,
                                                                   lizzieLet11_1_argbuf_d};
      2'd1:
        {srtarg_0_1_goMux_mux_onehot, srtarg_0_1_goMux_mux_mux} = {4'd2,
                                                                   contRet_0_1_1_argbuf_d};
      2'd2:
        {srtarg_0_1_goMux_mux_onehot, srtarg_0_1_goMux_mux_mux} = {4'd4,
                                                                   lizzieLet12_1_argbuf_d};
      2'd3:
        {srtarg_0_1_goMux_mux_onehot, srtarg_0_1_goMux_mux_mux} = {4'd8,
                                                                   lizzieLet13_1_argbuf_d};
      default:
        {srtarg_0_1_goMux_mux_onehot, srtarg_0_1_goMux_mux_mux} = {4'd0,
                                                                   {16'd0, 1'd0}};
    endcase
  assign srtarg_0_1_goMux_mux_d = {srtarg_0_1_goMux_mux_mux[16:1],
                                   (srtarg_0_1_goMux_mux_mux[0] && go_19_goMux_choice_1_d[0])};
  assign go_19_goMux_choice_1_r = (srtarg_0_1_goMux_mux_d[0] && srtarg_0_1_goMux_mux_r);
  assign {lizzieLet13_1_argbuf_r,
          lizzieLet12_1_argbuf_r,
          contRet_0_1_1_argbuf_r,
          lizzieLet11_1_argbuf_r} = (go_19_goMux_choice_1_r ? srtarg_0_1_goMux_mux_onehot :
                                     4'd0);
  
  /* mux (Ty C4,
     Ty Pointer_CTkron_kron_Int_Int_Int) : (go_19_goMux_choice_2,C4) [(lizzieLet6_7QNone_Int_1_argbuf,Pointer_CTkron_kron_Int_Int_Int),
                                                                      (sc_0_11_1_argbuf,Pointer_CTkron_kron_Int_Int_Int),
                                                                      (lizzieLet6_7QVal_Int_1_argbuf,Pointer_CTkron_kron_Int_Int_Int),
                                                                      (lizzieLet6_7QError_Int_1_argbuf,Pointer_CTkron_kron_Int_Int_Int)] > (scfarg_0_1_goMux_mux,Pointer_CTkron_kron_Int_Int_Int) */
  logic [16:0] scfarg_0_1_goMux_mux_mux;
  logic [3:0] scfarg_0_1_goMux_mux_onehot;
  always_comb
    unique case (go_19_goMux_choice_2_d[2:1])
      2'd0:
        {scfarg_0_1_goMux_mux_onehot, scfarg_0_1_goMux_mux_mux} = {4'd1,
                                                                   lizzieLet6_7QNone_Int_1_argbuf_d};
      2'd1:
        {scfarg_0_1_goMux_mux_onehot, scfarg_0_1_goMux_mux_mux} = {4'd2,
                                                                   sc_0_11_1_argbuf_d};
      2'd2:
        {scfarg_0_1_goMux_mux_onehot, scfarg_0_1_goMux_mux_mux} = {4'd4,
                                                                   lizzieLet6_7QVal_Int_1_argbuf_d};
      2'd3:
        {scfarg_0_1_goMux_mux_onehot, scfarg_0_1_goMux_mux_mux} = {4'd8,
                                                                   lizzieLet6_7QError_Int_1_argbuf_d};
      default:
        {scfarg_0_1_goMux_mux_onehot, scfarg_0_1_goMux_mux_mux} = {4'd0,
                                                                   {16'd0, 1'd0}};
    endcase
  assign scfarg_0_1_goMux_mux_d = {scfarg_0_1_goMux_mux_mux[16:1],
                                   (scfarg_0_1_goMux_mux_mux[0] && go_19_goMux_choice_2_d[0])};
  assign go_19_goMux_choice_2_r = (scfarg_0_1_goMux_mux_d[0] && scfarg_0_1_goMux_mux_r);
  assign {lizzieLet6_7QError_Int_1_argbuf_r,
          lizzieLet6_7QVal_Int_1_argbuf_r,
          sc_0_11_1_argbuf_r,
          lizzieLet6_7QNone_Int_1_argbuf_r} = (go_19_goMux_choice_2_r ? scfarg_0_1_goMux_mux_onehot :
                                               4'd0);
  
  /* dcon (Ty TupGo___Pointer_QTree_Int___Pointer_QTree_Int,
      Dcon TupGo___Pointer_QTree_Int___Pointer_QTree_Int) : [(go_1_argbuf,Go),
                                                             (wsvA_1_0,Pointer_QTree_Int),
                                                             (w1svB_1_1,Pointer_QTree_Int)] > ($wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Int_1,TupGo___Pointer_QTree_Int___Pointer_QTree_Int) */
  assign \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Int_1_d  = TupGo___Pointer_QTree_Int___Pointer_QTree_Int_dc((& {go_1_argbuf_d[0],
                                                                                                                          wsvA_1_0_d[0],
                                                                                                                          w1svB_1_1_d[0]}), go_1_argbuf_d, wsvA_1_0_d, w1svB_1_1_d);
  assign {go_1_argbuf_r,
          wsvA_1_0_r,
          w1svB_1_1_r} = {3 {(\$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Int_1_r  && \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Int_1_d [0])}};
  
  /* fork (Ty C5) : (go_20_goMux_choice,C5) > [(go_20_goMux_choice_1,C5),
                                          (go_20_goMux_choice_2,C5)] */
  logic [1:0] go_20_goMux_choice_emitted;
  logic [1:0] go_20_goMux_choice_done;
  assign go_20_goMux_choice_1_d = {go_20_goMux_choice_d[3:1],
                                   (go_20_goMux_choice_d[0] && (! go_20_goMux_choice_emitted[0]))};
  assign go_20_goMux_choice_2_d = {go_20_goMux_choice_d[3:1],
                                   (go_20_goMux_choice_d[0] && (! go_20_goMux_choice_emitted[1]))};
  assign go_20_goMux_choice_done = (go_20_goMux_choice_emitted | ({go_20_goMux_choice_2_d[0],
                                                                   go_20_goMux_choice_1_d[0]} & {go_20_goMux_choice_2_r,
                                                                                                 go_20_goMux_choice_1_r}));
  assign go_20_goMux_choice_r = (& go_20_goMux_choice_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_20_goMux_choice_emitted <= 2'd0;
    else
      go_20_goMux_choice_emitted <= (go_20_goMux_choice_r ? 2'd0 :
                                     go_20_goMux_choice_done);
  
  /* mux (Ty C5,
     Ty Pointer_QTree_Int) : (go_20_goMux_choice_1,C5) [(lizzieLet1_1_1_argbuf,Pointer_QTree_Int),
                                                        (contRet_0_2_1_argbuf,Pointer_QTree_Int),
                                                        (lizzieLet2_1_1_argbuf,Pointer_QTree_Int),
                                                        (lizzieLet3_1_1_argbuf,Pointer_QTree_Int),
                                                        (lizzieLet4_1_1_argbuf,Pointer_QTree_Int)] > (srtarg_0_2_goMux_mux,Pointer_QTree_Int) */
  logic [16:0] srtarg_0_2_goMux_mux_mux;
  logic [4:0] srtarg_0_2_goMux_mux_onehot;
  always_comb
    unique case (go_20_goMux_choice_1_d[3:1])
      3'd0:
        {srtarg_0_2_goMux_mux_onehot, srtarg_0_2_goMux_mux_mux} = {5'd1,
                                                                   lizzieLet1_1_1_argbuf_d};
      3'd1:
        {srtarg_0_2_goMux_mux_onehot, srtarg_0_2_goMux_mux_mux} = {5'd2,
                                                                   contRet_0_2_1_argbuf_d};
      3'd2:
        {srtarg_0_2_goMux_mux_onehot, srtarg_0_2_goMux_mux_mux} = {5'd4,
                                                                   lizzieLet2_1_1_argbuf_d};
      3'd3:
        {srtarg_0_2_goMux_mux_onehot, srtarg_0_2_goMux_mux_mux} = {5'd8,
                                                                   lizzieLet3_1_1_argbuf_d};
      3'd4:
        {srtarg_0_2_goMux_mux_onehot, srtarg_0_2_goMux_mux_mux} = {5'd16,
                                                                   lizzieLet4_1_1_argbuf_d};
      default:
        {srtarg_0_2_goMux_mux_onehot, srtarg_0_2_goMux_mux_mux} = {5'd0,
                                                                   {16'd0, 1'd0}};
    endcase
  assign srtarg_0_2_goMux_mux_d = {srtarg_0_2_goMux_mux_mux[16:1],
                                   (srtarg_0_2_goMux_mux_mux[0] && go_20_goMux_choice_1_d[0])};
  assign go_20_goMux_choice_1_r = (srtarg_0_2_goMux_mux_d[0] && srtarg_0_2_goMux_mux_r);
  assign {lizzieLet4_1_1_argbuf_r,
          lizzieLet3_1_1_argbuf_r,
          lizzieLet2_1_1_argbuf_r,
          contRet_0_2_1_argbuf_r,
          lizzieLet1_1_1_argbuf_r} = (go_20_goMux_choice_1_r ? srtarg_0_2_goMux_mux_onehot :
                                      5'd0);
  
  /* mux (Ty C5,
     Ty Pointer_CTmain_map'_Int_Int) : (go_20_goMux_choice_2,C5) [(lizzieLet10_6QNone_Int_1_argbuf,Pointer_CTmain_map'_Int_Int),
                                                                  (sc_0_15_1_argbuf,Pointer_CTmain_map'_Int_Int),
                                                                  (es_0_4_2MyFalse_1_argbuf,Pointer_CTmain_map'_Int_Int),
                                                                  (es_0_4_2MyTrue_1_argbuf,Pointer_CTmain_map'_Int_Int),
                                                                  (lizzieLet10_6QError_Int_1_argbuf,Pointer_CTmain_map'_Int_Int)] > (scfarg_0_2_goMux_mux,Pointer_CTmain_map'_Int_Int) */
  logic [16:0] scfarg_0_2_goMux_mux_mux;
  logic [4:0] scfarg_0_2_goMux_mux_onehot;
  always_comb
    unique case (go_20_goMux_choice_2_d[3:1])
      3'd0:
        {scfarg_0_2_goMux_mux_onehot, scfarg_0_2_goMux_mux_mux} = {5'd1,
                                                                   lizzieLet10_6QNone_Int_1_argbuf_d};
      3'd1:
        {scfarg_0_2_goMux_mux_onehot, scfarg_0_2_goMux_mux_mux} = {5'd2,
                                                                   sc_0_15_1_argbuf_d};
      3'd2:
        {scfarg_0_2_goMux_mux_onehot, scfarg_0_2_goMux_mux_mux} = {5'd4,
                                                                   es_0_4_2MyFalse_1_argbuf_d};
      3'd3:
        {scfarg_0_2_goMux_mux_onehot, scfarg_0_2_goMux_mux_mux} = {5'd8,
                                                                   es_0_4_2MyTrue_1_argbuf_d};
      3'd4:
        {scfarg_0_2_goMux_mux_onehot, scfarg_0_2_goMux_mux_mux} = {5'd16,
                                                                   lizzieLet10_6QError_Int_1_argbuf_d};
      default:
        {scfarg_0_2_goMux_mux_onehot, scfarg_0_2_goMux_mux_mux} = {5'd0,
                                                                   {16'd0, 1'd0}};
    endcase
  assign scfarg_0_2_goMux_mux_d = {scfarg_0_2_goMux_mux_mux[16:1],
                                   (scfarg_0_2_goMux_mux_mux[0] && go_20_goMux_choice_2_d[0])};
  assign go_20_goMux_choice_2_r = (scfarg_0_2_goMux_mux_d[0] && scfarg_0_2_goMux_mux_r);
  assign {lizzieLet10_6QError_Int_1_argbuf_r,
          es_0_4_2MyTrue_1_argbuf_r,
          es_0_4_2MyFalse_1_argbuf_r,
          sc_0_15_1_argbuf_r,
          lizzieLet10_6QNone_Int_1_argbuf_r} = (go_20_goMux_choice_2_r ? scfarg_0_2_goMux_mux_onehot :
                                                5'd0);
  
  /* fork (Ty C5) : (go_21_goMux_choice,C5) > [(go_21_goMux_choice_1,C5),
                                          (go_21_goMux_choice_2,C5)] */
  logic [1:0] go_21_goMux_choice_emitted;
  logic [1:0] go_21_goMux_choice_done;
  assign go_21_goMux_choice_1_d = {go_21_goMux_choice_d[3:1],
                                   (go_21_goMux_choice_d[0] && (! go_21_goMux_choice_emitted[0]))};
  assign go_21_goMux_choice_2_d = {go_21_goMux_choice_d[3:1],
                                   (go_21_goMux_choice_d[0] && (! go_21_goMux_choice_emitted[1]))};
  assign go_21_goMux_choice_done = (go_21_goMux_choice_emitted | ({go_21_goMux_choice_2_d[0],
                                                                   go_21_goMux_choice_1_d[0]} & {go_21_goMux_choice_2_r,
                                                                                                 go_21_goMux_choice_1_r}));
  assign go_21_goMux_choice_r = (& go_21_goMux_choice_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_21_goMux_choice_emitted <= 2'd0;
    else
      go_21_goMux_choice_emitted <= (go_21_goMux_choice_r ? 2'd0 :
                                     go_21_goMux_choice_done);
  
  /* mux (Ty C5,
     Ty Pointer_QTree_Int) : (go_21_goMux_choice_1,C5) [(lizzieLet6_1_1_argbuf,Pointer_QTree_Int),
                                                        (contRet_0_3_1_argbuf,Pointer_QTree_Int),
                                                        (lizzieLet7_1_1_argbuf,Pointer_QTree_Int),
                                                        (lizzieLet8_1_1_argbuf,Pointer_QTree_Int),
                                                        (lizzieLet9_1_1_argbuf,Pointer_QTree_Int)] > (srtarg_0_3_goMux_mux,Pointer_QTree_Int) */
  logic [16:0] srtarg_0_3_goMux_mux_mux;
  logic [4:0] srtarg_0_3_goMux_mux_onehot;
  always_comb
    unique case (go_21_goMux_choice_1_d[3:1])
      3'd0:
        {srtarg_0_3_goMux_mux_onehot, srtarg_0_3_goMux_mux_mux} = {5'd1,
                                                                   lizzieLet6_1_1_argbuf_d};
      3'd1:
        {srtarg_0_3_goMux_mux_onehot, srtarg_0_3_goMux_mux_mux} = {5'd2,
                                                                   contRet_0_3_1_argbuf_d};
      3'd2:
        {srtarg_0_3_goMux_mux_onehot, srtarg_0_3_goMux_mux_mux} = {5'd4,
                                                                   lizzieLet7_1_1_argbuf_d};
      3'd3:
        {srtarg_0_3_goMux_mux_onehot, srtarg_0_3_goMux_mux_mux} = {5'd8,
                                                                   lizzieLet8_1_1_argbuf_d};
      3'd4:
        {srtarg_0_3_goMux_mux_onehot, srtarg_0_3_goMux_mux_mux} = {5'd16,
                                                                   lizzieLet9_1_1_argbuf_d};
      default:
        {srtarg_0_3_goMux_mux_onehot, srtarg_0_3_goMux_mux_mux} = {5'd0,
                                                                   {16'd0, 1'd0}};
    endcase
  assign srtarg_0_3_goMux_mux_d = {srtarg_0_3_goMux_mux_mux[16:1],
                                   (srtarg_0_3_goMux_mux_mux[0] && go_21_goMux_choice_1_d[0])};
  assign go_21_goMux_choice_1_r = (srtarg_0_3_goMux_mux_d[0] && srtarg_0_3_goMux_mux_r);
  assign {lizzieLet9_1_1_argbuf_r,
          lizzieLet8_1_1_argbuf_r,
          lizzieLet7_1_1_argbuf_r,
          contRet_0_3_1_argbuf_r,
          lizzieLet6_1_1_argbuf_r} = (go_21_goMux_choice_1_r ? srtarg_0_3_goMux_mux_onehot :
                                      5'd0);
  
  /* mux (Ty C5,
     Ty Pointer_CTmap''_map''_Int_Int_Int) : (go_21_goMux_choice_2,C5) [(lizzieLet16_1_6QNone_Int_1_argbuf,Pointer_CTmap''_map''_Int_Int_Int),
                                                                        (sc_0_19_1_argbuf,Pointer_CTmap''_map''_Int_Int_Int),
                                                                        (es_0_5_2MyFalse_1_argbuf,Pointer_CTmap''_map''_Int_Int_Int),
                                                                        (es_0_5_2MyTrue_1_argbuf,Pointer_CTmap''_map''_Int_Int_Int),
                                                                        (lizzieLet16_1_6QError_Int_1_argbuf,Pointer_CTmap''_map''_Int_Int_Int)] > (scfarg_0_3_goMux_mux,Pointer_CTmap''_map''_Int_Int_Int) */
  logic [16:0] scfarg_0_3_goMux_mux_mux;
  logic [4:0] scfarg_0_3_goMux_mux_onehot;
  always_comb
    unique case (go_21_goMux_choice_2_d[3:1])
      3'd0:
        {scfarg_0_3_goMux_mux_onehot, scfarg_0_3_goMux_mux_mux} = {5'd1,
                                                                   lizzieLet16_1_6QNone_Int_1_argbuf_d};
      3'd1:
        {scfarg_0_3_goMux_mux_onehot, scfarg_0_3_goMux_mux_mux} = {5'd2,
                                                                   sc_0_19_1_argbuf_d};
      3'd2:
        {scfarg_0_3_goMux_mux_onehot, scfarg_0_3_goMux_mux_mux} = {5'd4,
                                                                   es_0_5_2MyFalse_1_argbuf_d};
      3'd3:
        {scfarg_0_3_goMux_mux_onehot, scfarg_0_3_goMux_mux_mux} = {5'd8,
                                                                   es_0_5_2MyTrue_1_argbuf_d};
      3'd4:
        {scfarg_0_3_goMux_mux_onehot, scfarg_0_3_goMux_mux_mux} = {5'd16,
                                                                   lizzieLet16_1_6QError_Int_1_argbuf_d};
      default:
        {scfarg_0_3_goMux_mux_onehot, scfarg_0_3_goMux_mux_mux} = {5'd0,
                                                                   {16'd0, 1'd0}};
    endcase
  assign scfarg_0_3_goMux_mux_d = {scfarg_0_3_goMux_mux_mux[16:1],
                                   (scfarg_0_3_goMux_mux_mux[0] && go_21_goMux_choice_2_d[0])};
  assign go_21_goMux_choice_2_r = (scfarg_0_3_goMux_mux_d[0] && scfarg_0_3_goMux_mux_r);
  assign {lizzieLet16_1_6QError_Int_1_argbuf_r,
          es_0_5_2MyTrue_1_argbuf_r,
          es_0_5_2MyFalse_1_argbuf_r,
          sc_0_19_1_argbuf_r,
          lizzieLet16_1_6QNone_Int_1_argbuf_r} = (go_21_goMux_choice_2_r ? scfarg_0_3_goMux_mux_onehot :
                                                  5'd0);
  
  /* dcon (Ty MyDTInt_Int,
      Dcon Dcon_main1) : [(go_7_1,Go)] > (go_7_1Dcon_main1,MyDTInt_Int) */
  assign go_7_1Dcon_main1_d = Dcon_main1_dc((& {go_7_1_d[0]}), go_7_1_d);
  assign {go_7_1_r} = {1 {(go_7_1Dcon_main1_r && go_7_1Dcon_main1_d[0])}};
  
  /* buf (Ty MyDTInt_Int) : (go_7_1Dcon_main1,MyDTInt_Int) > (es_2_1_argbuf,MyDTInt_Int) */
  MyDTInt_Int_t go_7_1Dcon_main1_bufchan_d;
  logic go_7_1Dcon_main1_bufchan_r;
  assign go_7_1Dcon_main1_r = ((! go_7_1Dcon_main1_bufchan_d[0]) || go_7_1Dcon_main1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_7_1Dcon_main1_bufchan_d <= 1'd0;
    else
      if (go_7_1Dcon_main1_r)
        go_7_1Dcon_main1_bufchan_d <= go_7_1Dcon_main1_d;
  MyDTInt_Int_t go_7_1Dcon_main1_bufchan_buf;
  assign go_7_1Dcon_main1_bufchan_r = (! go_7_1Dcon_main1_bufchan_buf[0]);
  assign es_2_1_argbuf_d = (go_7_1Dcon_main1_bufchan_buf[0] ? go_7_1Dcon_main1_bufchan_buf :
                            go_7_1Dcon_main1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_7_1Dcon_main1_bufchan_buf <= 1'd0;
    else
      if ((es_2_1_argbuf_r && go_7_1Dcon_main1_bufchan_buf[0]))
        go_7_1Dcon_main1_bufchan_buf <= 1'd0;
      else if (((! es_2_1_argbuf_r) && (! go_7_1Dcon_main1_bufchan_buf[0])))
        go_7_1Dcon_main1_bufchan_buf <= go_7_1Dcon_main1_bufchan_d;
  
  /* dcon (Ty MyDTInt_Bool,
      Dcon Dcon_eqZero) : [(go_7_2,Go)] > (go_7_2Dcon_eqZero,MyDTInt_Bool) */
  assign go_7_2Dcon_eqZero_d = Dcon_eqZero_dc((& {go_7_2_d[0]}), go_7_2_d);
  assign {go_7_2_r} = {1 {(go_7_2Dcon_eqZero_r && go_7_2Dcon_eqZero_d[0])}};
  
  /* buf (Ty MyDTInt_Bool) : (go_7_2Dcon_eqZero,MyDTInt_Bool) > (es_1_1_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t go_7_2Dcon_eqZero_bufchan_d;
  logic go_7_2Dcon_eqZero_bufchan_r;
  assign go_7_2Dcon_eqZero_r = ((! go_7_2Dcon_eqZero_bufchan_d[0]) || go_7_2Dcon_eqZero_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_7_2Dcon_eqZero_bufchan_d <= 1'd0;
    else
      if (go_7_2Dcon_eqZero_r)
        go_7_2Dcon_eqZero_bufchan_d <= go_7_2Dcon_eqZero_d;
  MyDTInt_Bool_t go_7_2Dcon_eqZero_bufchan_buf;
  assign go_7_2Dcon_eqZero_bufchan_r = (! go_7_2Dcon_eqZero_bufchan_buf[0]);
  assign es_1_1_argbuf_d = (go_7_2Dcon_eqZero_bufchan_buf[0] ? go_7_2Dcon_eqZero_bufchan_buf :
                            go_7_2Dcon_eqZero_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_7_2Dcon_eqZero_bufchan_buf <= 1'd0;
    else
      if ((es_1_1_argbuf_r && go_7_2Dcon_eqZero_bufchan_buf[0]))
        go_7_2Dcon_eqZero_bufchan_buf <= 1'd0;
      else if (((! es_1_1_argbuf_r) && (! go_7_2Dcon_eqZero_bufchan_buf[0])))
        go_7_2Dcon_eqZero_bufchan_buf <= go_7_2Dcon_eqZero_bufchan_d;
  
  /* dcon (Ty MyDTInt_Int_Int,
      Dcon Dcon_$fNumInt_$c*) : [(go_7_3,Go)] > (go_7_3Dcon_$fNumInt_$c*,MyDTInt_Int_Int) */
  assign \go_7_3Dcon_$fNumInt_$ctimes_d  = \Dcon_$fNumInt_$ctimes_dc ((& {go_7_3_d[0]}), go_7_3_d);
  assign {go_7_3_r} = {1 {(\go_7_3Dcon_$fNumInt_$ctimes_r  && \go_7_3Dcon_$fNumInt_$ctimes_d [0])}};
  
  /* buf (Ty MyDTInt_Int_Int) : (go_7_3Dcon_$fNumInt_$c*,MyDTInt_Int_Int) > (es_5_1_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t \go_7_3Dcon_$fNumInt_$ctimes_bufchan_d ;
  logic \go_7_3Dcon_$fNumInt_$ctimes_bufchan_r ;
  assign \go_7_3Dcon_$fNumInt_$ctimes_r  = ((! \go_7_3Dcon_$fNumInt_$ctimes_bufchan_d [0]) || \go_7_3Dcon_$fNumInt_$ctimes_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \go_7_3Dcon_$fNumInt_$ctimes_bufchan_d  <= 1'd0;
    else
      if (\go_7_3Dcon_$fNumInt_$ctimes_r )
        \go_7_3Dcon_$fNumInt_$ctimes_bufchan_d  <= \go_7_3Dcon_$fNumInt_$ctimes_d ;
  MyDTInt_Int_Int_t \go_7_3Dcon_$fNumInt_$ctimes_bufchan_buf ;
  assign \go_7_3Dcon_$fNumInt_$ctimes_bufchan_r  = (! \go_7_3Dcon_$fNumInt_$ctimes_bufchan_buf [0]);
  assign es_5_1_argbuf_d = (\go_7_3Dcon_$fNumInt_$ctimes_bufchan_buf [0] ? \go_7_3Dcon_$fNumInt_$ctimes_bufchan_buf  :
                            \go_7_3Dcon_$fNumInt_$ctimes_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \go_7_3Dcon_$fNumInt_$ctimes_bufchan_buf  <= 1'd0;
    else
      if ((es_5_1_argbuf_r && \go_7_3Dcon_$fNumInt_$ctimes_bufchan_buf [0]))
        \go_7_3Dcon_$fNumInt_$ctimes_bufchan_buf  <= 1'd0;
      else if (((! es_5_1_argbuf_r) && (! \go_7_3Dcon_$fNumInt_$ctimes_bufchan_buf [0])))
        \go_7_3Dcon_$fNumInt_$ctimes_bufchan_buf  <= \go_7_3Dcon_$fNumInt_$ctimes_bufchan_d ;
  
  /* dcon (Ty MyDTInt_Bool,
      Dcon Dcon_eqZero) : [(go_7_4,Go)] > (go_7_4Dcon_eqZero,MyDTInt_Bool) */
  assign go_7_4Dcon_eqZero_d = Dcon_eqZero_dc((& {go_7_4_d[0]}), go_7_4_d);
  assign {go_7_4_r} = {1 {(go_7_4Dcon_eqZero_r && go_7_4Dcon_eqZero_d[0])}};
  
  /* buf (Ty MyDTInt_Bool) : (go_7_4Dcon_eqZero,MyDTInt_Bool) > (es_4_1_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t go_7_4Dcon_eqZero_bufchan_d;
  logic go_7_4Dcon_eqZero_bufchan_r;
  assign go_7_4Dcon_eqZero_r = ((! go_7_4Dcon_eqZero_bufchan_d[0]) || go_7_4Dcon_eqZero_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_7_4Dcon_eqZero_bufchan_d <= 1'd0;
    else
      if (go_7_4Dcon_eqZero_r)
        go_7_4Dcon_eqZero_bufchan_d <= go_7_4Dcon_eqZero_d;
  MyDTInt_Bool_t go_7_4Dcon_eqZero_bufchan_buf;
  assign go_7_4Dcon_eqZero_bufchan_r = (! go_7_4Dcon_eqZero_bufchan_buf[0]);
  assign es_4_1_argbuf_d = (go_7_4Dcon_eqZero_bufchan_buf[0] ? go_7_4Dcon_eqZero_bufchan_buf :
                            go_7_4Dcon_eqZero_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_7_4Dcon_eqZero_bufchan_buf <= 1'd0;
    else
      if ((es_4_1_argbuf_r && go_7_4Dcon_eqZero_bufchan_buf[0]))
        go_7_4Dcon_eqZero_bufchan_buf <= 1'd0;
      else if (((! es_4_1_argbuf_r) && (! go_7_4Dcon_eqZero_bufchan_buf[0])))
        go_7_4Dcon_eqZero_bufchan_buf <= go_7_4Dcon_eqZero_bufchan_d;
  
  /* buf (Ty Go) : (go_7_5,Go) > (go_7_5_argbuf,Go) */
  Go_t go_7_5_bufchan_d;
  logic go_7_5_bufchan_r;
  assign go_7_5_r = ((! go_7_5_bufchan_d[0]) || go_7_5_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_7_5_bufchan_d <= 1'd0;
    else if (go_7_5_r) go_7_5_bufchan_d <= go_7_5_d;
  Go_t go_7_5_bufchan_buf;
  assign go_7_5_bufchan_r = (! go_7_5_bufchan_buf[0]);
  assign go_7_5_argbuf_d = (go_7_5_bufchan_buf[0] ? go_7_5_bufchan_buf :
                            go_7_5_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_7_5_bufchan_buf <= 1'd0;
    else
      if ((go_7_5_argbuf_r && go_7_5_bufchan_buf[0]))
        go_7_5_bufchan_buf <= 1'd0;
      else if (((! go_7_5_argbuf_r) && (! go_7_5_bufchan_buf[0])))
        go_7_5_bufchan_buf <= go_7_5_bufchan_d;
  
  /* dcon (Ty TupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int,
      Dcon TupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int) : [(go_7_5_argbuf,Go),
                                                                                              (es_4_1_argbuf,MyDTInt_Bool),
                                                                                              (es_5_1_argbuf,MyDTInt_Int_Int),
                                                                                              (wsvA_1_argbuf,Pointer_QTree_Int),
                                                                                              (w1svB_1_argbuf,Pointer_QTree_Int)] > (kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1,TupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int) */
  assign kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1_d = TupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_dc((& {go_7_5_argbuf_d[0],
                                                                                                                                                                                                         es_4_1_argbuf_d[0],
                                                                                                                                                                                                         es_5_1_argbuf_d[0],
                                                                                                                                                                                                         wsvA_1_argbuf_d[0],
                                                                                                                                                                                                         w1svB_1_argbuf_d[0]}), go_7_5_argbuf_d, es_4_1_argbuf_d, es_5_1_argbuf_d, wsvA_1_argbuf_d, w1svB_1_argbuf_d);
  assign {go_7_5_argbuf_r,
          es_4_1_argbuf_r,
          es_5_1_argbuf_r,
          wsvA_1_argbuf_r,
          w1svB_1_argbuf_r} = {5 {(kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1_r && kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1_d[0])}};
  
  /* buf (Ty Go) : (go_7_6,Go) > (go_7_6_argbuf,Go) */
  Go_t go_7_6_bufchan_d;
  logic go_7_6_bufchan_r;
  assign go_7_6_r = ((! go_7_6_bufchan_d[0]) || go_7_6_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_7_6_bufchan_d <= 1'd0;
    else if (go_7_6_r) go_7_6_bufchan_d <= go_7_6_d;
  Go_t go_7_6_bufchan_buf;
  assign go_7_6_bufchan_r = (! go_7_6_bufchan_buf[0]);
  assign go_7_6_argbuf_d = (go_7_6_bufchan_buf[0] ? go_7_6_bufchan_buf :
                            go_7_6_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_7_6_bufchan_buf <= 1'd0;
    else
      if ((go_7_6_argbuf_r && go_7_6_bufchan_buf[0]))
        go_7_6_bufchan_buf <= 1'd0;
      else if (((! go_7_6_argbuf_r) && (! go_7_6_bufchan_buf[0])))
        go_7_6_bufchan_buf <= go_7_6_bufchan_d;
  
  /* dcon (Ty TupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int,
      Dcon TupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int) : [(go_7_6_argbuf,Go),
                                                                      (es_1_1_argbuf,MyDTInt_Bool),
                                                                      (es_2_1_argbuf,MyDTInt_Int),
                                                                      (es_3_1_argbuf,Pointer_QTree_Int)] > (main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int_1,TupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int) */
  assign \main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int_1_d  = TupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int_dc((& {go_7_6_argbuf_d[0],
                                                                                                                                                       es_1_1_argbuf_d[0],
                                                                                                                                                       es_2_1_argbuf_d[0],
                                                                                                                                                       es_3_1_argbuf_d[0]}), go_7_6_argbuf_d, es_1_1_argbuf_d, es_2_1_argbuf_d, es_3_1_argbuf_d);
  assign {go_7_6_argbuf_r,
          es_1_1_argbuf_r,
          es_2_1_argbuf_r,
          es_3_1_argbuf_r} = {4 {(\main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int_1_r  && \main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int_1_d [0])}};
  
  /* buf (Ty Go) : (go_7_7,Go) > (go_7_7_argbuf,Go) */
  Go_t go_7_7_bufchan_d;
  logic go_7_7_bufchan_r;
  assign go_7_7_r = ((! go_7_7_bufchan_d[0]) || go_7_7_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_7_7_bufchan_d <= 1'd0;
    else if (go_7_7_r) go_7_7_bufchan_d <= go_7_7_d;
  Go_t go_7_7_bufchan_buf;
  assign go_7_7_bufchan_r = (! go_7_7_bufchan_buf[0]);
  assign go_7_7_argbuf_d = (go_7_7_bufchan_buf[0] ? go_7_7_bufchan_buf :
                            go_7_7_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_7_7_bufchan_buf <= 1'd0;
    else
      if ((go_7_7_argbuf_r && go_7_7_bufchan_buf[0]))
        go_7_7_bufchan_buf <= 1'd0;
      else if (((! go_7_7_argbuf_r) && (! go_7_7_bufchan_buf[0])))
        go_7_7_bufchan_buf <= go_7_7_bufchan_d;
  
  /* dcon (Ty TupGo___Pointer_QTree_Int,
      Dcon TupGo___Pointer_QTree_Int) : [(go_7_7_argbuf,Go),
                                         (es_0_1_1_argbuf,Pointer_QTree_Int)] > ($wnnz_IntTupGo___Pointer_QTree_Int_1,TupGo___Pointer_QTree_Int) */
  assign \$wnnz_IntTupGo___Pointer_QTree_Int_1_d  = TupGo___Pointer_QTree_Int_dc((& {go_7_7_argbuf_d[0],
                                                                                     es_0_1_1_argbuf_d[0]}), go_7_7_argbuf_d, es_0_1_1_argbuf_d);
  assign {go_7_7_argbuf_r,
          es_0_1_1_argbuf_r} = {2 {(\$wnnz_IntTupGo___Pointer_QTree_Int_1_r  && \$wnnz_IntTupGo___Pointer_QTree_Int_1_d [0])}};
  
  /* dcon (Ty CT$wnnz_Int,
      Dcon L$wnnz_Intsbos) : [(go_8_1,Go)] > (go_8_1L$wnnz_Intsbos,CT$wnnz_Int) */
  assign go_8_1L$wnnz_Intsbos_d = L$wnnz_Intsbos_dc((& {go_8_1_d[0]}), go_8_1_d);
  assign {go_8_1_r} = {1 {(go_8_1L$wnnz_Intsbos_r && go_8_1L$wnnz_Intsbos_d[0])}};
  
  /* buf (Ty CT$wnnz_Int) : (go_8_1L$wnnz_Intsbos,CT$wnnz_Int) > (lizzieLet0_1_argbuf,CT$wnnz_Int) */
  CT$wnnz_Int_t go_8_1L$wnnz_Intsbos_bufchan_d;
  logic go_8_1L$wnnz_Intsbos_bufchan_r;
  assign go_8_1L$wnnz_Intsbos_r = ((! go_8_1L$wnnz_Intsbos_bufchan_d[0]) || go_8_1L$wnnz_Intsbos_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      go_8_1L$wnnz_Intsbos_bufchan_d <= {115'd0, 1'd0};
    else
      if (go_8_1L$wnnz_Intsbos_r)
        go_8_1L$wnnz_Intsbos_bufchan_d <= go_8_1L$wnnz_Intsbos_d;
  CT$wnnz_Int_t go_8_1L$wnnz_Intsbos_bufchan_buf;
  assign go_8_1L$wnnz_Intsbos_bufchan_r = (! go_8_1L$wnnz_Intsbos_bufchan_buf[0]);
  assign lizzieLet0_1_argbuf_d = (go_8_1L$wnnz_Intsbos_bufchan_buf[0] ? go_8_1L$wnnz_Intsbos_bufchan_buf :
                                  go_8_1L$wnnz_Intsbos_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      go_8_1L$wnnz_Intsbos_bufchan_buf <= {115'd0, 1'd0};
    else
      if ((lizzieLet0_1_argbuf_r && go_8_1L$wnnz_Intsbos_bufchan_buf[0]))
        go_8_1L$wnnz_Intsbos_bufchan_buf <= {115'd0, 1'd0};
      else if (((! lizzieLet0_1_argbuf_r) && (! go_8_1L$wnnz_Intsbos_bufchan_buf[0])))
        go_8_1L$wnnz_Intsbos_bufchan_buf <= go_8_1L$wnnz_Intsbos_bufchan_d;
  
  /* buf (Ty Go) : (go_8_2,Go) > (go_8_2_argbuf,Go) */
  Go_t go_8_2_bufchan_d;
  logic go_8_2_bufchan_r;
  assign go_8_2_r = ((! go_8_2_bufchan_d[0]) || go_8_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_8_2_bufchan_d <= 1'd0;
    else if (go_8_2_r) go_8_2_bufchan_d <= go_8_2_d;
  Go_t go_8_2_bufchan_buf;
  assign go_8_2_bufchan_r = (! go_8_2_bufchan_buf[0]);
  assign go_8_2_argbuf_d = (go_8_2_bufchan_buf[0] ? go_8_2_bufchan_buf :
                            go_8_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_8_2_bufchan_buf <= 1'd0;
    else
      if ((go_8_2_argbuf_r && go_8_2_bufchan_buf[0]))
        go_8_2_bufchan_buf <= 1'd0;
      else if (((! go_8_2_argbuf_r) && (! go_8_2_bufchan_buf[0])))
        go_8_2_bufchan_buf <= go_8_2_bufchan_d;
  
  /* dcon (Ty TupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int,
      Dcon TupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int) : [(go_8_2_argbuf,Go),
                                                               (wsvt_1_argbuf,Pointer_QTree_Int),
                                                               (lizzieLet17_1_argbuf,Pointer_CT$wnnz_Int)] > (call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1,TupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int) */
  assign call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_d = TupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_dc((& {go_8_2_argbuf_d[0],
                                                                                                                                    wsvt_1_argbuf_d[0],
                                                                                                                                    lizzieLet17_1_argbuf_d[0]}), go_8_2_argbuf_d, wsvt_1_argbuf_d, lizzieLet17_1_argbuf_d);
  assign {go_8_2_argbuf_r,
          wsvt_1_argbuf_r,
          lizzieLet17_1_argbuf_r} = {3 {(call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_r && call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_d[0])}};
  
  /* buf (Ty MyDTInt_Bool) : (isZacL_2_2,MyDTInt_Bool) > (isZacL_2_2_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t isZacL_2_2_bufchan_d;
  logic isZacL_2_2_bufchan_r;
  assign isZacL_2_2_r = ((! isZacL_2_2_bufchan_d[0]) || isZacL_2_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) isZacL_2_2_bufchan_d <= 1'd0;
    else if (isZacL_2_2_r) isZacL_2_2_bufchan_d <= isZacL_2_2_d;
  MyDTInt_Bool_t isZacL_2_2_bufchan_buf;
  assign isZacL_2_2_bufchan_r = (! isZacL_2_2_bufchan_buf[0]);
  assign isZacL_2_2_argbuf_d = (isZacL_2_2_bufchan_buf[0] ? isZacL_2_2_bufchan_buf :
                                isZacL_2_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) isZacL_2_2_bufchan_buf <= 1'd0;
    else
      if ((isZacL_2_2_argbuf_r && isZacL_2_2_bufchan_buf[0]))
        isZacL_2_2_bufchan_buf <= 1'd0;
      else if (((! isZacL_2_2_argbuf_r) && (! isZacL_2_2_bufchan_buf[0])))
        isZacL_2_2_bufchan_buf <= isZacL_2_2_bufchan_d;
  
  /* fork (Ty MyDTInt_Bool) : (isZacL_2_destruct,MyDTInt_Bool) > [(isZacL_2_1,MyDTInt_Bool),
                                                             (isZacL_2_2,MyDTInt_Bool)] */
  logic [1:0] isZacL_2_destruct_emitted;
  logic [1:0] isZacL_2_destruct_done;
  assign isZacL_2_1_d = (isZacL_2_destruct_d[0] && (! isZacL_2_destruct_emitted[0]));
  assign isZacL_2_2_d = (isZacL_2_destruct_d[0] && (! isZacL_2_destruct_emitted[1]));
  assign isZacL_2_destruct_done = (isZacL_2_destruct_emitted | ({isZacL_2_2_d[0],
                                                                 isZacL_2_1_d[0]} & {isZacL_2_2_r,
                                                                                     isZacL_2_1_r}));
  assign isZacL_2_destruct_r = (& isZacL_2_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) isZacL_2_destruct_emitted <= 2'd0;
    else
      isZacL_2_destruct_emitted <= (isZacL_2_destruct_r ? 2'd0 :
                                    isZacL_2_destruct_done);
  
  /* buf (Ty MyDTInt_Bool) : (isZacL_3_2,MyDTInt_Bool) > (isZacL_3_2_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t isZacL_3_2_bufchan_d;
  logic isZacL_3_2_bufchan_r;
  assign isZacL_3_2_r = ((! isZacL_3_2_bufchan_d[0]) || isZacL_3_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) isZacL_3_2_bufchan_d <= 1'd0;
    else if (isZacL_3_2_r) isZacL_3_2_bufchan_d <= isZacL_3_2_d;
  MyDTInt_Bool_t isZacL_3_2_bufchan_buf;
  assign isZacL_3_2_bufchan_r = (! isZacL_3_2_bufchan_buf[0]);
  assign isZacL_3_2_argbuf_d = (isZacL_3_2_bufchan_buf[0] ? isZacL_3_2_bufchan_buf :
                                isZacL_3_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) isZacL_3_2_bufchan_buf <= 1'd0;
    else
      if ((isZacL_3_2_argbuf_r && isZacL_3_2_bufchan_buf[0]))
        isZacL_3_2_bufchan_buf <= 1'd0;
      else if (((! isZacL_3_2_argbuf_r) && (! isZacL_3_2_bufchan_buf[0])))
        isZacL_3_2_bufchan_buf <= isZacL_3_2_bufchan_d;
  
  /* fork (Ty MyDTInt_Bool) : (isZacL_3_destruct,MyDTInt_Bool) > [(isZacL_3_1,MyDTInt_Bool),
                                                             (isZacL_3_2,MyDTInt_Bool)] */
  logic [1:0] isZacL_3_destruct_emitted;
  logic [1:0] isZacL_3_destruct_done;
  assign isZacL_3_1_d = (isZacL_3_destruct_d[0] && (! isZacL_3_destruct_emitted[0]));
  assign isZacL_3_2_d = (isZacL_3_destruct_d[0] && (! isZacL_3_destruct_emitted[1]));
  assign isZacL_3_destruct_done = (isZacL_3_destruct_emitted | ({isZacL_3_2_d[0],
                                                                 isZacL_3_1_d[0]} & {isZacL_3_2_r,
                                                                                     isZacL_3_1_r}));
  assign isZacL_3_destruct_r = (& isZacL_3_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) isZacL_3_destruct_emitted <= 2'd0;
    else
      isZacL_3_destruct_emitted <= (isZacL_3_destruct_r ? 2'd0 :
                                    isZacL_3_destruct_done);
  
  /* buf (Ty MyDTInt_Bool) : (isZacL_4_destruct,MyDTInt_Bool) > (isZacL_4_1_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t isZacL_4_destruct_bufchan_d;
  logic isZacL_4_destruct_bufchan_r;
  assign isZacL_4_destruct_r = ((! isZacL_4_destruct_bufchan_d[0]) || isZacL_4_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) isZacL_4_destruct_bufchan_d <= 1'd0;
    else
      if (isZacL_4_destruct_r)
        isZacL_4_destruct_bufchan_d <= isZacL_4_destruct_d;
  MyDTInt_Bool_t isZacL_4_destruct_bufchan_buf;
  assign isZacL_4_destruct_bufchan_r = (! isZacL_4_destruct_bufchan_buf[0]);
  assign isZacL_4_1_argbuf_d = (isZacL_4_destruct_bufchan_buf[0] ? isZacL_4_destruct_bufchan_buf :
                                isZacL_4_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) isZacL_4_destruct_bufchan_buf <= 1'd0;
    else
      if ((isZacL_4_1_argbuf_r && isZacL_4_destruct_bufchan_buf[0]))
        isZacL_4_destruct_bufchan_buf <= 1'd0;
      else if (((! isZacL_4_1_argbuf_r) && (! isZacL_4_destruct_bufchan_buf[0])))
        isZacL_4_destruct_bufchan_buf <= isZacL_4_destruct_bufchan_d;
  
  /* buf (Ty MyDTInt_Bool) : (isZacT_2_2,MyDTInt_Bool) > (isZacT_2_2_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t isZacT_2_2_bufchan_d;
  logic isZacT_2_2_bufchan_r;
  assign isZacT_2_2_r = ((! isZacT_2_2_bufchan_d[0]) || isZacT_2_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) isZacT_2_2_bufchan_d <= 1'd0;
    else if (isZacT_2_2_r) isZacT_2_2_bufchan_d <= isZacT_2_2_d;
  MyDTInt_Bool_t isZacT_2_2_bufchan_buf;
  assign isZacT_2_2_bufchan_r = (! isZacT_2_2_bufchan_buf[0]);
  assign isZacT_2_2_argbuf_d = (isZacT_2_2_bufchan_buf[0] ? isZacT_2_2_bufchan_buf :
                                isZacT_2_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) isZacT_2_2_bufchan_buf <= 1'd0;
    else
      if ((isZacT_2_2_argbuf_r && isZacT_2_2_bufchan_buf[0]))
        isZacT_2_2_bufchan_buf <= 1'd0;
      else if (((! isZacT_2_2_argbuf_r) && (! isZacT_2_2_bufchan_buf[0])))
        isZacT_2_2_bufchan_buf <= isZacT_2_2_bufchan_d;
  
  /* fork (Ty MyDTInt_Bool) : (isZacT_2_destruct,MyDTInt_Bool) > [(isZacT_2_1,MyDTInt_Bool),
                                                             (isZacT_2_2,MyDTInt_Bool)] */
  logic [1:0] isZacT_2_destruct_emitted;
  logic [1:0] isZacT_2_destruct_done;
  assign isZacT_2_1_d = (isZacT_2_destruct_d[0] && (! isZacT_2_destruct_emitted[0]));
  assign isZacT_2_2_d = (isZacT_2_destruct_d[0] && (! isZacT_2_destruct_emitted[1]));
  assign isZacT_2_destruct_done = (isZacT_2_destruct_emitted | ({isZacT_2_2_d[0],
                                                                 isZacT_2_1_d[0]} & {isZacT_2_2_r,
                                                                                     isZacT_2_1_r}));
  assign isZacT_2_destruct_r = (& isZacT_2_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) isZacT_2_destruct_emitted <= 2'd0;
    else
      isZacT_2_destruct_emitted <= (isZacT_2_destruct_r ? 2'd0 :
                                    isZacT_2_destruct_done);
  
  /* buf (Ty MyDTInt_Bool) : (isZacT_3_2,MyDTInt_Bool) > (isZacT_3_2_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t isZacT_3_2_bufchan_d;
  logic isZacT_3_2_bufchan_r;
  assign isZacT_3_2_r = ((! isZacT_3_2_bufchan_d[0]) || isZacT_3_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) isZacT_3_2_bufchan_d <= 1'd0;
    else if (isZacT_3_2_r) isZacT_3_2_bufchan_d <= isZacT_3_2_d;
  MyDTInt_Bool_t isZacT_3_2_bufchan_buf;
  assign isZacT_3_2_bufchan_r = (! isZacT_3_2_bufchan_buf[0]);
  assign isZacT_3_2_argbuf_d = (isZacT_3_2_bufchan_buf[0] ? isZacT_3_2_bufchan_buf :
                                isZacT_3_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) isZacT_3_2_bufchan_buf <= 1'd0;
    else
      if ((isZacT_3_2_argbuf_r && isZacT_3_2_bufchan_buf[0]))
        isZacT_3_2_bufchan_buf <= 1'd0;
      else if (((! isZacT_3_2_argbuf_r) && (! isZacT_3_2_bufchan_buf[0])))
        isZacT_3_2_bufchan_buf <= isZacT_3_2_bufchan_d;
  
  /* fork (Ty MyDTInt_Bool) : (isZacT_3_destruct,MyDTInt_Bool) > [(isZacT_3_1,MyDTInt_Bool),
                                                             (isZacT_3_2,MyDTInt_Bool)] */
  logic [1:0] isZacT_3_destruct_emitted;
  logic [1:0] isZacT_3_destruct_done;
  assign isZacT_3_1_d = (isZacT_3_destruct_d[0] && (! isZacT_3_destruct_emitted[0]));
  assign isZacT_3_2_d = (isZacT_3_destruct_d[0] && (! isZacT_3_destruct_emitted[1]));
  assign isZacT_3_destruct_done = (isZacT_3_destruct_emitted | ({isZacT_3_2_d[0],
                                                                 isZacT_3_1_d[0]} & {isZacT_3_2_r,
                                                                                     isZacT_3_1_r}));
  assign isZacT_3_destruct_r = (& isZacT_3_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) isZacT_3_destruct_emitted <= 2'd0;
    else
      isZacT_3_destruct_emitted <= (isZacT_3_destruct_r ? 2'd0 :
                                    isZacT_3_destruct_done);
  
  /* buf (Ty MyDTInt_Bool) : (isZacT_4_destruct,MyDTInt_Bool) > (isZacT_4_1_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t isZacT_4_destruct_bufchan_d;
  logic isZacT_4_destruct_bufchan_r;
  assign isZacT_4_destruct_r = ((! isZacT_4_destruct_bufchan_d[0]) || isZacT_4_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) isZacT_4_destruct_bufchan_d <= 1'd0;
    else
      if (isZacT_4_destruct_r)
        isZacT_4_destruct_bufchan_d <= isZacT_4_destruct_d;
  MyDTInt_Bool_t isZacT_4_destruct_bufchan_buf;
  assign isZacT_4_destruct_bufchan_r = (! isZacT_4_destruct_bufchan_buf[0]);
  assign isZacT_4_1_argbuf_d = (isZacT_4_destruct_bufchan_buf[0] ? isZacT_4_destruct_bufchan_buf :
                                isZacT_4_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) isZacT_4_destruct_bufchan_buf <= 1'd0;
    else
      if ((isZacT_4_1_argbuf_r && isZacT_4_destruct_bufchan_buf[0]))
        isZacT_4_destruct_bufchan_buf <= 1'd0;
      else if (((! isZacT_4_1_argbuf_r) && (! isZacT_4_destruct_bufchan_buf[0])))
        isZacT_4_destruct_bufchan_buf <= isZacT_4_destruct_bufchan_d;
  
  /* buf (Ty MyDTInt_Bool) : (isZad2_2_2,MyDTInt_Bool) > (isZad2_2_2_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t isZad2_2_2_bufchan_d;
  logic isZad2_2_2_bufchan_r;
  assign isZad2_2_2_r = ((! isZad2_2_2_bufchan_d[0]) || isZad2_2_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) isZad2_2_2_bufchan_d <= 1'd0;
    else if (isZad2_2_2_r) isZad2_2_2_bufchan_d <= isZad2_2_2_d;
  MyDTInt_Bool_t isZad2_2_2_bufchan_buf;
  assign isZad2_2_2_bufchan_r = (! isZad2_2_2_bufchan_buf[0]);
  assign isZad2_2_2_argbuf_d = (isZad2_2_2_bufchan_buf[0] ? isZad2_2_2_bufchan_buf :
                                isZad2_2_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) isZad2_2_2_bufchan_buf <= 1'd0;
    else
      if ((isZad2_2_2_argbuf_r && isZad2_2_2_bufchan_buf[0]))
        isZad2_2_2_bufchan_buf <= 1'd0;
      else if (((! isZad2_2_2_argbuf_r) && (! isZad2_2_2_bufchan_buf[0])))
        isZad2_2_2_bufchan_buf <= isZad2_2_2_bufchan_d;
  
  /* fork (Ty MyDTInt_Bool) : (isZad2_2_destruct,MyDTInt_Bool) > [(isZad2_2_1,MyDTInt_Bool),
                                                             (isZad2_2_2,MyDTInt_Bool)] */
  logic [1:0] isZad2_2_destruct_emitted;
  logic [1:0] isZad2_2_destruct_done;
  assign isZad2_2_1_d = (isZad2_2_destruct_d[0] && (! isZad2_2_destruct_emitted[0]));
  assign isZad2_2_2_d = (isZad2_2_destruct_d[0] && (! isZad2_2_destruct_emitted[1]));
  assign isZad2_2_destruct_done = (isZad2_2_destruct_emitted | ({isZad2_2_2_d[0],
                                                                 isZad2_2_1_d[0]} & {isZad2_2_2_r,
                                                                                     isZad2_2_1_r}));
  assign isZad2_2_destruct_r = (& isZad2_2_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) isZad2_2_destruct_emitted <= 2'd0;
    else
      isZad2_2_destruct_emitted <= (isZad2_2_destruct_r ? 2'd0 :
                                    isZad2_2_destruct_done);
  
  /* buf (Ty MyDTInt_Bool) : (isZad2_3_2,MyDTInt_Bool) > (isZad2_3_2_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t isZad2_3_2_bufchan_d;
  logic isZad2_3_2_bufchan_r;
  assign isZad2_3_2_r = ((! isZad2_3_2_bufchan_d[0]) || isZad2_3_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) isZad2_3_2_bufchan_d <= 1'd0;
    else if (isZad2_3_2_r) isZad2_3_2_bufchan_d <= isZad2_3_2_d;
  MyDTInt_Bool_t isZad2_3_2_bufchan_buf;
  assign isZad2_3_2_bufchan_r = (! isZad2_3_2_bufchan_buf[0]);
  assign isZad2_3_2_argbuf_d = (isZad2_3_2_bufchan_buf[0] ? isZad2_3_2_bufchan_buf :
                                isZad2_3_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) isZad2_3_2_bufchan_buf <= 1'd0;
    else
      if ((isZad2_3_2_argbuf_r && isZad2_3_2_bufchan_buf[0]))
        isZad2_3_2_bufchan_buf <= 1'd0;
      else if (((! isZad2_3_2_argbuf_r) && (! isZad2_3_2_bufchan_buf[0])))
        isZad2_3_2_bufchan_buf <= isZad2_3_2_bufchan_d;
  
  /* fork (Ty MyDTInt_Bool) : (isZad2_3_destruct,MyDTInt_Bool) > [(isZad2_3_1,MyDTInt_Bool),
                                                             (isZad2_3_2,MyDTInt_Bool)] */
  logic [1:0] isZad2_3_destruct_emitted;
  logic [1:0] isZad2_3_destruct_done;
  assign isZad2_3_1_d = (isZad2_3_destruct_d[0] && (! isZad2_3_destruct_emitted[0]));
  assign isZad2_3_2_d = (isZad2_3_destruct_d[0] && (! isZad2_3_destruct_emitted[1]));
  assign isZad2_3_destruct_done = (isZad2_3_destruct_emitted | ({isZad2_3_2_d[0],
                                                                 isZad2_3_1_d[0]} & {isZad2_3_2_r,
                                                                                     isZad2_3_1_r}));
  assign isZad2_3_destruct_r = (& isZad2_3_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) isZad2_3_destruct_emitted <= 2'd0;
    else
      isZad2_3_destruct_emitted <= (isZad2_3_destruct_r ? 2'd0 :
                                    isZad2_3_destruct_done);
  
  /* buf (Ty MyDTInt_Bool) : (isZad2_4_destruct,MyDTInt_Bool) > (isZad2_4_1_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t isZad2_4_destruct_bufchan_d;
  logic isZad2_4_destruct_bufchan_r;
  assign isZad2_4_destruct_r = ((! isZad2_4_destruct_bufchan_d[0]) || isZad2_4_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) isZad2_4_destruct_bufchan_d <= 1'd0;
    else
      if (isZad2_4_destruct_r)
        isZad2_4_destruct_bufchan_d <= isZad2_4_destruct_d;
  MyDTInt_Bool_t isZad2_4_destruct_bufchan_buf;
  assign isZad2_4_destruct_bufchan_r = (! isZad2_4_destruct_bufchan_buf[0]);
  assign isZad2_4_1_argbuf_d = (isZad2_4_destruct_bufchan_buf[0] ? isZad2_4_destruct_bufchan_buf :
                                isZad2_4_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) isZad2_4_destruct_bufchan_buf <= 1'd0;
    else
      if ((isZad2_4_1_argbuf_r && isZad2_4_destruct_bufchan_buf[0]))
        isZad2_4_destruct_bufchan_buf <= 1'd0;
      else if (((! isZad2_4_1_argbuf_r) && (! isZad2_4_destruct_bufchan_buf[0])))
        isZad2_4_destruct_bufchan_buf <= isZad2_4_destruct_bufchan_d;
  
  /* destruct (Ty TupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int,
          Dcon TupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int) : (kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1,TupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int) > [(kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgo_15,Go),
                                                                                                                                                                                                                                                                                           (kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntisZad2_1,MyDTInt_Bool),
                                                                                                                                                                                                                                                                                           (kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgad3_1,MyDTInt_Int_Int),
                                                                                                                                                                                                                                                                                           (kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm1ad4_1,Pointer_QTree_Int),
                                                                                                                                                                                                                                                                                           (kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm2ad5_1,Pointer_QTree_Int)] */
  logic [4:0] kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1_emitted;
  logic [4:0] kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1_done;
  assign kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgo_15_d = (kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1_d[0] && (! kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1_emitted[0]));
  assign kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntisZad2_1_d = (kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1_d[0] && (! kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1_emitted[1]));
  assign kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgad3_1_d = (kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1_d[0] && (! kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1_emitted[2]));
  assign kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm1ad4_1_d = {kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1_d[16:1],
                                                                                                                         (kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1_d[0] && (! kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1_emitted[3]))};
  assign kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm2ad5_1_d = {kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1_d[32:17],
                                                                                                                         (kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1_d[0] && (! kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1_emitted[4]))};
  assign kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1_done = (kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1_emitted | ({kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm2ad5_1_d[0],
                                                                                                                                                                                                                                         kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm1ad4_1_d[0],
                                                                                                                                                                                                                                         kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgad3_1_d[0],
                                                                                                                                                                                                                                         kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntisZad2_1_d[0],
                                                                                                                                                                                                                                         kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgo_15_d[0]} & {kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm2ad5_1_r,
                                                                                                                                                                                                                                                                                                                                                           kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm1ad4_1_r,
                                                                                                                                                                                                                                                                                                                                                           kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgad3_1_r,
                                                                                                                                                                                                                                                                                                                                                           kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntisZad2_1_r,
                                                                                                                                                                                                                                                                                                                                                           kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgo_15_r}));
  assign kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1_r = (& kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1_emitted <= 5'd0;
    else
      kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1_emitted <= (kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1_r ? 5'd0 :
                                                                                                                        kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1_done);
  
  /* buf (Ty MyDTInt_Int_Int) : (kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgad3_1,MyDTInt_Int_Int) > (gad3_1_1_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgad3_1_bufchan_d;
  logic kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgad3_1_bufchan_r;
  assign kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgad3_1_r = ((! kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgad3_1_bufchan_d[0]) || kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgad3_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgad3_1_bufchan_d <= 1'd0;
    else
      if (kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgad3_1_r)
        kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgad3_1_bufchan_d <= kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgad3_1_d;
  MyDTInt_Int_Int_t kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgad3_1_bufchan_buf;
  assign kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgad3_1_bufchan_r = (! kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgad3_1_bufchan_buf[0]);
  assign gad3_1_1_argbuf_d = (kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgad3_1_bufchan_buf[0] ? kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgad3_1_bufchan_buf :
                              kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgad3_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgad3_1_bufchan_buf <= 1'd0;
    else
      if ((gad3_1_1_argbuf_r && kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgad3_1_bufchan_buf[0]))
        kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgad3_1_bufchan_buf <= 1'd0;
      else if (((! gad3_1_1_argbuf_r) && (! kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgad3_1_bufchan_buf[0])))
        kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgad3_1_bufchan_buf <= kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgad3_1_bufchan_d;
  
  /* fork (Ty Go) : (kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgo_15,Go) > [(go_15_1,Go),
                                                                                                                                (go_15_2,Go)] */
  logic [1:0] kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgo_15_emitted;
  logic [1:0] kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgo_15_done;
  assign go_15_1_d = (kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgo_15_d[0] && (! kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgo_15_emitted[0]));
  assign go_15_2_d = (kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgo_15_d[0] && (! kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgo_15_emitted[1]));
  assign kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgo_15_done = (kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgo_15_emitted | ({go_15_2_d[0],
                                                                                                                                                                                                                                               go_15_1_d[0]} & {go_15_2_r,
                                                                                                                                                                                                                                                                go_15_1_r}));
  assign kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgo_15_r = (& kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgo_15_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgo_15_emitted <= 2'd0;
    else
      kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgo_15_emitted <= (kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgo_15_r ? 2'd0 :
                                                                                                                           kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgo_15_done);
  
  /* buf (Ty MyDTInt_Bool) : (kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntisZad2_1,MyDTInt_Bool) > (isZad2_1_1_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntisZad2_1_bufchan_d;
  logic kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntisZad2_1_bufchan_r;
  assign kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntisZad2_1_r = ((! kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntisZad2_1_bufchan_d[0]) || kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntisZad2_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntisZad2_1_bufchan_d <= 1'd0;
    else
      if (kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntisZad2_1_r)
        kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntisZad2_1_bufchan_d <= kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntisZad2_1_d;
  MyDTInt_Bool_t kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntisZad2_1_bufchan_buf;
  assign kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntisZad2_1_bufchan_r = (! kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntisZad2_1_bufchan_buf[0]);
  assign isZad2_1_1_argbuf_d = (kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntisZad2_1_bufchan_buf[0] ? kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntisZad2_1_bufchan_buf :
                                kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntisZad2_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntisZad2_1_bufchan_buf <= 1'd0;
    else
      if ((isZad2_1_1_argbuf_r && kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntisZad2_1_bufchan_buf[0]))
        kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntisZad2_1_bufchan_buf <= 1'd0;
      else if (((! isZad2_1_1_argbuf_r) && (! kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntisZad2_1_bufchan_buf[0])))
        kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntisZad2_1_bufchan_buf <= kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntisZad2_1_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm1ad4_1,Pointer_QTree_Int) > (m1ad4_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm1ad4_1_bufchan_d;
  logic kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm1ad4_1_bufchan_r;
  assign kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm1ad4_1_r = ((! kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm1ad4_1_bufchan_d[0]) || kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm1ad4_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm1ad4_1_bufchan_d <= {16'd0,
                                                                                                                               1'd0};
    else
      if (kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm1ad4_1_r)
        kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm1ad4_1_bufchan_d <= kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm1ad4_1_d;
  Pointer_QTree_Int_t kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm1ad4_1_bufchan_buf;
  assign kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm1ad4_1_bufchan_r = (! kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm1ad4_1_bufchan_buf[0]);
  assign m1ad4_1_1_argbuf_d = (kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm1ad4_1_bufchan_buf[0] ? kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm1ad4_1_bufchan_buf :
                               kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm1ad4_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm1ad4_1_bufchan_buf <= {16'd0,
                                                                                                                                 1'd0};
    else
      if ((m1ad4_1_1_argbuf_r && kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm1ad4_1_bufchan_buf[0]))
        kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm1ad4_1_bufchan_buf <= {16'd0,
                                                                                                                                   1'd0};
      else if (((! m1ad4_1_1_argbuf_r) && (! kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm1ad4_1_bufchan_buf[0])))
        kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm1ad4_1_bufchan_buf <= kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm1ad4_1_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm2ad5_1,Pointer_QTree_Int) > (m2ad5_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm2ad5_1_bufchan_d;
  logic kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm2ad5_1_bufchan_r;
  assign kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm2ad5_1_r = ((! kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm2ad5_1_bufchan_d[0]) || kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm2ad5_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm2ad5_1_bufchan_d <= {16'd0,
                                                                                                                               1'd0};
    else
      if (kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm2ad5_1_r)
        kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm2ad5_1_bufchan_d <= kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm2ad5_1_d;
  Pointer_QTree_Int_t kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm2ad5_1_bufchan_buf;
  assign kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm2ad5_1_bufchan_r = (! kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm2ad5_1_bufchan_buf[0]);
  assign m2ad5_1_1_argbuf_d = (kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm2ad5_1_bufchan_buf[0] ? kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm2ad5_1_bufchan_buf :
                               kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm2ad5_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm2ad5_1_bufchan_buf <= {16'd0,
                                                                                                                                 1'd0};
    else
      if ((m2ad5_1_1_argbuf_r && kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm2ad5_1_bufchan_buf[0]))
        kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm2ad5_1_bufchan_buf <= {16'd0,
                                                                                                                                   1'd0};
      else if (((! m2ad5_1_1_argbuf_r) && (! kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm2ad5_1_bufchan_buf[0])))
        kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm2ad5_1_bufchan_buf <= kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm2ad5_1_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (kron_kron_Int_Int_Int_resbuf,Pointer_QTree_Int) > (es_3_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t kron_kron_Int_Int_Int_resbuf_bufchan_d;
  logic kron_kron_Int_Int_Int_resbuf_bufchan_r;
  assign kron_kron_Int_Int_Int_resbuf_r = ((! kron_kron_Int_Int_Int_resbuf_bufchan_d[0]) || kron_kron_Int_Int_Int_resbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      kron_kron_Int_Int_Int_resbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (kron_kron_Int_Int_Int_resbuf_r)
        kron_kron_Int_Int_Int_resbuf_bufchan_d <= kron_kron_Int_Int_Int_resbuf_d;
  Pointer_QTree_Int_t kron_kron_Int_Int_Int_resbuf_bufchan_buf;
  assign kron_kron_Int_Int_Int_resbuf_bufchan_r = (! kron_kron_Int_Int_Int_resbuf_bufchan_buf[0]);
  assign es_3_1_argbuf_d = (kron_kron_Int_Int_Int_resbuf_bufchan_buf[0] ? kron_kron_Int_Int_Int_resbuf_bufchan_buf :
                            kron_kron_Int_Int_Int_resbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      kron_kron_Int_Int_Int_resbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((es_3_1_argbuf_r && kron_kron_Int_Int_Int_resbuf_bufchan_buf[0]))
        kron_kron_Int_Int_Int_resbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! es_3_1_argbuf_r) && (! kron_kron_Int_Int_Int_resbuf_bufchan_buf[0])))
        kron_kron_Int_Int_Int_resbuf_bufchan_buf <= kron_kron_Int_Int_Int_resbuf_bufchan_d;
  
  /* destruct (Ty QTree_Int,
          Dcon QNode_Int) : (lizzieLet10_1QNode_Int,QTree_Int) > [(q1acP_destruct,Pointer_QTree_Int),
                                                                  (q2acQ_destruct,Pointer_QTree_Int),
                                                                  (q3acR_destruct,Pointer_QTree_Int),
                                                                  (q4acS_destruct,Pointer_QTree_Int)] */
  logic [3:0] lizzieLet10_1QNode_Int_emitted;
  logic [3:0] lizzieLet10_1QNode_Int_done;
  assign q1acP_destruct_d = {lizzieLet10_1QNode_Int_d[18:3],
                             (lizzieLet10_1QNode_Int_d[0] && (! lizzieLet10_1QNode_Int_emitted[0]))};
  assign q2acQ_destruct_d = {lizzieLet10_1QNode_Int_d[34:19],
                             (lizzieLet10_1QNode_Int_d[0] && (! lizzieLet10_1QNode_Int_emitted[1]))};
  assign q3acR_destruct_d = {lizzieLet10_1QNode_Int_d[50:35],
                             (lizzieLet10_1QNode_Int_d[0] && (! lizzieLet10_1QNode_Int_emitted[2]))};
  assign q4acS_destruct_d = {lizzieLet10_1QNode_Int_d[66:51],
                             (lizzieLet10_1QNode_Int_d[0] && (! lizzieLet10_1QNode_Int_emitted[3]))};
  assign lizzieLet10_1QNode_Int_done = (lizzieLet10_1QNode_Int_emitted | ({q4acS_destruct_d[0],
                                                                           q3acR_destruct_d[0],
                                                                           q2acQ_destruct_d[0],
                                                                           q1acP_destruct_d[0]} & {q4acS_destruct_r,
                                                                                                   q3acR_destruct_r,
                                                                                                   q2acQ_destruct_r,
                                                                                                   q1acP_destruct_r}));
  assign lizzieLet10_1QNode_Int_r = (& lizzieLet10_1QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet10_1QNode_Int_emitted <= 4'd0;
    else
      lizzieLet10_1QNode_Int_emitted <= (lizzieLet10_1QNode_Int_r ? 4'd0 :
                                         lizzieLet10_1QNode_Int_done);
  
  /* destruct (Ty QTree_Int,
          Dcon QVal_Int) : (lizzieLet10_1QVal_Int,QTree_Int) > [(vacO_destruct,Int)] */
  assign vacO_destruct_d = {lizzieLet10_1QVal_Int_d[34:3],
                            lizzieLet10_1QVal_Int_d[0]};
  assign lizzieLet10_1QVal_Int_r = vacO_destruct_r;
  
  /* demux (Ty QTree_Int,
       Ty QTree_Int) : (lizzieLet10_2,QTree_Int) (lizzieLet10_1,QTree_Int) > [(_32,QTree_Int),
                                                                              (lizzieLet10_1QVal_Int,QTree_Int),
                                                                              (lizzieLet10_1QNode_Int,QTree_Int),
                                                                              (_31,QTree_Int)] */
  logic [3:0] lizzieLet10_1_onehotd;
  always_comb
    if ((lizzieLet10_2_d[0] && lizzieLet10_1_d[0]))
      unique case (lizzieLet10_2_d[2:1])
        2'd0: lizzieLet10_1_onehotd = 4'd1;
        2'd1: lizzieLet10_1_onehotd = 4'd2;
        2'd2: lizzieLet10_1_onehotd = 4'd4;
        2'd3: lizzieLet10_1_onehotd = 4'd8;
        default: lizzieLet10_1_onehotd = 4'd0;
      endcase
    else lizzieLet10_1_onehotd = 4'd0;
  assign _32_d = {lizzieLet10_1_d[66:1], lizzieLet10_1_onehotd[0]};
  assign lizzieLet10_1QVal_Int_d = {lizzieLet10_1_d[66:1],
                                    lizzieLet10_1_onehotd[1]};
  assign lizzieLet10_1QNode_Int_d = {lizzieLet10_1_d[66:1],
                                     lizzieLet10_1_onehotd[2]};
  assign _31_d = {lizzieLet10_1_d[66:1], lizzieLet10_1_onehotd[3]};
  assign lizzieLet10_1_r = (| (lizzieLet10_1_onehotd & {_31_r,
                                                        lizzieLet10_1QNode_Int_r,
                                                        lizzieLet10_1QVal_Int_r,
                                                        _32_r}));
  assign lizzieLet10_2_r = lizzieLet10_1_r;
  
  /* demux (Ty QTree_Int,
       Ty MyDTInt_Int) : (lizzieLet10_3,QTree_Int) (gacM_goMux_mux,MyDTInt_Int) > [(_30,MyDTInt_Int),
                                                                                   (lizzieLet10_3QVal_Int,MyDTInt_Int),
                                                                                   (lizzieLet10_3QNode_Int,MyDTInt_Int),
                                                                                   (_29,MyDTInt_Int)] */
  logic [3:0] gacM_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet10_3_d[0] && gacM_goMux_mux_d[0]))
      unique case (lizzieLet10_3_d[2:1])
        2'd0: gacM_goMux_mux_onehotd = 4'd1;
        2'd1: gacM_goMux_mux_onehotd = 4'd2;
        2'd2: gacM_goMux_mux_onehotd = 4'd4;
        2'd3: gacM_goMux_mux_onehotd = 4'd8;
        default: gacM_goMux_mux_onehotd = 4'd0;
      endcase
    else gacM_goMux_mux_onehotd = 4'd0;
  assign _30_d = gacM_goMux_mux_onehotd[0];
  assign lizzieLet10_3QVal_Int_d = gacM_goMux_mux_onehotd[1];
  assign lizzieLet10_3QNode_Int_d = gacM_goMux_mux_onehotd[2];
  assign _29_d = gacM_goMux_mux_onehotd[3];
  assign gacM_goMux_mux_r = (| (gacM_goMux_mux_onehotd & {_29_r,
                                                          lizzieLet10_3QNode_Int_r,
                                                          lizzieLet10_3QVal_Int_r,
                                                          _30_r}));
  assign lizzieLet10_3_r = gacM_goMux_mux_r;
  
  /* fork (Ty MyDTInt_Int) : (lizzieLet10_3QNode_Int,MyDTInt_Int) > [(lizzieLet10_3QNode_Int_1,MyDTInt_Int),
                                                                (lizzieLet10_3QNode_Int_2,MyDTInt_Int)] */
  logic [1:0] lizzieLet10_3QNode_Int_emitted;
  logic [1:0] lizzieLet10_3QNode_Int_done;
  assign lizzieLet10_3QNode_Int_1_d = (lizzieLet10_3QNode_Int_d[0] && (! lizzieLet10_3QNode_Int_emitted[0]));
  assign lizzieLet10_3QNode_Int_2_d = (lizzieLet10_3QNode_Int_d[0] && (! lizzieLet10_3QNode_Int_emitted[1]));
  assign lizzieLet10_3QNode_Int_done = (lizzieLet10_3QNode_Int_emitted | ({lizzieLet10_3QNode_Int_2_d[0],
                                                                           lizzieLet10_3QNode_Int_1_d[0]} & {lizzieLet10_3QNode_Int_2_r,
                                                                                                             lizzieLet10_3QNode_Int_1_r}));
  assign lizzieLet10_3QNode_Int_r = (& lizzieLet10_3QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet10_3QNode_Int_emitted <= 2'd0;
    else
      lizzieLet10_3QNode_Int_emitted <= (lizzieLet10_3QNode_Int_r ? 2'd0 :
                                         lizzieLet10_3QNode_Int_done);
  
  /* buf (Ty MyDTInt_Int) : (lizzieLet10_3QNode_Int_2,MyDTInt_Int) > (lizzieLet10_3QNode_Int_2_argbuf,MyDTInt_Int) */
  MyDTInt_Int_t lizzieLet10_3QNode_Int_2_bufchan_d;
  logic lizzieLet10_3QNode_Int_2_bufchan_r;
  assign lizzieLet10_3QNode_Int_2_r = ((! lizzieLet10_3QNode_Int_2_bufchan_d[0]) || lizzieLet10_3QNode_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet10_3QNode_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet10_3QNode_Int_2_r)
        lizzieLet10_3QNode_Int_2_bufchan_d <= lizzieLet10_3QNode_Int_2_d;
  MyDTInt_Int_t lizzieLet10_3QNode_Int_2_bufchan_buf;
  assign lizzieLet10_3QNode_Int_2_bufchan_r = (! lizzieLet10_3QNode_Int_2_bufchan_buf[0]);
  assign lizzieLet10_3QNode_Int_2_argbuf_d = (lizzieLet10_3QNode_Int_2_bufchan_buf[0] ? lizzieLet10_3QNode_Int_2_bufchan_buf :
                                              lizzieLet10_3QNode_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet10_3QNode_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet10_3QNode_Int_2_argbuf_r && lizzieLet10_3QNode_Int_2_bufchan_buf[0]))
        lizzieLet10_3QNode_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet10_3QNode_Int_2_argbuf_r) && (! lizzieLet10_3QNode_Int_2_bufchan_buf[0])))
        lizzieLet10_3QNode_Int_2_bufchan_buf <= lizzieLet10_3QNode_Int_2_bufchan_d;
  
  /* buf (Ty MyDTInt_Int) : (lizzieLet10_3QVal_Int,MyDTInt_Int) > (lizzieLet10_3QVal_Int_1_argbuf,MyDTInt_Int) */
  MyDTInt_Int_t lizzieLet10_3QVal_Int_bufchan_d;
  logic lizzieLet10_3QVal_Int_bufchan_r;
  assign lizzieLet10_3QVal_Int_r = ((! lizzieLet10_3QVal_Int_bufchan_d[0]) || lizzieLet10_3QVal_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet10_3QVal_Int_bufchan_d <= 1'd0;
    else
      if (lizzieLet10_3QVal_Int_r)
        lizzieLet10_3QVal_Int_bufchan_d <= lizzieLet10_3QVal_Int_d;
  MyDTInt_Int_t lizzieLet10_3QVal_Int_bufchan_buf;
  assign lizzieLet10_3QVal_Int_bufchan_r = (! lizzieLet10_3QVal_Int_bufchan_buf[0]);
  assign lizzieLet10_3QVal_Int_1_argbuf_d = (lizzieLet10_3QVal_Int_bufchan_buf[0] ? lizzieLet10_3QVal_Int_bufchan_buf :
                                             lizzieLet10_3QVal_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet10_3QVal_Int_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet10_3QVal_Int_1_argbuf_r && lizzieLet10_3QVal_Int_bufchan_buf[0]))
        lizzieLet10_3QVal_Int_bufchan_buf <= 1'd0;
      else if (((! lizzieLet10_3QVal_Int_1_argbuf_r) && (! lizzieLet10_3QVal_Int_bufchan_buf[0])))
        lizzieLet10_3QVal_Int_bufchan_buf <= lizzieLet10_3QVal_Int_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Go) : (lizzieLet10_4,QTree_Int) (go_13_goMux_data,Go) > [(lizzieLet10_4QNone_Int,Go),
                                                                   (lizzieLet10_4QVal_Int,Go),
                                                                   (lizzieLet10_4QNode_Int,Go),
                                                                   (lizzieLet10_4QError_Int,Go)] */
  logic [3:0] go_13_goMux_data_onehotd;
  always_comb
    if ((lizzieLet10_4_d[0] && go_13_goMux_data_d[0]))
      unique case (lizzieLet10_4_d[2:1])
        2'd0: go_13_goMux_data_onehotd = 4'd1;
        2'd1: go_13_goMux_data_onehotd = 4'd2;
        2'd2: go_13_goMux_data_onehotd = 4'd4;
        2'd3: go_13_goMux_data_onehotd = 4'd8;
        default: go_13_goMux_data_onehotd = 4'd0;
      endcase
    else go_13_goMux_data_onehotd = 4'd0;
  assign lizzieLet10_4QNone_Int_d = go_13_goMux_data_onehotd[0];
  assign lizzieLet10_4QVal_Int_d = go_13_goMux_data_onehotd[1];
  assign lizzieLet10_4QNode_Int_d = go_13_goMux_data_onehotd[2];
  assign lizzieLet10_4QError_Int_d = go_13_goMux_data_onehotd[3];
  assign go_13_goMux_data_r = (| (go_13_goMux_data_onehotd & {lizzieLet10_4QError_Int_r,
                                                              lizzieLet10_4QNode_Int_r,
                                                              lizzieLet10_4QVal_Int_r,
                                                              lizzieLet10_4QNone_Int_r}));
  assign lizzieLet10_4_r = go_13_goMux_data_r;
  
  /* fork (Ty Go) : (lizzieLet10_4QError_Int,Go) > [(lizzieLet10_4QError_Int_1,Go),
                                               (lizzieLet10_4QError_Int_2,Go)] */
  logic [1:0] lizzieLet10_4QError_Int_emitted;
  logic [1:0] lizzieLet10_4QError_Int_done;
  assign lizzieLet10_4QError_Int_1_d = (lizzieLet10_4QError_Int_d[0] && (! lizzieLet10_4QError_Int_emitted[0]));
  assign lizzieLet10_4QError_Int_2_d = (lizzieLet10_4QError_Int_d[0] && (! lizzieLet10_4QError_Int_emitted[1]));
  assign lizzieLet10_4QError_Int_done = (lizzieLet10_4QError_Int_emitted | ({lizzieLet10_4QError_Int_2_d[0],
                                                                             lizzieLet10_4QError_Int_1_d[0]} & {lizzieLet10_4QError_Int_2_r,
                                                                                                                lizzieLet10_4QError_Int_1_r}));
  assign lizzieLet10_4QError_Int_r = (& lizzieLet10_4QError_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet10_4QError_Int_emitted <= 2'd0;
    else
      lizzieLet10_4QError_Int_emitted <= (lizzieLet10_4QError_Int_r ? 2'd0 :
                                          lizzieLet10_4QError_Int_done);
  
  /* dcon (Ty QTree_Int,
      Dcon QError_Int) : [(lizzieLet10_4QError_Int_1,Go)] > (lizzieLet10_4QError_Int_1QError_Int,QTree_Int) */
  assign lizzieLet10_4QError_Int_1QError_Int_d = QError_Int_dc((& {lizzieLet10_4QError_Int_1_d[0]}), lizzieLet10_4QError_Int_1_d);
  assign {lizzieLet10_4QError_Int_1_r} = {1 {(lizzieLet10_4QError_Int_1QError_Int_r && lizzieLet10_4QError_Int_1QError_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (lizzieLet10_4QError_Int_1QError_Int,QTree_Int) > (lizzieLet15_2_1_argbuf,QTree_Int) */
  QTree_Int_t lizzieLet10_4QError_Int_1QError_Int_bufchan_d;
  logic lizzieLet10_4QError_Int_1QError_Int_bufchan_r;
  assign lizzieLet10_4QError_Int_1QError_Int_r = ((! lizzieLet10_4QError_Int_1QError_Int_bufchan_d[0]) || lizzieLet10_4QError_Int_1QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet10_4QError_Int_1QError_Int_bufchan_d <= {66'd0, 1'd0};
    else
      if (lizzieLet10_4QError_Int_1QError_Int_r)
        lizzieLet10_4QError_Int_1QError_Int_bufchan_d <= lizzieLet10_4QError_Int_1QError_Int_d;
  QTree_Int_t lizzieLet10_4QError_Int_1QError_Int_bufchan_buf;
  assign lizzieLet10_4QError_Int_1QError_Int_bufchan_r = (! lizzieLet10_4QError_Int_1QError_Int_bufchan_buf[0]);
  assign lizzieLet15_2_1_argbuf_d = (lizzieLet10_4QError_Int_1QError_Int_bufchan_buf[0] ? lizzieLet10_4QError_Int_1QError_Int_bufchan_buf :
                                     lizzieLet10_4QError_Int_1QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet10_4QError_Int_1QError_Int_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((lizzieLet15_2_1_argbuf_r && lizzieLet10_4QError_Int_1QError_Int_bufchan_buf[0]))
        lizzieLet10_4QError_Int_1QError_Int_bufchan_buf <= {66'd0, 1'd0};
      else if (((! lizzieLet15_2_1_argbuf_r) && (! lizzieLet10_4QError_Int_1QError_Int_bufchan_buf[0])))
        lizzieLet10_4QError_Int_1QError_Int_bufchan_buf <= lizzieLet10_4QError_Int_1QError_Int_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet10_4QError_Int_2,Go) > (lizzieLet10_4QError_Int_2_argbuf,Go) */
  Go_t lizzieLet10_4QError_Int_2_bufchan_d;
  logic lizzieLet10_4QError_Int_2_bufchan_r;
  assign lizzieLet10_4QError_Int_2_r = ((! lizzieLet10_4QError_Int_2_bufchan_d[0]) || lizzieLet10_4QError_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet10_4QError_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet10_4QError_Int_2_r)
        lizzieLet10_4QError_Int_2_bufchan_d <= lizzieLet10_4QError_Int_2_d;
  Go_t lizzieLet10_4QError_Int_2_bufchan_buf;
  assign lizzieLet10_4QError_Int_2_bufchan_r = (! lizzieLet10_4QError_Int_2_bufchan_buf[0]);
  assign lizzieLet10_4QError_Int_2_argbuf_d = (lizzieLet10_4QError_Int_2_bufchan_buf[0] ? lizzieLet10_4QError_Int_2_bufchan_buf :
                                               lizzieLet10_4QError_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet10_4QError_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet10_4QError_Int_2_argbuf_r && lizzieLet10_4QError_Int_2_bufchan_buf[0]))
        lizzieLet10_4QError_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet10_4QError_Int_2_argbuf_r) && (! lizzieLet10_4QError_Int_2_bufchan_buf[0])))
        lizzieLet10_4QError_Int_2_bufchan_buf <= lizzieLet10_4QError_Int_2_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet10_4QNode_Int,Go) > (lizzieLet10_4QNode_Int_1_argbuf,Go) */
  Go_t lizzieLet10_4QNode_Int_bufchan_d;
  logic lizzieLet10_4QNode_Int_bufchan_r;
  assign lizzieLet10_4QNode_Int_r = ((! lizzieLet10_4QNode_Int_bufchan_d[0]) || lizzieLet10_4QNode_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet10_4QNode_Int_bufchan_d <= 1'd0;
    else
      if (lizzieLet10_4QNode_Int_r)
        lizzieLet10_4QNode_Int_bufchan_d <= lizzieLet10_4QNode_Int_d;
  Go_t lizzieLet10_4QNode_Int_bufchan_buf;
  assign lizzieLet10_4QNode_Int_bufchan_r = (! lizzieLet10_4QNode_Int_bufchan_buf[0]);
  assign lizzieLet10_4QNode_Int_1_argbuf_d = (lizzieLet10_4QNode_Int_bufchan_buf[0] ? lizzieLet10_4QNode_Int_bufchan_buf :
                                              lizzieLet10_4QNode_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet10_4QNode_Int_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet10_4QNode_Int_1_argbuf_r && lizzieLet10_4QNode_Int_bufchan_buf[0]))
        lizzieLet10_4QNode_Int_bufchan_buf <= 1'd0;
      else if (((! lizzieLet10_4QNode_Int_1_argbuf_r) && (! lizzieLet10_4QNode_Int_bufchan_buf[0])))
        lizzieLet10_4QNode_Int_bufchan_buf <= lizzieLet10_4QNode_Int_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet10_4QNone_Int,Go) > [(lizzieLet10_4QNone_Int_1,Go),
                                              (lizzieLet10_4QNone_Int_2,Go)] */
  logic [1:0] lizzieLet10_4QNone_Int_emitted;
  logic [1:0] lizzieLet10_4QNone_Int_done;
  assign lizzieLet10_4QNone_Int_1_d = (lizzieLet10_4QNone_Int_d[0] && (! lizzieLet10_4QNone_Int_emitted[0]));
  assign lizzieLet10_4QNone_Int_2_d = (lizzieLet10_4QNone_Int_d[0] && (! lizzieLet10_4QNone_Int_emitted[1]));
  assign lizzieLet10_4QNone_Int_done = (lizzieLet10_4QNone_Int_emitted | ({lizzieLet10_4QNone_Int_2_d[0],
                                                                           lizzieLet10_4QNone_Int_1_d[0]} & {lizzieLet10_4QNone_Int_2_r,
                                                                                                             lizzieLet10_4QNone_Int_1_r}));
  assign lizzieLet10_4QNone_Int_r = (& lizzieLet10_4QNone_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet10_4QNone_Int_emitted <= 2'd0;
    else
      lizzieLet10_4QNone_Int_emitted <= (lizzieLet10_4QNone_Int_r ? 2'd0 :
                                         lizzieLet10_4QNone_Int_done);
  
  /* dcon (Ty QTree_Int,
      Dcon QNone_Int) : [(lizzieLet10_4QNone_Int_1,Go)] > (lizzieLet10_4QNone_Int_1QNone_Int,QTree_Int) */
  assign lizzieLet10_4QNone_Int_1QNone_Int_d = QNone_Int_dc((& {lizzieLet10_4QNone_Int_1_d[0]}), lizzieLet10_4QNone_Int_1_d);
  assign {lizzieLet10_4QNone_Int_1_r} = {1 {(lizzieLet10_4QNone_Int_1QNone_Int_r && lizzieLet10_4QNone_Int_1QNone_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (lizzieLet10_4QNone_Int_1QNone_Int,QTree_Int) > (lizzieLet11_1_1_argbuf,QTree_Int) */
  QTree_Int_t lizzieLet10_4QNone_Int_1QNone_Int_bufchan_d;
  logic lizzieLet10_4QNone_Int_1QNone_Int_bufchan_r;
  assign lizzieLet10_4QNone_Int_1QNone_Int_r = ((! lizzieLet10_4QNone_Int_1QNone_Int_bufchan_d[0]) || lizzieLet10_4QNone_Int_1QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet10_4QNone_Int_1QNone_Int_bufchan_d <= {66'd0, 1'd0};
    else
      if (lizzieLet10_4QNone_Int_1QNone_Int_r)
        lizzieLet10_4QNone_Int_1QNone_Int_bufchan_d <= lizzieLet10_4QNone_Int_1QNone_Int_d;
  QTree_Int_t lizzieLet10_4QNone_Int_1QNone_Int_bufchan_buf;
  assign lizzieLet10_4QNone_Int_1QNone_Int_bufchan_r = (! lizzieLet10_4QNone_Int_1QNone_Int_bufchan_buf[0]);
  assign lizzieLet11_1_1_argbuf_d = (lizzieLet10_4QNone_Int_1QNone_Int_bufchan_buf[0] ? lizzieLet10_4QNone_Int_1QNone_Int_bufchan_buf :
                                     lizzieLet10_4QNone_Int_1QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet10_4QNone_Int_1QNone_Int_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((lizzieLet11_1_1_argbuf_r && lizzieLet10_4QNone_Int_1QNone_Int_bufchan_buf[0]))
        lizzieLet10_4QNone_Int_1QNone_Int_bufchan_buf <= {66'd0, 1'd0};
      else if (((! lizzieLet11_1_1_argbuf_r) && (! lizzieLet10_4QNone_Int_1QNone_Int_bufchan_buf[0])))
        lizzieLet10_4QNone_Int_1QNone_Int_bufchan_buf <= lizzieLet10_4QNone_Int_1QNone_Int_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet10_4QNone_Int_2,Go) > (lizzieLet10_4QNone_Int_2_argbuf,Go) */
  Go_t lizzieLet10_4QNone_Int_2_bufchan_d;
  logic lizzieLet10_4QNone_Int_2_bufchan_r;
  assign lizzieLet10_4QNone_Int_2_r = ((! lizzieLet10_4QNone_Int_2_bufchan_d[0]) || lizzieLet10_4QNone_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet10_4QNone_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet10_4QNone_Int_2_r)
        lizzieLet10_4QNone_Int_2_bufchan_d <= lizzieLet10_4QNone_Int_2_d;
  Go_t lizzieLet10_4QNone_Int_2_bufchan_buf;
  assign lizzieLet10_4QNone_Int_2_bufchan_r = (! lizzieLet10_4QNone_Int_2_bufchan_buf[0]);
  assign lizzieLet10_4QNone_Int_2_argbuf_d = (lizzieLet10_4QNone_Int_2_bufchan_buf[0] ? lizzieLet10_4QNone_Int_2_bufchan_buf :
                                              lizzieLet10_4QNone_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet10_4QNone_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet10_4QNone_Int_2_argbuf_r && lizzieLet10_4QNone_Int_2_bufchan_buf[0]))
        lizzieLet10_4QNone_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet10_4QNone_Int_2_argbuf_r) && (! lizzieLet10_4QNone_Int_2_bufchan_buf[0])))
        lizzieLet10_4QNone_Int_2_bufchan_buf <= lizzieLet10_4QNone_Int_2_bufchan_d;
  
  /* mergectrl (Ty C5,Ty Go) : [(lizzieLet10_4QNone_Int_2_argbuf,Go),
                           (lizzieLet34_3Lcall_main_map'_Int_Int0_1_argbuf,Go),
                           (es_0_4_1MyFalse_1_argbuf,Go),
                           (es_0_4_1MyTrue_2_argbuf,Go),
                           (lizzieLet10_4QError_Int_2_argbuf,Go)] > (go_20_goMux_choice,C5) (go_20_goMux_data,Go) */
  logic [4:0] lizzieLet10_4QNone_Int_2_argbuf_select_d;
  assign lizzieLet10_4QNone_Int_2_argbuf_select_d = ((| lizzieLet10_4QNone_Int_2_argbuf_select_q) ? lizzieLet10_4QNone_Int_2_argbuf_select_q :
                                                     (lizzieLet10_4QNone_Int_2_argbuf_d[0] ? 5'd1 :
                                                      (\lizzieLet34_3Lcall_main_map'_Int_Int0_1_argbuf_d [0] ? 5'd2 :
                                                       (es_0_4_1MyFalse_1_argbuf_d[0] ? 5'd4 :
                                                        (es_0_4_1MyTrue_2_argbuf_d[0] ? 5'd8 :
                                                         (lizzieLet10_4QError_Int_2_argbuf_d[0] ? 5'd16 :
                                                          5'd0))))));
  logic [4:0] lizzieLet10_4QNone_Int_2_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet10_4QNone_Int_2_argbuf_select_q <= 5'd0;
    else
      lizzieLet10_4QNone_Int_2_argbuf_select_q <= (lizzieLet10_4QNone_Int_2_argbuf_done ? 5'd0 :
                                                   lizzieLet10_4QNone_Int_2_argbuf_select_d);
  logic [1:0] lizzieLet10_4QNone_Int_2_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet10_4QNone_Int_2_argbuf_emit_q <= 2'd0;
    else
      lizzieLet10_4QNone_Int_2_argbuf_emit_q <= (lizzieLet10_4QNone_Int_2_argbuf_done ? 2'd0 :
                                                 lizzieLet10_4QNone_Int_2_argbuf_emit_d);
  logic [1:0] lizzieLet10_4QNone_Int_2_argbuf_emit_d;
  assign lizzieLet10_4QNone_Int_2_argbuf_emit_d = (lizzieLet10_4QNone_Int_2_argbuf_emit_q | ({go_20_goMux_choice_d[0],
                                                                                              go_20_goMux_data_d[0]} & {go_20_goMux_choice_r,
                                                                                                                        go_20_goMux_data_r}));
  logic lizzieLet10_4QNone_Int_2_argbuf_done;
  assign lizzieLet10_4QNone_Int_2_argbuf_done = (& lizzieLet10_4QNone_Int_2_argbuf_emit_d);
  assign {lizzieLet10_4QError_Int_2_argbuf_r,
          es_0_4_1MyTrue_2_argbuf_r,
          es_0_4_1MyFalse_1_argbuf_r,
          \lizzieLet34_3Lcall_main_map'_Int_Int0_1_argbuf_r ,
          lizzieLet10_4QNone_Int_2_argbuf_r} = (lizzieLet10_4QNone_Int_2_argbuf_done ? lizzieLet10_4QNone_Int_2_argbuf_select_d :
                                                5'd0);
  assign go_20_goMux_data_d = ((lizzieLet10_4QNone_Int_2_argbuf_select_d[0] && (! lizzieLet10_4QNone_Int_2_argbuf_emit_q[0])) ? lizzieLet10_4QNone_Int_2_argbuf_d :
                               ((lizzieLet10_4QNone_Int_2_argbuf_select_d[1] && (! lizzieLet10_4QNone_Int_2_argbuf_emit_q[0])) ? \lizzieLet34_3Lcall_main_map'_Int_Int0_1_argbuf_d  :
                                ((lizzieLet10_4QNone_Int_2_argbuf_select_d[2] && (! lizzieLet10_4QNone_Int_2_argbuf_emit_q[0])) ? es_0_4_1MyFalse_1_argbuf_d :
                                 ((lizzieLet10_4QNone_Int_2_argbuf_select_d[3] && (! lizzieLet10_4QNone_Int_2_argbuf_emit_q[0])) ? es_0_4_1MyTrue_2_argbuf_d :
                                  ((lizzieLet10_4QNone_Int_2_argbuf_select_d[4] && (! lizzieLet10_4QNone_Int_2_argbuf_emit_q[0])) ? lizzieLet10_4QError_Int_2_argbuf_d :
                                   1'd0)))));
  assign go_20_goMux_choice_d = ((lizzieLet10_4QNone_Int_2_argbuf_select_d[0] && (! lizzieLet10_4QNone_Int_2_argbuf_emit_q[1])) ? C1_5_dc(1'd1) :
                                 ((lizzieLet10_4QNone_Int_2_argbuf_select_d[1] && (! lizzieLet10_4QNone_Int_2_argbuf_emit_q[1])) ? C2_5_dc(1'd1) :
                                  ((lizzieLet10_4QNone_Int_2_argbuf_select_d[2] && (! lizzieLet10_4QNone_Int_2_argbuf_emit_q[1])) ? C3_5_dc(1'd1) :
                                   ((lizzieLet10_4QNone_Int_2_argbuf_select_d[3] && (! lizzieLet10_4QNone_Int_2_argbuf_emit_q[1])) ? C4_5_dc(1'd1) :
                                    ((lizzieLet10_4QNone_Int_2_argbuf_select_d[4] && (! lizzieLet10_4QNone_Int_2_argbuf_emit_q[1])) ? C5_5_dc(1'd1) :
                                     {3'd0, 1'd0})))));
  
  /* fork (Ty Go) : (lizzieLet10_4QVal_Int,Go) > [(lizzieLet10_4QVal_Int_1,Go),
                                             (lizzieLet10_4QVal_Int_2,Go),
                                             (lizzieLet10_4QVal_Int_3,Go)] */
  logic [2:0] lizzieLet10_4QVal_Int_emitted;
  logic [2:0] lizzieLet10_4QVal_Int_done;
  assign lizzieLet10_4QVal_Int_1_d = (lizzieLet10_4QVal_Int_d[0] && (! lizzieLet10_4QVal_Int_emitted[0]));
  assign lizzieLet10_4QVal_Int_2_d = (lizzieLet10_4QVal_Int_d[0] && (! lizzieLet10_4QVal_Int_emitted[1]));
  assign lizzieLet10_4QVal_Int_3_d = (lizzieLet10_4QVal_Int_d[0] && (! lizzieLet10_4QVal_Int_emitted[2]));
  assign lizzieLet10_4QVal_Int_done = (lizzieLet10_4QVal_Int_emitted | ({lizzieLet10_4QVal_Int_3_d[0],
                                                                         lizzieLet10_4QVal_Int_2_d[0],
                                                                         lizzieLet10_4QVal_Int_1_d[0]} & {lizzieLet10_4QVal_Int_3_r,
                                                                                                          lizzieLet10_4QVal_Int_2_r,
                                                                                                          lizzieLet10_4QVal_Int_1_r}));
  assign lizzieLet10_4QVal_Int_r = (& lizzieLet10_4QVal_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet10_4QVal_Int_emitted <= 3'd0;
    else
      lizzieLet10_4QVal_Int_emitted <= (lizzieLet10_4QVal_Int_r ? 3'd0 :
                                        lizzieLet10_4QVal_Int_done);
  
  /* buf (Ty Go) : (lizzieLet10_4QVal_Int_1,Go) > (lizzieLet10_4QVal_Int_1_argbuf,Go) */
  Go_t lizzieLet10_4QVal_Int_1_bufchan_d;
  logic lizzieLet10_4QVal_Int_1_bufchan_r;
  assign lizzieLet10_4QVal_Int_1_r = ((! lizzieLet10_4QVal_Int_1_bufchan_d[0]) || lizzieLet10_4QVal_Int_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet10_4QVal_Int_1_bufchan_d <= 1'd0;
    else
      if (lizzieLet10_4QVal_Int_1_r)
        lizzieLet10_4QVal_Int_1_bufchan_d <= lizzieLet10_4QVal_Int_1_d;
  Go_t lizzieLet10_4QVal_Int_1_bufchan_buf;
  assign lizzieLet10_4QVal_Int_1_bufchan_r = (! lizzieLet10_4QVal_Int_1_bufchan_buf[0]);
  assign lizzieLet10_4QVal_Int_1_argbuf_d = (lizzieLet10_4QVal_Int_1_bufchan_buf[0] ? lizzieLet10_4QVal_Int_1_bufchan_buf :
                                             lizzieLet10_4QVal_Int_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet10_4QVal_Int_1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet10_4QVal_Int_1_argbuf_r && lizzieLet10_4QVal_Int_1_bufchan_buf[0]))
        lizzieLet10_4QVal_Int_1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet10_4QVal_Int_1_argbuf_r) && (! lizzieLet10_4QVal_Int_1_bufchan_buf[0])))
        lizzieLet10_4QVal_Int_1_bufchan_buf <= lizzieLet10_4QVal_Int_1_bufchan_d;
  
  /* dcon (Ty TupGo___MyDTInt_Int___Int,
      Dcon TupGo___MyDTInt_Int___Int) : [(lizzieLet10_4QVal_Int_1_argbuf,Go),
                                         (lizzieLet10_3QVal_Int_1_argbuf,MyDTInt_Int),
                                         (vacO_1_argbuf,Int)] > (applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1,TupGo___MyDTInt_Int___Int) */
  assign applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_d = TupGo___MyDTInt_Int___Int_dc((& {lizzieLet10_4QVal_Int_1_argbuf_d[0],
                                                                                          lizzieLet10_3QVal_Int_1_argbuf_d[0],
                                                                                          vacO_1_argbuf_d[0]}), lizzieLet10_4QVal_Int_1_argbuf_d, lizzieLet10_3QVal_Int_1_argbuf_d, vacO_1_argbuf_d);
  assign {lizzieLet10_4QVal_Int_1_argbuf_r,
          lizzieLet10_3QVal_Int_1_argbuf_r,
          vacO_1_argbuf_r} = {3 {(applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_r && applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_d[0])}};
  
  /* buf (Ty Go) : (lizzieLet10_4QVal_Int_2,Go) > (lizzieLet10_4QVal_Int_2_argbuf,Go) */
  Go_t lizzieLet10_4QVal_Int_2_bufchan_d;
  logic lizzieLet10_4QVal_Int_2_bufchan_r;
  assign lizzieLet10_4QVal_Int_2_r = ((! lizzieLet10_4QVal_Int_2_bufchan_d[0]) || lizzieLet10_4QVal_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet10_4QVal_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet10_4QVal_Int_2_r)
        lizzieLet10_4QVal_Int_2_bufchan_d <= lizzieLet10_4QVal_Int_2_d;
  Go_t lizzieLet10_4QVal_Int_2_bufchan_buf;
  assign lizzieLet10_4QVal_Int_2_bufchan_r = (! lizzieLet10_4QVal_Int_2_bufchan_buf[0]);
  assign lizzieLet10_4QVal_Int_2_argbuf_d = (lizzieLet10_4QVal_Int_2_bufchan_buf[0] ? lizzieLet10_4QVal_Int_2_bufchan_buf :
                                             lizzieLet10_4QVal_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet10_4QVal_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet10_4QVal_Int_2_argbuf_r && lizzieLet10_4QVal_Int_2_bufchan_buf[0]))
        lizzieLet10_4QVal_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet10_4QVal_Int_2_argbuf_r) && (! lizzieLet10_4QVal_Int_2_bufchan_buf[0])))
        lizzieLet10_4QVal_Int_2_bufchan_buf <= lizzieLet10_4QVal_Int_2_bufchan_d;
  
  /* dcon (Ty TupGo___MyDTInt_Bool___Int,
      Dcon TupGo___MyDTInt_Bool___Int) : [(lizzieLet10_4QVal_Int_2_argbuf,Go),
                                          (lizzieLet10_5QVal_Int_1_argbuf,MyDTInt_Bool),
                                          (xacr_1_argbuf,Int)] > (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int2,TupGo___MyDTInt_Bool___Int) */
  assign applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int2_d = TupGo___MyDTInt_Bool___Int_dc((& {lizzieLet10_4QVal_Int_2_argbuf_d[0],
                                                                                            lizzieLet10_5QVal_Int_1_argbuf_d[0],
                                                                                            xacr_1_argbuf_d[0]}), lizzieLet10_4QVal_Int_2_argbuf_d, lizzieLet10_5QVal_Int_1_argbuf_d, xacr_1_argbuf_d);
  assign {lizzieLet10_4QVal_Int_2_argbuf_r,
          lizzieLet10_5QVal_Int_1_argbuf_r,
          xacr_1_argbuf_r} = {3 {(applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int2_r && applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int2_d[0])}};
  
  /* demux (Ty QTree_Int,
       Ty MyDTInt_Bool) : (lizzieLet10_5,QTree_Int) (isZacL_goMux_mux,MyDTInt_Bool) > [(_28,MyDTInt_Bool),
                                                                                       (lizzieLet10_5QVal_Int,MyDTInt_Bool),
                                                                                       (lizzieLet10_5QNode_Int,MyDTInt_Bool),
                                                                                       (_27,MyDTInt_Bool)] */
  logic [3:0] isZacL_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet10_5_d[0] && isZacL_goMux_mux_d[0]))
      unique case (lizzieLet10_5_d[2:1])
        2'd0: isZacL_goMux_mux_onehotd = 4'd1;
        2'd1: isZacL_goMux_mux_onehotd = 4'd2;
        2'd2: isZacL_goMux_mux_onehotd = 4'd4;
        2'd3: isZacL_goMux_mux_onehotd = 4'd8;
        default: isZacL_goMux_mux_onehotd = 4'd0;
      endcase
    else isZacL_goMux_mux_onehotd = 4'd0;
  assign _28_d = isZacL_goMux_mux_onehotd[0];
  assign lizzieLet10_5QVal_Int_d = isZacL_goMux_mux_onehotd[1];
  assign lizzieLet10_5QNode_Int_d = isZacL_goMux_mux_onehotd[2];
  assign _27_d = isZacL_goMux_mux_onehotd[3];
  assign isZacL_goMux_mux_r = (| (isZacL_goMux_mux_onehotd & {_27_r,
                                                              lizzieLet10_5QNode_Int_r,
                                                              lizzieLet10_5QVal_Int_r,
                                                              _28_r}));
  assign lizzieLet10_5_r = isZacL_goMux_mux_r;
  
  /* fork (Ty MyDTInt_Bool) : (lizzieLet10_5QNode_Int,MyDTInt_Bool) > [(lizzieLet10_5QNode_Int_1,MyDTInt_Bool),
                                                                  (lizzieLet10_5QNode_Int_2,MyDTInt_Bool)] */
  logic [1:0] lizzieLet10_5QNode_Int_emitted;
  logic [1:0] lizzieLet10_5QNode_Int_done;
  assign lizzieLet10_5QNode_Int_1_d = (lizzieLet10_5QNode_Int_d[0] && (! lizzieLet10_5QNode_Int_emitted[0]));
  assign lizzieLet10_5QNode_Int_2_d = (lizzieLet10_5QNode_Int_d[0] && (! lizzieLet10_5QNode_Int_emitted[1]));
  assign lizzieLet10_5QNode_Int_done = (lizzieLet10_5QNode_Int_emitted | ({lizzieLet10_5QNode_Int_2_d[0],
                                                                           lizzieLet10_5QNode_Int_1_d[0]} & {lizzieLet10_5QNode_Int_2_r,
                                                                                                             lizzieLet10_5QNode_Int_1_r}));
  assign lizzieLet10_5QNode_Int_r = (& lizzieLet10_5QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet10_5QNode_Int_emitted <= 2'd0;
    else
      lizzieLet10_5QNode_Int_emitted <= (lizzieLet10_5QNode_Int_r ? 2'd0 :
                                         lizzieLet10_5QNode_Int_done);
  
  /* buf (Ty MyDTInt_Bool) : (lizzieLet10_5QNode_Int_2,MyDTInt_Bool) > (lizzieLet10_5QNode_Int_2_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t lizzieLet10_5QNode_Int_2_bufchan_d;
  logic lizzieLet10_5QNode_Int_2_bufchan_r;
  assign lizzieLet10_5QNode_Int_2_r = ((! lizzieLet10_5QNode_Int_2_bufchan_d[0]) || lizzieLet10_5QNode_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet10_5QNode_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet10_5QNode_Int_2_r)
        lizzieLet10_5QNode_Int_2_bufchan_d <= lizzieLet10_5QNode_Int_2_d;
  MyDTInt_Bool_t lizzieLet10_5QNode_Int_2_bufchan_buf;
  assign lizzieLet10_5QNode_Int_2_bufchan_r = (! lizzieLet10_5QNode_Int_2_bufchan_buf[0]);
  assign lizzieLet10_5QNode_Int_2_argbuf_d = (lizzieLet10_5QNode_Int_2_bufchan_buf[0] ? lizzieLet10_5QNode_Int_2_bufchan_buf :
                                              lizzieLet10_5QNode_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet10_5QNode_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet10_5QNode_Int_2_argbuf_r && lizzieLet10_5QNode_Int_2_bufchan_buf[0]))
        lizzieLet10_5QNode_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet10_5QNode_Int_2_argbuf_r) && (! lizzieLet10_5QNode_Int_2_bufchan_buf[0])))
        lizzieLet10_5QNode_Int_2_bufchan_buf <= lizzieLet10_5QNode_Int_2_bufchan_d;
  
  /* buf (Ty MyDTInt_Bool) : (lizzieLet10_5QVal_Int,MyDTInt_Bool) > (lizzieLet10_5QVal_Int_1_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t lizzieLet10_5QVal_Int_bufchan_d;
  logic lizzieLet10_5QVal_Int_bufchan_r;
  assign lizzieLet10_5QVal_Int_r = ((! lizzieLet10_5QVal_Int_bufchan_d[0]) || lizzieLet10_5QVal_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet10_5QVal_Int_bufchan_d <= 1'd0;
    else
      if (lizzieLet10_5QVal_Int_r)
        lizzieLet10_5QVal_Int_bufchan_d <= lizzieLet10_5QVal_Int_d;
  MyDTInt_Bool_t lizzieLet10_5QVal_Int_bufchan_buf;
  assign lizzieLet10_5QVal_Int_bufchan_r = (! lizzieLet10_5QVal_Int_bufchan_buf[0]);
  assign lizzieLet10_5QVal_Int_1_argbuf_d = (lizzieLet10_5QVal_Int_bufchan_buf[0] ? lizzieLet10_5QVal_Int_bufchan_buf :
                                             lizzieLet10_5QVal_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet10_5QVal_Int_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet10_5QVal_Int_1_argbuf_r && lizzieLet10_5QVal_Int_bufchan_buf[0]))
        lizzieLet10_5QVal_Int_bufchan_buf <= 1'd0;
      else if (((! lizzieLet10_5QVal_Int_1_argbuf_r) && (! lizzieLet10_5QVal_Int_bufchan_buf[0])))
        lizzieLet10_5QVal_Int_bufchan_buf <= lizzieLet10_5QVal_Int_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_CTmain_map'_Int_Int) : (lizzieLet10_6,QTree_Int) (sc_0_2_goMux_mux,Pointer_CTmain_map'_Int_Int) > [(lizzieLet10_6QNone_Int,Pointer_CTmain_map'_Int_Int),
                                                                                                                     (lizzieLet10_6QVal_Int,Pointer_CTmain_map'_Int_Int),
                                                                                                                     (lizzieLet10_6QNode_Int,Pointer_CTmain_map'_Int_Int),
                                                                                                                     (lizzieLet10_6QError_Int,Pointer_CTmain_map'_Int_Int)] */
  logic [3:0] sc_0_2_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet10_6_d[0] && sc_0_2_goMux_mux_d[0]))
      unique case (lizzieLet10_6_d[2:1])
        2'd0: sc_0_2_goMux_mux_onehotd = 4'd1;
        2'd1: sc_0_2_goMux_mux_onehotd = 4'd2;
        2'd2: sc_0_2_goMux_mux_onehotd = 4'd4;
        2'd3: sc_0_2_goMux_mux_onehotd = 4'd8;
        default: sc_0_2_goMux_mux_onehotd = 4'd0;
      endcase
    else sc_0_2_goMux_mux_onehotd = 4'd0;
  assign lizzieLet10_6QNone_Int_d = {sc_0_2_goMux_mux_d[16:1],
                                     sc_0_2_goMux_mux_onehotd[0]};
  assign lizzieLet10_6QVal_Int_d = {sc_0_2_goMux_mux_d[16:1],
                                    sc_0_2_goMux_mux_onehotd[1]};
  assign lizzieLet10_6QNode_Int_d = {sc_0_2_goMux_mux_d[16:1],
                                     sc_0_2_goMux_mux_onehotd[2]};
  assign lizzieLet10_6QError_Int_d = {sc_0_2_goMux_mux_d[16:1],
                                      sc_0_2_goMux_mux_onehotd[3]};
  assign sc_0_2_goMux_mux_r = (| (sc_0_2_goMux_mux_onehotd & {lizzieLet10_6QError_Int_r,
                                                              lizzieLet10_6QNode_Int_r,
                                                              lizzieLet10_6QVal_Int_r,
                                                              lizzieLet10_6QNone_Int_r}));
  assign lizzieLet10_6_r = sc_0_2_goMux_mux_r;
  
  /* buf (Ty Pointer_CTmain_map'_Int_Int) : (lizzieLet10_6QError_Int,Pointer_CTmain_map'_Int_Int) > (lizzieLet10_6QError_Int_1_argbuf,Pointer_CTmain_map'_Int_Int) */
  \Pointer_CTmain_map'_Int_Int_t  lizzieLet10_6QError_Int_bufchan_d;
  logic lizzieLet10_6QError_Int_bufchan_r;
  assign lizzieLet10_6QError_Int_r = ((! lizzieLet10_6QError_Int_bufchan_d[0]) || lizzieLet10_6QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet10_6QError_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet10_6QError_Int_r)
        lizzieLet10_6QError_Int_bufchan_d <= lizzieLet10_6QError_Int_d;
  \Pointer_CTmain_map'_Int_Int_t  lizzieLet10_6QError_Int_bufchan_buf;
  assign lizzieLet10_6QError_Int_bufchan_r = (! lizzieLet10_6QError_Int_bufchan_buf[0]);
  assign lizzieLet10_6QError_Int_1_argbuf_d = (lizzieLet10_6QError_Int_bufchan_buf[0] ? lizzieLet10_6QError_Int_bufchan_buf :
                                               lizzieLet10_6QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet10_6QError_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet10_6QError_Int_1_argbuf_r && lizzieLet10_6QError_Int_bufchan_buf[0]))
        lizzieLet10_6QError_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet10_6QError_Int_1_argbuf_r) && (! lizzieLet10_6QError_Int_bufchan_buf[0])))
        lizzieLet10_6QError_Int_bufchan_buf <= lizzieLet10_6QError_Int_bufchan_d;
  
  /* dcon (Ty CTmain_map'_Int_Int,
      Dcon Lcall_main_map'_Int_Int3) : [(lizzieLet10_6QNode_Int,Pointer_CTmain_map'_Int_Int),
                                        (lizzieLet10_5QNode_Int_1,MyDTInt_Bool),
                                        (lizzieLet10_3QNode_Int_1,MyDTInt_Int),
                                        (q1acP_destruct,Pointer_QTree_Int),
                                        (q2acQ_destruct,Pointer_QTree_Int),
                                        (q3acR_destruct,Pointer_QTree_Int)] > (lizzieLet10_6QNode_Int_1lizzieLet10_5QNode_Int_1lizzieLet10_3QNode_Int_1q1acP_1q2acQ_1q3acR_1Lcall_main_map'_Int_Int3,CTmain_map'_Int_Int) */
  assign \lizzieLet10_6QNode_Int_1lizzieLet10_5QNode_Int_1lizzieLet10_3QNode_Int_1q1acP_1q2acQ_1q3acR_1Lcall_main_map'_Int_Int3_d  = \Lcall_main_map'_Int_Int3_dc ((& {lizzieLet10_6QNode_Int_d[0],
                                                                                                                                                                       lizzieLet10_5QNode_Int_1_d[0],
                                                                                                                                                                       lizzieLet10_3QNode_Int_1_d[0],
                                                                                                                                                                       q1acP_destruct_d[0],
                                                                                                                                                                       q2acQ_destruct_d[0],
                                                                                                                                                                       q3acR_destruct_d[0]}), lizzieLet10_6QNode_Int_d, lizzieLet10_5QNode_Int_1_d, lizzieLet10_3QNode_Int_1_d, q1acP_destruct_d, q2acQ_destruct_d, q3acR_destruct_d);
  assign {lizzieLet10_6QNode_Int_r,
          lizzieLet10_5QNode_Int_1_r,
          lizzieLet10_3QNode_Int_1_r,
          q1acP_destruct_r,
          q2acQ_destruct_r,
          q3acR_destruct_r} = {6 {(\lizzieLet10_6QNode_Int_1lizzieLet10_5QNode_Int_1lizzieLet10_3QNode_Int_1q1acP_1q2acQ_1q3acR_1Lcall_main_map'_Int_Int3_r  && \lizzieLet10_6QNode_Int_1lizzieLet10_5QNode_Int_1lizzieLet10_3QNode_Int_1q1acP_1q2acQ_1q3acR_1Lcall_main_map'_Int_Int3_d [0])}};
  
  /* buf (Ty CTmain_map'_Int_Int) : (lizzieLet10_6QNode_Int_1lizzieLet10_5QNode_Int_1lizzieLet10_3QNode_Int_1q1acP_1q2acQ_1q3acR_1Lcall_main_map'_Int_Int3,CTmain_map'_Int_Int) > (lizzieLet14_1_argbuf,CTmain_map'_Int_Int) */
  \CTmain_map'_Int_Int_t  \lizzieLet10_6QNode_Int_1lizzieLet10_5QNode_Int_1lizzieLet10_3QNode_Int_1q1acP_1q2acQ_1q3acR_1Lcall_main_map'_Int_Int3_bufchan_d ;
  logic \lizzieLet10_6QNode_Int_1lizzieLet10_5QNode_Int_1lizzieLet10_3QNode_Int_1q1acP_1q2acQ_1q3acR_1Lcall_main_map'_Int_Int3_bufchan_r ;
  assign \lizzieLet10_6QNode_Int_1lizzieLet10_5QNode_Int_1lizzieLet10_3QNode_Int_1q1acP_1q2acQ_1q3acR_1Lcall_main_map'_Int_Int3_r  = ((! \lizzieLet10_6QNode_Int_1lizzieLet10_5QNode_Int_1lizzieLet10_3QNode_Int_1q1acP_1q2acQ_1q3acR_1Lcall_main_map'_Int_Int3_bufchan_d [0]) || \lizzieLet10_6QNode_Int_1lizzieLet10_5QNode_Int_1lizzieLet10_3QNode_Int_1q1acP_1q2acQ_1q3acR_1Lcall_main_map'_Int_Int3_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet10_6QNode_Int_1lizzieLet10_5QNode_Int_1lizzieLet10_3QNode_Int_1q1acP_1q2acQ_1q3acR_1Lcall_main_map'_Int_Int3_bufchan_d  <= {67'd0,
                                                                                                                                            1'd0};
    else
      if (\lizzieLet10_6QNode_Int_1lizzieLet10_5QNode_Int_1lizzieLet10_3QNode_Int_1q1acP_1q2acQ_1q3acR_1Lcall_main_map'_Int_Int3_r )
        \lizzieLet10_6QNode_Int_1lizzieLet10_5QNode_Int_1lizzieLet10_3QNode_Int_1q1acP_1q2acQ_1q3acR_1Lcall_main_map'_Int_Int3_bufchan_d  <= \lizzieLet10_6QNode_Int_1lizzieLet10_5QNode_Int_1lizzieLet10_3QNode_Int_1q1acP_1q2acQ_1q3acR_1Lcall_main_map'_Int_Int3_d ;
  \CTmain_map'_Int_Int_t  \lizzieLet10_6QNode_Int_1lizzieLet10_5QNode_Int_1lizzieLet10_3QNode_Int_1q1acP_1q2acQ_1q3acR_1Lcall_main_map'_Int_Int3_bufchan_buf ;
  assign \lizzieLet10_6QNode_Int_1lizzieLet10_5QNode_Int_1lizzieLet10_3QNode_Int_1q1acP_1q2acQ_1q3acR_1Lcall_main_map'_Int_Int3_bufchan_r  = (! \lizzieLet10_6QNode_Int_1lizzieLet10_5QNode_Int_1lizzieLet10_3QNode_Int_1q1acP_1q2acQ_1q3acR_1Lcall_main_map'_Int_Int3_bufchan_buf [0]);
  assign lizzieLet14_1_argbuf_d = (\lizzieLet10_6QNode_Int_1lizzieLet10_5QNode_Int_1lizzieLet10_3QNode_Int_1q1acP_1q2acQ_1q3acR_1Lcall_main_map'_Int_Int3_bufchan_buf [0] ? \lizzieLet10_6QNode_Int_1lizzieLet10_5QNode_Int_1lizzieLet10_3QNode_Int_1q1acP_1q2acQ_1q3acR_1Lcall_main_map'_Int_Int3_bufchan_buf  :
                                   \lizzieLet10_6QNode_Int_1lizzieLet10_5QNode_Int_1lizzieLet10_3QNode_Int_1q1acP_1q2acQ_1q3acR_1Lcall_main_map'_Int_Int3_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet10_6QNode_Int_1lizzieLet10_5QNode_Int_1lizzieLet10_3QNode_Int_1q1acP_1q2acQ_1q3acR_1Lcall_main_map'_Int_Int3_bufchan_buf  <= {67'd0,
                                                                                                                                              1'd0};
    else
      if ((lizzieLet14_1_argbuf_r && \lizzieLet10_6QNode_Int_1lizzieLet10_5QNode_Int_1lizzieLet10_3QNode_Int_1q1acP_1q2acQ_1q3acR_1Lcall_main_map'_Int_Int3_bufchan_buf [0]))
        \lizzieLet10_6QNode_Int_1lizzieLet10_5QNode_Int_1lizzieLet10_3QNode_Int_1q1acP_1q2acQ_1q3acR_1Lcall_main_map'_Int_Int3_bufchan_buf  <= {67'd0,
                                                                                                                                                1'd0};
      else if (((! lizzieLet14_1_argbuf_r) && (! \lizzieLet10_6QNode_Int_1lizzieLet10_5QNode_Int_1lizzieLet10_3QNode_Int_1q1acP_1q2acQ_1q3acR_1Lcall_main_map'_Int_Int3_bufchan_buf [0])))
        \lizzieLet10_6QNode_Int_1lizzieLet10_5QNode_Int_1lizzieLet10_3QNode_Int_1q1acP_1q2acQ_1q3acR_1Lcall_main_map'_Int_Int3_bufchan_buf  <= \lizzieLet10_6QNode_Int_1lizzieLet10_5QNode_Int_1lizzieLet10_3QNode_Int_1q1acP_1q2acQ_1q3acR_1Lcall_main_map'_Int_Int3_bufchan_d ;
  
  /* buf (Ty Pointer_CTmain_map'_Int_Int) : (lizzieLet10_6QNone_Int,Pointer_CTmain_map'_Int_Int) > (lizzieLet10_6QNone_Int_1_argbuf,Pointer_CTmain_map'_Int_Int) */
  \Pointer_CTmain_map'_Int_Int_t  lizzieLet10_6QNone_Int_bufchan_d;
  logic lizzieLet10_6QNone_Int_bufchan_r;
  assign lizzieLet10_6QNone_Int_r = ((! lizzieLet10_6QNone_Int_bufchan_d[0]) || lizzieLet10_6QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet10_6QNone_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet10_6QNone_Int_r)
        lizzieLet10_6QNone_Int_bufchan_d <= lizzieLet10_6QNone_Int_d;
  \Pointer_CTmain_map'_Int_Int_t  lizzieLet10_6QNone_Int_bufchan_buf;
  assign lizzieLet10_6QNone_Int_bufchan_r = (! lizzieLet10_6QNone_Int_bufchan_buf[0]);
  assign lizzieLet10_6QNone_Int_1_argbuf_d = (lizzieLet10_6QNone_Int_bufchan_buf[0] ? lizzieLet10_6QNone_Int_bufchan_buf :
                                              lizzieLet10_6QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet10_6QNone_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet10_6QNone_Int_1_argbuf_r && lizzieLet10_6QNone_Int_bufchan_buf[0]))
        lizzieLet10_6QNone_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet10_6QNone_Int_1_argbuf_r) && (! lizzieLet10_6QNone_Int_bufchan_buf[0])))
        lizzieLet10_6QNone_Int_bufchan_buf <= lizzieLet10_6QNone_Int_bufchan_d;
  
  /* destruct (Ty QTree_Int,
          Dcon QNode_Int) : (lizzieLet16_1_1QNode_Int,QTree_Int) > [(q1acY_destruct,Pointer_QTree_Int),
                                                                    (q2acZ_destruct,Pointer_QTree_Int),
                                                                    (q3ad0_destruct,Pointer_QTree_Int),
                                                                    (q4ad1_destruct,Pointer_QTree_Int)] */
  logic [3:0] lizzieLet16_1_1QNode_Int_emitted;
  logic [3:0] lizzieLet16_1_1QNode_Int_done;
  assign q1acY_destruct_d = {lizzieLet16_1_1QNode_Int_d[18:3],
                             (lizzieLet16_1_1QNode_Int_d[0] && (! lizzieLet16_1_1QNode_Int_emitted[0]))};
  assign q2acZ_destruct_d = {lizzieLet16_1_1QNode_Int_d[34:19],
                             (lizzieLet16_1_1QNode_Int_d[0] && (! lizzieLet16_1_1QNode_Int_emitted[1]))};
  assign q3ad0_destruct_d = {lizzieLet16_1_1QNode_Int_d[50:35],
                             (lizzieLet16_1_1QNode_Int_d[0] && (! lizzieLet16_1_1QNode_Int_emitted[2]))};
  assign q4ad1_destruct_d = {lizzieLet16_1_1QNode_Int_d[66:51],
                             (lizzieLet16_1_1QNode_Int_d[0] && (! lizzieLet16_1_1QNode_Int_emitted[3]))};
  assign lizzieLet16_1_1QNode_Int_done = (lizzieLet16_1_1QNode_Int_emitted | ({q4ad1_destruct_d[0],
                                                                               q3ad0_destruct_d[0],
                                                                               q2acZ_destruct_d[0],
                                                                               q1acY_destruct_d[0]} & {q4ad1_destruct_r,
                                                                                                       q3ad0_destruct_r,
                                                                                                       q2acZ_destruct_r,
                                                                                                       q1acY_destruct_r}));
  assign lizzieLet16_1_1QNode_Int_r = (& lizzieLet16_1_1QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet16_1_1QNode_Int_emitted <= 4'd0;
    else
      lizzieLet16_1_1QNode_Int_emitted <= (lizzieLet16_1_1QNode_Int_r ? 4'd0 :
                                           lizzieLet16_1_1QNode_Int_done);
  
  /* destruct (Ty QTree_Int,
          Dcon QVal_Int) : (lizzieLet16_1_1QVal_Int,QTree_Int) > [(vacX_destruct,Int)] */
  assign vacX_destruct_d = {lizzieLet16_1_1QVal_Int_d[34:3],
                            lizzieLet16_1_1QVal_Int_d[0]};
  assign lizzieLet16_1_1QVal_Int_r = vacX_destruct_r;
  
  /* demux (Ty QTree_Int,
       Ty QTree_Int) : (lizzieLet16_1_2,QTree_Int) (lizzieLet16_1_1,QTree_Int) > [(_26,QTree_Int),
                                                                                  (lizzieLet16_1_1QVal_Int,QTree_Int),
                                                                                  (lizzieLet16_1_1QNode_Int,QTree_Int),
                                                                                  (_25,QTree_Int)] */
  logic [3:0] lizzieLet16_1_1_onehotd;
  always_comb
    if ((lizzieLet16_1_2_d[0] && lizzieLet16_1_1_d[0]))
      unique case (lizzieLet16_1_2_d[2:1])
        2'd0: lizzieLet16_1_1_onehotd = 4'd1;
        2'd1: lizzieLet16_1_1_onehotd = 4'd2;
        2'd2: lizzieLet16_1_1_onehotd = 4'd4;
        2'd3: lizzieLet16_1_1_onehotd = 4'd8;
        default: lizzieLet16_1_1_onehotd = 4'd0;
      endcase
    else lizzieLet16_1_1_onehotd = 4'd0;
  assign _26_d = {lizzieLet16_1_1_d[66:1],
                  lizzieLet16_1_1_onehotd[0]};
  assign lizzieLet16_1_1QVal_Int_d = {lizzieLet16_1_1_d[66:1],
                                      lizzieLet16_1_1_onehotd[1]};
  assign lizzieLet16_1_1QNode_Int_d = {lizzieLet16_1_1_d[66:1],
                                       lizzieLet16_1_1_onehotd[2]};
  assign _25_d = {lizzieLet16_1_1_d[66:1],
                  lizzieLet16_1_1_onehotd[3]};
  assign lizzieLet16_1_1_r = (| (lizzieLet16_1_1_onehotd & {_25_r,
                                                            lizzieLet16_1_1QNode_Int_r,
                                                            lizzieLet16_1_1QVal_Int_r,
                                                            _26_r}));
  assign lizzieLet16_1_2_r = lizzieLet16_1_1_r;
  
  /* demux (Ty QTree_Int,
       Ty MyDTInt_Int_Int) : (lizzieLet16_1_3,QTree_Int) (gacU_goMux_mux,MyDTInt_Int_Int) > [(_24,MyDTInt_Int_Int),
                                                                                             (lizzieLet16_1_3QVal_Int,MyDTInt_Int_Int),
                                                                                             (lizzieLet16_1_3QNode_Int,MyDTInt_Int_Int),
                                                                                             (_23,MyDTInt_Int_Int)] */
  logic [3:0] gacU_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet16_1_3_d[0] && gacU_goMux_mux_d[0]))
      unique case (lizzieLet16_1_3_d[2:1])
        2'd0: gacU_goMux_mux_onehotd = 4'd1;
        2'd1: gacU_goMux_mux_onehotd = 4'd2;
        2'd2: gacU_goMux_mux_onehotd = 4'd4;
        2'd3: gacU_goMux_mux_onehotd = 4'd8;
        default: gacU_goMux_mux_onehotd = 4'd0;
      endcase
    else gacU_goMux_mux_onehotd = 4'd0;
  assign _24_d = gacU_goMux_mux_onehotd[0];
  assign lizzieLet16_1_3QVal_Int_d = gacU_goMux_mux_onehotd[1];
  assign lizzieLet16_1_3QNode_Int_d = gacU_goMux_mux_onehotd[2];
  assign _23_d = gacU_goMux_mux_onehotd[3];
  assign gacU_goMux_mux_r = (| (gacU_goMux_mux_onehotd & {_23_r,
                                                          lizzieLet16_1_3QNode_Int_r,
                                                          lizzieLet16_1_3QVal_Int_r,
                                                          _24_r}));
  assign lizzieLet16_1_3_r = gacU_goMux_mux_r;
  
  /* fork (Ty MyDTInt_Int_Int) : (lizzieLet16_1_3QNode_Int,MyDTInt_Int_Int) > [(lizzieLet16_1_3QNode_Int_1,MyDTInt_Int_Int),
                                                                          (lizzieLet16_1_3QNode_Int_2,MyDTInt_Int_Int)] */
  logic [1:0] lizzieLet16_1_3QNode_Int_emitted;
  logic [1:0] lizzieLet16_1_3QNode_Int_done;
  assign lizzieLet16_1_3QNode_Int_1_d = (lizzieLet16_1_3QNode_Int_d[0] && (! lizzieLet16_1_3QNode_Int_emitted[0]));
  assign lizzieLet16_1_3QNode_Int_2_d = (lizzieLet16_1_3QNode_Int_d[0] && (! lizzieLet16_1_3QNode_Int_emitted[1]));
  assign lizzieLet16_1_3QNode_Int_done = (lizzieLet16_1_3QNode_Int_emitted | ({lizzieLet16_1_3QNode_Int_2_d[0],
                                                                               lizzieLet16_1_3QNode_Int_1_d[0]} & {lizzieLet16_1_3QNode_Int_2_r,
                                                                                                                   lizzieLet16_1_3QNode_Int_1_r}));
  assign lizzieLet16_1_3QNode_Int_r = (& lizzieLet16_1_3QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet16_1_3QNode_Int_emitted <= 2'd0;
    else
      lizzieLet16_1_3QNode_Int_emitted <= (lizzieLet16_1_3QNode_Int_r ? 2'd0 :
                                           lizzieLet16_1_3QNode_Int_done);
  
  /* buf (Ty MyDTInt_Int_Int) : (lizzieLet16_1_3QNode_Int_2,MyDTInt_Int_Int) > (lizzieLet16_1_3QNode_Int_2_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t lizzieLet16_1_3QNode_Int_2_bufchan_d;
  logic lizzieLet16_1_3QNode_Int_2_bufchan_r;
  assign lizzieLet16_1_3QNode_Int_2_r = ((! lizzieLet16_1_3QNode_Int_2_bufchan_d[0]) || lizzieLet16_1_3QNode_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet16_1_3QNode_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet16_1_3QNode_Int_2_r)
        lizzieLet16_1_3QNode_Int_2_bufchan_d <= lizzieLet16_1_3QNode_Int_2_d;
  MyDTInt_Int_Int_t lizzieLet16_1_3QNode_Int_2_bufchan_buf;
  assign lizzieLet16_1_3QNode_Int_2_bufchan_r = (! lizzieLet16_1_3QNode_Int_2_bufchan_buf[0]);
  assign lizzieLet16_1_3QNode_Int_2_argbuf_d = (lizzieLet16_1_3QNode_Int_2_bufchan_buf[0] ? lizzieLet16_1_3QNode_Int_2_bufchan_buf :
                                                lizzieLet16_1_3QNode_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet16_1_3QNode_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet16_1_3QNode_Int_2_argbuf_r && lizzieLet16_1_3QNode_Int_2_bufchan_buf[0]))
        lizzieLet16_1_3QNode_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet16_1_3QNode_Int_2_argbuf_r) && (! lizzieLet16_1_3QNode_Int_2_bufchan_buf[0])))
        lizzieLet16_1_3QNode_Int_2_bufchan_buf <= lizzieLet16_1_3QNode_Int_2_bufchan_d;
  
  /* buf (Ty MyDTInt_Int_Int) : (lizzieLet16_1_3QVal_Int,MyDTInt_Int_Int) > (lizzieLet16_1_3QVal_Int_1_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t lizzieLet16_1_3QVal_Int_bufchan_d;
  logic lizzieLet16_1_3QVal_Int_bufchan_r;
  assign lizzieLet16_1_3QVal_Int_r = ((! lizzieLet16_1_3QVal_Int_bufchan_d[0]) || lizzieLet16_1_3QVal_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet16_1_3QVal_Int_bufchan_d <= 1'd0;
    else
      if (lizzieLet16_1_3QVal_Int_r)
        lizzieLet16_1_3QVal_Int_bufchan_d <= lizzieLet16_1_3QVal_Int_d;
  MyDTInt_Int_Int_t lizzieLet16_1_3QVal_Int_bufchan_buf;
  assign lizzieLet16_1_3QVal_Int_bufchan_r = (! lizzieLet16_1_3QVal_Int_bufchan_buf[0]);
  assign lizzieLet16_1_3QVal_Int_1_argbuf_d = (lizzieLet16_1_3QVal_Int_bufchan_buf[0] ? lizzieLet16_1_3QVal_Int_bufchan_buf :
                                               lizzieLet16_1_3QVal_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet16_1_3QVal_Int_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet16_1_3QVal_Int_1_argbuf_r && lizzieLet16_1_3QVal_Int_bufchan_buf[0]))
        lizzieLet16_1_3QVal_Int_bufchan_buf <= 1'd0;
      else if (((! lizzieLet16_1_3QVal_Int_1_argbuf_r) && (! lizzieLet16_1_3QVal_Int_bufchan_buf[0])))
        lizzieLet16_1_3QVal_Int_bufchan_buf <= lizzieLet16_1_3QVal_Int_bufchan_d;
  
  /* dcon (Ty TupMyDTInt_Int_Int___Int___Int,
      Dcon TupMyDTInt_Int_Int___Int___Int) : [(lizzieLet16_1_3QVal_Int_1_argbuf,MyDTInt_Int_Int),
                                              (lizzieLet16_1_7QVal_Int_1_argbuf,Int),
                                              (vacX_1_argbuf,Int)] > (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1,TupMyDTInt_Int_Int___Int___Int) */
  assign applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_d = TupMyDTInt_Int_Int___Int___Int_dc((& {lizzieLet16_1_3QVal_Int_1_argbuf_d[0],
                                                                                                        lizzieLet16_1_7QVal_Int_1_argbuf_d[0],
                                                                                                        vacX_1_argbuf_d[0]}), lizzieLet16_1_3QVal_Int_1_argbuf_d, lizzieLet16_1_7QVal_Int_1_argbuf_d, vacX_1_argbuf_d);
  assign {lizzieLet16_1_3QVal_Int_1_argbuf_r,
          lizzieLet16_1_7QVal_Int_1_argbuf_r,
          vacX_1_argbuf_r} = {3 {(applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_r && applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_d[0])}};
  
  /* demux (Ty QTree_Int,
       Ty Go) : (lizzieLet16_1_4,QTree_Int) (go_14_goMux_data,Go) > [(lizzieLet16_1_4QNone_Int,Go),
                                                                     (lizzieLet16_1_4QVal_Int,Go),
                                                                     (lizzieLet16_1_4QNode_Int,Go),
                                                                     (lizzieLet16_1_4QError_Int,Go)] */
  logic [3:0] go_14_goMux_data_onehotd;
  always_comb
    if ((lizzieLet16_1_4_d[0] && go_14_goMux_data_d[0]))
      unique case (lizzieLet16_1_4_d[2:1])
        2'd0: go_14_goMux_data_onehotd = 4'd1;
        2'd1: go_14_goMux_data_onehotd = 4'd2;
        2'd2: go_14_goMux_data_onehotd = 4'd4;
        2'd3: go_14_goMux_data_onehotd = 4'd8;
        default: go_14_goMux_data_onehotd = 4'd0;
      endcase
    else go_14_goMux_data_onehotd = 4'd0;
  assign lizzieLet16_1_4QNone_Int_d = go_14_goMux_data_onehotd[0];
  assign lizzieLet16_1_4QVal_Int_d = go_14_goMux_data_onehotd[1];
  assign lizzieLet16_1_4QNode_Int_d = go_14_goMux_data_onehotd[2];
  assign lizzieLet16_1_4QError_Int_d = go_14_goMux_data_onehotd[3];
  assign go_14_goMux_data_r = (| (go_14_goMux_data_onehotd & {lizzieLet16_1_4QError_Int_r,
                                                              lizzieLet16_1_4QNode_Int_r,
                                                              lizzieLet16_1_4QVal_Int_r,
                                                              lizzieLet16_1_4QNone_Int_r}));
  assign lizzieLet16_1_4_r = go_14_goMux_data_r;
  
  /* fork (Ty Go) : (lizzieLet16_1_4QError_Int,Go) > [(lizzieLet16_1_4QError_Int_1,Go),
                                                 (lizzieLet16_1_4QError_Int_2,Go)] */
  logic [1:0] lizzieLet16_1_4QError_Int_emitted;
  logic [1:0] lizzieLet16_1_4QError_Int_done;
  assign lizzieLet16_1_4QError_Int_1_d = (lizzieLet16_1_4QError_Int_d[0] && (! lizzieLet16_1_4QError_Int_emitted[0]));
  assign lizzieLet16_1_4QError_Int_2_d = (lizzieLet16_1_4QError_Int_d[0] && (! lizzieLet16_1_4QError_Int_emitted[1]));
  assign lizzieLet16_1_4QError_Int_done = (lizzieLet16_1_4QError_Int_emitted | ({lizzieLet16_1_4QError_Int_2_d[0],
                                                                                 lizzieLet16_1_4QError_Int_1_d[0]} & {lizzieLet16_1_4QError_Int_2_r,
                                                                                                                      lizzieLet16_1_4QError_Int_1_r}));
  assign lizzieLet16_1_4QError_Int_r = (& lizzieLet16_1_4QError_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet16_1_4QError_Int_emitted <= 2'd0;
    else
      lizzieLet16_1_4QError_Int_emitted <= (lizzieLet16_1_4QError_Int_r ? 2'd0 :
                                            lizzieLet16_1_4QError_Int_done);
  
  /* dcon (Ty QTree_Int,
      Dcon QError_Int) : [(lizzieLet16_1_4QError_Int_1,Go)] > (lizzieLet16_1_4QError_Int_1QError_Int,QTree_Int) */
  assign lizzieLet16_1_4QError_Int_1QError_Int_d = QError_Int_dc((& {lizzieLet16_1_4QError_Int_1_d[0]}), lizzieLet16_1_4QError_Int_1_d);
  assign {lizzieLet16_1_4QError_Int_1_r} = {1 {(lizzieLet16_1_4QError_Int_1QError_Int_r && lizzieLet16_1_4QError_Int_1QError_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (lizzieLet16_1_4QError_Int_1QError_Int,QTree_Int) > (lizzieLet21_1_argbuf,QTree_Int) */
  QTree_Int_t lizzieLet16_1_4QError_Int_1QError_Int_bufchan_d;
  logic lizzieLet16_1_4QError_Int_1QError_Int_bufchan_r;
  assign lizzieLet16_1_4QError_Int_1QError_Int_r = ((! lizzieLet16_1_4QError_Int_1QError_Int_bufchan_d[0]) || lizzieLet16_1_4QError_Int_1QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet16_1_4QError_Int_1QError_Int_bufchan_d <= {66'd0, 1'd0};
    else
      if (lizzieLet16_1_4QError_Int_1QError_Int_r)
        lizzieLet16_1_4QError_Int_1QError_Int_bufchan_d <= lizzieLet16_1_4QError_Int_1QError_Int_d;
  QTree_Int_t lizzieLet16_1_4QError_Int_1QError_Int_bufchan_buf;
  assign lizzieLet16_1_4QError_Int_1QError_Int_bufchan_r = (! lizzieLet16_1_4QError_Int_1QError_Int_bufchan_buf[0]);
  assign lizzieLet21_1_argbuf_d = (lizzieLet16_1_4QError_Int_1QError_Int_bufchan_buf[0] ? lizzieLet16_1_4QError_Int_1QError_Int_bufchan_buf :
                                   lizzieLet16_1_4QError_Int_1QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet16_1_4QError_Int_1QError_Int_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((lizzieLet21_1_argbuf_r && lizzieLet16_1_4QError_Int_1QError_Int_bufchan_buf[0]))
        lizzieLet16_1_4QError_Int_1QError_Int_bufchan_buf <= {66'd0, 1'd0};
      else if (((! lizzieLet21_1_argbuf_r) && (! lizzieLet16_1_4QError_Int_1QError_Int_bufchan_buf[0])))
        lizzieLet16_1_4QError_Int_1QError_Int_bufchan_buf <= lizzieLet16_1_4QError_Int_1QError_Int_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet16_1_4QError_Int_2,Go) > (lizzieLet16_1_4QError_Int_2_argbuf,Go) */
  Go_t lizzieLet16_1_4QError_Int_2_bufchan_d;
  logic lizzieLet16_1_4QError_Int_2_bufchan_r;
  assign lizzieLet16_1_4QError_Int_2_r = ((! lizzieLet16_1_4QError_Int_2_bufchan_d[0]) || lizzieLet16_1_4QError_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet16_1_4QError_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet16_1_4QError_Int_2_r)
        lizzieLet16_1_4QError_Int_2_bufchan_d <= lizzieLet16_1_4QError_Int_2_d;
  Go_t lizzieLet16_1_4QError_Int_2_bufchan_buf;
  assign lizzieLet16_1_4QError_Int_2_bufchan_r = (! lizzieLet16_1_4QError_Int_2_bufchan_buf[0]);
  assign lizzieLet16_1_4QError_Int_2_argbuf_d = (lizzieLet16_1_4QError_Int_2_bufchan_buf[0] ? lizzieLet16_1_4QError_Int_2_bufchan_buf :
                                                 lizzieLet16_1_4QError_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet16_1_4QError_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet16_1_4QError_Int_2_argbuf_r && lizzieLet16_1_4QError_Int_2_bufchan_buf[0]))
        lizzieLet16_1_4QError_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet16_1_4QError_Int_2_argbuf_r) && (! lizzieLet16_1_4QError_Int_2_bufchan_buf[0])))
        lizzieLet16_1_4QError_Int_2_bufchan_buf <= lizzieLet16_1_4QError_Int_2_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet16_1_4QNode_Int,Go) > (lizzieLet16_1_4QNode_Int_1_argbuf,Go) */
  Go_t lizzieLet16_1_4QNode_Int_bufchan_d;
  logic lizzieLet16_1_4QNode_Int_bufchan_r;
  assign lizzieLet16_1_4QNode_Int_r = ((! lizzieLet16_1_4QNode_Int_bufchan_d[0]) || lizzieLet16_1_4QNode_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet16_1_4QNode_Int_bufchan_d <= 1'd0;
    else
      if (lizzieLet16_1_4QNode_Int_r)
        lizzieLet16_1_4QNode_Int_bufchan_d <= lizzieLet16_1_4QNode_Int_d;
  Go_t lizzieLet16_1_4QNode_Int_bufchan_buf;
  assign lizzieLet16_1_4QNode_Int_bufchan_r = (! lizzieLet16_1_4QNode_Int_bufchan_buf[0]);
  assign lizzieLet16_1_4QNode_Int_1_argbuf_d = (lizzieLet16_1_4QNode_Int_bufchan_buf[0] ? lizzieLet16_1_4QNode_Int_bufchan_buf :
                                                lizzieLet16_1_4QNode_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet16_1_4QNode_Int_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet16_1_4QNode_Int_1_argbuf_r && lizzieLet16_1_4QNode_Int_bufchan_buf[0]))
        lizzieLet16_1_4QNode_Int_bufchan_buf <= 1'd0;
      else if (((! lizzieLet16_1_4QNode_Int_1_argbuf_r) && (! lizzieLet16_1_4QNode_Int_bufchan_buf[0])))
        lizzieLet16_1_4QNode_Int_bufchan_buf <= lizzieLet16_1_4QNode_Int_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet16_1_4QNone_Int,Go) > [(lizzieLet16_1_4QNone_Int_1,Go),
                                                (lizzieLet16_1_4QNone_Int_2,Go)] */
  logic [1:0] lizzieLet16_1_4QNone_Int_emitted;
  logic [1:0] lizzieLet16_1_4QNone_Int_done;
  assign lizzieLet16_1_4QNone_Int_1_d = (lizzieLet16_1_4QNone_Int_d[0] && (! lizzieLet16_1_4QNone_Int_emitted[0]));
  assign lizzieLet16_1_4QNone_Int_2_d = (lizzieLet16_1_4QNone_Int_d[0] && (! lizzieLet16_1_4QNone_Int_emitted[1]));
  assign lizzieLet16_1_4QNone_Int_done = (lizzieLet16_1_4QNone_Int_emitted | ({lizzieLet16_1_4QNone_Int_2_d[0],
                                                                               lizzieLet16_1_4QNone_Int_1_d[0]} & {lizzieLet16_1_4QNone_Int_2_r,
                                                                                                                   lizzieLet16_1_4QNone_Int_1_r}));
  assign lizzieLet16_1_4QNone_Int_r = (& lizzieLet16_1_4QNone_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet16_1_4QNone_Int_emitted <= 2'd0;
    else
      lizzieLet16_1_4QNone_Int_emitted <= (lizzieLet16_1_4QNone_Int_r ? 2'd0 :
                                           lizzieLet16_1_4QNone_Int_done);
  
  /* dcon (Ty QTree_Int,
      Dcon QNone_Int) : [(lizzieLet16_1_4QNone_Int_1,Go)] > (lizzieLet16_1_4QNone_Int_1QNone_Int,QTree_Int) */
  assign lizzieLet16_1_4QNone_Int_1QNone_Int_d = QNone_Int_dc((& {lizzieLet16_1_4QNone_Int_1_d[0]}), lizzieLet16_1_4QNone_Int_1_d);
  assign {lizzieLet16_1_4QNone_Int_1_r} = {1 {(lizzieLet16_1_4QNone_Int_1QNone_Int_r && lizzieLet16_1_4QNone_Int_1QNone_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (lizzieLet16_1_4QNone_Int_1QNone_Int,QTree_Int) > (lizzieLet17_1_1_argbuf,QTree_Int) */
  QTree_Int_t lizzieLet16_1_4QNone_Int_1QNone_Int_bufchan_d;
  logic lizzieLet16_1_4QNone_Int_1QNone_Int_bufchan_r;
  assign lizzieLet16_1_4QNone_Int_1QNone_Int_r = ((! lizzieLet16_1_4QNone_Int_1QNone_Int_bufchan_d[0]) || lizzieLet16_1_4QNone_Int_1QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet16_1_4QNone_Int_1QNone_Int_bufchan_d <= {66'd0, 1'd0};
    else
      if (lizzieLet16_1_4QNone_Int_1QNone_Int_r)
        lizzieLet16_1_4QNone_Int_1QNone_Int_bufchan_d <= lizzieLet16_1_4QNone_Int_1QNone_Int_d;
  QTree_Int_t lizzieLet16_1_4QNone_Int_1QNone_Int_bufchan_buf;
  assign lizzieLet16_1_4QNone_Int_1QNone_Int_bufchan_r = (! lizzieLet16_1_4QNone_Int_1QNone_Int_bufchan_buf[0]);
  assign lizzieLet17_1_1_argbuf_d = (lizzieLet16_1_4QNone_Int_1QNone_Int_bufchan_buf[0] ? lizzieLet16_1_4QNone_Int_1QNone_Int_bufchan_buf :
                                     lizzieLet16_1_4QNone_Int_1QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet16_1_4QNone_Int_1QNone_Int_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((lizzieLet17_1_1_argbuf_r && lizzieLet16_1_4QNone_Int_1QNone_Int_bufchan_buf[0]))
        lizzieLet16_1_4QNone_Int_1QNone_Int_bufchan_buf <= {66'd0, 1'd0};
      else if (((! lizzieLet17_1_1_argbuf_r) && (! lizzieLet16_1_4QNone_Int_1QNone_Int_bufchan_buf[0])))
        lizzieLet16_1_4QNone_Int_1QNone_Int_bufchan_buf <= lizzieLet16_1_4QNone_Int_1QNone_Int_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet16_1_4QNone_Int_2,Go) > (lizzieLet16_1_4QNone_Int_2_argbuf,Go) */
  Go_t lizzieLet16_1_4QNone_Int_2_bufchan_d;
  logic lizzieLet16_1_4QNone_Int_2_bufchan_r;
  assign lizzieLet16_1_4QNone_Int_2_r = ((! lizzieLet16_1_4QNone_Int_2_bufchan_d[0]) || lizzieLet16_1_4QNone_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet16_1_4QNone_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet16_1_4QNone_Int_2_r)
        lizzieLet16_1_4QNone_Int_2_bufchan_d <= lizzieLet16_1_4QNone_Int_2_d;
  Go_t lizzieLet16_1_4QNone_Int_2_bufchan_buf;
  assign lizzieLet16_1_4QNone_Int_2_bufchan_r = (! lizzieLet16_1_4QNone_Int_2_bufchan_buf[0]);
  assign lizzieLet16_1_4QNone_Int_2_argbuf_d = (lizzieLet16_1_4QNone_Int_2_bufchan_buf[0] ? lizzieLet16_1_4QNone_Int_2_bufchan_buf :
                                                lizzieLet16_1_4QNone_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet16_1_4QNone_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet16_1_4QNone_Int_2_argbuf_r && lizzieLet16_1_4QNone_Int_2_bufchan_buf[0]))
        lizzieLet16_1_4QNone_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet16_1_4QNone_Int_2_argbuf_r) && (! lizzieLet16_1_4QNone_Int_2_bufchan_buf[0])))
        lizzieLet16_1_4QNone_Int_2_bufchan_buf <= lizzieLet16_1_4QNone_Int_2_bufchan_d;
  
  /* mergectrl (Ty C5,Ty Go) : [(lizzieLet16_1_4QNone_Int_2_argbuf,Go),
                           (lizzieLet39_3Lcall_map''_map''_Int_Int_Int0_1_argbuf,Go),
                           (es_0_5_1MyFalse_1_argbuf,Go),
                           (es_0_5_1MyTrue_2_argbuf,Go),
                           (lizzieLet16_1_4QError_Int_2_argbuf,Go)] > (go_21_goMux_choice,C5) (go_21_goMux_data,Go) */
  logic [4:0] lizzieLet16_1_4QNone_Int_2_argbuf_select_d;
  assign lizzieLet16_1_4QNone_Int_2_argbuf_select_d = ((| lizzieLet16_1_4QNone_Int_2_argbuf_select_q) ? lizzieLet16_1_4QNone_Int_2_argbuf_select_q :
                                                       (lizzieLet16_1_4QNone_Int_2_argbuf_d[0] ? 5'd1 :
                                                        (\lizzieLet39_3Lcall_map''_map''_Int_Int_Int0_1_argbuf_d [0] ? 5'd2 :
                                                         (es_0_5_1MyFalse_1_argbuf_d[0] ? 5'd4 :
                                                          (es_0_5_1MyTrue_2_argbuf_d[0] ? 5'd8 :
                                                           (lizzieLet16_1_4QError_Int_2_argbuf_d[0] ? 5'd16 :
                                                            5'd0))))));
  logic [4:0] lizzieLet16_1_4QNone_Int_2_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet16_1_4QNone_Int_2_argbuf_select_q <= 5'd0;
    else
      lizzieLet16_1_4QNone_Int_2_argbuf_select_q <= (lizzieLet16_1_4QNone_Int_2_argbuf_done ? 5'd0 :
                                                     lizzieLet16_1_4QNone_Int_2_argbuf_select_d);
  logic [1:0] lizzieLet16_1_4QNone_Int_2_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet16_1_4QNone_Int_2_argbuf_emit_q <= 2'd0;
    else
      lizzieLet16_1_4QNone_Int_2_argbuf_emit_q <= (lizzieLet16_1_4QNone_Int_2_argbuf_done ? 2'd0 :
                                                   lizzieLet16_1_4QNone_Int_2_argbuf_emit_d);
  logic [1:0] lizzieLet16_1_4QNone_Int_2_argbuf_emit_d;
  assign lizzieLet16_1_4QNone_Int_2_argbuf_emit_d = (lizzieLet16_1_4QNone_Int_2_argbuf_emit_q | ({go_21_goMux_choice_d[0],
                                                                                                  go_21_goMux_data_d[0]} & {go_21_goMux_choice_r,
                                                                                                                            go_21_goMux_data_r}));
  logic lizzieLet16_1_4QNone_Int_2_argbuf_done;
  assign lizzieLet16_1_4QNone_Int_2_argbuf_done = (& lizzieLet16_1_4QNone_Int_2_argbuf_emit_d);
  assign {lizzieLet16_1_4QError_Int_2_argbuf_r,
          es_0_5_1MyTrue_2_argbuf_r,
          es_0_5_1MyFalse_1_argbuf_r,
          \lizzieLet39_3Lcall_map''_map''_Int_Int_Int0_1_argbuf_r ,
          lizzieLet16_1_4QNone_Int_2_argbuf_r} = (lizzieLet16_1_4QNone_Int_2_argbuf_done ? lizzieLet16_1_4QNone_Int_2_argbuf_select_d :
                                                  5'd0);
  assign go_21_goMux_data_d = ((lizzieLet16_1_4QNone_Int_2_argbuf_select_d[0] && (! lizzieLet16_1_4QNone_Int_2_argbuf_emit_q[0])) ? lizzieLet16_1_4QNone_Int_2_argbuf_d :
                               ((lizzieLet16_1_4QNone_Int_2_argbuf_select_d[1] && (! lizzieLet16_1_4QNone_Int_2_argbuf_emit_q[0])) ? \lizzieLet39_3Lcall_map''_map''_Int_Int_Int0_1_argbuf_d  :
                                ((lizzieLet16_1_4QNone_Int_2_argbuf_select_d[2] && (! lizzieLet16_1_4QNone_Int_2_argbuf_emit_q[0])) ? es_0_5_1MyFalse_1_argbuf_d :
                                 ((lizzieLet16_1_4QNone_Int_2_argbuf_select_d[3] && (! lizzieLet16_1_4QNone_Int_2_argbuf_emit_q[0])) ? es_0_5_1MyTrue_2_argbuf_d :
                                  ((lizzieLet16_1_4QNone_Int_2_argbuf_select_d[4] && (! lizzieLet16_1_4QNone_Int_2_argbuf_emit_q[0])) ? lizzieLet16_1_4QError_Int_2_argbuf_d :
                                   1'd0)))));
  assign go_21_goMux_choice_d = ((lizzieLet16_1_4QNone_Int_2_argbuf_select_d[0] && (! lizzieLet16_1_4QNone_Int_2_argbuf_emit_q[1])) ? C1_5_dc(1'd1) :
                                 ((lizzieLet16_1_4QNone_Int_2_argbuf_select_d[1] && (! lizzieLet16_1_4QNone_Int_2_argbuf_emit_q[1])) ? C2_5_dc(1'd1) :
                                  ((lizzieLet16_1_4QNone_Int_2_argbuf_select_d[2] && (! lizzieLet16_1_4QNone_Int_2_argbuf_emit_q[1])) ? C3_5_dc(1'd1) :
                                   ((lizzieLet16_1_4QNone_Int_2_argbuf_select_d[3] && (! lizzieLet16_1_4QNone_Int_2_argbuf_emit_q[1])) ? C4_5_dc(1'd1) :
                                    ((lizzieLet16_1_4QNone_Int_2_argbuf_select_d[4] && (! lizzieLet16_1_4QNone_Int_2_argbuf_emit_q[1])) ? C5_5_dc(1'd1) :
                                     {3'd0, 1'd0})))));
  
  /* fork (Ty Go) : (lizzieLet16_1_4QVal_Int,Go) > [(lizzieLet16_1_4QVal_Int_1,Go),
                                               (lizzieLet16_1_4QVal_Int_2,Go)] */
  logic [1:0] lizzieLet16_1_4QVal_Int_emitted;
  logic [1:0] lizzieLet16_1_4QVal_Int_done;
  assign lizzieLet16_1_4QVal_Int_1_d = (lizzieLet16_1_4QVal_Int_d[0] && (! lizzieLet16_1_4QVal_Int_emitted[0]));
  assign lizzieLet16_1_4QVal_Int_2_d = (lizzieLet16_1_4QVal_Int_d[0] && (! lizzieLet16_1_4QVal_Int_emitted[1]));
  assign lizzieLet16_1_4QVal_Int_done = (lizzieLet16_1_4QVal_Int_emitted | ({lizzieLet16_1_4QVal_Int_2_d[0],
                                                                             lizzieLet16_1_4QVal_Int_1_d[0]} & {lizzieLet16_1_4QVal_Int_2_r,
                                                                                                                lizzieLet16_1_4QVal_Int_1_r}));
  assign lizzieLet16_1_4QVal_Int_r = (& lizzieLet16_1_4QVal_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet16_1_4QVal_Int_emitted <= 2'd0;
    else
      lizzieLet16_1_4QVal_Int_emitted <= (lizzieLet16_1_4QVal_Int_r ? 2'd0 :
                                          lizzieLet16_1_4QVal_Int_done);
  
  /* buf (Ty Go) : (lizzieLet16_1_4QVal_Int_1,Go) > (lizzieLet16_1_4QVal_Int_1_argbuf,Go) */
  Go_t lizzieLet16_1_4QVal_Int_1_bufchan_d;
  logic lizzieLet16_1_4QVal_Int_1_bufchan_r;
  assign lizzieLet16_1_4QVal_Int_1_r = ((! lizzieLet16_1_4QVal_Int_1_bufchan_d[0]) || lizzieLet16_1_4QVal_Int_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet16_1_4QVal_Int_1_bufchan_d <= 1'd0;
    else
      if (lizzieLet16_1_4QVal_Int_1_r)
        lizzieLet16_1_4QVal_Int_1_bufchan_d <= lizzieLet16_1_4QVal_Int_1_d;
  Go_t lizzieLet16_1_4QVal_Int_1_bufchan_buf;
  assign lizzieLet16_1_4QVal_Int_1_bufchan_r = (! lizzieLet16_1_4QVal_Int_1_bufchan_buf[0]);
  assign lizzieLet16_1_4QVal_Int_1_argbuf_d = (lizzieLet16_1_4QVal_Int_1_bufchan_buf[0] ? lizzieLet16_1_4QVal_Int_1_bufchan_buf :
                                               lizzieLet16_1_4QVal_Int_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet16_1_4QVal_Int_1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet16_1_4QVal_Int_1_argbuf_r && lizzieLet16_1_4QVal_Int_1_bufchan_buf[0]))
        lizzieLet16_1_4QVal_Int_1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet16_1_4QVal_Int_1_argbuf_r) && (! lizzieLet16_1_4QVal_Int_1_bufchan_buf[0])))
        lizzieLet16_1_4QVal_Int_1_bufchan_buf <= lizzieLet16_1_4QVal_Int_1_bufchan_d;
  
  /* dcon (Ty TupGo___MyDTInt_Bool___Int,
      Dcon TupGo___MyDTInt_Bool___Int) : [(lizzieLet16_1_4QVal_Int_1_argbuf,Go),
                                          (lizzieLet16_1_5QVal_Int_1_argbuf,MyDTInt_Bool),
                                          (xacr_1_1_argbuf,Int)] > (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1,TupGo___MyDTInt_Bool___Int) */
  assign applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_d = TupGo___MyDTInt_Bool___Int_dc((& {lizzieLet16_1_4QVal_Int_1_argbuf_d[0],
                                                                                             lizzieLet16_1_5QVal_Int_1_argbuf_d[0],
                                                                                             xacr_1_1_argbuf_d[0]}), lizzieLet16_1_4QVal_Int_1_argbuf_d, lizzieLet16_1_5QVal_Int_1_argbuf_d, xacr_1_1_argbuf_d);
  assign {lizzieLet16_1_4QVal_Int_1_argbuf_r,
          lizzieLet16_1_5QVal_Int_1_argbuf_r,
          xacr_1_1_argbuf_r} = {3 {(applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_r && applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_d[0])}};
  
  /* demux (Ty QTree_Int,
       Ty MyDTInt_Bool) : (lizzieLet16_1_5,QTree_Int) (isZacT_goMux_mux,MyDTInt_Bool) > [(_22,MyDTInt_Bool),
                                                                                         (lizzieLet16_1_5QVal_Int,MyDTInt_Bool),
                                                                                         (lizzieLet16_1_5QNode_Int,MyDTInt_Bool),
                                                                                         (_21,MyDTInt_Bool)] */
  logic [3:0] isZacT_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet16_1_5_d[0] && isZacT_goMux_mux_d[0]))
      unique case (lizzieLet16_1_5_d[2:1])
        2'd0: isZacT_goMux_mux_onehotd = 4'd1;
        2'd1: isZacT_goMux_mux_onehotd = 4'd2;
        2'd2: isZacT_goMux_mux_onehotd = 4'd4;
        2'd3: isZacT_goMux_mux_onehotd = 4'd8;
        default: isZacT_goMux_mux_onehotd = 4'd0;
      endcase
    else isZacT_goMux_mux_onehotd = 4'd0;
  assign _22_d = isZacT_goMux_mux_onehotd[0];
  assign lizzieLet16_1_5QVal_Int_d = isZacT_goMux_mux_onehotd[1];
  assign lizzieLet16_1_5QNode_Int_d = isZacT_goMux_mux_onehotd[2];
  assign _21_d = isZacT_goMux_mux_onehotd[3];
  assign isZacT_goMux_mux_r = (| (isZacT_goMux_mux_onehotd & {_21_r,
                                                              lizzieLet16_1_5QNode_Int_r,
                                                              lizzieLet16_1_5QVal_Int_r,
                                                              _22_r}));
  assign lizzieLet16_1_5_r = isZacT_goMux_mux_r;
  
  /* fork (Ty MyDTInt_Bool) : (lizzieLet16_1_5QNode_Int,MyDTInt_Bool) > [(lizzieLet16_1_5QNode_Int_1,MyDTInt_Bool),
                                                                    (lizzieLet16_1_5QNode_Int_2,MyDTInt_Bool)] */
  logic [1:0] lizzieLet16_1_5QNode_Int_emitted;
  logic [1:0] lizzieLet16_1_5QNode_Int_done;
  assign lizzieLet16_1_5QNode_Int_1_d = (lizzieLet16_1_5QNode_Int_d[0] && (! lizzieLet16_1_5QNode_Int_emitted[0]));
  assign lizzieLet16_1_5QNode_Int_2_d = (lizzieLet16_1_5QNode_Int_d[0] && (! lizzieLet16_1_5QNode_Int_emitted[1]));
  assign lizzieLet16_1_5QNode_Int_done = (lizzieLet16_1_5QNode_Int_emitted | ({lizzieLet16_1_5QNode_Int_2_d[0],
                                                                               lizzieLet16_1_5QNode_Int_1_d[0]} & {lizzieLet16_1_5QNode_Int_2_r,
                                                                                                                   lizzieLet16_1_5QNode_Int_1_r}));
  assign lizzieLet16_1_5QNode_Int_r = (& lizzieLet16_1_5QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet16_1_5QNode_Int_emitted <= 2'd0;
    else
      lizzieLet16_1_5QNode_Int_emitted <= (lizzieLet16_1_5QNode_Int_r ? 2'd0 :
                                           lizzieLet16_1_5QNode_Int_done);
  
  /* buf (Ty MyDTInt_Bool) : (lizzieLet16_1_5QNode_Int_2,MyDTInt_Bool) > (lizzieLet16_1_5QNode_Int_2_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t lizzieLet16_1_5QNode_Int_2_bufchan_d;
  logic lizzieLet16_1_5QNode_Int_2_bufchan_r;
  assign lizzieLet16_1_5QNode_Int_2_r = ((! lizzieLet16_1_5QNode_Int_2_bufchan_d[0]) || lizzieLet16_1_5QNode_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet16_1_5QNode_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet16_1_5QNode_Int_2_r)
        lizzieLet16_1_5QNode_Int_2_bufchan_d <= lizzieLet16_1_5QNode_Int_2_d;
  MyDTInt_Bool_t lizzieLet16_1_5QNode_Int_2_bufchan_buf;
  assign lizzieLet16_1_5QNode_Int_2_bufchan_r = (! lizzieLet16_1_5QNode_Int_2_bufchan_buf[0]);
  assign lizzieLet16_1_5QNode_Int_2_argbuf_d = (lizzieLet16_1_5QNode_Int_2_bufchan_buf[0] ? lizzieLet16_1_5QNode_Int_2_bufchan_buf :
                                                lizzieLet16_1_5QNode_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet16_1_5QNode_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet16_1_5QNode_Int_2_argbuf_r && lizzieLet16_1_5QNode_Int_2_bufchan_buf[0]))
        lizzieLet16_1_5QNode_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet16_1_5QNode_Int_2_argbuf_r) && (! lizzieLet16_1_5QNode_Int_2_bufchan_buf[0])))
        lizzieLet16_1_5QNode_Int_2_bufchan_buf <= lizzieLet16_1_5QNode_Int_2_bufchan_d;
  
  /* buf (Ty MyDTInt_Bool) : (lizzieLet16_1_5QVal_Int,MyDTInt_Bool) > (lizzieLet16_1_5QVal_Int_1_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t lizzieLet16_1_5QVal_Int_bufchan_d;
  logic lizzieLet16_1_5QVal_Int_bufchan_r;
  assign lizzieLet16_1_5QVal_Int_r = ((! lizzieLet16_1_5QVal_Int_bufchan_d[0]) || lizzieLet16_1_5QVal_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet16_1_5QVal_Int_bufchan_d <= 1'd0;
    else
      if (lizzieLet16_1_5QVal_Int_r)
        lizzieLet16_1_5QVal_Int_bufchan_d <= lizzieLet16_1_5QVal_Int_d;
  MyDTInt_Bool_t lizzieLet16_1_5QVal_Int_bufchan_buf;
  assign lizzieLet16_1_5QVal_Int_bufchan_r = (! lizzieLet16_1_5QVal_Int_bufchan_buf[0]);
  assign lizzieLet16_1_5QVal_Int_1_argbuf_d = (lizzieLet16_1_5QVal_Int_bufchan_buf[0] ? lizzieLet16_1_5QVal_Int_bufchan_buf :
                                               lizzieLet16_1_5QVal_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet16_1_5QVal_Int_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet16_1_5QVal_Int_1_argbuf_r && lizzieLet16_1_5QVal_Int_bufchan_buf[0]))
        lizzieLet16_1_5QVal_Int_bufchan_buf <= 1'd0;
      else if (((! lizzieLet16_1_5QVal_Int_1_argbuf_r) && (! lizzieLet16_1_5QVal_Int_bufchan_buf[0])))
        lizzieLet16_1_5QVal_Int_bufchan_buf <= lizzieLet16_1_5QVal_Int_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_CTmap''_map''_Int_Int_Int) : (lizzieLet16_1_6,QTree_Int) (sc_0_3_goMux_mux,Pointer_CTmap''_map''_Int_Int_Int) > [(lizzieLet16_1_6QNone_Int,Pointer_CTmap''_map''_Int_Int_Int),
                                                                                                                                   (lizzieLet16_1_6QVal_Int,Pointer_CTmap''_map''_Int_Int_Int),
                                                                                                                                   (lizzieLet16_1_6QNode_Int,Pointer_CTmap''_map''_Int_Int_Int),
                                                                                                                                   (lizzieLet16_1_6QError_Int,Pointer_CTmap''_map''_Int_Int_Int)] */
  logic [3:0] sc_0_3_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet16_1_6_d[0] && sc_0_3_goMux_mux_d[0]))
      unique case (lizzieLet16_1_6_d[2:1])
        2'd0: sc_0_3_goMux_mux_onehotd = 4'd1;
        2'd1: sc_0_3_goMux_mux_onehotd = 4'd2;
        2'd2: sc_0_3_goMux_mux_onehotd = 4'd4;
        2'd3: sc_0_3_goMux_mux_onehotd = 4'd8;
        default: sc_0_3_goMux_mux_onehotd = 4'd0;
      endcase
    else sc_0_3_goMux_mux_onehotd = 4'd0;
  assign lizzieLet16_1_6QNone_Int_d = {sc_0_3_goMux_mux_d[16:1],
                                       sc_0_3_goMux_mux_onehotd[0]};
  assign lizzieLet16_1_6QVal_Int_d = {sc_0_3_goMux_mux_d[16:1],
                                      sc_0_3_goMux_mux_onehotd[1]};
  assign lizzieLet16_1_6QNode_Int_d = {sc_0_3_goMux_mux_d[16:1],
                                       sc_0_3_goMux_mux_onehotd[2]};
  assign lizzieLet16_1_6QError_Int_d = {sc_0_3_goMux_mux_d[16:1],
                                        sc_0_3_goMux_mux_onehotd[3]};
  assign sc_0_3_goMux_mux_r = (| (sc_0_3_goMux_mux_onehotd & {lizzieLet16_1_6QError_Int_r,
                                                              lizzieLet16_1_6QNode_Int_r,
                                                              lizzieLet16_1_6QVal_Int_r,
                                                              lizzieLet16_1_6QNone_Int_r}));
  assign lizzieLet16_1_6_r = sc_0_3_goMux_mux_r;
  
  /* buf (Ty Pointer_CTmap''_map''_Int_Int_Int) : (lizzieLet16_1_6QError_Int,Pointer_CTmap''_map''_Int_Int_Int) > (lizzieLet16_1_6QError_Int_1_argbuf,Pointer_CTmap''_map''_Int_Int_Int) */
  \Pointer_CTmap''_map''_Int_Int_Int_t  lizzieLet16_1_6QError_Int_bufchan_d;
  logic lizzieLet16_1_6QError_Int_bufchan_r;
  assign lizzieLet16_1_6QError_Int_r = ((! lizzieLet16_1_6QError_Int_bufchan_d[0]) || lizzieLet16_1_6QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet16_1_6QError_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet16_1_6QError_Int_r)
        lizzieLet16_1_6QError_Int_bufchan_d <= lizzieLet16_1_6QError_Int_d;
  \Pointer_CTmap''_map''_Int_Int_Int_t  lizzieLet16_1_6QError_Int_bufchan_buf;
  assign lizzieLet16_1_6QError_Int_bufchan_r = (! lizzieLet16_1_6QError_Int_bufchan_buf[0]);
  assign lizzieLet16_1_6QError_Int_1_argbuf_d = (lizzieLet16_1_6QError_Int_bufchan_buf[0] ? lizzieLet16_1_6QError_Int_bufchan_buf :
                                                 lizzieLet16_1_6QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet16_1_6QError_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet16_1_6QError_Int_1_argbuf_r && lizzieLet16_1_6QError_Int_bufchan_buf[0]))
        lizzieLet16_1_6QError_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet16_1_6QError_Int_1_argbuf_r) && (! lizzieLet16_1_6QError_Int_bufchan_buf[0])))
        lizzieLet16_1_6QError_Int_bufchan_buf <= lizzieLet16_1_6QError_Int_bufchan_d;
  
  /* dcon (Ty CTmap''_map''_Int_Int_Int,
      Dcon Lcall_map''_map''_Int_Int_Int3) : [(lizzieLet16_1_6QNode_Int,Pointer_CTmap''_map''_Int_Int_Int),
                                              (lizzieLet16_1_5QNode_Int_1,MyDTInt_Bool),
                                              (lizzieLet16_1_3QNode_Int_1,MyDTInt_Int_Int),
                                              (lizzieLet16_1_7QNode_Int_1,Int),
                                              (q1acY_destruct,Pointer_QTree_Int),
                                              (q2acZ_destruct,Pointer_QTree_Int),
                                              (q3ad0_destruct,Pointer_QTree_Int)] > (lizzieLet16_1_6QNode_Int_1lizzieLet16_1_5QNode_Int_1lizzieLet16_1_3QNode_Int_1lizzieLet16_1_7QNode_Int_1q1acY_1q2acZ_1q3ad0_1Lcall_map''_map''_Int_Int_Int3,CTmap''_map''_Int_Int_Int) */
  assign \lizzieLet16_1_6QNode_Int_1lizzieLet16_1_5QNode_Int_1lizzieLet16_1_3QNode_Int_1lizzieLet16_1_7QNode_Int_1q1acY_1q2acZ_1q3ad0_1Lcall_map''_map''_Int_Int_Int3_d  = \Lcall_map''_map''_Int_Int_Int3_dc ((& {lizzieLet16_1_6QNode_Int_d[0],
                                                                                                                                                                                                                   lizzieLet16_1_5QNode_Int_1_d[0],
                                                                                                                                                                                                                   lizzieLet16_1_3QNode_Int_1_d[0],
                                                                                                                                                                                                                   lizzieLet16_1_7QNode_Int_1_d[0],
                                                                                                                                                                                                                   q1acY_destruct_d[0],
                                                                                                                                                                                                                   q2acZ_destruct_d[0],
                                                                                                                                                                                                                   q3ad0_destruct_d[0]}), lizzieLet16_1_6QNode_Int_d, lizzieLet16_1_5QNode_Int_1_d, lizzieLet16_1_3QNode_Int_1_d, lizzieLet16_1_7QNode_Int_1_d, q1acY_destruct_d, q2acZ_destruct_d, q3ad0_destruct_d);
  assign {lizzieLet16_1_6QNode_Int_r,
          lizzieLet16_1_5QNode_Int_1_r,
          lizzieLet16_1_3QNode_Int_1_r,
          lizzieLet16_1_7QNode_Int_1_r,
          q1acY_destruct_r,
          q2acZ_destruct_r,
          q3ad0_destruct_r} = {7 {(\lizzieLet16_1_6QNode_Int_1lizzieLet16_1_5QNode_Int_1lizzieLet16_1_3QNode_Int_1lizzieLet16_1_7QNode_Int_1q1acY_1q2acZ_1q3ad0_1Lcall_map''_map''_Int_Int_Int3_r  && \lizzieLet16_1_6QNode_Int_1lizzieLet16_1_5QNode_Int_1lizzieLet16_1_3QNode_Int_1lizzieLet16_1_7QNode_Int_1q1acY_1q2acZ_1q3ad0_1Lcall_map''_map''_Int_Int_Int3_d [0])}};
  
  /* buf (Ty CTmap''_map''_Int_Int_Int) : (lizzieLet16_1_6QNode_Int_1lizzieLet16_1_5QNode_Int_1lizzieLet16_1_3QNode_Int_1lizzieLet16_1_7QNode_Int_1q1acY_1q2acZ_1q3ad0_1Lcall_map''_map''_Int_Int_Int3,CTmap''_map''_Int_Int_Int) > (lizzieLet20_1_argbuf,CTmap''_map''_Int_Int_Int) */
  \CTmap''_map''_Int_Int_Int_t  \lizzieLet16_1_6QNode_Int_1lizzieLet16_1_5QNode_Int_1lizzieLet16_1_3QNode_Int_1lizzieLet16_1_7QNode_Int_1q1acY_1q2acZ_1q3ad0_1Lcall_map''_map''_Int_Int_Int3_bufchan_d ;
  logic \lizzieLet16_1_6QNode_Int_1lizzieLet16_1_5QNode_Int_1lizzieLet16_1_3QNode_Int_1lizzieLet16_1_7QNode_Int_1q1acY_1q2acZ_1q3ad0_1Lcall_map''_map''_Int_Int_Int3_bufchan_r ;
  assign \lizzieLet16_1_6QNode_Int_1lizzieLet16_1_5QNode_Int_1lizzieLet16_1_3QNode_Int_1lizzieLet16_1_7QNode_Int_1q1acY_1q2acZ_1q3ad0_1Lcall_map''_map''_Int_Int_Int3_r  = ((! \lizzieLet16_1_6QNode_Int_1lizzieLet16_1_5QNode_Int_1lizzieLet16_1_3QNode_Int_1lizzieLet16_1_7QNode_Int_1q1acY_1q2acZ_1q3ad0_1Lcall_map''_map''_Int_Int_Int3_bufchan_d [0]) || \lizzieLet16_1_6QNode_Int_1lizzieLet16_1_5QNode_Int_1lizzieLet16_1_3QNode_Int_1lizzieLet16_1_7QNode_Int_1q1acY_1q2acZ_1q3ad0_1Lcall_map''_map''_Int_Int_Int3_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet16_1_6QNode_Int_1lizzieLet16_1_5QNode_Int_1lizzieLet16_1_3QNode_Int_1lizzieLet16_1_7QNode_Int_1q1acY_1q2acZ_1q3ad0_1Lcall_map''_map''_Int_Int_Int3_bufchan_d  <= {99'd0,
                                                                                                                                                                                  1'd0};
    else
      if (\lizzieLet16_1_6QNode_Int_1lizzieLet16_1_5QNode_Int_1lizzieLet16_1_3QNode_Int_1lizzieLet16_1_7QNode_Int_1q1acY_1q2acZ_1q3ad0_1Lcall_map''_map''_Int_Int_Int3_r )
        \lizzieLet16_1_6QNode_Int_1lizzieLet16_1_5QNode_Int_1lizzieLet16_1_3QNode_Int_1lizzieLet16_1_7QNode_Int_1q1acY_1q2acZ_1q3ad0_1Lcall_map''_map''_Int_Int_Int3_bufchan_d  <= \lizzieLet16_1_6QNode_Int_1lizzieLet16_1_5QNode_Int_1lizzieLet16_1_3QNode_Int_1lizzieLet16_1_7QNode_Int_1q1acY_1q2acZ_1q3ad0_1Lcall_map''_map''_Int_Int_Int3_d ;
  \CTmap''_map''_Int_Int_Int_t  \lizzieLet16_1_6QNode_Int_1lizzieLet16_1_5QNode_Int_1lizzieLet16_1_3QNode_Int_1lizzieLet16_1_7QNode_Int_1q1acY_1q2acZ_1q3ad0_1Lcall_map''_map''_Int_Int_Int3_bufchan_buf ;
  assign \lizzieLet16_1_6QNode_Int_1lizzieLet16_1_5QNode_Int_1lizzieLet16_1_3QNode_Int_1lizzieLet16_1_7QNode_Int_1q1acY_1q2acZ_1q3ad0_1Lcall_map''_map''_Int_Int_Int3_bufchan_r  = (! \lizzieLet16_1_6QNode_Int_1lizzieLet16_1_5QNode_Int_1lizzieLet16_1_3QNode_Int_1lizzieLet16_1_7QNode_Int_1q1acY_1q2acZ_1q3ad0_1Lcall_map''_map''_Int_Int_Int3_bufchan_buf [0]);
  assign lizzieLet20_1_argbuf_d = (\lizzieLet16_1_6QNode_Int_1lizzieLet16_1_5QNode_Int_1lizzieLet16_1_3QNode_Int_1lizzieLet16_1_7QNode_Int_1q1acY_1q2acZ_1q3ad0_1Lcall_map''_map''_Int_Int_Int3_bufchan_buf [0] ? \lizzieLet16_1_6QNode_Int_1lizzieLet16_1_5QNode_Int_1lizzieLet16_1_3QNode_Int_1lizzieLet16_1_7QNode_Int_1q1acY_1q2acZ_1q3ad0_1Lcall_map''_map''_Int_Int_Int3_bufchan_buf  :
                                   \lizzieLet16_1_6QNode_Int_1lizzieLet16_1_5QNode_Int_1lizzieLet16_1_3QNode_Int_1lizzieLet16_1_7QNode_Int_1q1acY_1q2acZ_1q3ad0_1Lcall_map''_map''_Int_Int_Int3_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet16_1_6QNode_Int_1lizzieLet16_1_5QNode_Int_1lizzieLet16_1_3QNode_Int_1lizzieLet16_1_7QNode_Int_1q1acY_1q2acZ_1q3ad0_1Lcall_map''_map''_Int_Int_Int3_bufchan_buf  <= {99'd0,
                                                                                                                                                                                    1'd0};
    else
      if ((lizzieLet20_1_argbuf_r && \lizzieLet16_1_6QNode_Int_1lizzieLet16_1_5QNode_Int_1lizzieLet16_1_3QNode_Int_1lizzieLet16_1_7QNode_Int_1q1acY_1q2acZ_1q3ad0_1Lcall_map''_map''_Int_Int_Int3_bufchan_buf [0]))
        \lizzieLet16_1_6QNode_Int_1lizzieLet16_1_5QNode_Int_1lizzieLet16_1_3QNode_Int_1lizzieLet16_1_7QNode_Int_1q1acY_1q2acZ_1q3ad0_1Lcall_map''_map''_Int_Int_Int3_bufchan_buf  <= {99'd0,
                                                                                                                                                                                      1'd0};
      else if (((! lizzieLet20_1_argbuf_r) && (! \lizzieLet16_1_6QNode_Int_1lizzieLet16_1_5QNode_Int_1lizzieLet16_1_3QNode_Int_1lizzieLet16_1_7QNode_Int_1q1acY_1q2acZ_1q3ad0_1Lcall_map''_map''_Int_Int_Int3_bufchan_buf [0])))
        \lizzieLet16_1_6QNode_Int_1lizzieLet16_1_5QNode_Int_1lizzieLet16_1_3QNode_Int_1lizzieLet16_1_7QNode_Int_1q1acY_1q2acZ_1q3ad0_1Lcall_map''_map''_Int_Int_Int3_bufchan_buf  <= \lizzieLet16_1_6QNode_Int_1lizzieLet16_1_5QNode_Int_1lizzieLet16_1_3QNode_Int_1lizzieLet16_1_7QNode_Int_1q1acY_1q2acZ_1q3ad0_1Lcall_map''_map''_Int_Int_Int3_bufchan_d ;
  
  /* buf (Ty Pointer_CTmap''_map''_Int_Int_Int) : (lizzieLet16_1_6QNone_Int,Pointer_CTmap''_map''_Int_Int_Int) > (lizzieLet16_1_6QNone_Int_1_argbuf,Pointer_CTmap''_map''_Int_Int_Int) */
  \Pointer_CTmap''_map''_Int_Int_Int_t  lizzieLet16_1_6QNone_Int_bufchan_d;
  logic lizzieLet16_1_6QNone_Int_bufchan_r;
  assign lizzieLet16_1_6QNone_Int_r = ((! lizzieLet16_1_6QNone_Int_bufchan_d[0]) || lizzieLet16_1_6QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet16_1_6QNone_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet16_1_6QNone_Int_r)
        lizzieLet16_1_6QNone_Int_bufchan_d <= lizzieLet16_1_6QNone_Int_d;
  \Pointer_CTmap''_map''_Int_Int_Int_t  lizzieLet16_1_6QNone_Int_bufchan_buf;
  assign lizzieLet16_1_6QNone_Int_bufchan_r = (! lizzieLet16_1_6QNone_Int_bufchan_buf[0]);
  assign lizzieLet16_1_6QNone_Int_1_argbuf_d = (lizzieLet16_1_6QNone_Int_bufchan_buf[0] ? lizzieLet16_1_6QNone_Int_bufchan_buf :
                                                lizzieLet16_1_6QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet16_1_6QNone_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet16_1_6QNone_Int_1_argbuf_r && lizzieLet16_1_6QNone_Int_bufchan_buf[0]))
        lizzieLet16_1_6QNone_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet16_1_6QNone_Int_1_argbuf_r) && (! lizzieLet16_1_6QNone_Int_bufchan_buf[0])))
        lizzieLet16_1_6QNone_Int_bufchan_buf <= lizzieLet16_1_6QNone_Int_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Int) : (lizzieLet16_1_7,QTree_Int) (v'acV_goMux_mux,Int) > [(_20,Int),
                                                                      (lizzieLet16_1_7QVal_Int,Int),
                                                                      (lizzieLet16_1_7QNode_Int,Int),
                                                                      (_19,Int)] */
  logic [3:0] \v'acV_goMux_mux_onehotd ;
  always_comb
    if ((lizzieLet16_1_7_d[0] && \v'acV_goMux_mux_d [0]))
      unique case (lizzieLet16_1_7_d[2:1])
        2'd0: \v'acV_goMux_mux_onehotd  = 4'd1;
        2'd1: \v'acV_goMux_mux_onehotd  = 4'd2;
        2'd2: \v'acV_goMux_mux_onehotd  = 4'd4;
        2'd3: \v'acV_goMux_mux_onehotd  = 4'd8;
        default: \v'acV_goMux_mux_onehotd  = 4'd0;
      endcase
    else \v'acV_goMux_mux_onehotd  = 4'd0;
  assign _20_d = {\v'acV_goMux_mux_d [32:1],
                  \v'acV_goMux_mux_onehotd [0]};
  assign lizzieLet16_1_7QVal_Int_d = {\v'acV_goMux_mux_d [32:1],
                                      \v'acV_goMux_mux_onehotd [1]};
  assign lizzieLet16_1_7QNode_Int_d = {\v'acV_goMux_mux_d [32:1],
                                       \v'acV_goMux_mux_onehotd [2]};
  assign _19_d = {\v'acV_goMux_mux_d [32:1],
                  \v'acV_goMux_mux_onehotd [3]};
  assign \v'acV_goMux_mux_r  = (| (\v'acV_goMux_mux_onehotd  & {_19_r,
                                                                lizzieLet16_1_7QNode_Int_r,
                                                                lizzieLet16_1_7QVal_Int_r,
                                                                _20_r}));
  assign lizzieLet16_1_7_r = \v'acV_goMux_mux_r ;
  
  /* fork (Ty Int) : (lizzieLet16_1_7QNode_Int,Int) > [(lizzieLet16_1_7QNode_Int_1,Int),
                                                  (lizzieLet16_1_7QNode_Int_2,Int)] */
  logic [1:0] lizzieLet16_1_7QNode_Int_emitted;
  logic [1:0] lizzieLet16_1_7QNode_Int_done;
  assign lizzieLet16_1_7QNode_Int_1_d = {lizzieLet16_1_7QNode_Int_d[32:1],
                                         (lizzieLet16_1_7QNode_Int_d[0] && (! lizzieLet16_1_7QNode_Int_emitted[0]))};
  assign lizzieLet16_1_7QNode_Int_2_d = {lizzieLet16_1_7QNode_Int_d[32:1],
                                         (lizzieLet16_1_7QNode_Int_d[0] && (! lizzieLet16_1_7QNode_Int_emitted[1]))};
  assign lizzieLet16_1_7QNode_Int_done = (lizzieLet16_1_7QNode_Int_emitted | ({lizzieLet16_1_7QNode_Int_2_d[0],
                                                                               lizzieLet16_1_7QNode_Int_1_d[0]} & {lizzieLet16_1_7QNode_Int_2_r,
                                                                                                                   lizzieLet16_1_7QNode_Int_1_r}));
  assign lizzieLet16_1_7QNode_Int_r = (& lizzieLet16_1_7QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet16_1_7QNode_Int_emitted <= 2'd0;
    else
      lizzieLet16_1_7QNode_Int_emitted <= (lizzieLet16_1_7QNode_Int_r ? 2'd0 :
                                           lizzieLet16_1_7QNode_Int_done);
  
  /* buf (Ty Int) : (lizzieLet16_1_7QNode_Int_2,Int) > (lizzieLet16_1_7QNode_Int_2_argbuf,Int) */
  Int_t lizzieLet16_1_7QNode_Int_2_bufchan_d;
  logic lizzieLet16_1_7QNode_Int_2_bufchan_r;
  assign lizzieLet16_1_7QNode_Int_2_r = ((! lizzieLet16_1_7QNode_Int_2_bufchan_d[0]) || lizzieLet16_1_7QNode_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet16_1_7QNode_Int_2_bufchan_d <= {32'd0, 1'd0};
    else
      if (lizzieLet16_1_7QNode_Int_2_r)
        lizzieLet16_1_7QNode_Int_2_bufchan_d <= lizzieLet16_1_7QNode_Int_2_d;
  Int_t lizzieLet16_1_7QNode_Int_2_bufchan_buf;
  assign lizzieLet16_1_7QNode_Int_2_bufchan_r = (! lizzieLet16_1_7QNode_Int_2_bufchan_buf[0]);
  assign lizzieLet16_1_7QNode_Int_2_argbuf_d = (lizzieLet16_1_7QNode_Int_2_bufchan_buf[0] ? lizzieLet16_1_7QNode_Int_2_bufchan_buf :
                                                lizzieLet16_1_7QNode_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet16_1_7QNode_Int_2_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((lizzieLet16_1_7QNode_Int_2_argbuf_r && lizzieLet16_1_7QNode_Int_2_bufchan_buf[0]))
        lizzieLet16_1_7QNode_Int_2_bufchan_buf <= {32'd0, 1'd0};
      else if (((! lizzieLet16_1_7QNode_Int_2_argbuf_r) && (! lizzieLet16_1_7QNode_Int_2_bufchan_buf[0])))
        lizzieLet16_1_7QNode_Int_2_bufchan_buf <= lizzieLet16_1_7QNode_Int_2_bufchan_d;
  
  /* buf (Ty Int) : (lizzieLet16_1_7QVal_Int,Int) > (lizzieLet16_1_7QVal_Int_1_argbuf,Int) */
  Int_t lizzieLet16_1_7QVal_Int_bufchan_d;
  logic lizzieLet16_1_7QVal_Int_bufchan_r;
  assign lizzieLet16_1_7QVal_Int_r = ((! lizzieLet16_1_7QVal_Int_bufchan_d[0]) || lizzieLet16_1_7QVal_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet16_1_7QVal_Int_bufchan_d <= {32'd0, 1'd0};
    else
      if (lizzieLet16_1_7QVal_Int_r)
        lizzieLet16_1_7QVal_Int_bufchan_d <= lizzieLet16_1_7QVal_Int_d;
  Int_t lizzieLet16_1_7QVal_Int_bufchan_buf;
  assign lizzieLet16_1_7QVal_Int_bufchan_r = (! lizzieLet16_1_7QVal_Int_bufchan_buf[0]);
  assign lizzieLet16_1_7QVal_Int_1_argbuf_d = (lizzieLet16_1_7QVal_Int_bufchan_buf[0] ? lizzieLet16_1_7QVal_Int_bufchan_buf :
                                               lizzieLet16_1_7QVal_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet16_1_7QVal_Int_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((lizzieLet16_1_7QVal_Int_1_argbuf_r && lizzieLet16_1_7QVal_Int_bufchan_buf[0]))
        lizzieLet16_1_7QVal_Int_bufchan_buf <= {32'd0, 1'd0};
      else if (((! lizzieLet16_1_7QVal_Int_1_argbuf_r) && (! lizzieLet16_1_7QVal_Int_bufchan_buf[0])))
        lizzieLet16_1_7QVal_Int_bufchan_buf <= lizzieLet16_1_7QVal_Int_bufchan_d;
  
  /* buf (Ty Bool) : (lizzieLet1_1wild1X1h_1_Eq,Bool) > (lizzieLet2_1_argbuf,Bool) */
  Bool_t lizzieLet1_1wild1X1h_1_Eq_bufchan_d;
  logic lizzieLet1_1wild1X1h_1_Eq_bufchan_r;
  assign lizzieLet1_1wild1X1h_1_Eq_r = ((! lizzieLet1_1wild1X1h_1_Eq_bufchan_d[0]) || lizzieLet1_1wild1X1h_1_Eq_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet1_1wild1X1h_1_Eq_bufchan_d <= {1'd0, 1'd0};
    else
      if (lizzieLet1_1wild1X1h_1_Eq_r)
        lizzieLet1_1wild1X1h_1_Eq_bufchan_d <= lizzieLet1_1wild1X1h_1_Eq_d;
  Bool_t lizzieLet1_1wild1X1h_1_Eq_bufchan_buf;
  assign lizzieLet1_1wild1X1h_1_Eq_bufchan_r = (! lizzieLet1_1wild1X1h_1_Eq_bufchan_buf[0]);
  assign lizzieLet2_1_argbuf_d = (lizzieLet1_1wild1X1h_1_Eq_bufchan_buf[0] ? lizzieLet1_1wild1X1h_1_Eq_bufchan_buf :
                                  lizzieLet1_1wild1X1h_1_Eq_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet1_1wild1X1h_1_Eq_bufchan_buf <= {1'd0, 1'd0};
    else
      if ((lizzieLet2_1_argbuf_r && lizzieLet1_1wild1X1h_1_Eq_bufchan_buf[0]))
        lizzieLet1_1wild1X1h_1_Eq_bufchan_buf <= {1'd0, 1'd0};
      else if (((! lizzieLet2_1_argbuf_r) && (! lizzieLet1_1wild1X1h_1_Eq_bufchan_buf[0])))
        lizzieLet1_1wild1X1h_1_Eq_bufchan_buf <= lizzieLet1_1wild1X1h_1_Eq_bufchan_d;
  
  /* destruct (Ty CT$wnnz_Int,
          Dcon Lcall_$wnnz_Int0) : (lizzieLet25_1Lcall_$wnnz_Int0,CT$wnnz_Int) > [(wwsvw_3_destruct,Int#),
                                                                                  (ww1XwI_2_destruct,Int#),
                                                                                  (ww2XwL_1_destruct,Int#),
                                                                                  (sc_0_7_destruct,Pointer_CT$wnnz_Int)] */
  logic [3:0] lizzieLet25_1Lcall_$wnnz_Int0_emitted;
  logic [3:0] lizzieLet25_1Lcall_$wnnz_Int0_done;
  assign wwsvw_3_destruct_d = {lizzieLet25_1Lcall_$wnnz_Int0_d[35:4],
                               (lizzieLet25_1Lcall_$wnnz_Int0_d[0] && (! lizzieLet25_1Lcall_$wnnz_Int0_emitted[0]))};
  assign ww1XwI_2_destruct_d = {lizzieLet25_1Lcall_$wnnz_Int0_d[67:36],
                                (lizzieLet25_1Lcall_$wnnz_Int0_d[0] && (! lizzieLet25_1Lcall_$wnnz_Int0_emitted[1]))};
  assign ww2XwL_1_destruct_d = {lizzieLet25_1Lcall_$wnnz_Int0_d[99:68],
                                (lizzieLet25_1Lcall_$wnnz_Int0_d[0] && (! lizzieLet25_1Lcall_$wnnz_Int0_emitted[2]))};
  assign sc_0_7_destruct_d = {lizzieLet25_1Lcall_$wnnz_Int0_d[115:100],
                              (lizzieLet25_1Lcall_$wnnz_Int0_d[0] && (! lizzieLet25_1Lcall_$wnnz_Int0_emitted[3]))};
  assign lizzieLet25_1Lcall_$wnnz_Int0_done = (lizzieLet25_1Lcall_$wnnz_Int0_emitted | ({sc_0_7_destruct_d[0],
                                                                                         ww2XwL_1_destruct_d[0],
                                                                                         ww1XwI_2_destruct_d[0],
                                                                                         wwsvw_3_destruct_d[0]} & {sc_0_7_destruct_r,
                                                                                                                   ww2XwL_1_destruct_r,
                                                                                                                   ww1XwI_2_destruct_r,
                                                                                                                   wwsvw_3_destruct_r}));
  assign lizzieLet25_1Lcall_$wnnz_Int0_r = (& lizzieLet25_1Lcall_$wnnz_Int0_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet25_1Lcall_$wnnz_Int0_emitted <= 4'd0;
    else
      lizzieLet25_1Lcall_$wnnz_Int0_emitted <= (lizzieLet25_1Lcall_$wnnz_Int0_r ? 4'd0 :
                                                lizzieLet25_1Lcall_$wnnz_Int0_done);
  
  /* destruct (Ty CT$wnnz_Int,
          Dcon Lcall_$wnnz_Int1) : (lizzieLet25_1Lcall_$wnnz_Int1,CT$wnnz_Int) > [(wwsvw_2_destruct,Int#),
                                                                                  (ww1XwI_1_destruct,Int#),
                                                                                  (sc_0_6_destruct,Pointer_CT$wnnz_Int),
                                                                                  (q4ac3_3_destruct,Pointer_QTree_Int)] */
  logic [3:0] lizzieLet25_1Lcall_$wnnz_Int1_emitted;
  logic [3:0] lizzieLet25_1Lcall_$wnnz_Int1_done;
  assign wwsvw_2_destruct_d = {lizzieLet25_1Lcall_$wnnz_Int1_d[35:4],
                               (lizzieLet25_1Lcall_$wnnz_Int1_d[0] && (! lizzieLet25_1Lcall_$wnnz_Int1_emitted[0]))};
  assign ww1XwI_1_destruct_d = {lizzieLet25_1Lcall_$wnnz_Int1_d[67:36],
                                (lizzieLet25_1Lcall_$wnnz_Int1_d[0] && (! lizzieLet25_1Lcall_$wnnz_Int1_emitted[1]))};
  assign sc_0_6_destruct_d = {lizzieLet25_1Lcall_$wnnz_Int1_d[83:68],
                              (lizzieLet25_1Lcall_$wnnz_Int1_d[0] && (! lizzieLet25_1Lcall_$wnnz_Int1_emitted[2]))};
  assign q4ac3_3_destruct_d = {lizzieLet25_1Lcall_$wnnz_Int1_d[99:84],
                               (lizzieLet25_1Lcall_$wnnz_Int1_d[0] && (! lizzieLet25_1Lcall_$wnnz_Int1_emitted[3]))};
  assign lizzieLet25_1Lcall_$wnnz_Int1_done = (lizzieLet25_1Lcall_$wnnz_Int1_emitted | ({q4ac3_3_destruct_d[0],
                                                                                         sc_0_6_destruct_d[0],
                                                                                         ww1XwI_1_destruct_d[0],
                                                                                         wwsvw_2_destruct_d[0]} & {q4ac3_3_destruct_r,
                                                                                                                   sc_0_6_destruct_r,
                                                                                                                   ww1XwI_1_destruct_r,
                                                                                                                   wwsvw_2_destruct_r}));
  assign lizzieLet25_1Lcall_$wnnz_Int1_r = (& lizzieLet25_1Lcall_$wnnz_Int1_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet25_1Lcall_$wnnz_Int1_emitted <= 4'd0;
    else
      lizzieLet25_1Lcall_$wnnz_Int1_emitted <= (lizzieLet25_1Lcall_$wnnz_Int1_r ? 4'd0 :
                                                lizzieLet25_1Lcall_$wnnz_Int1_done);
  
  /* destruct (Ty CT$wnnz_Int,
          Dcon Lcall_$wnnz_Int2) : (lizzieLet25_1Lcall_$wnnz_Int2,CT$wnnz_Int) > [(wwsvw_1_destruct,Int#),
                                                                                  (sc_0_5_destruct,Pointer_CT$wnnz_Int),
                                                                                  (q4ac3_2_destruct,Pointer_QTree_Int),
                                                                                  (q3ac2_2_destruct,Pointer_QTree_Int)] */
  logic [3:0] lizzieLet25_1Lcall_$wnnz_Int2_emitted;
  logic [3:0] lizzieLet25_1Lcall_$wnnz_Int2_done;
  assign wwsvw_1_destruct_d = {lizzieLet25_1Lcall_$wnnz_Int2_d[35:4],
                               (lizzieLet25_1Lcall_$wnnz_Int2_d[0] && (! lizzieLet25_1Lcall_$wnnz_Int2_emitted[0]))};
  assign sc_0_5_destruct_d = {lizzieLet25_1Lcall_$wnnz_Int2_d[51:36],
                              (lizzieLet25_1Lcall_$wnnz_Int2_d[0] && (! lizzieLet25_1Lcall_$wnnz_Int2_emitted[1]))};
  assign q4ac3_2_destruct_d = {lizzieLet25_1Lcall_$wnnz_Int2_d[67:52],
                               (lizzieLet25_1Lcall_$wnnz_Int2_d[0] && (! lizzieLet25_1Lcall_$wnnz_Int2_emitted[2]))};
  assign q3ac2_2_destruct_d = {lizzieLet25_1Lcall_$wnnz_Int2_d[83:68],
                               (lizzieLet25_1Lcall_$wnnz_Int2_d[0] && (! lizzieLet25_1Lcall_$wnnz_Int2_emitted[3]))};
  assign lizzieLet25_1Lcall_$wnnz_Int2_done = (lizzieLet25_1Lcall_$wnnz_Int2_emitted | ({q3ac2_2_destruct_d[0],
                                                                                         q4ac3_2_destruct_d[0],
                                                                                         sc_0_5_destruct_d[0],
                                                                                         wwsvw_1_destruct_d[0]} & {q3ac2_2_destruct_r,
                                                                                                                   q4ac3_2_destruct_r,
                                                                                                                   sc_0_5_destruct_r,
                                                                                                                   wwsvw_1_destruct_r}));
  assign lizzieLet25_1Lcall_$wnnz_Int2_r = (& lizzieLet25_1Lcall_$wnnz_Int2_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet25_1Lcall_$wnnz_Int2_emitted <= 4'd0;
    else
      lizzieLet25_1Lcall_$wnnz_Int2_emitted <= (lizzieLet25_1Lcall_$wnnz_Int2_r ? 4'd0 :
                                                lizzieLet25_1Lcall_$wnnz_Int2_done);
  
  /* destruct (Ty CT$wnnz_Int,
          Dcon Lcall_$wnnz_Int3) : (lizzieLet25_1Lcall_$wnnz_Int3,CT$wnnz_Int) > [(sc_0_4_destruct,Pointer_CT$wnnz_Int),
                                                                                  (q4ac3_1_destruct,Pointer_QTree_Int),
                                                                                  (q3ac2_1_destruct,Pointer_QTree_Int),
                                                                                  (q2ac1_1_destruct,Pointer_QTree_Int)] */
  logic [3:0] lizzieLet25_1Lcall_$wnnz_Int3_emitted;
  logic [3:0] lizzieLet25_1Lcall_$wnnz_Int3_done;
  assign sc_0_4_destruct_d = {lizzieLet25_1Lcall_$wnnz_Int3_d[19:4],
                              (lizzieLet25_1Lcall_$wnnz_Int3_d[0] && (! lizzieLet25_1Lcall_$wnnz_Int3_emitted[0]))};
  assign q4ac3_1_destruct_d = {lizzieLet25_1Lcall_$wnnz_Int3_d[35:20],
                               (lizzieLet25_1Lcall_$wnnz_Int3_d[0] && (! lizzieLet25_1Lcall_$wnnz_Int3_emitted[1]))};
  assign q3ac2_1_destruct_d = {lizzieLet25_1Lcall_$wnnz_Int3_d[51:36],
                               (lizzieLet25_1Lcall_$wnnz_Int3_d[0] && (! lizzieLet25_1Lcall_$wnnz_Int3_emitted[2]))};
  assign q2ac1_1_destruct_d = {lizzieLet25_1Lcall_$wnnz_Int3_d[67:52],
                               (lizzieLet25_1Lcall_$wnnz_Int3_d[0] && (! lizzieLet25_1Lcall_$wnnz_Int3_emitted[3]))};
  assign lizzieLet25_1Lcall_$wnnz_Int3_done = (lizzieLet25_1Lcall_$wnnz_Int3_emitted | ({q2ac1_1_destruct_d[0],
                                                                                         q3ac2_1_destruct_d[0],
                                                                                         q4ac3_1_destruct_d[0],
                                                                                         sc_0_4_destruct_d[0]} & {q2ac1_1_destruct_r,
                                                                                                                  q3ac2_1_destruct_r,
                                                                                                                  q4ac3_1_destruct_r,
                                                                                                                  sc_0_4_destruct_r}));
  assign lizzieLet25_1Lcall_$wnnz_Int3_r = (& lizzieLet25_1Lcall_$wnnz_Int3_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet25_1Lcall_$wnnz_Int3_emitted <= 4'd0;
    else
      lizzieLet25_1Lcall_$wnnz_Int3_emitted <= (lizzieLet25_1Lcall_$wnnz_Int3_r ? 4'd0 :
                                                lizzieLet25_1Lcall_$wnnz_Int3_done);
  
  /* demux (Ty CT$wnnz_Int,
       Ty CT$wnnz_Int) : (lizzieLet25_2,CT$wnnz_Int) (lizzieLet25_1,CT$wnnz_Int) > [(_18,CT$wnnz_Int),
                                                                                    (lizzieLet25_1Lcall_$wnnz_Int3,CT$wnnz_Int),
                                                                                    (lizzieLet25_1Lcall_$wnnz_Int2,CT$wnnz_Int),
                                                                                    (lizzieLet25_1Lcall_$wnnz_Int1,CT$wnnz_Int),
                                                                                    (lizzieLet25_1Lcall_$wnnz_Int0,CT$wnnz_Int)] */
  logic [4:0] lizzieLet25_1_onehotd;
  always_comb
    if ((lizzieLet25_2_d[0] && lizzieLet25_1_d[0]))
      unique case (lizzieLet25_2_d[3:1])
        3'd0: lizzieLet25_1_onehotd = 5'd1;
        3'd1: lizzieLet25_1_onehotd = 5'd2;
        3'd2: lizzieLet25_1_onehotd = 5'd4;
        3'd3: lizzieLet25_1_onehotd = 5'd8;
        3'd4: lizzieLet25_1_onehotd = 5'd16;
        default: lizzieLet25_1_onehotd = 5'd0;
      endcase
    else lizzieLet25_1_onehotd = 5'd0;
  assign _18_d = {lizzieLet25_1_d[115:1], lizzieLet25_1_onehotd[0]};
  assign lizzieLet25_1Lcall_$wnnz_Int3_d = {lizzieLet25_1_d[115:1],
                                            lizzieLet25_1_onehotd[1]};
  assign lizzieLet25_1Lcall_$wnnz_Int2_d = {lizzieLet25_1_d[115:1],
                                            lizzieLet25_1_onehotd[2]};
  assign lizzieLet25_1Lcall_$wnnz_Int1_d = {lizzieLet25_1_d[115:1],
                                            lizzieLet25_1_onehotd[3]};
  assign lizzieLet25_1Lcall_$wnnz_Int0_d = {lizzieLet25_1_d[115:1],
                                            lizzieLet25_1_onehotd[4]};
  assign lizzieLet25_1_r = (| (lizzieLet25_1_onehotd & {lizzieLet25_1Lcall_$wnnz_Int0_r,
                                                        lizzieLet25_1Lcall_$wnnz_Int1_r,
                                                        lizzieLet25_1Lcall_$wnnz_Int2_r,
                                                        lizzieLet25_1Lcall_$wnnz_Int3_r,
                                                        _18_r}));
  assign lizzieLet25_2_r = lizzieLet25_1_r;
  
  /* demux (Ty CT$wnnz_Int,
       Ty Go) : (lizzieLet25_3,CT$wnnz_Int) (go_18_goMux_data,Go) > [(_17,Go),
                                                                     (lizzieLet25_3Lcall_$wnnz_Int3,Go),
                                                                     (lizzieLet25_3Lcall_$wnnz_Int2,Go),
                                                                     (lizzieLet25_3Lcall_$wnnz_Int1,Go),
                                                                     (lizzieLet25_3Lcall_$wnnz_Int0,Go)] */
  logic [4:0] go_18_goMux_data_onehotd;
  always_comb
    if ((lizzieLet25_3_d[0] && go_18_goMux_data_d[0]))
      unique case (lizzieLet25_3_d[3:1])
        3'd0: go_18_goMux_data_onehotd = 5'd1;
        3'd1: go_18_goMux_data_onehotd = 5'd2;
        3'd2: go_18_goMux_data_onehotd = 5'd4;
        3'd3: go_18_goMux_data_onehotd = 5'd8;
        3'd4: go_18_goMux_data_onehotd = 5'd16;
        default: go_18_goMux_data_onehotd = 5'd0;
      endcase
    else go_18_goMux_data_onehotd = 5'd0;
  assign _17_d = go_18_goMux_data_onehotd[0];
  assign lizzieLet25_3Lcall_$wnnz_Int3_d = go_18_goMux_data_onehotd[1];
  assign lizzieLet25_3Lcall_$wnnz_Int2_d = go_18_goMux_data_onehotd[2];
  assign lizzieLet25_3Lcall_$wnnz_Int1_d = go_18_goMux_data_onehotd[3];
  assign lizzieLet25_3Lcall_$wnnz_Int0_d = go_18_goMux_data_onehotd[4];
  assign go_18_goMux_data_r = (| (go_18_goMux_data_onehotd & {lizzieLet25_3Lcall_$wnnz_Int0_r,
                                                              lizzieLet25_3Lcall_$wnnz_Int1_r,
                                                              lizzieLet25_3Lcall_$wnnz_Int2_r,
                                                              lizzieLet25_3Lcall_$wnnz_Int3_r,
                                                              _17_r}));
  assign lizzieLet25_3_r = go_18_goMux_data_r;
  
  /* buf (Ty Go) : (lizzieLet25_3Lcall_$wnnz_Int0,Go) > (lizzieLet25_3Lcall_$wnnz_Int0_1_argbuf,Go) */
  Go_t lizzieLet25_3Lcall_$wnnz_Int0_bufchan_d;
  logic lizzieLet25_3Lcall_$wnnz_Int0_bufchan_r;
  assign lizzieLet25_3Lcall_$wnnz_Int0_r = ((! lizzieLet25_3Lcall_$wnnz_Int0_bufchan_d[0]) || lizzieLet25_3Lcall_$wnnz_Int0_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet25_3Lcall_$wnnz_Int0_bufchan_d <= 1'd0;
    else
      if (lizzieLet25_3Lcall_$wnnz_Int0_r)
        lizzieLet25_3Lcall_$wnnz_Int0_bufchan_d <= lizzieLet25_3Lcall_$wnnz_Int0_d;
  Go_t lizzieLet25_3Lcall_$wnnz_Int0_bufchan_buf;
  assign lizzieLet25_3Lcall_$wnnz_Int0_bufchan_r = (! lizzieLet25_3Lcall_$wnnz_Int0_bufchan_buf[0]);
  assign lizzieLet25_3Lcall_$wnnz_Int0_1_argbuf_d = (lizzieLet25_3Lcall_$wnnz_Int0_bufchan_buf[0] ? lizzieLet25_3Lcall_$wnnz_Int0_bufchan_buf :
                                                     lizzieLet25_3Lcall_$wnnz_Int0_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet25_3Lcall_$wnnz_Int0_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet25_3Lcall_$wnnz_Int0_1_argbuf_r && lizzieLet25_3Lcall_$wnnz_Int0_bufchan_buf[0]))
        lizzieLet25_3Lcall_$wnnz_Int0_bufchan_buf <= 1'd0;
      else if (((! lizzieLet25_3Lcall_$wnnz_Int0_1_argbuf_r) && (! lizzieLet25_3Lcall_$wnnz_Int0_bufchan_buf[0])))
        lizzieLet25_3Lcall_$wnnz_Int0_bufchan_buf <= lizzieLet25_3Lcall_$wnnz_Int0_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet25_3Lcall_$wnnz_Int1,Go) > (lizzieLet25_3Lcall_$wnnz_Int1_1_argbuf,Go) */
  Go_t lizzieLet25_3Lcall_$wnnz_Int1_bufchan_d;
  logic lizzieLet25_3Lcall_$wnnz_Int1_bufchan_r;
  assign lizzieLet25_3Lcall_$wnnz_Int1_r = ((! lizzieLet25_3Lcall_$wnnz_Int1_bufchan_d[0]) || lizzieLet25_3Lcall_$wnnz_Int1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet25_3Lcall_$wnnz_Int1_bufchan_d <= 1'd0;
    else
      if (lizzieLet25_3Lcall_$wnnz_Int1_r)
        lizzieLet25_3Lcall_$wnnz_Int1_bufchan_d <= lizzieLet25_3Lcall_$wnnz_Int1_d;
  Go_t lizzieLet25_3Lcall_$wnnz_Int1_bufchan_buf;
  assign lizzieLet25_3Lcall_$wnnz_Int1_bufchan_r = (! lizzieLet25_3Lcall_$wnnz_Int1_bufchan_buf[0]);
  assign lizzieLet25_3Lcall_$wnnz_Int1_1_argbuf_d = (lizzieLet25_3Lcall_$wnnz_Int1_bufchan_buf[0] ? lizzieLet25_3Lcall_$wnnz_Int1_bufchan_buf :
                                                     lizzieLet25_3Lcall_$wnnz_Int1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet25_3Lcall_$wnnz_Int1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet25_3Lcall_$wnnz_Int1_1_argbuf_r && lizzieLet25_3Lcall_$wnnz_Int1_bufchan_buf[0]))
        lizzieLet25_3Lcall_$wnnz_Int1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet25_3Lcall_$wnnz_Int1_1_argbuf_r) && (! lizzieLet25_3Lcall_$wnnz_Int1_bufchan_buf[0])))
        lizzieLet25_3Lcall_$wnnz_Int1_bufchan_buf <= lizzieLet25_3Lcall_$wnnz_Int1_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet25_3Lcall_$wnnz_Int2,Go) > (lizzieLet25_3Lcall_$wnnz_Int2_1_argbuf,Go) */
  Go_t lizzieLet25_3Lcall_$wnnz_Int2_bufchan_d;
  logic lizzieLet25_3Lcall_$wnnz_Int2_bufchan_r;
  assign lizzieLet25_3Lcall_$wnnz_Int2_r = ((! lizzieLet25_3Lcall_$wnnz_Int2_bufchan_d[0]) || lizzieLet25_3Lcall_$wnnz_Int2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet25_3Lcall_$wnnz_Int2_bufchan_d <= 1'd0;
    else
      if (lizzieLet25_3Lcall_$wnnz_Int2_r)
        lizzieLet25_3Lcall_$wnnz_Int2_bufchan_d <= lizzieLet25_3Lcall_$wnnz_Int2_d;
  Go_t lizzieLet25_3Lcall_$wnnz_Int2_bufchan_buf;
  assign lizzieLet25_3Lcall_$wnnz_Int2_bufchan_r = (! lizzieLet25_3Lcall_$wnnz_Int2_bufchan_buf[0]);
  assign lizzieLet25_3Lcall_$wnnz_Int2_1_argbuf_d = (lizzieLet25_3Lcall_$wnnz_Int2_bufchan_buf[0] ? lizzieLet25_3Lcall_$wnnz_Int2_bufchan_buf :
                                                     lizzieLet25_3Lcall_$wnnz_Int2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet25_3Lcall_$wnnz_Int2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet25_3Lcall_$wnnz_Int2_1_argbuf_r && lizzieLet25_3Lcall_$wnnz_Int2_bufchan_buf[0]))
        lizzieLet25_3Lcall_$wnnz_Int2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet25_3Lcall_$wnnz_Int2_1_argbuf_r) && (! lizzieLet25_3Lcall_$wnnz_Int2_bufchan_buf[0])))
        lizzieLet25_3Lcall_$wnnz_Int2_bufchan_buf <= lizzieLet25_3Lcall_$wnnz_Int2_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet25_3Lcall_$wnnz_Int3,Go) > (lizzieLet25_3Lcall_$wnnz_Int3_1_argbuf,Go) */
  Go_t lizzieLet25_3Lcall_$wnnz_Int3_bufchan_d;
  logic lizzieLet25_3Lcall_$wnnz_Int3_bufchan_r;
  assign lizzieLet25_3Lcall_$wnnz_Int3_r = ((! lizzieLet25_3Lcall_$wnnz_Int3_bufchan_d[0]) || lizzieLet25_3Lcall_$wnnz_Int3_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet25_3Lcall_$wnnz_Int3_bufchan_d <= 1'd0;
    else
      if (lizzieLet25_3Lcall_$wnnz_Int3_r)
        lizzieLet25_3Lcall_$wnnz_Int3_bufchan_d <= lizzieLet25_3Lcall_$wnnz_Int3_d;
  Go_t lizzieLet25_3Lcall_$wnnz_Int3_bufchan_buf;
  assign lizzieLet25_3Lcall_$wnnz_Int3_bufchan_r = (! lizzieLet25_3Lcall_$wnnz_Int3_bufchan_buf[0]);
  assign lizzieLet25_3Lcall_$wnnz_Int3_1_argbuf_d = (lizzieLet25_3Lcall_$wnnz_Int3_bufchan_buf[0] ? lizzieLet25_3Lcall_$wnnz_Int3_bufchan_buf :
                                                     lizzieLet25_3Lcall_$wnnz_Int3_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet25_3Lcall_$wnnz_Int3_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet25_3Lcall_$wnnz_Int3_1_argbuf_r && lizzieLet25_3Lcall_$wnnz_Int3_bufchan_buf[0]))
        lizzieLet25_3Lcall_$wnnz_Int3_bufchan_buf <= 1'd0;
      else if (((! lizzieLet25_3Lcall_$wnnz_Int3_1_argbuf_r) && (! lizzieLet25_3Lcall_$wnnz_Int3_bufchan_buf[0])))
        lizzieLet25_3Lcall_$wnnz_Int3_bufchan_buf <= lizzieLet25_3Lcall_$wnnz_Int3_bufchan_d;
  
  /* demux (Ty CT$wnnz_Int,
       Ty Int#) : (lizzieLet25_4,CT$wnnz_Int) (srtarg_0_goMux_mux,Int#) > [(lizzieLet25_4L$wnnz_Intsbos,Int#),
                                                                           (lizzieLet25_4Lcall_$wnnz_Int3,Int#),
                                                                           (lizzieLet25_4Lcall_$wnnz_Int2,Int#),
                                                                           (lizzieLet25_4Lcall_$wnnz_Int1,Int#),
                                                                           (lizzieLet25_4Lcall_$wnnz_Int0,Int#)] */
  logic [4:0] srtarg_0_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet25_4_d[0] && srtarg_0_goMux_mux_d[0]))
      unique case (lizzieLet25_4_d[3:1])
        3'd0: srtarg_0_goMux_mux_onehotd = 5'd1;
        3'd1: srtarg_0_goMux_mux_onehotd = 5'd2;
        3'd2: srtarg_0_goMux_mux_onehotd = 5'd4;
        3'd3: srtarg_0_goMux_mux_onehotd = 5'd8;
        3'd4: srtarg_0_goMux_mux_onehotd = 5'd16;
        default: srtarg_0_goMux_mux_onehotd = 5'd0;
      endcase
    else srtarg_0_goMux_mux_onehotd = 5'd0;
  assign lizzieLet25_4L$wnnz_Intsbos_d = {srtarg_0_goMux_mux_d[32:1],
                                          srtarg_0_goMux_mux_onehotd[0]};
  assign lizzieLet25_4Lcall_$wnnz_Int3_d = {srtarg_0_goMux_mux_d[32:1],
                                            srtarg_0_goMux_mux_onehotd[1]};
  assign lizzieLet25_4Lcall_$wnnz_Int2_d = {srtarg_0_goMux_mux_d[32:1],
                                            srtarg_0_goMux_mux_onehotd[2]};
  assign lizzieLet25_4Lcall_$wnnz_Int1_d = {srtarg_0_goMux_mux_d[32:1],
                                            srtarg_0_goMux_mux_onehotd[3]};
  assign lizzieLet25_4Lcall_$wnnz_Int0_d = {srtarg_0_goMux_mux_d[32:1],
                                            srtarg_0_goMux_mux_onehotd[4]};
  assign srtarg_0_goMux_mux_r = (| (srtarg_0_goMux_mux_onehotd & {lizzieLet25_4Lcall_$wnnz_Int0_r,
                                                                  lizzieLet25_4Lcall_$wnnz_Int1_r,
                                                                  lizzieLet25_4Lcall_$wnnz_Int2_r,
                                                                  lizzieLet25_4Lcall_$wnnz_Int3_r,
                                                                  lizzieLet25_4L$wnnz_Intsbos_r}));
  assign lizzieLet25_4_r = srtarg_0_goMux_mux_r;
  
  /* fork (Ty Int#) : (lizzieLet25_4L$wnnz_Intsbos,Int#) > [(lizzieLet25_4L$wnnz_Intsbos_1_merge_merge_fork_1,Int#),
                                                       (lizzieLet25_4L$wnnz_Intsbos_1_merge_merge_fork_2,Int#)] */
  logic [1:0] lizzieLet25_4L$wnnz_Intsbos_emitted;
  logic [1:0] lizzieLet25_4L$wnnz_Intsbos_done;
  assign lizzieLet25_4L$wnnz_Intsbos_1_merge_merge_fork_1_d = {lizzieLet25_4L$wnnz_Intsbos_d[32:1],
                                                               (lizzieLet25_4L$wnnz_Intsbos_d[0] && (! lizzieLet25_4L$wnnz_Intsbos_emitted[0]))};
  assign lizzieLet25_4L$wnnz_Intsbos_1_merge_merge_fork_2_d = {lizzieLet25_4L$wnnz_Intsbos_d[32:1],
                                                               (lizzieLet25_4L$wnnz_Intsbos_d[0] && (! lizzieLet25_4L$wnnz_Intsbos_emitted[1]))};
  assign lizzieLet25_4L$wnnz_Intsbos_done = (lizzieLet25_4L$wnnz_Intsbos_emitted | ({lizzieLet25_4L$wnnz_Intsbos_1_merge_merge_fork_2_d[0],
                                                                                     lizzieLet25_4L$wnnz_Intsbos_1_merge_merge_fork_1_d[0]} & {lizzieLet25_4L$wnnz_Intsbos_1_merge_merge_fork_2_r,
                                                                                                                                               lizzieLet25_4L$wnnz_Intsbos_1_merge_merge_fork_1_r}));
  assign lizzieLet25_4L$wnnz_Intsbos_r = (& lizzieLet25_4L$wnnz_Intsbos_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet25_4L$wnnz_Intsbos_emitted <= 2'd0;
    else
      lizzieLet25_4L$wnnz_Intsbos_emitted <= (lizzieLet25_4L$wnnz_Intsbos_r ? 2'd0 :
                                              lizzieLet25_4L$wnnz_Intsbos_done);
  
  /* togo (Ty Int#) : (lizzieLet25_4L$wnnz_Intsbos_1_merge_merge_fork_1,Int#) > (call_$wnnz_Int_goConst,Go) */
  assign call_$wnnz_Int_goConst_d = lizzieLet25_4L$wnnz_Intsbos_1_merge_merge_fork_1_d[0];
  assign lizzieLet25_4L$wnnz_Intsbos_1_merge_merge_fork_1_r = call_$wnnz_Int_goConst_r;
  
  /* buf (Ty Int#) : (lizzieLet25_4L$wnnz_Intsbos_1_merge_merge_fork_2,Int#) > ($wnnz_Int_resbuf,Int#) */
  \Int#_t  lizzieLet25_4L$wnnz_Intsbos_1_merge_merge_fork_2_bufchan_d;
  logic lizzieLet25_4L$wnnz_Intsbos_1_merge_merge_fork_2_bufchan_r;
  assign lizzieLet25_4L$wnnz_Intsbos_1_merge_merge_fork_2_r = ((! lizzieLet25_4L$wnnz_Intsbos_1_merge_merge_fork_2_bufchan_d[0]) || lizzieLet25_4L$wnnz_Intsbos_1_merge_merge_fork_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet25_4L$wnnz_Intsbos_1_merge_merge_fork_2_bufchan_d <= {32'd0,
                                                                     1'd0};
    else
      if (lizzieLet25_4L$wnnz_Intsbos_1_merge_merge_fork_2_r)
        lizzieLet25_4L$wnnz_Intsbos_1_merge_merge_fork_2_bufchan_d <= lizzieLet25_4L$wnnz_Intsbos_1_merge_merge_fork_2_d;
  \Int#_t  lizzieLet25_4L$wnnz_Intsbos_1_merge_merge_fork_2_bufchan_buf;
  assign lizzieLet25_4L$wnnz_Intsbos_1_merge_merge_fork_2_bufchan_r = (! lizzieLet25_4L$wnnz_Intsbos_1_merge_merge_fork_2_bufchan_buf[0]);
  assign \$wnnz_Int_resbuf_d  = (lizzieLet25_4L$wnnz_Intsbos_1_merge_merge_fork_2_bufchan_buf[0] ? lizzieLet25_4L$wnnz_Intsbos_1_merge_merge_fork_2_bufchan_buf :
                                 lizzieLet25_4L$wnnz_Intsbos_1_merge_merge_fork_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet25_4L$wnnz_Intsbos_1_merge_merge_fork_2_bufchan_buf <= {32'd0,
                                                                       1'd0};
    else
      if ((\$wnnz_Int_resbuf_r  && lizzieLet25_4L$wnnz_Intsbos_1_merge_merge_fork_2_bufchan_buf[0]))
        lizzieLet25_4L$wnnz_Intsbos_1_merge_merge_fork_2_bufchan_buf <= {32'd0,
                                                                         1'd0};
      else if (((! \$wnnz_Int_resbuf_r ) && (! lizzieLet25_4L$wnnz_Intsbos_1_merge_merge_fork_2_bufchan_buf[0])))
        lizzieLet25_4L$wnnz_Intsbos_1_merge_merge_fork_2_bufchan_buf <= lizzieLet25_4L$wnnz_Intsbos_1_merge_merge_fork_2_bufchan_d;
  
  /* dcon (Ty CT$wnnz_Int,
      Dcon Lcall_$wnnz_Int2) : [(lizzieLet25_4Lcall_$wnnz_Int3,Int#),
                                (sc_0_4_destruct,Pointer_CT$wnnz_Int),
                                (q4ac3_1_destruct,Pointer_QTree_Int),
                                (q3ac2_1_destruct,Pointer_QTree_Int)] > (lizzieLet25_4Lcall_$wnnz_Int3_1sc_0_4_1q4ac3_1_1q3ac2_1_1Lcall_$wnnz_Int2,CT$wnnz_Int) */
  assign lizzieLet25_4Lcall_$wnnz_Int3_1sc_0_4_1q4ac3_1_1q3ac2_1_1Lcall_$wnnz_Int2_d = Lcall_$wnnz_Int2_dc((& {lizzieLet25_4Lcall_$wnnz_Int3_d[0],
                                                                                                               sc_0_4_destruct_d[0],
                                                                                                               q4ac3_1_destruct_d[0],
                                                                                                               q3ac2_1_destruct_d[0]}), lizzieLet25_4Lcall_$wnnz_Int3_d, sc_0_4_destruct_d, q4ac3_1_destruct_d, q3ac2_1_destruct_d);
  assign {lizzieLet25_4Lcall_$wnnz_Int3_r,
          sc_0_4_destruct_r,
          q4ac3_1_destruct_r,
          q3ac2_1_destruct_r} = {4 {(lizzieLet25_4Lcall_$wnnz_Int3_1sc_0_4_1q4ac3_1_1q3ac2_1_1Lcall_$wnnz_Int2_r && lizzieLet25_4Lcall_$wnnz_Int3_1sc_0_4_1q4ac3_1_1q3ac2_1_1Lcall_$wnnz_Int2_d[0])}};
  
  /* buf (Ty CT$wnnz_Int) : (lizzieLet25_4Lcall_$wnnz_Int3_1sc_0_4_1q4ac3_1_1q3ac2_1_1Lcall_$wnnz_Int2,CT$wnnz_Int) > (lizzieLet26_1_argbuf,CT$wnnz_Int) */
  CT$wnnz_Int_t lizzieLet25_4Lcall_$wnnz_Int3_1sc_0_4_1q4ac3_1_1q3ac2_1_1Lcall_$wnnz_Int2_bufchan_d;
  logic lizzieLet25_4Lcall_$wnnz_Int3_1sc_0_4_1q4ac3_1_1q3ac2_1_1Lcall_$wnnz_Int2_bufchan_r;
  assign lizzieLet25_4Lcall_$wnnz_Int3_1sc_0_4_1q4ac3_1_1q3ac2_1_1Lcall_$wnnz_Int2_r = ((! lizzieLet25_4Lcall_$wnnz_Int3_1sc_0_4_1q4ac3_1_1q3ac2_1_1Lcall_$wnnz_Int2_bufchan_d[0]) || lizzieLet25_4Lcall_$wnnz_Int3_1sc_0_4_1q4ac3_1_1q3ac2_1_1Lcall_$wnnz_Int2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet25_4Lcall_$wnnz_Int3_1sc_0_4_1q4ac3_1_1q3ac2_1_1Lcall_$wnnz_Int2_bufchan_d <= {115'd0,
                                                                                              1'd0};
    else
      if (lizzieLet25_4Lcall_$wnnz_Int3_1sc_0_4_1q4ac3_1_1q3ac2_1_1Lcall_$wnnz_Int2_r)
        lizzieLet25_4Lcall_$wnnz_Int3_1sc_0_4_1q4ac3_1_1q3ac2_1_1Lcall_$wnnz_Int2_bufchan_d <= lizzieLet25_4Lcall_$wnnz_Int3_1sc_0_4_1q4ac3_1_1q3ac2_1_1Lcall_$wnnz_Int2_d;
  CT$wnnz_Int_t lizzieLet25_4Lcall_$wnnz_Int3_1sc_0_4_1q4ac3_1_1q3ac2_1_1Lcall_$wnnz_Int2_bufchan_buf;
  assign lizzieLet25_4Lcall_$wnnz_Int3_1sc_0_4_1q4ac3_1_1q3ac2_1_1Lcall_$wnnz_Int2_bufchan_r = (! lizzieLet25_4Lcall_$wnnz_Int3_1sc_0_4_1q4ac3_1_1q3ac2_1_1Lcall_$wnnz_Int2_bufchan_buf[0]);
  assign lizzieLet26_1_argbuf_d = (lizzieLet25_4Lcall_$wnnz_Int3_1sc_0_4_1q4ac3_1_1q3ac2_1_1Lcall_$wnnz_Int2_bufchan_buf[0] ? lizzieLet25_4Lcall_$wnnz_Int3_1sc_0_4_1q4ac3_1_1q3ac2_1_1Lcall_$wnnz_Int2_bufchan_buf :
                                   lizzieLet25_4Lcall_$wnnz_Int3_1sc_0_4_1q4ac3_1_1q3ac2_1_1Lcall_$wnnz_Int2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet25_4Lcall_$wnnz_Int3_1sc_0_4_1q4ac3_1_1q3ac2_1_1Lcall_$wnnz_Int2_bufchan_buf <= {115'd0,
                                                                                                1'd0};
    else
      if ((lizzieLet26_1_argbuf_r && lizzieLet25_4Lcall_$wnnz_Int3_1sc_0_4_1q4ac3_1_1q3ac2_1_1Lcall_$wnnz_Int2_bufchan_buf[0]))
        lizzieLet25_4Lcall_$wnnz_Int3_1sc_0_4_1q4ac3_1_1q3ac2_1_1Lcall_$wnnz_Int2_bufchan_buf <= {115'd0,
                                                                                                  1'd0};
      else if (((! lizzieLet26_1_argbuf_r) && (! lizzieLet25_4Lcall_$wnnz_Int3_1sc_0_4_1q4ac3_1_1q3ac2_1_1Lcall_$wnnz_Int2_bufchan_buf[0])))
        lizzieLet25_4Lcall_$wnnz_Int3_1sc_0_4_1q4ac3_1_1q3ac2_1_1Lcall_$wnnz_Int2_bufchan_buf <= lizzieLet25_4Lcall_$wnnz_Int3_1sc_0_4_1q4ac3_1_1q3ac2_1_1Lcall_$wnnz_Int2_bufchan_d;
  
  /* destruct (Ty CTkron_kron_Int_Int_Int,
          Dcon Lcall_kron_kron_Int_Int_Int0) : (lizzieLet29_1Lcall_kron_kron_Int_Int_Int0,CTkron_kron_Int_Int_Int) > [(es_1_1_destruct,Pointer_QTree_Int),
                                                                                                                      (es_2_2_destruct,Pointer_QTree_Int),
                                                                                                                      (es_3_3_destruct,Pointer_QTree_Int),
                                                                                                                      (sc_0_11_destruct,Pointer_CTkron_kron_Int_Int_Int)] */
  logic [3:0] lizzieLet29_1Lcall_kron_kron_Int_Int_Int0_emitted;
  logic [3:0] lizzieLet29_1Lcall_kron_kron_Int_Int_Int0_done;
  assign es_1_1_destruct_d = {lizzieLet29_1Lcall_kron_kron_Int_Int_Int0_d[19:4],
                              (lizzieLet29_1Lcall_kron_kron_Int_Int_Int0_d[0] && (! lizzieLet29_1Lcall_kron_kron_Int_Int_Int0_emitted[0]))};
  assign es_2_2_destruct_d = {lizzieLet29_1Lcall_kron_kron_Int_Int_Int0_d[35:20],
                              (lizzieLet29_1Lcall_kron_kron_Int_Int_Int0_d[0] && (! lizzieLet29_1Lcall_kron_kron_Int_Int_Int0_emitted[1]))};
  assign es_3_3_destruct_d = {lizzieLet29_1Lcall_kron_kron_Int_Int_Int0_d[51:36],
                              (lizzieLet29_1Lcall_kron_kron_Int_Int_Int0_d[0] && (! lizzieLet29_1Lcall_kron_kron_Int_Int_Int0_emitted[2]))};
  assign sc_0_11_destruct_d = {lizzieLet29_1Lcall_kron_kron_Int_Int_Int0_d[67:52],
                               (lizzieLet29_1Lcall_kron_kron_Int_Int_Int0_d[0] && (! lizzieLet29_1Lcall_kron_kron_Int_Int_Int0_emitted[3]))};
  assign lizzieLet29_1Lcall_kron_kron_Int_Int_Int0_done = (lizzieLet29_1Lcall_kron_kron_Int_Int_Int0_emitted | ({sc_0_11_destruct_d[0],
                                                                                                                 es_3_3_destruct_d[0],
                                                                                                                 es_2_2_destruct_d[0],
                                                                                                                 es_1_1_destruct_d[0]} & {sc_0_11_destruct_r,
                                                                                                                                          es_3_3_destruct_r,
                                                                                                                                          es_2_2_destruct_r,
                                                                                                                                          es_1_1_destruct_r}));
  assign lizzieLet29_1Lcall_kron_kron_Int_Int_Int0_r = (& lizzieLet29_1Lcall_kron_kron_Int_Int_Int0_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet29_1Lcall_kron_kron_Int_Int_Int0_emitted <= 4'd0;
    else
      lizzieLet29_1Lcall_kron_kron_Int_Int_Int0_emitted <= (lizzieLet29_1Lcall_kron_kron_Int_Int_Int0_r ? 4'd0 :
                                                            lizzieLet29_1Lcall_kron_kron_Int_Int_Int0_done);
  
  /* destruct (Ty CTkron_kron_Int_Int_Int,
          Dcon Lcall_kron_kron_Int_Int_Int1) : (lizzieLet29_1Lcall_kron_kron_Int_Int_Int1,CTkron_kron_Int_Int_Int) > [(es_2_1_destruct,Pointer_QTree_Int),
                                                                                                                      (es_3_2_destruct,Pointer_QTree_Int),
                                                                                                                      (sc_0_10_destruct,Pointer_CTkron_kron_Int_Int_Int),
                                                                                                                      (isZad2_4_destruct,MyDTInt_Bool),
                                                                                                                      (gad3_4_destruct,MyDTInt_Int_Int),
                                                                                                                      (q1ad7_3_destruct,Pointer_QTree_Int),
                                                                                                                      (m2ad5_4_destruct,Pointer_QTree_Int)] */
  logic [6:0] lizzieLet29_1Lcall_kron_kron_Int_Int_Int1_emitted;
  logic [6:0] lizzieLet29_1Lcall_kron_kron_Int_Int_Int1_done;
  assign es_2_1_destruct_d = {lizzieLet29_1Lcall_kron_kron_Int_Int_Int1_d[19:4],
                              (lizzieLet29_1Lcall_kron_kron_Int_Int_Int1_d[0] && (! lizzieLet29_1Lcall_kron_kron_Int_Int_Int1_emitted[0]))};
  assign es_3_2_destruct_d = {lizzieLet29_1Lcall_kron_kron_Int_Int_Int1_d[35:20],
                              (lizzieLet29_1Lcall_kron_kron_Int_Int_Int1_d[0] && (! lizzieLet29_1Lcall_kron_kron_Int_Int_Int1_emitted[1]))};
  assign sc_0_10_destruct_d = {lizzieLet29_1Lcall_kron_kron_Int_Int_Int1_d[51:36],
                               (lizzieLet29_1Lcall_kron_kron_Int_Int_Int1_d[0] && (! lizzieLet29_1Lcall_kron_kron_Int_Int_Int1_emitted[2]))};
  assign isZad2_4_destruct_d = (lizzieLet29_1Lcall_kron_kron_Int_Int_Int1_d[0] && (! lizzieLet29_1Lcall_kron_kron_Int_Int_Int1_emitted[3]));
  assign gad3_4_destruct_d = (lizzieLet29_1Lcall_kron_kron_Int_Int_Int1_d[0] && (! lizzieLet29_1Lcall_kron_kron_Int_Int_Int1_emitted[4]));
  assign q1ad7_3_destruct_d = {lizzieLet29_1Lcall_kron_kron_Int_Int_Int1_d[67:52],
                               (lizzieLet29_1Lcall_kron_kron_Int_Int_Int1_d[0] && (! lizzieLet29_1Lcall_kron_kron_Int_Int_Int1_emitted[5]))};
  assign m2ad5_4_destruct_d = {lizzieLet29_1Lcall_kron_kron_Int_Int_Int1_d[83:68],
                               (lizzieLet29_1Lcall_kron_kron_Int_Int_Int1_d[0] && (! lizzieLet29_1Lcall_kron_kron_Int_Int_Int1_emitted[6]))};
  assign lizzieLet29_1Lcall_kron_kron_Int_Int_Int1_done = (lizzieLet29_1Lcall_kron_kron_Int_Int_Int1_emitted | ({m2ad5_4_destruct_d[0],
                                                                                                                 q1ad7_3_destruct_d[0],
                                                                                                                 gad3_4_destruct_d[0],
                                                                                                                 isZad2_4_destruct_d[0],
                                                                                                                 sc_0_10_destruct_d[0],
                                                                                                                 es_3_2_destruct_d[0],
                                                                                                                 es_2_1_destruct_d[0]} & {m2ad5_4_destruct_r,
                                                                                                                                          q1ad7_3_destruct_r,
                                                                                                                                          gad3_4_destruct_r,
                                                                                                                                          isZad2_4_destruct_r,
                                                                                                                                          sc_0_10_destruct_r,
                                                                                                                                          es_3_2_destruct_r,
                                                                                                                                          es_2_1_destruct_r}));
  assign lizzieLet29_1Lcall_kron_kron_Int_Int_Int1_r = (& lizzieLet29_1Lcall_kron_kron_Int_Int_Int1_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet29_1Lcall_kron_kron_Int_Int_Int1_emitted <= 7'd0;
    else
      lizzieLet29_1Lcall_kron_kron_Int_Int_Int1_emitted <= (lizzieLet29_1Lcall_kron_kron_Int_Int_Int1_r ? 7'd0 :
                                                            lizzieLet29_1Lcall_kron_kron_Int_Int_Int1_done);
  
  /* destruct (Ty CTkron_kron_Int_Int_Int,
          Dcon Lcall_kron_kron_Int_Int_Int2) : (lizzieLet29_1Lcall_kron_kron_Int_Int_Int2,CTkron_kron_Int_Int_Int) > [(es_3_1_destruct,Pointer_QTree_Int),
                                                                                                                      (sc_0_9_destruct,Pointer_CTkron_kron_Int_Int_Int),
                                                                                                                      (isZad2_3_destruct,MyDTInt_Bool),
                                                                                                                      (gad3_3_destruct,MyDTInt_Int_Int),
                                                                                                                      (q1ad7_2_destruct,Pointer_QTree_Int),
                                                                                                                      (m2ad5_3_destruct,Pointer_QTree_Int),
                                                                                                                      (q2ad8_2_destruct,Pointer_QTree_Int)] */
  logic [6:0] lizzieLet29_1Lcall_kron_kron_Int_Int_Int2_emitted;
  logic [6:0] lizzieLet29_1Lcall_kron_kron_Int_Int_Int2_done;
  assign es_3_1_destruct_d = {lizzieLet29_1Lcall_kron_kron_Int_Int_Int2_d[19:4],
                              (lizzieLet29_1Lcall_kron_kron_Int_Int_Int2_d[0] && (! lizzieLet29_1Lcall_kron_kron_Int_Int_Int2_emitted[0]))};
  assign sc_0_9_destruct_d = {lizzieLet29_1Lcall_kron_kron_Int_Int_Int2_d[35:20],
                              (lizzieLet29_1Lcall_kron_kron_Int_Int_Int2_d[0] && (! lizzieLet29_1Lcall_kron_kron_Int_Int_Int2_emitted[1]))};
  assign isZad2_3_destruct_d = (lizzieLet29_1Lcall_kron_kron_Int_Int_Int2_d[0] && (! lizzieLet29_1Lcall_kron_kron_Int_Int_Int2_emitted[2]));
  assign gad3_3_destruct_d = (lizzieLet29_1Lcall_kron_kron_Int_Int_Int2_d[0] && (! lizzieLet29_1Lcall_kron_kron_Int_Int_Int2_emitted[3]));
  assign q1ad7_2_destruct_d = {lizzieLet29_1Lcall_kron_kron_Int_Int_Int2_d[51:36],
                               (lizzieLet29_1Lcall_kron_kron_Int_Int_Int2_d[0] && (! lizzieLet29_1Lcall_kron_kron_Int_Int_Int2_emitted[4]))};
  assign m2ad5_3_destruct_d = {lizzieLet29_1Lcall_kron_kron_Int_Int_Int2_d[67:52],
                               (lizzieLet29_1Lcall_kron_kron_Int_Int_Int2_d[0] && (! lizzieLet29_1Lcall_kron_kron_Int_Int_Int2_emitted[5]))};
  assign q2ad8_2_destruct_d = {lizzieLet29_1Lcall_kron_kron_Int_Int_Int2_d[83:68],
                               (lizzieLet29_1Lcall_kron_kron_Int_Int_Int2_d[0] && (! lizzieLet29_1Lcall_kron_kron_Int_Int_Int2_emitted[6]))};
  assign lizzieLet29_1Lcall_kron_kron_Int_Int_Int2_done = (lizzieLet29_1Lcall_kron_kron_Int_Int_Int2_emitted | ({q2ad8_2_destruct_d[0],
                                                                                                                 m2ad5_3_destruct_d[0],
                                                                                                                 q1ad7_2_destruct_d[0],
                                                                                                                 gad3_3_destruct_d[0],
                                                                                                                 isZad2_3_destruct_d[0],
                                                                                                                 sc_0_9_destruct_d[0],
                                                                                                                 es_3_1_destruct_d[0]} & {q2ad8_2_destruct_r,
                                                                                                                                          m2ad5_3_destruct_r,
                                                                                                                                          q1ad7_2_destruct_r,
                                                                                                                                          gad3_3_destruct_r,
                                                                                                                                          isZad2_3_destruct_r,
                                                                                                                                          sc_0_9_destruct_r,
                                                                                                                                          es_3_1_destruct_r}));
  assign lizzieLet29_1Lcall_kron_kron_Int_Int_Int2_r = (& lizzieLet29_1Lcall_kron_kron_Int_Int_Int2_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet29_1Lcall_kron_kron_Int_Int_Int2_emitted <= 7'd0;
    else
      lizzieLet29_1Lcall_kron_kron_Int_Int_Int2_emitted <= (lizzieLet29_1Lcall_kron_kron_Int_Int_Int2_r ? 7'd0 :
                                                            lizzieLet29_1Lcall_kron_kron_Int_Int_Int2_done);
  
  /* destruct (Ty CTkron_kron_Int_Int_Int,
          Dcon Lcall_kron_kron_Int_Int_Int3) : (lizzieLet29_1Lcall_kron_kron_Int_Int_Int3,CTkron_kron_Int_Int_Int) > [(sc_0_8_destruct,Pointer_CTkron_kron_Int_Int_Int),
                                                                                                                      (isZad2_2_destruct,MyDTInt_Bool),
                                                                                                                      (gad3_2_destruct,MyDTInt_Int_Int),
                                                                                                                      (q1ad7_1_destruct,Pointer_QTree_Int),
                                                                                                                      (m2ad5_2_destruct,Pointer_QTree_Int),
                                                                                                                      (q2ad8_1_destruct,Pointer_QTree_Int),
                                                                                                                      (q3ad9_1_destruct,Pointer_QTree_Int)] */
  logic [6:0] lizzieLet29_1Lcall_kron_kron_Int_Int_Int3_emitted;
  logic [6:0] lizzieLet29_1Lcall_kron_kron_Int_Int_Int3_done;
  assign sc_0_8_destruct_d = {lizzieLet29_1Lcall_kron_kron_Int_Int_Int3_d[19:4],
                              (lizzieLet29_1Lcall_kron_kron_Int_Int_Int3_d[0] && (! lizzieLet29_1Lcall_kron_kron_Int_Int_Int3_emitted[0]))};
  assign isZad2_2_destruct_d = (lizzieLet29_1Lcall_kron_kron_Int_Int_Int3_d[0] && (! lizzieLet29_1Lcall_kron_kron_Int_Int_Int3_emitted[1]));
  assign gad3_2_destruct_d = (lizzieLet29_1Lcall_kron_kron_Int_Int_Int3_d[0] && (! lizzieLet29_1Lcall_kron_kron_Int_Int_Int3_emitted[2]));
  assign q1ad7_1_destruct_d = {lizzieLet29_1Lcall_kron_kron_Int_Int_Int3_d[35:20],
                               (lizzieLet29_1Lcall_kron_kron_Int_Int_Int3_d[0] && (! lizzieLet29_1Lcall_kron_kron_Int_Int_Int3_emitted[3]))};
  assign m2ad5_2_destruct_d = {lizzieLet29_1Lcall_kron_kron_Int_Int_Int3_d[51:36],
                               (lizzieLet29_1Lcall_kron_kron_Int_Int_Int3_d[0] && (! lizzieLet29_1Lcall_kron_kron_Int_Int_Int3_emitted[4]))};
  assign q2ad8_1_destruct_d = {lizzieLet29_1Lcall_kron_kron_Int_Int_Int3_d[67:52],
                               (lizzieLet29_1Lcall_kron_kron_Int_Int_Int3_d[0] && (! lizzieLet29_1Lcall_kron_kron_Int_Int_Int3_emitted[5]))};
  assign q3ad9_1_destruct_d = {lizzieLet29_1Lcall_kron_kron_Int_Int_Int3_d[83:68],
                               (lizzieLet29_1Lcall_kron_kron_Int_Int_Int3_d[0] && (! lizzieLet29_1Lcall_kron_kron_Int_Int_Int3_emitted[6]))};
  assign lizzieLet29_1Lcall_kron_kron_Int_Int_Int3_done = (lizzieLet29_1Lcall_kron_kron_Int_Int_Int3_emitted | ({q3ad9_1_destruct_d[0],
                                                                                                                 q2ad8_1_destruct_d[0],
                                                                                                                 m2ad5_2_destruct_d[0],
                                                                                                                 q1ad7_1_destruct_d[0],
                                                                                                                 gad3_2_destruct_d[0],
                                                                                                                 isZad2_2_destruct_d[0],
                                                                                                                 sc_0_8_destruct_d[0]} & {q3ad9_1_destruct_r,
                                                                                                                                          q2ad8_1_destruct_r,
                                                                                                                                          m2ad5_2_destruct_r,
                                                                                                                                          q1ad7_1_destruct_r,
                                                                                                                                          gad3_2_destruct_r,
                                                                                                                                          isZad2_2_destruct_r,
                                                                                                                                          sc_0_8_destruct_r}));
  assign lizzieLet29_1Lcall_kron_kron_Int_Int_Int3_r = (& lizzieLet29_1Lcall_kron_kron_Int_Int_Int3_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet29_1Lcall_kron_kron_Int_Int_Int3_emitted <= 7'd0;
    else
      lizzieLet29_1Lcall_kron_kron_Int_Int_Int3_emitted <= (lizzieLet29_1Lcall_kron_kron_Int_Int_Int3_r ? 7'd0 :
                                                            lizzieLet29_1Lcall_kron_kron_Int_Int_Int3_done);
  
  /* demux (Ty CTkron_kron_Int_Int_Int,
       Ty CTkron_kron_Int_Int_Int) : (lizzieLet29_2,CTkron_kron_Int_Int_Int) (lizzieLet29_1,CTkron_kron_Int_Int_Int) > [(_16,CTkron_kron_Int_Int_Int),
                                                                                                                        (lizzieLet29_1Lcall_kron_kron_Int_Int_Int3,CTkron_kron_Int_Int_Int),
                                                                                                                        (lizzieLet29_1Lcall_kron_kron_Int_Int_Int2,CTkron_kron_Int_Int_Int),
                                                                                                                        (lizzieLet29_1Lcall_kron_kron_Int_Int_Int1,CTkron_kron_Int_Int_Int),
                                                                                                                        (lizzieLet29_1Lcall_kron_kron_Int_Int_Int0,CTkron_kron_Int_Int_Int)] */
  logic [4:0] lizzieLet29_1_onehotd;
  always_comb
    if ((lizzieLet29_2_d[0] && lizzieLet29_1_d[0]))
      unique case (lizzieLet29_2_d[3:1])
        3'd0: lizzieLet29_1_onehotd = 5'd1;
        3'd1: lizzieLet29_1_onehotd = 5'd2;
        3'd2: lizzieLet29_1_onehotd = 5'd4;
        3'd3: lizzieLet29_1_onehotd = 5'd8;
        3'd4: lizzieLet29_1_onehotd = 5'd16;
        default: lizzieLet29_1_onehotd = 5'd0;
      endcase
    else lizzieLet29_1_onehotd = 5'd0;
  assign _16_d = {lizzieLet29_1_d[83:1], lizzieLet29_1_onehotd[0]};
  assign lizzieLet29_1Lcall_kron_kron_Int_Int_Int3_d = {lizzieLet29_1_d[83:1],
                                                        lizzieLet29_1_onehotd[1]};
  assign lizzieLet29_1Lcall_kron_kron_Int_Int_Int2_d = {lizzieLet29_1_d[83:1],
                                                        lizzieLet29_1_onehotd[2]};
  assign lizzieLet29_1Lcall_kron_kron_Int_Int_Int1_d = {lizzieLet29_1_d[83:1],
                                                        lizzieLet29_1_onehotd[3]};
  assign lizzieLet29_1Lcall_kron_kron_Int_Int_Int0_d = {lizzieLet29_1_d[83:1],
                                                        lizzieLet29_1_onehotd[4]};
  assign lizzieLet29_1_r = (| (lizzieLet29_1_onehotd & {lizzieLet29_1Lcall_kron_kron_Int_Int_Int0_r,
                                                        lizzieLet29_1Lcall_kron_kron_Int_Int_Int1_r,
                                                        lizzieLet29_1Lcall_kron_kron_Int_Int_Int2_r,
                                                        lizzieLet29_1Lcall_kron_kron_Int_Int_Int3_r,
                                                        _16_r}));
  assign lizzieLet29_2_r = lizzieLet29_1_r;
  
  /* demux (Ty CTkron_kron_Int_Int_Int,
       Ty Go) : (lizzieLet29_3,CTkron_kron_Int_Int_Int) (go_19_goMux_data,Go) > [(_15,Go),
                                                                                 (lizzieLet29_3Lcall_kron_kron_Int_Int_Int3,Go),
                                                                                 (lizzieLet29_3Lcall_kron_kron_Int_Int_Int2,Go),
                                                                                 (lizzieLet29_3Lcall_kron_kron_Int_Int_Int1,Go),
                                                                                 (lizzieLet29_3Lcall_kron_kron_Int_Int_Int0,Go)] */
  logic [4:0] go_19_goMux_data_onehotd;
  always_comb
    if ((lizzieLet29_3_d[0] && go_19_goMux_data_d[0]))
      unique case (lizzieLet29_3_d[3:1])
        3'd0: go_19_goMux_data_onehotd = 5'd1;
        3'd1: go_19_goMux_data_onehotd = 5'd2;
        3'd2: go_19_goMux_data_onehotd = 5'd4;
        3'd3: go_19_goMux_data_onehotd = 5'd8;
        3'd4: go_19_goMux_data_onehotd = 5'd16;
        default: go_19_goMux_data_onehotd = 5'd0;
      endcase
    else go_19_goMux_data_onehotd = 5'd0;
  assign _15_d = go_19_goMux_data_onehotd[0];
  assign lizzieLet29_3Lcall_kron_kron_Int_Int_Int3_d = go_19_goMux_data_onehotd[1];
  assign lizzieLet29_3Lcall_kron_kron_Int_Int_Int2_d = go_19_goMux_data_onehotd[2];
  assign lizzieLet29_3Lcall_kron_kron_Int_Int_Int1_d = go_19_goMux_data_onehotd[3];
  assign lizzieLet29_3Lcall_kron_kron_Int_Int_Int0_d = go_19_goMux_data_onehotd[4];
  assign go_19_goMux_data_r = (| (go_19_goMux_data_onehotd & {lizzieLet29_3Lcall_kron_kron_Int_Int_Int0_r,
                                                              lizzieLet29_3Lcall_kron_kron_Int_Int_Int1_r,
                                                              lizzieLet29_3Lcall_kron_kron_Int_Int_Int2_r,
                                                              lizzieLet29_3Lcall_kron_kron_Int_Int_Int3_r,
                                                              _15_r}));
  assign lizzieLet29_3_r = go_19_goMux_data_r;
  
  /* buf (Ty Go) : (lizzieLet29_3Lcall_kron_kron_Int_Int_Int0,Go) > (lizzieLet29_3Lcall_kron_kron_Int_Int_Int0_1_argbuf,Go) */
  Go_t lizzieLet29_3Lcall_kron_kron_Int_Int_Int0_bufchan_d;
  logic lizzieLet29_3Lcall_kron_kron_Int_Int_Int0_bufchan_r;
  assign lizzieLet29_3Lcall_kron_kron_Int_Int_Int0_r = ((! lizzieLet29_3Lcall_kron_kron_Int_Int_Int0_bufchan_d[0]) || lizzieLet29_3Lcall_kron_kron_Int_Int_Int0_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet29_3Lcall_kron_kron_Int_Int_Int0_bufchan_d <= 1'd0;
    else
      if (lizzieLet29_3Lcall_kron_kron_Int_Int_Int0_r)
        lizzieLet29_3Lcall_kron_kron_Int_Int_Int0_bufchan_d <= lizzieLet29_3Lcall_kron_kron_Int_Int_Int0_d;
  Go_t lizzieLet29_3Lcall_kron_kron_Int_Int_Int0_bufchan_buf;
  assign lizzieLet29_3Lcall_kron_kron_Int_Int_Int0_bufchan_r = (! lizzieLet29_3Lcall_kron_kron_Int_Int_Int0_bufchan_buf[0]);
  assign lizzieLet29_3Lcall_kron_kron_Int_Int_Int0_1_argbuf_d = (lizzieLet29_3Lcall_kron_kron_Int_Int_Int0_bufchan_buf[0] ? lizzieLet29_3Lcall_kron_kron_Int_Int_Int0_bufchan_buf :
                                                                 lizzieLet29_3Lcall_kron_kron_Int_Int_Int0_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet29_3Lcall_kron_kron_Int_Int_Int0_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet29_3Lcall_kron_kron_Int_Int_Int0_1_argbuf_r && lizzieLet29_3Lcall_kron_kron_Int_Int_Int0_bufchan_buf[0]))
        lizzieLet29_3Lcall_kron_kron_Int_Int_Int0_bufchan_buf <= 1'd0;
      else if (((! lizzieLet29_3Lcall_kron_kron_Int_Int_Int0_1_argbuf_r) && (! lizzieLet29_3Lcall_kron_kron_Int_Int_Int0_bufchan_buf[0])))
        lizzieLet29_3Lcall_kron_kron_Int_Int_Int0_bufchan_buf <= lizzieLet29_3Lcall_kron_kron_Int_Int_Int0_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet29_3Lcall_kron_kron_Int_Int_Int1,Go) > (lizzieLet29_3Lcall_kron_kron_Int_Int_Int1_1_argbuf,Go) */
  Go_t lizzieLet29_3Lcall_kron_kron_Int_Int_Int1_bufchan_d;
  logic lizzieLet29_3Lcall_kron_kron_Int_Int_Int1_bufchan_r;
  assign lizzieLet29_3Lcall_kron_kron_Int_Int_Int1_r = ((! lizzieLet29_3Lcall_kron_kron_Int_Int_Int1_bufchan_d[0]) || lizzieLet29_3Lcall_kron_kron_Int_Int_Int1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet29_3Lcall_kron_kron_Int_Int_Int1_bufchan_d <= 1'd0;
    else
      if (lizzieLet29_3Lcall_kron_kron_Int_Int_Int1_r)
        lizzieLet29_3Lcall_kron_kron_Int_Int_Int1_bufchan_d <= lizzieLet29_3Lcall_kron_kron_Int_Int_Int1_d;
  Go_t lizzieLet29_3Lcall_kron_kron_Int_Int_Int1_bufchan_buf;
  assign lizzieLet29_3Lcall_kron_kron_Int_Int_Int1_bufchan_r = (! lizzieLet29_3Lcall_kron_kron_Int_Int_Int1_bufchan_buf[0]);
  assign lizzieLet29_3Lcall_kron_kron_Int_Int_Int1_1_argbuf_d = (lizzieLet29_3Lcall_kron_kron_Int_Int_Int1_bufchan_buf[0] ? lizzieLet29_3Lcall_kron_kron_Int_Int_Int1_bufchan_buf :
                                                                 lizzieLet29_3Lcall_kron_kron_Int_Int_Int1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet29_3Lcall_kron_kron_Int_Int_Int1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet29_3Lcall_kron_kron_Int_Int_Int1_1_argbuf_r && lizzieLet29_3Lcall_kron_kron_Int_Int_Int1_bufchan_buf[0]))
        lizzieLet29_3Lcall_kron_kron_Int_Int_Int1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet29_3Lcall_kron_kron_Int_Int_Int1_1_argbuf_r) && (! lizzieLet29_3Lcall_kron_kron_Int_Int_Int1_bufchan_buf[0])))
        lizzieLet29_3Lcall_kron_kron_Int_Int_Int1_bufchan_buf <= lizzieLet29_3Lcall_kron_kron_Int_Int_Int1_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet29_3Lcall_kron_kron_Int_Int_Int2,Go) > (lizzieLet29_3Lcall_kron_kron_Int_Int_Int2_1_argbuf,Go) */
  Go_t lizzieLet29_3Lcall_kron_kron_Int_Int_Int2_bufchan_d;
  logic lizzieLet29_3Lcall_kron_kron_Int_Int_Int2_bufchan_r;
  assign lizzieLet29_3Lcall_kron_kron_Int_Int_Int2_r = ((! lizzieLet29_3Lcall_kron_kron_Int_Int_Int2_bufchan_d[0]) || lizzieLet29_3Lcall_kron_kron_Int_Int_Int2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet29_3Lcall_kron_kron_Int_Int_Int2_bufchan_d <= 1'd0;
    else
      if (lizzieLet29_3Lcall_kron_kron_Int_Int_Int2_r)
        lizzieLet29_3Lcall_kron_kron_Int_Int_Int2_bufchan_d <= lizzieLet29_3Lcall_kron_kron_Int_Int_Int2_d;
  Go_t lizzieLet29_3Lcall_kron_kron_Int_Int_Int2_bufchan_buf;
  assign lizzieLet29_3Lcall_kron_kron_Int_Int_Int2_bufchan_r = (! lizzieLet29_3Lcall_kron_kron_Int_Int_Int2_bufchan_buf[0]);
  assign lizzieLet29_3Lcall_kron_kron_Int_Int_Int2_1_argbuf_d = (lizzieLet29_3Lcall_kron_kron_Int_Int_Int2_bufchan_buf[0] ? lizzieLet29_3Lcall_kron_kron_Int_Int_Int2_bufchan_buf :
                                                                 lizzieLet29_3Lcall_kron_kron_Int_Int_Int2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet29_3Lcall_kron_kron_Int_Int_Int2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet29_3Lcall_kron_kron_Int_Int_Int2_1_argbuf_r && lizzieLet29_3Lcall_kron_kron_Int_Int_Int2_bufchan_buf[0]))
        lizzieLet29_3Lcall_kron_kron_Int_Int_Int2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet29_3Lcall_kron_kron_Int_Int_Int2_1_argbuf_r) && (! lizzieLet29_3Lcall_kron_kron_Int_Int_Int2_bufchan_buf[0])))
        lizzieLet29_3Lcall_kron_kron_Int_Int_Int2_bufchan_buf <= lizzieLet29_3Lcall_kron_kron_Int_Int_Int2_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet29_3Lcall_kron_kron_Int_Int_Int3,Go) > (lizzieLet29_3Lcall_kron_kron_Int_Int_Int3_1_argbuf,Go) */
  Go_t lizzieLet29_3Lcall_kron_kron_Int_Int_Int3_bufchan_d;
  logic lizzieLet29_3Lcall_kron_kron_Int_Int_Int3_bufchan_r;
  assign lizzieLet29_3Lcall_kron_kron_Int_Int_Int3_r = ((! lizzieLet29_3Lcall_kron_kron_Int_Int_Int3_bufchan_d[0]) || lizzieLet29_3Lcall_kron_kron_Int_Int_Int3_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet29_3Lcall_kron_kron_Int_Int_Int3_bufchan_d <= 1'd0;
    else
      if (lizzieLet29_3Lcall_kron_kron_Int_Int_Int3_r)
        lizzieLet29_3Lcall_kron_kron_Int_Int_Int3_bufchan_d <= lizzieLet29_3Lcall_kron_kron_Int_Int_Int3_d;
  Go_t lizzieLet29_3Lcall_kron_kron_Int_Int_Int3_bufchan_buf;
  assign lizzieLet29_3Lcall_kron_kron_Int_Int_Int3_bufchan_r = (! lizzieLet29_3Lcall_kron_kron_Int_Int_Int3_bufchan_buf[0]);
  assign lizzieLet29_3Lcall_kron_kron_Int_Int_Int3_1_argbuf_d = (lizzieLet29_3Lcall_kron_kron_Int_Int_Int3_bufchan_buf[0] ? lizzieLet29_3Lcall_kron_kron_Int_Int_Int3_bufchan_buf :
                                                                 lizzieLet29_3Lcall_kron_kron_Int_Int_Int3_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet29_3Lcall_kron_kron_Int_Int_Int3_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet29_3Lcall_kron_kron_Int_Int_Int3_1_argbuf_r && lizzieLet29_3Lcall_kron_kron_Int_Int_Int3_bufchan_buf[0]))
        lizzieLet29_3Lcall_kron_kron_Int_Int_Int3_bufchan_buf <= 1'd0;
      else if (((! lizzieLet29_3Lcall_kron_kron_Int_Int_Int3_1_argbuf_r) && (! lizzieLet29_3Lcall_kron_kron_Int_Int_Int3_bufchan_buf[0])))
        lizzieLet29_3Lcall_kron_kron_Int_Int_Int3_bufchan_buf <= lizzieLet29_3Lcall_kron_kron_Int_Int_Int3_bufchan_d;
  
  /* demux (Ty CTkron_kron_Int_Int_Int,
       Ty Pointer_QTree_Int) : (lizzieLet29_4,CTkron_kron_Int_Int_Int) (srtarg_0_1_goMux_mux,Pointer_QTree_Int) > [(lizzieLet29_4Lkron_kron_Int_Int_Intsbos,Pointer_QTree_Int),
                                                                                                                   (lizzieLet29_4Lcall_kron_kron_Int_Int_Int3,Pointer_QTree_Int),
                                                                                                                   (lizzieLet29_4Lcall_kron_kron_Int_Int_Int2,Pointer_QTree_Int),
                                                                                                                   (lizzieLet29_4Lcall_kron_kron_Int_Int_Int1,Pointer_QTree_Int),
                                                                                                                   (lizzieLet29_4Lcall_kron_kron_Int_Int_Int0,Pointer_QTree_Int)] */
  logic [4:0] srtarg_0_1_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet29_4_d[0] && srtarg_0_1_goMux_mux_d[0]))
      unique case (lizzieLet29_4_d[3:1])
        3'd0: srtarg_0_1_goMux_mux_onehotd = 5'd1;
        3'd1: srtarg_0_1_goMux_mux_onehotd = 5'd2;
        3'd2: srtarg_0_1_goMux_mux_onehotd = 5'd4;
        3'd3: srtarg_0_1_goMux_mux_onehotd = 5'd8;
        3'd4: srtarg_0_1_goMux_mux_onehotd = 5'd16;
        default: srtarg_0_1_goMux_mux_onehotd = 5'd0;
      endcase
    else srtarg_0_1_goMux_mux_onehotd = 5'd0;
  assign lizzieLet29_4Lkron_kron_Int_Int_Intsbos_d = {srtarg_0_1_goMux_mux_d[16:1],
                                                      srtarg_0_1_goMux_mux_onehotd[0]};
  assign lizzieLet29_4Lcall_kron_kron_Int_Int_Int3_d = {srtarg_0_1_goMux_mux_d[16:1],
                                                        srtarg_0_1_goMux_mux_onehotd[1]};
  assign lizzieLet29_4Lcall_kron_kron_Int_Int_Int2_d = {srtarg_0_1_goMux_mux_d[16:1],
                                                        srtarg_0_1_goMux_mux_onehotd[2]};
  assign lizzieLet29_4Lcall_kron_kron_Int_Int_Int1_d = {srtarg_0_1_goMux_mux_d[16:1],
                                                        srtarg_0_1_goMux_mux_onehotd[3]};
  assign lizzieLet29_4Lcall_kron_kron_Int_Int_Int0_d = {srtarg_0_1_goMux_mux_d[16:1],
                                                        srtarg_0_1_goMux_mux_onehotd[4]};
  assign srtarg_0_1_goMux_mux_r = (| (srtarg_0_1_goMux_mux_onehotd & {lizzieLet29_4Lcall_kron_kron_Int_Int_Int0_r,
                                                                      lizzieLet29_4Lcall_kron_kron_Int_Int_Int1_r,
                                                                      lizzieLet29_4Lcall_kron_kron_Int_Int_Int2_r,
                                                                      lizzieLet29_4Lcall_kron_kron_Int_Int_Int3_r,
                                                                      lizzieLet29_4Lkron_kron_Int_Int_Intsbos_r}));
  assign lizzieLet29_4_r = srtarg_0_1_goMux_mux_r;
  
  /* dcon (Ty QTree_Int,
      Dcon QNode_Int) : [(lizzieLet29_4Lcall_kron_kron_Int_Int_Int0,Pointer_QTree_Int),
                         (es_1_1_destruct,Pointer_QTree_Int),
                         (es_2_2_destruct,Pointer_QTree_Int),
                         (es_3_3_destruct,Pointer_QTree_Int)] > (lizzieLet29_4Lcall_kron_kron_Int_Int_Int0_1es_1_1_1es_2_2_1es_3_3_1QNode_Int,QTree_Int) */
  assign lizzieLet29_4Lcall_kron_kron_Int_Int_Int0_1es_1_1_1es_2_2_1es_3_3_1QNode_Int_d = QNode_Int_dc((& {lizzieLet29_4Lcall_kron_kron_Int_Int_Int0_d[0],
                                                                                                           es_1_1_destruct_d[0],
                                                                                                           es_2_2_destruct_d[0],
                                                                                                           es_3_3_destruct_d[0]}), lizzieLet29_4Lcall_kron_kron_Int_Int_Int0_d, es_1_1_destruct_d, es_2_2_destruct_d, es_3_3_destruct_d);
  assign {lizzieLet29_4Lcall_kron_kron_Int_Int_Int0_r,
          es_1_1_destruct_r,
          es_2_2_destruct_r,
          es_3_3_destruct_r} = {4 {(lizzieLet29_4Lcall_kron_kron_Int_Int_Int0_1es_1_1_1es_2_2_1es_3_3_1QNode_Int_r && lizzieLet29_4Lcall_kron_kron_Int_Int_Int0_1es_1_1_1es_2_2_1es_3_3_1QNode_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (lizzieLet29_4Lcall_kron_kron_Int_Int_Int0_1es_1_1_1es_2_2_1es_3_3_1QNode_Int,QTree_Int) > (lizzieLet33_1_argbuf,QTree_Int) */
  QTree_Int_t lizzieLet29_4Lcall_kron_kron_Int_Int_Int0_1es_1_1_1es_2_2_1es_3_3_1QNode_Int_bufchan_d;
  logic lizzieLet29_4Lcall_kron_kron_Int_Int_Int0_1es_1_1_1es_2_2_1es_3_3_1QNode_Int_bufchan_r;
  assign lizzieLet29_4Lcall_kron_kron_Int_Int_Int0_1es_1_1_1es_2_2_1es_3_3_1QNode_Int_r = ((! lizzieLet29_4Lcall_kron_kron_Int_Int_Int0_1es_1_1_1es_2_2_1es_3_3_1QNode_Int_bufchan_d[0]) || lizzieLet29_4Lcall_kron_kron_Int_Int_Int0_1es_1_1_1es_2_2_1es_3_3_1QNode_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet29_4Lcall_kron_kron_Int_Int_Int0_1es_1_1_1es_2_2_1es_3_3_1QNode_Int_bufchan_d <= {66'd0,
                                                                                                 1'd0};
    else
      if (lizzieLet29_4Lcall_kron_kron_Int_Int_Int0_1es_1_1_1es_2_2_1es_3_3_1QNode_Int_r)
        lizzieLet29_4Lcall_kron_kron_Int_Int_Int0_1es_1_1_1es_2_2_1es_3_3_1QNode_Int_bufchan_d <= lizzieLet29_4Lcall_kron_kron_Int_Int_Int0_1es_1_1_1es_2_2_1es_3_3_1QNode_Int_d;
  QTree_Int_t lizzieLet29_4Lcall_kron_kron_Int_Int_Int0_1es_1_1_1es_2_2_1es_3_3_1QNode_Int_bufchan_buf;
  assign lizzieLet29_4Lcall_kron_kron_Int_Int_Int0_1es_1_1_1es_2_2_1es_3_3_1QNode_Int_bufchan_r = (! lizzieLet29_4Lcall_kron_kron_Int_Int_Int0_1es_1_1_1es_2_2_1es_3_3_1QNode_Int_bufchan_buf[0]);
  assign lizzieLet33_1_argbuf_d = (lizzieLet29_4Lcall_kron_kron_Int_Int_Int0_1es_1_1_1es_2_2_1es_3_3_1QNode_Int_bufchan_buf[0] ? lizzieLet29_4Lcall_kron_kron_Int_Int_Int0_1es_1_1_1es_2_2_1es_3_3_1QNode_Int_bufchan_buf :
                                   lizzieLet29_4Lcall_kron_kron_Int_Int_Int0_1es_1_1_1es_2_2_1es_3_3_1QNode_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet29_4Lcall_kron_kron_Int_Int_Int0_1es_1_1_1es_2_2_1es_3_3_1QNode_Int_bufchan_buf <= {66'd0,
                                                                                                   1'd0};
    else
      if ((lizzieLet33_1_argbuf_r && lizzieLet29_4Lcall_kron_kron_Int_Int_Int0_1es_1_1_1es_2_2_1es_3_3_1QNode_Int_bufchan_buf[0]))
        lizzieLet29_4Lcall_kron_kron_Int_Int_Int0_1es_1_1_1es_2_2_1es_3_3_1QNode_Int_bufchan_buf <= {66'd0,
                                                                                                     1'd0};
      else if (((! lizzieLet33_1_argbuf_r) && (! lizzieLet29_4Lcall_kron_kron_Int_Int_Int0_1es_1_1_1es_2_2_1es_3_3_1QNode_Int_bufchan_buf[0])))
        lizzieLet29_4Lcall_kron_kron_Int_Int_Int0_1es_1_1_1es_2_2_1es_3_3_1QNode_Int_bufchan_buf <= lizzieLet29_4Lcall_kron_kron_Int_Int_Int0_1es_1_1_1es_2_2_1es_3_3_1QNode_Int_bufchan_d;
  
  /* dcon (Ty CTkron_kron_Int_Int_Int,
      Dcon Lcall_kron_kron_Int_Int_Int0) : [(lizzieLet29_4Lcall_kron_kron_Int_Int_Int1,Pointer_QTree_Int),
                                            (es_2_1_destruct,Pointer_QTree_Int),
                                            (es_3_2_destruct,Pointer_QTree_Int),
                                            (sc_0_10_destruct,Pointer_CTkron_kron_Int_Int_Int)] > (lizzieLet29_4Lcall_kron_kron_Int_Int_Int1_1es_2_1_1es_3_2_1sc_0_10_1Lcall_kron_kron_Int_Int_Int0,CTkron_kron_Int_Int_Int) */
  assign lizzieLet29_4Lcall_kron_kron_Int_Int_Int1_1es_2_1_1es_3_2_1sc_0_10_1Lcall_kron_kron_Int_Int_Int0_d = Lcall_kron_kron_Int_Int_Int0_dc((& {lizzieLet29_4Lcall_kron_kron_Int_Int_Int1_d[0],
                                                                                                                                                  es_2_1_destruct_d[0],
                                                                                                                                                  es_3_2_destruct_d[0],
                                                                                                                                                  sc_0_10_destruct_d[0]}), lizzieLet29_4Lcall_kron_kron_Int_Int_Int1_d, es_2_1_destruct_d, es_3_2_destruct_d, sc_0_10_destruct_d);
  assign {lizzieLet29_4Lcall_kron_kron_Int_Int_Int1_r,
          es_2_1_destruct_r,
          es_3_2_destruct_r,
          sc_0_10_destruct_r} = {4 {(lizzieLet29_4Lcall_kron_kron_Int_Int_Int1_1es_2_1_1es_3_2_1sc_0_10_1Lcall_kron_kron_Int_Int_Int0_r && lizzieLet29_4Lcall_kron_kron_Int_Int_Int1_1es_2_1_1es_3_2_1sc_0_10_1Lcall_kron_kron_Int_Int_Int0_d[0])}};
  
  /* buf (Ty CTkron_kron_Int_Int_Int) : (lizzieLet29_4Lcall_kron_kron_Int_Int_Int1_1es_2_1_1es_3_2_1sc_0_10_1Lcall_kron_kron_Int_Int_Int0,CTkron_kron_Int_Int_Int) > (lizzieLet32_1_argbuf,CTkron_kron_Int_Int_Int) */
  CTkron_kron_Int_Int_Int_t lizzieLet29_4Lcall_kron_kron_Int_Int_Int1_1es_2_1_1es_3_2_1sc_0_10_1Lcall_kron_kron_Int_Int_Int0_bufchan_d;
  logic lizzieLet29_4Lcall_kron_kron_Int_Int_Int1_1es_2_1_1es_3_2_1sc_0_10_1Lcall_kron_kron_Int_Int_Int0_bufchan_r;
  assign lizzieLet29_4Lcall_kron_kron_Int_Int_Int1_1es_2_1_1es_3_2_1sc_0_10_1Lcall_kron_kron_Int_Int_Int0_r = ((! lizzieLet29_4Lcall_kron_kron_Int_Int_Int1_1es_2_1_1es_3_2_1sc_0_10_1Lcall_kron_kron_Int_Int_Int0_bufchan_d[0]) || lizzieLet29_4Lcall_kron_kron_Int_Int_Int1_1es_2_1_1es_3_2_1sc_0_10_1Lcall_kron_kron_Int_Int_Int0_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet29_4Lcall_kron_kron_Int_Int_Int1_1es_2_1_1es_3_2_1sc_0_10_1Lcall_kron_kron_Int_Int_Int0_bufchan_d <= {83'd0,
                                                                                                                     1'd0};
    else
      if (lizzieLet29_4Lcall_kron_kron_Int_Int_Int1_1es_2_1_1es_3_2_1sc_0_10_1Lcall_kron_kron_Int_Int_Int0_r)
        lizzieLet29_4Lcall_kron_kron_Int_Int_Int1_1es_2_1_1es_3_2_1sc_0_10_1Lcall_kron_kron_Int_Int_Int0_bufchan_d <= lizzieLet29_4Lcall_kron_kron_Int_Int_Int1_1es_2_1_1es_3_2_1sc_0_10_1Lcall_kron_kron_Int_Int_Int0_d;
  CTkron_kron_Int_Int_Int_t lizzieLet29_4Lcall_kron_kron_Int_Int_Int1_1es_2_1_1es_3_2_1sc_0_10_1Lcall_kron_kron_Int_Int_Int0_bufchan_buf;
  assign lizzieLet29_4Lcall_kron_kron_Int_Int_Int1_1es_2_1_1es_3_2_1sc_0_10_1Lcall_kron_kron_Int_Int_Int0_bufchan_r = (! lizzieLet29_4Lcall_kron_kron_Int_Int_Int1_1es_2_1_1es_3_2_1sc_0_10_1Lcall_kron_kron_Int_Int_Int0_bufchan_buf[0]);
  assign lizzieLet32_1_argbuf_d = (lizzieLet29_4Lcall_kron_kron_Int_Int_Int1_1es_2_1_1es_3_2_1sc_0_10_1Lcall_kron_kron_Int_Int_Int0_bufchan_buf[0] ? lizzieLet29_4Lcall_kron_kron_Int_Int_Int1_1es_2_1_1es_3_2_1sc_0_10_1Lcall_kron_kron_Int_Int_Int0_bufchan_buf :
                                   lizzieLet29_4Lcall_kron_kron_Int_Int_Int1_1es_2_1_1es_3_2_1sc_0_10_1Lcall_kron_kron_Int_Int_Int0_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet29_4Lcall_kron_kron_Int_Int_Int1_1es_2_1_1es_3_2_1sc_0_10_1Lcall_kron_kron_Int_Int_Int0_bufchan_buf <= {83'd0,
                                                                                                                       1'd0};
    else
      if ((lizzieLet32_1_argbuf_r && lizzieLet29_4Lcall_kron_kron_Int_Int_Int1_1es_2_1_1es_3_2_1sc_0_10_1Lcall_kron_kron_Int_Int_Int0_bufchan_buf[0]))
        lizzieLet29_4Lcall_kron_kron_Int_Int_Int1_1es_2_1_1es_3_2_1sc_0_10_1Lcall_kron_kron_Int_Int_Int0_bufchan_buf <= {83'd0,
                                                                                                                         1'd0};
      else if (((! lizzieLet32_1_argbuf_r) && (! lizzieLet29_4Lcall_kron_kron_Int_Int_Int1_1es_2_1_1es_3_2_1sc_0_10_1Lcall_kron_kron_Int_Int_Int0_bufchan_buf[0])))
        lizzieLet29_4Lcall_kron_kron_Int_Int_Int1_1es_2_1_1es_3_2_1sc_0_10_1Lcall_kron_kron_Int_Int_Int0_bufchan_buf <= lizzieLet29_4Lcall_kron_kron_Int_Int_Int1_1es_2_1_1es_3_2_1sc_0_10_1Lcall_kron_kron_Int_Int_Int0_bufchan_d;
  
  /* dcon (Ty CTkron_kron_Int_Int_Int,
      Dcon Lcall_kron_kron_Int_Int_Int1) : [(lizzieLet29_4Lcall_kron_kron_Int_Int_Int2,Pointer_QTree_Int),
                                            (es_3_1_destruct,Pointer_QTree_Int),
                                            (sc_0_9_destruct,Pointer_CTkron_kron_Int_Int_Int),
                                            (isZad2_3_1,MyDTInt_Bool),
                                            (gad3_3_1,MyDTInt_Int_Int),
                                            (q1ad7_2_destruct,Pointer_QTree_Int),
                                            (m2ad5_3_1,Pointer_QTree_Int)] > (lizzieLet29_4Lcall_kron_kron_Int_Int_Int2_1es_3_1_1sc_0_9_1isZad2_3_1gad3_3_1q1ad7_2_1m2ad5_3_1Lcall_kron_kron_Int_Int_Int1,CTkron_kron_Int_Int_Int) */
  assign lizzieLet29_4Lcall_kron_kron_Int_Int_Int2_1es_3_1_1sc_0_9_1isZad2_3_1gad3_3_1q1ad7_2_1m2ad5_3_1Lcall_kron_kron_Int_Int_Int1_d = Lcall_kron_kron_Int_Int_Int1_dc((& {lizzieLet29_4Lcall_kron_kron_Int_Int_Int2_d[0],
                                                                                                                                                                             es_3_1_destruct_d[0],
                                                                                                                                                                             sc_0_9_destruct_d[0],
                                                                                                                                                                             isZad2_3_1_d[0],
                                                                                                                                                                             gad3_3_1_d[0],
                                                                                                                                                                             q1ad7_2_destruct_d[0],
                                                                                                                                                                             m2ad5_3_1_d[0]}), lizzieLet29_4Lcall_kron_kron_Int_Int_Int2_d, es_3_1_destruct_d, sc_0_9_destruct_d, isZad2_3_1_d, gad3_3_1_d, q1ad7_2_destruct_d, m2ad5_3_1_d);
  assign {lizzieLet29_4Lcall_kron_kron_Int_Int_Int2_r,
          es_3_1_destruct_r,
          sc_0_9_destruct_r,
          isZad2_3_1_r,
          gad3_3_1_r,
          q1ad7_2_destruct_r,
          m2ad5_3_1_r} = {7 {(lizzieLet29_4Lcall_kron_kron_Int_Int_Int2_1es_3_1_1sc_0_9_1isZad2_3_1gad3_3_1q1ad7_2_1m2ad5_3_1Lcall_kron_kron_Int_Int_Int1_r && lizzieLet29_4Lcall_kron_kron_Int_Int_Int2_1es_3_1_1sc_0_9_1isZad2_3_1gad3_3_1q1ad7_2_1m2ad5_3_1Lcall_kron_kron_Int_Int_Int1_d[0])}};
  
  /* buf (Ty CTkron_kron_Int_Int_Int) : (lizzieLet29_4Lcall_kron_kron_Int_Int_Int2_1es_3_1_1sc_0_9_1isZad2_3_1gad3_3_1q1ad7_2_1m2ad5_3_1Lcall_kron_kron_Int_Int_Int1,CTkron_kron_Int_Int_Int) > (lizzieLet31_1_argbuf,CTkron_kron_Int_Int_Int) */
  CTkron_kron_Int_Int_Int_t lizzieLet29_4Lcall_kron_kron_Int_Int_Int2_1es_3_1_1sc_0_9_1isZad2_3_1gad3_3_1q1ad7_2_1m2ad5_3_1Lcall_kron_kron_Int_Int_Int1_bufchan_d;
  logic lizzieLet29_4Lcall_kron_kron_Int_Int_Int2_1es_3_1_1sc_0_9_1isZad2_3_1gad3_3_1q1ad7_2_1m2ad5_3_1Lcall_kron_kron_Int_Int_Int1_bufchan_r;
  assign lizzieLet29_4Lcall_kron_kron_Int_Int_Int2_1es_3_1_1sc_0_9_1isZad2_3_1gad3_3_1q1ad7_2_1m2ad5_3_1Lcall_kron_kron_Int_Int_Int1_r = ((! lizzieLet29_4Lcall_kron_kron_Int_Int_Int2_1es_3_1_1sc_0_9_1isZad2_3_1gad3_3_1q1ad7_2_1m2ad5_3_1Lcall_kron_kron_Int_Int_Int1_bufchan_d[0]) || lizzieLet29_4Lcall_kron_kron_Int_Int_Int2_1es_3_1_1sc_0_9_1isZad2_3_1gad3_3_1q1ad7_2_1m2ad5_3_1Lcall_kron_kron_Int_Int_Int1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet29_4Lcall_kron_kron_Int_Int_Int2_1es_3_1_1sc_0_9_1isZad2_3_1gad3_3_1q1ad7_2_1m2ad5_3_1Lcall_kron_kron_Int_Int_Int1_bufchan_d <= {83'd0,
                                                                                                                                                1'd0};
    else
      if (lizzieLet29_4Lcall_kron_kron_Int_Int_Int2_1es_3_1_1sc_0_9_1isZad2_3_1gad3_3_1q1ad7_2_1m2ad5_3_1Lcall_kron_kron_Int_Int_Int1_r)
        lizzieLet29_4Lcall_kron_kron_Int_Int_Int2_1es_3_1_1sc_0_9_1isZad2_3_1gad3_3_1q1ad7_2_1m2ad5_3_1Lcall_kron_kron_Int_Int_Int1_bufchan_d <= lizzieLet29_4Lcall_kron_kron_Int_Int_Int2_1es_3_1_1sc_0_9_1isZad2_3_1gad3_3_1q1ad7_2_1m2ad5_3_1Lcall_kron_kron_Int_Int_Int1_d;
  CTkron_kron_Int_Int_Int_t lizzieLet29_4Lcall_kron_kron_Int_Int_Int2_1es_3_1_1sc_0_9_1isZad2_3_1gad3_3_1q1ad7_2_1m2ad5_3_1Lcall_kron_kron_Int_Int_Int1_bufchan_buf;
  assign lizzieLet29_4Lcall_kron_kron_Int_Int_Int2_1es_3_1_1sc_0_9_1isZad2_3_1gad3_3_1q1ad7_2_1m2ad5_3_1Lcall_kron_kron_Int_Int_Int1_bufchan_r = (! lizzieLet29_4Lcall_kron_kron_Int_Int_Int2_1es_3_1_1sc_0_9_1isZad2_3_1gad3_3_1q1ad7_2_1m2ad5_3_1Lcall_kron_kron_Int_Int_Int1_bufchan_buf[0]);
  assign lizzieLet31_1_argbuf_d = (lizzieLet29_4Lcall_kron_kron_Int_Int_Int2_1es_3_1_1sc_0_9_1isZad2_3_1gad3_3_1q1ad7_2_1m2ad5_3_1Lcall_kron_kron_Int_Int_Int1_bufchan_buf[0] ? lizzieLet29_4Lcall_kron_kron_Int_Int_Int2_1es_3_1_1sc_0_9_1isZad2_3_1gad3_3_1q1ad7_2_1m2ad5_3_1Lcall_kron_kron_Int_Int_Int1_bufchan_buf :
                                   lizzieLet29_4Lcall_kron_kron_Int_Int_Int2_1es_3_1_1sc_0_9_1isZad2_3_1gad3_3_1q1ad7_2_1m2ad5_3_1Lcall_kron_kron_Int_Int_Int1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet29_4Lcall_kron_kron_Int_Int_Int2_1es_3_1_1sc_0_9_1isZad2_3_1gad3_3_1q1ad7_2_1m2ad5_3_1Lcall_kron_kron_Int_Int_Int1_bufchan_buf <= {83'd0,
                                                                                                                                                  1'd0};
    else
      if ((lizzieLet31_1_argbuf_r && lizzieLet29_4Lcall_kron_kron_Int_Int_Int2_1es_3_1_1sc_0_9_1isZad2_3_1gad3_3_1q1ad7_2_1m2ad5_3_1Lcall_kron_kron_Int_Int_Int1_bufchan_buf[0]))
        lizzieLet29_4Lcall_kron_kron_Int_Int_Int2_1es_3_1_1sc_0_9_1isZad2_3_1gad3_3_1q1ad7_2_1m2ad5_3_1Lcall_kron_kron_Int_Int_Int1_bufchan_buf <= {83'd0,
                                                                                                                                                    1'd0};
      else if (((! lizzieLet31_1_argbuf_r) && (! lizzieLet29_4Lcall_kron_kron_Int_Int_Int2_1es_3_1_1sc_0_9_1isZad2_3_1gad3_3_1q1ad7_2_1m2ad5_3_1Lcall_kron_kron_Int_Int_Int1_bufchan_buf[0])))
        lizzieLet29_4Lcall_kron_kron_Int_Int_Int2_1es_3_1_1sc_0_9_1isZad2_3_1gad3_3_1q1ad7_2_1m2ad5_3_1Lcall_kron_kron_Int_Int_Int1_bufchan_buf <= lizzieLet29_4Lcall_kron_kron_Int_Int_Int2_1es_3_1_1sc_0_9_1isZad2_3_1gad3_3_1q1ad7_2_1m2ad5_3_1Lcall_kron_kron_Int_Int_Int1_bufchan_d;
  
  /* dcon (Ty CTkron_kron_Int_Int_Int,
      Dcon Lcall_kron_kron_Int_Int_Int2) : [(lizzieLet29_4Lcall_kron_kron_Int_Int_Int3,Pointer_QTree_Int),
                                            (sc_0_8_destruct,Pointer_CTkron_kron_Int_Int_Int),
                                            (isZad2_2_1,MyDTInt_Bool),
                                            (gad3_2_1,MyDTInt_Int_Int),
                                            (q1ad7_1_destruct,Pointer_QTree_Int),
                                            (m2ad5_2_1,Pointer_QTree_Int),
                                            (q2ad8_1_destruct,Pointer_QTree_Int)] > (lizzieLet29_4Lcall_kron_kron_Int_Int_Int3_1sc_0_8_1isZad2_2_1gad3_2_1q1ad7_1_1m2ad5_2_1q2ad8_1_1Lcall_kron_kron_Int_Int_Int2,CTkron_kron_Int_Int_Int) */
  assign lizzieLet29_4Lcall_kron_kron_Int_Int_Int3_1sc_0_8_1isZad2_2_1gad3_2_1q1ad7_1_1m2ad5_2_1q2ad8_1_1Lcall_kron_kron_Int_Int_Int2_d = Lcall_kron_kron_Int_Int_Int2_dc((& {lizzieLet29_4Lcall_kron_kron_Int_Int_Int3_d[0],
                                                                                                                                                                              sc_0_8_destruct_d[0],
                                                                                                                                                                              isZad2_2_1_d[0],
                                                                                                                                                                              gad3_2_1_d[0],
                                                                                                                                                                              q1ad7_1_destruct_d[0],
                                                                                                                                                                              m2ad5_2_1_d[0],
                                                                                                                                                                              q2ad8_1_destruct_d[0]}), lizzieLet29_4Lcall_kron_kron_Int_Int_Int3_d, sc_0_8_destruct_d, isZad2_2_1_d, gad3_2_1_d, q1ad7_1_destruct_d, m2ad5_2_1_d, q2ad8_1_destruct_d);
  assign {lizzieLet29_4Lcall_kron_kron_Int_Int_Int3_r,
          sc_0_8_destruct_r,
          isZad2_2_1_r,
          gad3_2_1_r,
          q1ad7_1_destruct_r,
          m2ad5_2_1_r,
          q2ad8_1_destruct_r} = {7 {(lizzieLet29_4Lcall_kron_kron_Int_Int_Int3_1sc_0_8_1isZad2_2_1gad3_2_1q1ad7_1_1m2ad5_2_1q2ad8_1_1Lcall_kron_kron_Int_Int_Int2_r && lizzieLet29_4Lcall_kron_kron_Int_Int_Int3_1sc_0_8_1isZad2_2_1gad3_2_1q1ad7_1_1m2ad5_2_1q2ad8_1_1Lcall_kron_kron_Int_Int_Int2_d[0])}};
  
  /* buf (Ty CTkron_kron_Int_Int_Int) : (lizzieLet29_4Lcall_kron_kron_Int_Int_Int3_1sc_0_8_1isZad2_2_1gad3_2_1q1ad7_1_1m2ad5_2_1q2ad8_1_1Lcall_kron_kron_Int_Int_Int2,CTkron_kron_Int_Int_Int) > (lizzieLet30_1_argbuf,CTkron_kron_Int_Int_Int) */
  CTkron_kron_Int_Int_Int_t lizzieLet29_4Lcall_kron_kron_Int_Int_Int3_1sc_0_8_1isZad2_2_1gad3_2_1q1ad7_1_1m2ad5_2_1q2ad8_1_1Lcall_kron_kron_Int_Int_Int2_bufchan_d;
  logic lizzieLet29_4Lcall_kron_kron_Int_Int_Int3_1sc_0_8_1isZad2_2_1gad3_2_1q1ad7_1_1m2ad5_2_1q2ad8_1_1Lcall_kron_kron_Int_Int_Int2_bufchan_r;
  assign lizzieLet29_4Lcall_kron_kron_Int_Int_Int3_1sc_0_8_1isZad2_2_1gad3_2_1q1ad7_1_1m2ad5_2_1q2ad8_1_1Lcall_kron_kron_Int_Int_Int2_r = ((! lizzieLet29_4Lcall_kron_kron_Int_Int_Int3_1sc_0_8_1isZad2_2_1gad3_2_1q1ad7_1_1m2ad5_2_1q2ad8_1_1Lcall_kron_kron_Int_Int_Int2_bufchan_d[0]) || lizzieLet29_4Lcall_kron_kron_Int_Int_Int3_1sc_0_8_1isZad2_2_1gad3_2_1q1ad7_1_1m2ad5_2_1q2ad8_1_1Lcall_kron_kron_Int_Int_Int2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet29_4Lcall_kron_kron_Int_Int_Int3_1sc_0_8_1isZad2_2_1gad3_2_1q1ad7_1_1m2ad5_2_1q2ad8_1_1Lcall_kron_kron_Int_Int_Int2_bufchan_d <= {83'd0,
                                                                                                                                                 1'd0};
    else
      if (lizzieLet29_4Lcall_kron_kron_Int_Int_Int3_1sc_0_8_1isZad2_2_1gad3_2_1q1ad7_1_1m2ad5_2_1q2ad8_1_1Lcall_kron_kron_Int_Int_Int2_r)
        lizzieLet29_4Lcall_kron_kron_Int_Int_Int3_1sc_0_8_1isZad2_2_1gad3_2_1q1ad7_1_1m2ad5_2_1q2ad8_1_1Lcall_kron_kron_Int_Int_Int2_bufchan_d <= lizzieLet29_4Lcall_kron_kron_Int_Int_Int3_1sc_0_8_1isZad2_2_1gad3_2_1q1ad7_1_1m2ad5_2_1q2ad8_1_1Lcall_kron_kron_Int_Int_Int2_d;
  CTkron_kron_Int_Int_Int_t lizzieLet29_4Lcall_kron_kron_Int_Int_Int3_1sc_0_8_1isZad2_2_1gad3_2_1q1ad7_1_1m2ad5_2_1q2ad8_1_1Lcall_kron_kron_Int_Int_Int2_bufchan_buf;
  assign lizzieLet29_4Lcall_kron_kron_Int_Int_Int3_1sc_0_8_1isZad2_2_1gad3_2_1q1ad7_1_1m2ad5_2_1q2ad8_1_1Lcall_kron_kron_Int_Int_Int2_bufchan_r = (! lizzieLet29_4Lcall_kron_kron_Int_Int_Int3_1sc_0_8_1isZad2_2_1gad3_2_1q1ad7_1_1m2ad5_2_1q2ad8_1_1Lcall_kron_kron_Int_Int_Int2_bufchan_buf[0]);
  assign lizzieLet30_1_argbuf_d = (lizzieLet29_4Lcall_kron_kron_Int_Int_Int3_1sc_0_8_1isZad2_2_1gad3_2_1q1ad7_1_1m2ad5_2_1q2ad8_1_1Lcall_kron_kron_Int_Int_Int2_bufchan_buf[0] ? lizzieLet29_4Lcall_kron_kron_Int_Int_Int3_1sc_0_8_1isZad2_2_1gad3_2_1q1ad7_1_1m2ad5_2_1q2ad8_1_1Lcall_kron_kron_Int_Int_Int2_bufchan_buf :
                                   lizzieLet29_4Lcall_kron_kron_Int_Int_Int3_1sc_0_8_1isZad2_2_1gad3_2_1q1ad7_1_1m2ad5_2_1q2ad8_1_1Lcall_kron_kron_Int_Int_Int2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet29_4Lcall_kron_kron_Int_Int_Int3_1sc_0_8_1isZad2_2_1gad3_2_1q1ad7_1_1m2ad5_2_1q2ad8_1_1Lcall_kron_kron_Int_Int_Int2_bufchan_buf <= {83'd0,
                                                                                                                                                   1'd0};
    else
      if ((lizzieLet30_1_argbuf_r && lizzieLet29_4Lcall_kron_kron_Int_Int_Int3_1sc_0_8_1isZad2_2_1gad3_2_1q1ad7_1_1m2ad5_2_1q2ad8_1_1Lcall_kron_kron_Int_Int_Int2_bufchan_buf[0]))
        lizzieLet29_4Lcall_kron_kron_Int_Int_Int3_1sc_0_8_1isZad2_2_1gad3_2_1q1ad7_1_1m2ad5_2_1q2ad8_1_1Lcall_kron_kron_Int_Int_Int2_bufchan_buf <= {83'd0,
                                                                                                                                                     1'd0};
      else if (((! lizzieLet30_1_argbuf_r) && (! lizzieLet29_4Lcall_kron_kron_Int_Int_Int3_1sc_0_8_1isZad2_2_1gad3_2_1q1ad7_1_1m2ad5_2_1q2ad8_1_1Lcall_kron_kron_Int_Int_Int2_bufchan_buf[0])))
        lizzieLet29_4Lcall_kron_kron_Int_Int_Int3_1sc_0_8_1isZad2_2_1gad3_2_1q1ad7_1_1m2ad5_2_1q2ad8_1_1Lcall_kron_kron_Int_Int_Int2_bufchan_buf <= lizzieLet29_4Lcall_kron_kron_Int_Int_Int3_1sc_0_8_1isZad2_2_1gad3_2_1q1ad7_1_1m2ad5_2_1q2ad8_1_1Lcall_kron_kron_Int_Int_Int2_bufchan_d;
  
  /* fork (Ty Pointer_QTree_Int) : (lizzieLet29_4Lkron_kron_Int_Int_Intsbos,Pointer_QTree_Int) > [(lizzieLet29_4Lkron_kron_Int_Int_Intsbos_1_merge_merge_fork_1,Pointer_QTree_Int),
                                                                                             (lizzieLet29_4Lkron_kron_Int_Int_Intsbos_1_merge_merge_fork_2,Pointer_QTree_Int)] */
  logic [1:0] lizzieLet29_4Lkron_kron_Int_Int_Intsbos_emitted;
  logic [1:0] lizzieLet29_4Lkron_kron_Int_Int_Intsbos_done;
  assign lizzieLet29_4Lkron_kron_Int_Int_Intsbos_1_merge_merge_fork_1_d = {lizzieLet29_4Lkron_kron_Int_Int_Intsbos_d[16:1],
                                                                           (lizzieLet29_4Lkron_kron_Int_Int_Intsbos_d[0] && (! lizzieLet29_4Lkron_kron_Int_Int_Intsbos_emitted[0]))};
  assign lizzieLet29_4Lkron_kron_Int_Int_Intsbos_1_merge_merge_fork_2_d = {lizzieLet29_4Lkron_kron_Int_Int_Intsbos_d[16:1],
                                                                           (lizzieLet29_4Lkron_kron_Int_Int_Intsbos_d[0] && (! lizzieLet29_4Lkron_kron_Int_Int_Intsbos_emitted[1]))};
  assign lizzieLet29_4Lkron_kron_Int_Int_Intsbos_done = (lizzieLet29_4Lkron_kron_Int_Int_Intsbos_emitted | ({lizzieLet29_4Lkron_kron_Int_Int_Intsbos_1_merge_merge_fork_2_d[0],
                                                                                                             lizzieLet29_4Lkron_kron_Int_Int_Intsbos_1_merge_merge_fork_1_d[0]} & {lizzieLet29_4Lkron_kron_Int_Int_Intsbos_1_merge_merge_fork_2_r,
                                                                                                                                                                                   lizzieLet29_4Lkron_kron_Int_Int_Intsbos_1_merge_merge_fork_1_r}));
  assign lizzieLet29_4Lkron_kron_Int_Int_Intsbos_r = (& lizzieLet29_4Lkron_kron_Int_Int_Intsbos_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet29_4Lkron_kron_Int_Int_Intsbos_emitted <= 2'd0;
    else
      lizzieLet29_4Lkron_kron_Int_Int_Intsbos_emitted <= (lizzieLet29_4Lkron_kron_Int_Int_Intsbos_r ? 2'd0 :
                                                          lizzieLet29_4Lkron_kron_Int_Int_Intsbos_done);
  
  /* togo (Ty Pointer_QTree_Int) : (lizzieLet29_4Lkron_kron_Int_Int_Intsbos_1_merge_merge_fork_1,Pointer_QTree_Int) > (call_kron_kron_Int_Int_Int_goConst,Go) */
  assign call_kron_kron_Int_Int_Int_goConst_d = lizzieLet29_4Lkron_kron_Int_Int_Intsbos_1_merge_merge_fork_1_d[0];
  assign lizzieLet29_4Lkron_kron_Int_Int_Intsbos_1_merge_merge_fork_1_r = call_kron_kron_Int_Int_Int_goConst_r;
  
  /* buf (Ty Pointer_QTree_Int) : (lizzieLet29_4Lkron_kron_Int_Int_Intsbos_1_merge_merge_fork_2,Pointer_QTree_Int) > (kron_kron_Int_Int_Int_resbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t lizzieLet29_4Lkron_kron_Int_Int_Intsbos_1_merge_merge_fork_2_bufchan_d;
  logic lizzieLet29_4Lkron_kron_Int_Int_Intsbos_1_merge_merge_fork_2_bufchan_r;
  assign lizzieLet29_4Lkron_kron_Int_Int_Intsbos_1_merge_merge_fork_2_r = ((! lizzieLet29_4Lkron_kron_Int_Int_Intsbos_1_merge_merge_fork_2_bufchan_d[0]) || lizzieLet29_4Lkron_kron_Int_Int_Intsbos_1_merge_merge_fork_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet29_4Lkron_kron_Int_Int_Intsbos_1_merge_merge_fork_2_bufchan_d <= {16'd0,
                                                                                 1'd0};
    else
      if (lizzieLet29_4Lkron_kron_Int_Int_Intsbos_1_merge_merge_fork_2_r)
        lizzieLet29_4Lkron_kron_Int_Int_Intsbos_1_merge_merge_fork_2_bufchan_d <= lizzieLet29_4Lkron_kron_Int_Int_Intsbos_1_merge_merge_fork_2_d;
  Pointer_QTree_Int_t lizzieLet29_4Lkron_kron_Int_Int_Intsbos_1_merge_merge_fork_2_bufchan_buf;
  assign lizzieLet29_4Lkron_kron_Int_Int_Intsbos_1_merge_merge_fork_2_bufchan_r = (! lizzieLet29_4Lkron_kron_Int_Int_Intsbos_1_merge_merge_fork_2_bufchan_buf[0]);
  assign kron_kron_Int_Int_Int_resbuf_d = (lizzieLet29_4Lkron_kron_Int_Int_Intsbos_1_merge_merge_fork_2_bufchan_buf[0] ? lizzieLet29_4Lkron_kron_Int_Int_Intsbos_1_merge_merge_fork_2_bufchan_buf :
                                           lizzieLet29_4Lkron_kron_Int_Int_Intsbos_1_merge_merge_fork_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet29_4Lkron_kron_Int_Int_Intsbos_1_merge_merge_fork_2_bufchan_buf <= {16'd0,
                                                                                   1'd0};
    else
      if ((kron_kron_Int_Int_Int_resbuf_r && lizzieLet29_4Lkron_kron_Int_Int_Intsbos_1_merge_merge_fork_2_bufchan_buf[0]))
        lizzieLet29_4Lkron_kron_Int_Int_Intsbos_1_merge_merge_fork_2_bufchan_buf <= {16'd0,
                                                                                     1'd0};
      else if (((! kron_kron_Int_Int_Int_resbuf_r) && (! lizzieLet29_4Lkron_kron_Int_Int_Intsbos_1_merge_merge_fork_2_bufchan_buf[0])))
        lizzieLet29_4Lkron_kron_Int_Int_Intsbos_1_merge_merge_fork_2_bufchan_buf <= lizzieLet29_4Lkron_kron_Int_Int_Intsbos_1_merge_merge_fork_2_bufchan_d;
  
  /* destruct (Ty CTmain_map'_Int_Int,
          Dcon Lcall_main_map'_Int_Int0) : (lizzieLet34_1Lcall_main_map'_Int_Int0,CTmain_map'_Int_Int) > [(es_2_3_destruct,Pointer_QTree_Int),
                                                                                                          (es_3_5_destruct,Pointer_QTree_Int),
                                                                                                          (es_4_4_destruct,Pointer_QTree_Int),
                                                                                                          (sc_0_15_destruct,Pointer_CTmain_map'_Int_Int)] */
  logic [3:0] \lizzieLet34_1Lcall_main_map'_Int_Int0_emitted ;
  logic [3:0] \lizzieLet34_1Lcall_main_map'_Int_Int0_done ;
  assign es_2_3_destruct_d = {\lizzieLet34_1Lcall_main_map'_Int_Int0_d [19:4],
                              (\lizzieLet34_1Lcall_main_map'_Int_Int0_d [0] && (! \lizzieLet34_1Lcall_main_map'_Int_Int0_emitted [0]))};
  assign es_3_5_destruct_d = {\lizzieLet34_1Lcall_main_map'_Int_Int0_d [35:20],
                              (\lizzieLet34_1Lcall_main_map'_Int_Int0_d [0] && (! \lizzieLet34_1Lcall_main_map'_Int_Int0_emitted [1]))};
  assign es_4_4_destruct_d = {\lizzieLet34_1Lcall_main_map'_Int_Int0_d [51:36],
                              (\lizzieLet34_1Lcall_main_map'_Int_Int0_d [0] && (! \lizzieLet34_1Lcall_main_map'_Int_Int0_emitted [2]))};
  assign sc_0_15_destruct_d = {\lizzieLet34_1Lcall_main_map'_Int_Int0_d [67:52],
                               (\lizzieLet34_1Lcall_main_map'_Int_Int0_d [0] && (! \lizzieLet34_1Lcall_main_map'_Int_Int0_emitted [3]))};
  assign \lizzieLet34_1Lcall_main_map'_Int_Int0_done  = (\lizzieLet34_1Lcall_main_map'_Int_Int0_emitted  | ({sc_0_15_destruct_d[0],
                                                                                                             es_4_4_destruct_d[0],
                                                                                                             es_3_5_destruct_d[0],
                                                                                                             es_2_3_destruct_d[0]} & {sc_0_15_destruct_r,
                                                                                                                                      es_4_4_destruct_r,
                                                                                                                                      es_3_5_destruct_r,
                                                                                                                                      es_2_3_destruct_r}));
  assign \lizzieLet34_1Lcall_main_map'_Int_Int0_r  = (& \lizzieLet34_1Lcall_main_map'_Int_Int0_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet34_1Lcall_main_map'_Int_Int0_emitted  <= 4'd0;
    else
      \lizzieLet34_1Lcall_main_map'_Int_Int0_emitted  <= (\lizzieLet34_1Lcall_main_map'_Int_Int0_r  ? 4'd0 :
                                                          \lizzieLet34_1Lcall_main_map'_Int_Int0_done );
  
  /* destruct (Ty CTmain_map'_Int_Int,
          Dcon Lcall_main_map'_Int_Int1) : (lizzieLet34_1Lcall_main_map'_Int_Int1,CTmain_map'_Int_Int) > [(es_3_4_destruct,Pointer_QTree_Int),
                                                                                                          (es_4_3_destruct,Pointer_QTree_Int),
                                                                                                          (sc_0_14_destruct,Pointer_CTmain_map'_Int_Int),
                                                                                                          (isZacL_4_destruct,MyDTInt_Bool),
                                                                                                          (gacM_4_destruct,MyDTInt_Int),
                                                                                                          (q1acP_3_destruct,Pointer_QTree_Int)] */
  logic [5:0] \lizzieLet34_1Lcall_main_map'_Int_Int1_emitted ;
  logic [5:0] \lizzieLet34_1Lcall_main_map'_Int_Int1_done ;
  assign es_3_4_destruct_d = {\lizzieLet34_1Lcall_main_map'_Int_Int1_d [19:4],
                              (\lizzieLet34_1Lcall_main_map'_Int_Int1_d [0] && (! \lizzieLet34_1Lcall_main_map'_Int_Int1_emitted [0]))};
  assign es_4_3_destruct_d = {\lizzieLet34_1Lcall_main_map'_Int_Int1_d [35:20],
                              (\lizzieLet34_1Lcall_main_map'_Int_Int1_d [0] && (! \lizzieLet34_1Lcall_main_map'_Int_Int1_emitted [1]))};
  assign sc_0_14_destruct_d = {\lizzieLet34_1Lcall_main_map'_Int_Int1_d [51:36],
                               (\lizzieLet34_1Lcall_main_map'_Int_Int1_d [0] && (! \lizzieLet34_1Lcall_main_map'_Int_Int1_emitted [2]))};
  assign isZacL_4_destruct_d = (\lizzieLet34_1Lcall_main_map'_Int_Int1_d [0] && (! \lizzieLet34_1Lcall_main_map'_Int_Int1_emitted [3]));
  assign gacM_4_destruct_d = (\lizzieLet34_1Lcall_main_map'_Int_Int1_d [0] && (! \lizzieLet34_1Lcall_main_map'_Int_Int1_emitted [4]));
  assign q1acP_3_destruct_d = {\lizzieLet34_1Lcall_main_map'_Int_Int1_d [67:52],
                               (\lizzieLet34_1Lcall_main_map'_Int_Int1_d [0] && (! \lizzieLet34_1Lcall_main_map'_Int_Int1_emitted [5]))};
  assign \lizzieLet34_1Lcall_main_map'_Int_Int1_done  = (\lizzieLet34_1Lcall_main_map'_Int_Int1_emitted  | ({q1acP_3_destruct_d[0],
                                                                                                             gacM_4_destruct_d[0],
                                                                                                             isZacL_4_destruct_d[0],
                                                                                                             sc_0_14_destruct_d[0],
                                                                                                             es_4_3_destruct_d[0],
                                                                                                             es_3_4_destruct_d[0]} & {q1acP_3_destruct_r,
                                                                                                                                      gacM_4_destruct_r,
                                                                                                                                      isZacL_4_destruct_r,
                                                                                                                                      sc_0_14_destruct_r,
                                                                                                                                      es_4_3_destruct_r,
                                                                                                                                      es_3_4_destruct_r}));
  assign \lizzieLet34_1Lcall_main_map'_Int_Int1_r  = (& \lizzieLet34_1Lcall_main_map'_Int_Int1_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet34_1Lcall_main_map'_Int_Int1_emitted  <= 6'd0;
    else
      \lizzieLet34_1Lcall_main_map'_Int_Int1_emitted  <= (\lizzieLet34_1Lcall_main_map'_Int_Int1_r  ? 6'd0 :
                                                          \lizzieLet34_1Lcall_main_map'_Int_Int1_done );
  
  /* destruct (Ty CTmain_map'_Int_Int,
          Dcon Lcall_main_map'_Int_Int2) : (lizzieLet34_1Lcall_main_map'_Int_Int2,CTmain_map'_Int_Int) > [(es_4_2_destruct,Pointer_QTree_Int),
                                                                                                          (sc_0_13_destruct,Pointer_CTmain_map'_Int_Int),
                                                                                                          (isZacL_3_destruct,MyDTInt_Bool),
                                                                                                          (gacM_3_destruct,MyDTInt_Int),
                                                                                                          (q1acP_2_destruct,Pointer_QTree_Int),
                                                                                                          (q2acQ_2_destruct,Pointer_QTree_Int)] */
  logic [5:0] \lizzieLet34_1Lcall_main_map'_Int_Int2_emitted ;
  logic [5:0] \lizzieLet34_1Lcall_main_map'_Int_Int2_done ;
  assign es_4_2_destruct_d = {\lizzieLet34_1Lcall_main_map'_Int_Int2_d [19:4],
                              (\lizzieLet34_1Lcall_main_map'_Int_Int2_d [0] && (! \lizzieLet34_1Lcall_main_map'_Int_Int2_emitted [0]))};
  assign sc_0_13_destruct_d = {\lizzieLet34_1Lcall_main_map'_Int_Int2_d [35:20],
                               (\lizzieLet34_1Lcall_main_map'_Int_Int2_d [0] && (! \lizzieLet34_1Lcall_main_map'_Int_Int2_emitted [1]))};
  assign isZacL_3_destruct_d = (\lizzieLet34_1Lcall_main_map'_Int_Int2_d [0] && (! \lizzieLet34_1Lcall_main_map'_Int_Int2_emitted [2]));
  assign gacM_3_destruct_d = (\lizzieLet34_1Lcall_main_map'_Int_Int2_d [0] && (! \lizzieLet34_1Lcall_main_map'_Int_Int2_emitted [3]));
  assign q1acP_2_destruct_d = {\lizzieLet34_1Lcall_main_map'_Int_Int2_d [51:36],
                               (\lizzieLet34_1Lcall_main_map'_Int_Int2_d [0] && (! \lizzieLet34_1Lcall_main_map'_Int_Int2_emitted [4]))};
  assign q2acQ_2_destruct_d = {\lizzieLet34_1Lcall_main_map'_Int_Int2_d [67:52],
                               (\lizzieLet34_1Lcall_main_map'_Int_Int2_d [0] && (! \lizzieLet34_1Lcall_main_map'_Int_Int2_emitted [5]))};
  assign \lizzieLet34_1Lcall_main_map'_Int_Int2_done  = (\lizzieLet34_1Lcall_main_map'_Int_Int2_emitted  | ({q2acQ_2_destruct_d[0],
                                                                                                             q1acP_2_destruct_d[0],
                                                                                                             gacM_3_destruct_d[0],
                                                                                                             isZacL_3_destruct_d[0],
                                                                                                             sc_0_13_destruct_d[0],
                                                                                                             es_4_2_destruct_d[0]} & {q2acQ_2_destruct_r,
                                                                                                                                      q1acP_2_destruct_r,
                                                                                                                                      gacM_3_destruct_r,
                                                                                                                                      isZacL_3_destruct_r,
                                                                                                                                      sc_0_13_destruct_r,
                                                                                                                                      es_4_2_destruct_r}));
  assign \lizzieLet34_1Lcall_main_map'_Int_Int2_r  = (& \lizzieLet34_1Lcall_main_map'_Int_Int2_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet34_1Lcall_main_map'_Int_Int2_emitted  <= 6'd0;
    else
      \lizzieLet34_1Lcall_main_map'_Int_Int2_emitted  <= (\lizzieLet34_1Lcall_main_map'_Int_Int2_r  ? 6'd0 :
                                                          \lizzieLet34_1Lcall_main_map'_Int_Int2_done );
  
  /* destruct (Ty CTmain_map'_Int_Int,
          Dcon Lcall_main_map'_Int_Int3) : (lizzieLet34_1Lcall_main_map'_Int_Int3,CTmain_map'_Int_Int) > [(sc_0_12_destruct,Pointer_CTmain_map'_Int_Int),
                                                                                                          (isZacL_2_destruct,MyDTInt_Bool),
                                                                                                          (gacM_2_destruct,MyDTInt_Int),
                                                                                                          (q1acP_1_destruct,Pointer_QTree_Int),
                                                                                                          (q2acQ_1_destruct,Pointer_QTree_Int),
                                                                                                          (q3acR_1_destruct,Pointer_QTree_Int)] */
  logic [5:0] \lizzieLet34_1Lcall_main_map'_Int_Int3_emitted ;
  logic [5:0] \lizzieLet34_1Lcall_main_map'_Int_Int3_done ;
  assign sc_0_12_destruct_d = {\lizzieLet34_1Lcall_main_map'_Int_Int3_d [19:4],
                               (\lizzieLet34_1Lcall_main_map'_Int_Int3_d [0] && (! \lizzieLet34_1Lcall_main_map'_Int_Int3_emitted [0]))};
  assign isZacL_2_destruct_d = (\lizzieLet34_1Lcall_main_map'_Int_Int3_d [0] && (! \lizzieLet34_1Lcall_main_map'_Int_Int3_emitted [1]));
  assign gacM_2_destruct_d = (\lizzieLet34_1Lcall_main_map'_Int_Int3_d [0] && (! \lizzieLet34_1Lcall_main_map'_Int_Int3_emitted [2]));
  assign q1acP_1_destruct_d = {\lizzieLet34_1Lcall_main_map'_Int_Int3_d [35:20],
                               (\lizzieLet34_1Lcall_main_map'_Int_Int3_d [0] && (! \lizzieLet34_1Lcall_main_map'_Int_Int3_emitted [3]))};
  assign q2acQ_1_destruct_d = {\lizzieLet34_1Lcall_main_map'_Int_Int3_d [51:36],
                               (\lizzieLet34_1Lcall_main_map'_Int_Int3_d [0] && (! \lizzieLet34_1Lcall_main_map'_Int_Int3_emitted [4]))};
  assign q3acR_1_destruct_d = {\lizzieLet34_1Lcall_main_map'_Int_Int3_d [67:52],
                               (\lizzieLet34_1Lcall_main_map'_Int_Int3_d [0] && (! \lizzieLet34_1Lcall_main_map'_Int_Int3_emitted [5]))};
  assign \lizzieLet34_1Lcall_main_map'_Int_Int3_done  = (\lizzieLet34_1Lcall_main_map'_Int_Int3_emitted  | ({q3acR_1_destruct_d[0],
                                                                                                             q2acQ_1_destruct_d[0],
                                                                                                             q1acP_1_destruct_d[0],
                                                                                                             gacM_2_destruct_d[0],
                                                                                                             isZacL_2_destruct_d[0],
                                                                                                             sc_0_12_destruct_d[0]} & {q3acR_1_destruct_r,
                                                                                                                                       q2acQ_1_destruct_r,
                                                                                                                                       q1acP_1_destruct_r,
                                                                                                                                       gacM_2_destruct_r,
                                                                                                                                       isZacL_2_destruct_r,
                                                                                                                                       sc_0_12_destruct_r}));
  assign \lizzieLet34_1Lcall_main_map'_Int_Int3_r  = (& \lizzieLet34_1Lcall_main_map'_Int_Int3_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet34_1Lcall_main_map'_Int_Int3_emitted  <= 6'd0;
    else
      \lizzieLet34_1Lcall_main_map'_Int_Int3_emitted  <= (\lizzieLet34_1Lcall_main_map'_Int_Int3_r  ? 6'd0 :
                                                          \lizzieLet34_1Lcall_main_map'_Int_Int3_done );
  
  /* demux (Ty CTmain_map'_Int_Int,
       Ty CTmain_map'_Int_Int) : (lizzieLet34_2,CTmain_map'_Int_Int) (lizzieLet34_1,CTmain_map'_Int_Int) > [(_14,CTmain_map'_Int_Int),
                                                                                                            (lizzieLet34_1Lcall_main_map'_Int_Int3,CTmain_map'_Int_Int),
                                                                                                            (lizzieLet34_1Lcall_main_map'_Int_Int2,CTmain_map'_Int_Int),
                                                                                                            (lizzieLet34_1Lcall_main_map'_Int_Int1,CTmain_map'_Int_Int),
                                                                                                            (lizzieLet34_1Lcall_main_map'_Int_Int0,CTmain_map'_Int_Int)] */
  logic [4:0] lizzieLet34_1_onehotd;
  always_comb
    if ((lizzieLet34_2_d[0] && lizzieLet34_1_d[0]))
      unique case (lizzieLet34_2_d[3:1])
        3'd0: lizzieLet34_1_onehotd = 5'd1;
        3'd1: lizzieLet34_1_onehotd = 5'd2;
        3'd2: lizzieLet34_1_onehotd = 5'd4;
        3'd3: lizzieLet34_1_onehotd = 5'd8;
        3'd4: lizzieLet34_1_onehotd = 5'd16;
        default: lizzieLet34_1_onehotd = 5'd0;
      endcase
    else lizzieLet34_1_onehotd = 5'd0;
  assign _14_d = {lizzieLet34_1_d[67:1], lizzieLet34_1_onehotd[0]};
  assign \lizzieLet34_1Lcall_main_map'_Int_Int3_d  = {lizzieLet34_1_d[67:1],
                                                      lizzieLet34_1_onehotd[1]};
  assign \lizzieLet34_1Lcall_main_map'_Int_Int2_d  = {lizzieLet34_1_d[67:1],
                                                      lizzieLet34_1_onehotd[2]};
  assign \lizzieLet34_1Lcall_main_map'_Int_Int1_d  = {lizzieLet34_1_d[67:1],
                                                      lizzieLet34_1_onehotd[3]};
  assign \lizzieLet34_1Lcall_main_map'_Int_Int0_d  = {lizzieLet34_1_d[67:1],
                                                      lizzieLet34_1_onehotd[4]};
  assign lizzieLet34_1_r = (| (lizzieLet34_1_onehotd & {\lizzieLet34_1Lcall_main_map'_Int_Int0_r ,
                                                        \lizzieLet34_1Lcall_main_map'_Int_Int1_r ,
                                                        \lizzieLet34_1Lcall_main_map'_Int_Int2_r ,
                                                        \lizzieLet34_1Lcall_main_map'_Int_Int3_r ,
                                                        _14_r}));
  assign lizzieLet34_2_r = lizzieLet34_1_r;
  
  /* demux (Ty CTmain_map'_Int_Int,
       Ty Go) : (lizzieLet34_3,CTmain_map'_Int_Int) (go_20_goMux_data,Go) > [(_13,Go),
                                                                             (lizzieLet34_3Lcall_main_map'_Int_Int3,Go),
                                                                             (lizzieLet34_3Lcall_main_map'_Int_Int2,Go),
                                                                             (lizzieLet34_3Lcall_main_map'_Int_Int1,Go),
                                                                             (lizzieLet34_3Lcall_main_map'_Int_Int0,Go)] */
  logic [4:0] go_20_goMux_data_onehotd;
  always_comb
    if ((lizzieLet34_3_d[0] && go_20_goMux_data_d[0]))
      unique case (lizzieLet34_3_d[3:1])
        3'd0: go_20_goMux_data_onehotd = 5'd1;
        3'd1: go_20_goMux_data_onehotd = 5'd2;
        3'd2: go_20_goMux_data_onehotd = 5'd4;
        3'd3: go_20_goMux_data_onehotd = 5'd8;
        3'd4: go_20_goMux_data_onehotd = 5'd16;
        default: go_20_goMux_data_onehotd = 5'd0;
      endcase
    else go_20_goMux_data_onehotd = 5'd0;
  assign _13_d = go_20_goMux_data_onehotd[0];
  assign \lizzieLet34_3Lcall_main_map'_Int_Int3_d  = go_20_goMux_data_onehotd[1];
  assign \lizzieLet34_3Lcall_main_map'_Int_Int2_d  = go_20_goMux_data_onehotd[2];
  assign \lizzieLet34_3Lcall_main_map'_Int_Int1_d  = go_20_goMux_data_onehotd[3];
  assign \lizzieLet34_3Lcall_main_map'_Int_Int0_d  = go_20_goMux_data_onehotd[4];
  assign go_20_goMux_data_r = (| (go_20_goMux_data_onehotd & {\lizzieLet34_3Lcall_main_map'_Int_Int0_r ,
                                                              \lizzieLet34_3Lcall_main_map'_Int_Int1_r ,
                                                              \lizzieLet34_3Lcall_main_map'_Int_Int2_r ,
                                                              \lizzieLet34_3Lcall_main_map'_Int_Int3_r ,
                                                              _13_r}));
  assign lizzieLet34_3_r = go_20_goMux_data_r;
  
  /* buf (Ty Go) : (lizzieLet34_3Lcall_main_map'_Int_Int0,Go) > (lizzieLet34_3Lcall_main_map'_Int_Int0_1_argbuf,Go) */
  Go_t \lizzieLet34_3Lcall_main_map'_Int_Int0_bufchan_d ;
  logic \lizzieLet34_3Lcall_main_map'_Int_Int0_bufchan_r ;
  assign \lizzieLet34_3Lcall_main_map'_Int_Int0_r  = ((! \lizzieLet34_3Lcall_main_map'_Int_Int0_bufchan_d [0]) || \lizzieLet34_3Lcall_main_map'_Int_Int0_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet34_3Lcall_main_map'_Int_Int0_bufchan_d  <= 1'd0;
    else
      if (\lizzieLet34_3Lcall_main_map'_Int_Int0_r )
        \lizzieLet34_3Lcall_main_map'_Int_Int0_bufchan_d  <= \lizzieLet34_3Lcall_main_map'_Int_Int0_d ;
  Go_t \lizzieLet34_3Lcall_main_map'_Int_Int0_bufchan_buf ;
  assign \lizzieLet34_3Lcall_main_map'_Int_Int0_bufchan_r  = (! \lizzieLet34_3Lcall_main_map'_Int_Int0_bufchan_buf [0]);
  assign \lizzieLet34_3Lcall_main_map'_Int_Int0_1_argbuf_d  = (\lizzieLet34_3Lcall_main_map'_Int_Int0_bufchan_buf [0] ? \lizzieLet34_3Lcall_main_map'_Int_Int0_bufchan_buf  :
                                                               \lizzieLet34_3Lcall_main_map'_Int_Int0_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet34_3Lcall_main_map'_Int_Int0_bufchan_buf  <= 1'd0;
    else
      if ((\lizzieLet34_3Lcall_main_map'_Int_Int0_1_argbuf_r  && \lizzieLet34_3Lcall_main_map'_Int_Int0_bufchan_buf [0]))
        \lizzieLet34_3Lcall_main_map'_Int_Int0_bufchan_buf  <= 1'd0;
      else if (((! \lizzieLet34_3Lcall_main_map'_Int_Int0_1_argbuf_r ) && (! \lizzieLet34_3Lcall_main_map'_Int_Int0_bufchan_buf [0])))
        \lizzieLet34_3Lcall_main_map'_Int_Int0_bufchan_buf  <= \lizzieLet34_3Lcall_main_map'_Int_Int0_bufchan_d ;
  
  /* buf (Ty Go) : (lizzieLet34_3Lcall_main_map'_Int_Int1,Go) > (lizzieLet34_3Lcall_main_map'_Int_Int1_1_argbuf,Go) */
  Go_t \lizzieLet34_3Lcall_main_map'_Int_Int1_bufchan_d ;
  logic \lizzieLet34_3Lcall_main_map'_Int_Int1_bufchan_r ;
  assign \lizzieLet34_3Lcall_main_map'_Int_Int1_r  = ((! \lizzieLet34_3Lcall_main_map'_Int_Int1_bufchan_d [0]) || \lizzieLet34_3Lcall_main_map'_Int_Int1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet34_3Lcall_main_map'_Int_Int1_bufchan_d  <= 1'd0;
    else
      if (\lizzieLet34_3Lcall_main_map'_Int_Int1_r )
        \lizzieLet34_3Lcall_main_map'_Int_Int1_bufchan_d  <= \lizzieLet34_3Lcall_main_map'_Int_Int1_d ;
  Go_t \lizzieLet34_3Lcall_main_map'_Int_Int1_bufchan_buf ;
  assign \lizzieLet34_3Lcall_main_map'_Int_Int1_bufchan_r  = (! \lizzieLet34_3Lcall_main_map'_Int_Int1_bufchan_buf [0]);
  assign \lizzieLet34_3Lcall_main_map'_Int_Int1_1_argbuf_d  = (\lizzieLet34_3Lcall_main_map'_Int_Int1_bufchan_buf [0] ? \lizzieLet34_3Lcall_main_map'_Int_Int1_bufchan_buf  :
                                                               \lizzieLet34_3Lcall_main_map'_Int_Int1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet34_3Lcall_main_map'_Int_Int1_bufchan_buf  <= 1'd0;
    else
      if ((\lizzieLet34_3Lcall_main_map'_Int_Int1_1_argbuf_r  && \lizzieLet34_3Lcall_main_map'_Int_Int1_bufchan_buf [0]))
        \lizzieLet34_3Lcall_main_map'_Int_Int1_bufchan_buf  <= 1'd0;
      else if (((! \lizzieLet34_3Lcall_main_map'_Int_Int1_1_argbuf_r ) && (! \lizzieLet34_3Lcall_main_map'_Int_Int1_bufchan_buf [0])))
        \lizzieLet34_3Lcall_main_map'_Int_Int1_bufchan_buf  <= \lizzieLet34_3Lcall_main_map'_Int_Int1_bufchan_d ;
  
  /* buf (Ty Go) : (lizzieLet34_3Lcall_main_map'_Int_Int2,Go) > (lizzieLet34_3Lcall_main_map'_Int_Int2_1_argbuf,Go) */
  Go_t \lizzieLet34_3Lcall_main_map'_Int_Int2_bufchan_d ;
  logic \lizzieLet34_3Lcall_main_map'_Int_Int2_bufchan_r ;
  assign \lizzieLet34_3Lcall_main_map'_Int_Int2_r  = ((! \lizzieLet34_3Lcall_main_map'_Int_Int2_bufchan_d [0]) || \lizzieLet34_3Lcall_main_map'_Int_Int2_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet34_3Lcall_main_map'_Int_Int2_bufchan_d  <= 1'd0;
    else
      if (\lizzieLet34_3Lcall_main_map'_Int_Int2_r )
        \lizzieLet34_3Lcall_main_map'_Int_Int2_bufchan_d  <= \lizzieLet34_3Lcall_main_map'_Int_Int2_d ;
  Go_t \lizzieLet34_3Lcall_main_map'_Int_Int2_bufchan_buf ;
  assign \lizzieLet34_3Lcall_main_map'_Int_Int2_bufchan_r  = (! \lizzieLet34_3Lcall_main_map'_Int_Int2_bufchan_buf [0]);
  assign \lizzieLet34_3Lcall_main_map'_Int_Int2_1_argbuf_d  = (\lizzieLet34_3Lcall_main_map'_Int_Int2_bufchan_buf [0] ? \lizzieLet34_3Lcall_main_map'_Int_Int2_bufchan_buf  :
                                                               \lizzieLet34_3Lcall_main_map'_Int_Int2_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet34_3Lcall_main_map'_Int_Int2_bufchan_buf  <= 1'd0;
    else
      if ((\lizzieLet34_3Lcall_main_map'_Int_Int2_1_argbuf_r  && \lizzieLet34_3Lcall_main_map'_Int_Int2_bufchan_buf [0]))
        \lizzieLet34_3Lcall_main_map'_Int_Int2_bufchan_buf  <= 1'd0;
      else if (((! \lizzieLet34_3Lcall_main_map'_Int_Int2_1_argbuf_r ) && (! \lizzieLet34_3Lcall_main_map'_Int_Int2_bufchan_buf [0])))
        \lizzieLet34_3Lcall_main_map'_Int_Int2_bufchan_buf  <= \lizzieLet34_3Lcall_main_map'_Int_Int2_bufchan_d ;
  
  /* buf (Ty Go) : (lizzieLet34_3Lcall_main_map'_Int_Int3,Go) > (lizzieLet34_3Lcall_main_map'_Int_Int3_1_argbuf,Go) */
  Go_t \lizzieLet34_3Lcall_main_map'_Int_Int3_bufchan_d ;
  logic \lizzieLet34_3Lcall_main_map'_Int_Int3_bufchan_r ;
  assign \lizzieLet34_3Lcall_main_map'_Int_Int3_r  = ((! \lizzieLet34_3Lcall_main_map'_Int_Int3_bufchan_d [0]) || \lizzieLet34_3Lcall_main_map'_Int_Int3_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet34_3Lcall_main_map'_Int_Int3_bufchan_d  <= 1'd0;
    else
      if (\lizzieLet34_3Lcall_main_map'_Int_Int3_r )
        \lizzieLet34_3Lcall_main_map'_Int_Int3_bufchan_d  <= \lizzieLet34_3Lcall_main_map'_Int_Int3_d ;
  Go_t \lizzieLet34_3Lcall_main_map'_Int_Int3_bufchan_buf ;
  assign \lizzieLet34_3Lcall_main_map'_Int_Int3_bufchan_r  = (! \lizzieLet34_3Lcall_main_map'_Int_Int3_bufchan_buf [0]);
  assign \lizzieLet34_3Lcall_main_map'_Int_Int3_1_argbuf_d  = (\lizzieLet34_3Lcall_main_map'_Int_Int3_bufchan_buf [0] ? \lizzieLet34_3Lcall_main_map'_Int_Int3_bufchan_buf  :
                                                               \lizzieLet34_3Lcall_main_map'_Int_Int3_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet34_3Lcall_main_map'_Int_Int3_bufchan_buf  <= 1'd0;
    else
      if ((\lizzieLet34_3Lcall_main_map'_Int_Int3_1_argbuf_r  && \lizzieLet34_3Lcall_main_map'_Int_Int3_bufchan_buf [0]))
        \lizzieLet34_3Lcall_main_map'_Int_Int3_bufchan_buf  <= 1'd0;
      else if (((! \lizzieLet34_3Lcall_main_map'_Int_Int3_1_argbuf_r ) && (! \lizzieLet34_3Lcall_main_map'_Int_Int3_bufchan_buf [0])))
        \lizzieLet34_3Lcall_main_map'_Int_Int3_bufchan_buf  <= \lizzieLet34_3Lcall_main_map'_Int_Int3_bufchan_d ;
  
  /* demux (Ty CTmain_map'_Int_Int,
       Ty Pointer_QTree_Int) : (lizzieLet34_4,CTmain_map'_Int_Int) (srtarg_0_2_goMux_mux,Pointer_QTree_Int) > [(lizzieLet34_4Lmain_map'_Int_Intsbos,Pointer_QTree_Int),
                                                                                                               (lizzieLet34_4Lcall_main_map'_Int_Int3,Pointer_QTree_Int),
                                                                                                               (lizzieLet34_4Lcall_main_map'_Int_Int2,Pointer_QTree_Int),
                                                                                                               (lizzieLet34_4Lcall_main_map'_Int_Int1,Pointer_QTree_Int),
                                                                                                               (lizzieLet34_4Lcall_main_map'_Int_Int0,Pointer_QTree_Int)] */
  logic [4:0] srtarg_0_2_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet34_4_d[0] && srtarg_0_2_goMux_mux_d[0]))
      unique case (lizzieLet34_4_d[3:1])
        3'd0: srtarg_0_2_goMux_mux_onehotd = 5'd1;
        3'd1: srtarg_0_2_goMux_mux_onehotd = 5'd2;
        3'd2: srtarg_0_2_goMux_mux_onehotd = 5'd4;
        3'd3: srtarg_0_2_goMux_mux_onehotd = 5'd8;
        3'd4: srtarg_0_2_goMux_mux_onehotd = 5'd16;
        default: srtarg_0_2_goMux_mux_onehotd = 5'd0;
      endcase
    else srtarg_0_2_goMux_mux_onehotd = 5'd0;
  assign \lizzieLet34_4Lmain_map'_Int_Intsbos_d  = {srtarg_0_2_goMux_mux_d[16:1],
                                                    srtarg_0_2_goMux_mux_onehotd[0]};
  assign \lizzieLet34_4Lcall_main_map'_Int_Int3_d  = {srtarg_0_2_goMux_mux_d[16:1],
                                                      srtarg_0_2_goMux_mux_onehotd[1]};
  assign \lizzieLet34_4Lcall_main_map'_Int_Int2_d  = {srtarg_0_2_goMux_mux_d[16:1],
                                                      srtarg_0_2_goMux_mux_onehotd[2]};
  assign \lizzieLet34_4Lcall_main_map'_Int_Int1_d  = {srtarg_0_2_goMux_mux_d[16:1],
                                                      srtarg_0_2_goMux_mux_onehotd[3]};
  assign \lizzieLet34_4Lcall_main_map'_Int_Int0_d  = {srtarg_0_2_goMux_mux_d[16:1],
                                                      srtarg_0_2_goMux_mux_onehotd[4]};
  assign srtarg_0_2_goMux_mux_r = (| (srtarg_0_2_goMux_mux_onehotd & {\lizzieLet34_4Lcall_main_map'_Int_Int0_r ,
                                                                      \lizzieLet34_4Lcall_main_map'_Int_Int1_r ,
                                                                      \lizzieLet34_4Lcall_main_map'_Int_Int2_r ,
                                                                      \lizzieLet34_4Lcall_main_map'_Int_Int3_r ,
                                                                      \lizzieLet34_4Lmain_map'_Int_Intsbos_r }));
  assign lizzieLet34_4_r = srtarg_0_2_goMux_mux_r;
  
  /* dcon (Ty QTree_Int,
      Dcon QNode_Int) : [(lizzieLet34_4Lcall_main_map'_Int_Int0,Pointer_QTree_Int),
                         (es_2_3_destruct,Pointer_QTree_Int),
                         (es_3_5_destruct,Pointer_QTree_Int),
                         (es_4_4_destruct,Pointer_QTree_Int)] > (lizzieLet34_4Lcall_main_map'_Int_Int0_1es_2_3_1es_3_5_1es_4_4_1QNode_Int,QTree_Int) */
  assign \lizzieLet34_4Lcall_main_map'_Int_Int0_1es_2_3_1es_3_5_1es_4_4_1QNode_Int_d  = QNode_Int_dc((& {\lizzieLet34_4Lcall_main_map'_Int_Int0_d [0],
                                                                                                         es_2_3_destruct_d[0],
                                                                                                         es_3_5_destruct_d[0],
                                                                                                         es_4_4_destruct_d[0]}), \lizzieLet34_4Lcall_main_map'_Int_Int0_d , es_2_3_destruct_d, es_3_5_destruct_d, es_4_4_destruct_d);
  assign {\lizzieLet34_4Lcall_main_map'_Int_Int0_r ,
          es_2_3_destruct_r,
          es_3_5_destruct_r,
          es_4_4_destruct_r} = {4 {(\lizzieLet34_4Lcall_main_map'_Int_Int0_1es_2_3_1es_3_5_1es_4_4_1QNode_Int_r  && \lizzieLet34_4Lcall_main_map'_Int_Int0_1es_2_3_1es_3_5_1es_4_4_1QNode_Int_d [0])}};
  
  /* buf (Ty QTree_Int) : (lizzieLet34_4Lcall_main_map'_Int_Int0_1es_2_3_1es_3_5_1es_4_4_1QNode_Int,QTree_Int) > (lizzieLet38_1_argbuf,QTree_Int) */
  QTree_Int_t \lizzieLet34_4Lcall_main_map'_Int_Int0_1es_2_3_1es_3_5_1es_4_4_1QNode_Int_bufchan_d ;
  logic \lizzieLet34_4Lcall_main_map'_Int_Int0_1es_2_3_1es_3_5_1es_4_4_1QNode_Int_bufchan_r ;
  assign \lizzieLet34_4Lcall_main_map'_Int_Int0_1es_2_3_1es_3_5_1es_4_4_1QNode_Int_r  = ((! \lizzieLet34_4Lcall_main_map'_Int_Int0_1es_2_3_1es_3_5_1es_4_4_1QNode_Int_bufchan_d [0]) || \lizzieLet34_4Lcall_main_map'_Int_Int0_1es_2_3_1es_3_5_1es_4_4_1QNode_Int_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet34_4Lcall_main_map'_Int_Int0_1es_2_3_1es_3_5_1es_4_4_1QNode_Int_bufchan_d  <= {66'd0,
                                                                                               1'd0};
    else
      if (\lizzieLet34_4Lcall_main_map'_Int_Int0_1es_2_3_1es_3_5_1es_4_4_1QNode_Int_r )
        \lizzieLet34_4Lcall_main_map'_Int_Int0_1es_2_3_1es_3_5_1es_4_4_1QNode_Int_bufchan_d  <= \lizzieLet34_4Lcall_main_map'_Int_Int0_1es_2_3_1es_3_5_1es_4_4_1QNode_Int_d ;
  QTree_Int_t \lizzieLet34_4Lcall_main_map'_Int_Int0_1es_2_3_1es_3_5_1es_4_4_1QNode_Int_bufchan_buf ;
  assign \lizzieLet34_4Lcall_main_map'_Int_Int0_1es_2_3_1es_3_5_1es_4_4_1QNode_Int_bufchan_r  = (! \lizzieLet34_4Lcall_main_map'_Int_Int0_1es_2_3_1es_3_5_1es_4_4_1QNode_Int_bufchan_buf [0]);
  assign lizzieLet38_1_argbuf_d = (\lizzieLet34_4Lcall_main_map'_Int_Int0_1es_2_3_1es_3_5_1es_4_4_1QNode_Int_bufchan_buf [0] ? \lizzieLet34_4Lcall_main_map'_Int_Int0_1es_2_3_1es_3_5_1es_4_4_1QNode_Int_bufchan_buf  :
                                   \lizzieLet34_4Lcall_main_map'_Int_Int0_1es_2_3_1es_3_5_1es_4_4_1QNode_Int_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet34_4Lcall_main_map'_Int_Int0_1es_2_3_1es_3_5_1es_4_4_1QNode_Int_bufchan_buf  <= {66'd0,
                                                                                                 1'd0};
    else
      if ((lizzieLet38_1_argbuf_r && \lizzieLet34_4Lcall_main_map'_Int_Int0_1es_2_3_1es_3_5_1es_4_4_1QNode_Int_bufchan_buf [0]))
        \lizzieLet34_4Lcall_main_map'_Int_Int0_1es_2_3_1es_3_5_1es_4_4_1QNode_Int_bufchan_buf  <= {66'd0,
                                                                                                   1'd0};
      else if (((! lizzieLet38_1_argbuf_r) && (! \lizzieLet34_4Lcall_main_map'_Int_Int0_1es_2_3_1es_3_5_1es_4_4_1QNode_Int_bufchan_buf [0])))
        \lizzieLet34_4Lcall_main_map'_Int_Int0_1es_2_3_1es_3_5_1es_4_4_1QNode_Int_bufchan_buf  <= \lizzieLet34_4Lcall_main_map'_Int_Int0_1es_2_3_1es_3_5_1es_4_4_1QNode_Int_bufchan_d ;
  
  /* dcon (Ty CTmain_map'_Int_Int,
      Dcon Lcall_main_map'_Int_Int0) : [(lizzieLet34_4Lcall_main_map'_Int_Int1,Pointer_QTree_Int),
                                        (es_3_4_destruct,Pointer_QTree_Int),
                                        (es_4_3_destruct,Pointer_QTree_Int),
                                        (sc_0_14_destruct,Pointer_CTmain_map'_Int_Int)] > (lizzieLet34_4Lcall_main_map'_Int_Int1_1es_3_4_1es_4_3_1sc_0_14_1Lcall_main_map'_Int_Int0,CTmain_map'_Int_Int) */
  assign \lizzieLet34_4Lcall_main_map'_Int_Int1_1es_3_4_1es_4_3_1sc_0_14_1Lcall_main_map'_Int_Int0_d  = \Lcall_main_map'_Int_Int0_dc ((& {\lizzieLet34_4Lcall_main_map'_Int_Int1_d [0],
                                                                                                                                          es_3_4_destruct_d[0],
                                                                                                                                          es_4_3_destruct_d[0],
                                                                                                                                          sc_0_14_destruct_d[0]}), \lizzieLet34_4Lcall_main_map'_Int_Int1_d , es_3_4_destruct_d, es_4_3_destruct_d, sc_0_14_destruct_d);
  assign {\lizzieLet34_4Lcall_main_map'_Int_Int1_r ,
          es_3_4_destruct_r,
          es_4_3_destruct_r,
          sc_0_14_destruct_r} = {4 {(\lizzieLet34_4Lcall_main_map'_Int_Int1_1es_3_4_1es_4_3_1sc_0_14_1Lcall_main_map'_Int_Int0_r  && \lizzieLet34_4Lcall_main_map'_Int_Int1_1es_3_4_1es_4_3_1sc_0_14_1Lcall_main_map'_Int_Int0_d [0])}};
  
  /* buf (Ty CTmain_map'_Int_Int) : (lizzieLet34_4Lcall_main_map'_Int_Int1_1es_3_4_1es_4_3_1sc_0_14_1Lcall_main_map'_Int_Int0,CTmain_map'_Int_Int) > (lizzieLet37_1_argbuf,CTmain_map'_Int_Int) */
  \CTmain_map'_Int_Int_t  \lizzieLet34_4Lcall_main_map'_Int_Int1_1es_3_4_1es_4_3_1sc_0_14_1Lcall_main_map'_Int_Int0_bufchan_d ;
  logic \lizzieLet34_4Lcall_main_map'_Int_Int1_1es_3_4_1es_4_3_1sc_0_14_1Lcall_main_map'_Int_Int0_bufchan_r ;
  assign \lizzieLet34_4Lcall_main_map'_Int_Int1_1es_3_4_1es_4_3_1sc_0_14_1Lcall_main_map'_Int_Int0_r  = ((! \lizzieLet34_4Lcall_main_map'_Int_Int1_1es_3_4_1es_4_3_1sc_0_14_1Lcall_main_map'_Int_Int0_bufchan_d [0]) || \lizzieLet34_4Lcall_main_map'_Int_Int1_1es_3_4_1es_4_3_1sc_0_14_1Lcall_main_map'_Int_Int0_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet34_4Lcall_main_map'_Int_Int1_1es_3_4_1es_4_3_1sc_0_14_1Lcall_main_map'_Int_Int0_bufchan_d  <= {67'd0,
                                                                                                               1'd0};
    else
      if (\lizzieLet34_4Lcall_main_map'_Int_Int1_1es_3_4_1es_4_3_1sc_0_14_1Lcall_main_map'_Int_Int0_r )
        \lizzieLet34_4Lcall_main_map'_Int_Int1_1es_3_4_1es_4_3_1sc_0_14_1Lcall_main_map'_Int_Int0_bufchan_d  <= \lizzieLet34_4Lcall_main_map'_Int_Int1_1es_3_4_1es_4_3_1sc_0_14_1Lcall_main_map'_Int_Int0_d ;
  \CTmain_map'_Int_Int_t  \lizzieLet34_4Lcall_main_map'_Int_Int1_1es_3_4_1es_4_3_1sc_0_14_1Lcall_main_map'_Int_Int0_bufchan_buf ;
  assign \lizzieLet34_4Lcall_main_map'_Int_Int1_1es_3_4_1es_4_3_1sc_0_14_1Lcall_main_map'_Int_Int0_bufchan_r  = (! \lizzieLet34_4Lcall_main_map'_Int_Int1_1es_3_4_1es_4_3_1sc_0_14_1Lcall_main_map'_Int_Int0_bufchan_buf [0]);
  assign lizzieLet37_1_argbuf_d = (\lizzieLet34_4Lcall_main_map'_Int_Int1_1es_3_4_1es_4_3_1sc_0_14_1Lcall_main_map'_Int_Int0_bufchan_buf [0] ? \lizzieLet34_4Lcall_main_map'_Int_Int1_1es_3_4_1es_4_3_1sc_0_14_1Lcall_main_map'_Int_Int0_bufchan_buf  :
                                   \lizzieLet34_4Lcall_main_map'_Int_Int1_1es_3_4_1es_4_3_1sc_0_14_1Lcall_main_map'_Int_Int0_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet34_4Lcall_main_map'_Int_Int1_1es_3_4_1es_4_3_1sc_0_14_1Lcall_main_map'_Int_Int0_bufchan_buf  <= {67'd0,
                                                                                                                 1'd0};
    else
      if ((lizzieLet37_1_argbuf_r && \lizzieLet34_4Lcall_main_map'_Int_Int1_1es_3_4_1es_4_3_1sc_0_14_1Lcall_main_map'_Int_Int0_bufchan_buf [0]))
        \lizzieLet34_4Lcall_main_map'_Int_Int1_1es_3_4_1es_4_3_1sc_0_14_1Lcall_main_map'_Int_Int0_bufchan_buf  <= {67'd0,
                                                                                                                   1'd0};
      else if (((! lizzieLet37_1_argbuf_r) && (! \lizzieLet34_4Lcall_main_map'_Int_Int1_1es_3_4_1es_4_3_1sc_0_14_1Lcall_main_map'_Int_Int0_bufchan_buf [0])))
        \lizzieLet34_4Lcall_main_map'_Int_Int1_1es_3_4_1es_4_3_1sc_0_14_1Lcall_main_map'_Int_Int0_bufchan_buf  <= \lizzieLet34_4Lcall_main_map'_Int_Int1_1es_3_4_1es_4_3_1sc_0_14_1Lcall_main_map'_Int_Int0_bufchan_d ;
  
  /* dcon (Ty CTmain_map'_Int_Int,
      Dcon Lcall_main_map'_Int_Int1) : [(lizzieLet34_4Lcall_main_map'_Int_Int2,Pointer_QTree_Int),
                                        (es_4_2_destruct,Pointer_QTree_Int),
                                        (sc_0_13_destruct,Pointer_CTmain_map'_Int_Int),
                                        (isZacL_3_1,MyDTInt_Bool),
                                        (gacM_3_1,MyDTInt_Int),
                                        (q1acP_2_destruct,Pointer_QTree_Int)] > (lizzieLet34_4Lcall_main_map'_Int_Int2_1es_4_2_1sc_0_13_1isZacL_3_1gacM_3_1q1acP_2_1Lcall_main_map'_Int_Int1,CTmain_map'_Int_Int) */
  assign \lizzieLet34_4Lcall_main_map'_Int_Int2_1es_4_2_1sc_0_13_1isZacL_3_1gacM_3_1q1acP_2_1Lcall_main_map'_Int_Int1_d  = \Lcall_main_map'_Int_Int1_dc ((& {\lizzieLet34_4Lcall_main_map'_Int_Int2_d [0],
                                                                                                                                                             es_4_2_destruct_d[0],
                                                                                                                                                             sc_0_13_destruct_d[0],
                                                                                                                                                             isZacL_3_1_d[0],
                                                                                                                                                             gacM_3_1_d[0],
                                                                                                                                                             q1acP_2_destruct_d[0]}), \lizzieLet34_4Lcall_main_map'_Int_Int2_d , es_4_2_destruct_d, sc_0_13_destruct_d, isZacL_3_1_d, gacM_3_1_d, q1acP_2_destruct_d);
  assign {\lizzieLet34_4Lcall_main_map'_Int_Int2_r ,
          es_4_2_destruct_r,
          sc_0_13_destruct_r,
          isZacL_3_1_r,
          gacM_3_1_r,
          q1acP_2_destruct_r} = {6 {(\lizzieLet34_4Lcall_main_map'_Int_Int2_1es_4_2_1sc_0_13_1isZacL_3_1gacM_3_1q1acP_2_1Lcall_main_map'_Int_Int1_r  && \lizzieLet34_4Lcall_main_map'_Int_Int2_1es_4_2_1sc_0_13_1isZacL_3_1gacM_3_1q1acP_2_1Lcall_main_map'_Int_Int1_d [0])}};
  
  /* buf (Ty CTmain_map'_Int_Int) : (lizzieLet34_4Lcall_main_map'_Int_Int2_1es_4_2_1sc_0_13_1isZacL_3_1gacM_3_1q1acP_2_1Lcall_main_map'_Int_Int1,CTmain_map'_Int_Int) > (lizzieLet36_1_argbuf,CTmain_map'_Int_Int) */
  \CTmain_map'_Int_Int_t  \lizzieLet34_4Lcall_main_map'_Int_Int2_1es_4_2_1sc_0_13_1isZacL_3_1gacM_3_1q1acP_2_1Lcall_main_map'_Int_Int1_bufchan_d ;
  logic \lizzieLet34_4Lcall_main_map'_Int_Int2_1es_4_2_1sc_0_13_1isZacL_3_1gacM_3_1q1acP_2_1Lcall_main_map'_Int_Int1_bufchan_r ;
  assign \lizzieLet34_4Lcall_main_map'_Int_Int2_1es_4_2_1sc_0_13_1isZacL_3_1gacM_3_1q1acP_2_1Lcall_main_map'_Int_Int1_r  = ((! \lizzieLet34_4Lcall_main_map'_Int_Int2_1es_4_2_1sc_0_13_1isZacL_3_1gacM_3_1q1acP_2_1Lcall_main_map'_Int_Int1_bufchan_d [0]) || \lizzieLet34_4Lcall_main_map'_Int_Int2_1es_4_2_1sc_0_13_1isZacL_3_1gacM_3_1q1acP_2_1Lcall_main_map'_Int_Int1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet34_4Lcall_main_map'_Int_Int2_1es_4_2_1sc_0_13_1isZacL_3_1gacM_3_1q1acP_2_1Lcall_main_map'_Int_Int1_bufchan_d  <= {67'd0,
                                                                                                                                  1'd0};
    else
      if (\lizzieLet34_4Lcall_main_map'_Int_Int2_1es_4_2_1sc_0_13_1isZacL_3_1gacM_3_1q1acP_2_1Lcall_main_map'_Int_Int1_r )
        \lizzieLet34_4Lcall_main_map'_Int_Int2_1es_4_2_1sc_0_13_1isZacL_3_1gacM_3_1q1acP_2_1Lcall_main_map'_Int_Int1_bufchan_d  <= \lizzieLet34_4Lcall_main_map'_Int_Int2_1es_4_2_1sc_0_13_1isZacL_3_1gacM_3_1q1acP_2_1Lcall_main_map'_Int_Int1_d ;
  \CTmain_map'_Int_Int_t  \lizzieLet34_4Lcall_main_map'_Int_Int2_1es_4_2_1sc_0_13_1isZacL_3_1gacM_3_1q1acP_2_1Lcall_main_map'_Int_Int1_bufchan_buf ;
  assign \lizzieLet34_4Lcall_main_map'_Int_Int2_1es_4_2_1sc_0_13_1isZacL_3_1gacM_3_1q1acP_2_1Lcall_main_map'_Int_Int1_bufchan_r  = (! \lizzieLet34_4Lcall_main_map'_Int_Int2_1es_4_2_1sc_0_13_1isZacL_3_1gacM_3_1q1acP_2_1Lcall_main_map'_Int_Int1_bufchan_buf [0]);
  assign lizzieLet36_1_argbuf_d = (\lizzieLet34_4Lcall_main_map'_Int_Int2_1es_4_2_1sc_0_13_1isZacL_3_1gacM_3_1q1acP_2_1Lcall_main_map'_Int_Int1_bufchan_buf [0] ? \lizzieLet34_4Lcall_main_map'_Int_Int2_1es_4_2_1sc_0_13_1isZacL_3_1gacM_3_1q1acP_2_1Lcall_main_map'_Int_Int1_bufchan_buf  :
                                   \lizzieLet34_4Lcall_main_map'_Int_Int2_1es_4_2_1sc_0_13_1isZacL_3_1gacM_3_1q1acP_2_1Lcall_main_map'_Int_Int1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet34_4Lcall_main_map'_Int_Int2_1es_4_2_1sc_0_13_1isZacL_3_1gacM_3_1q1acP_2_1Lcall_main_map'_Int_Int1_bufchan_buf  <= {67'd0,
                                                                                                                                    1'd0};
    else
      if ((lizzieLet36_1_argbuf_r && \lizzieLet34_4Lcall_main_map'_Int_Int2_1es_4_2_1sc_0_13_1isZacL_3_1gacM_3_1q1acP_2_1Lcall_main_map'_Int_Int1_bufchan_buf [0]))
        \lizzieLet34_4Lcall_main_map'_Int_Int2_1es_4_2_1sc_0_13_1isZacL_3_1gacM_3_1q1acP_2_1Lcall_main_map'_Int_Int1_bufchan_buf  <= {67'd0,
                                                                                                                                      1'd0};
      else if (((! lizzieLet36_1_argbuf_r) && (! \lizzieLet34_4Lcall_main_map'_Int_Int2_1es_4_2_1sc_0_13_1isZacL_3_1gacM_3_1q1acP_2_1Lcall_main_map'_Int_Int1_bufchan_buf [0])))
        \lizzieLet34_4Lcall_main_map'_Int_Int2_1es_4_2_1sc_0_13_1isZacL_3_1gacM_3_1q1acP_2_1Lcall_main_map'_Int_Int1_bufchan_buf  <= \lizzieLet34_4Lcall_main_map'_Int_Int2_1es_4_2_1sc_0_13_1isZacL_3_1gacM_3_1q1acP_2_1Lcall_main_map'_Int_Int1_bufchan_d ;
  
  /* dcon (Ty CTmain_map'_Int_Int,
      Dcon Lcall_main_map'_Int_Int2) : [(lizzieLet34_4Lcall_main_map'_Int_Int3,Pointer_QTree_Int),
                                        (sc_0_12_destruct,Pointer_CTmain_map'_Int_Int),
                                        (isZacL_2_1,MyDTInt_Bool),
                                        (gacM_2_1,MyDTInt_Int),
                                        (q1acP_1_destruct,Pointer_QTree_Int),
                                        (q2acQ_1_destruct,Pointer_QTree_Int)] > (lizzieLet34_4Lcall_main_map'_Int_Int3_1sc_0_12_1isZacL_2_1gacM_2_1q1acP_1_1q2acQ_1_1Lcall_main_map'_Int_Int2,CTmain_map'_Int_Int) */
  assign \lizzieLet34_4Lcall_main_map'_Int_Int3_1sc_0_12_1isZacL_2_1gacM_2_1q1acP_1_1q2acQ_1_1Lcall_main_map'_Int_Int2_d  = \Lcall_main_map'_Int_Int2_dc ((& {\lizzieLet34_4Lcall_main_map'_Int_Int3_d [0],
                                                                                                                                                              sc_0_12_destruct_d[0],
                                                                                                                                                              isZacL_2_1_d[0],
                                                                                                                                                              gacM_2_1_d[0],
                                                                                                                                                              q1acP_1_destruct_d[0],
                                                                                                                                                              q2acQ_1_destruct_d[0]}), \lizzieLet34_4Lcall_main_map'_Int_Int3_d , sc_0_12_destruct_d, isZacL_2_1_d, gacM_2_1_d, q1acP_1_destruct_d, q2acQ_1_destruct_d);
  assign {\lizzieLet34_4Lcall_main_map'_Int_Int3_r ,
          sc_0_12_destruct_r,
          isZacL_2_1_r,
          gacM_2_1_r,
          q1acP_1_destruct_r,
          q2acQ_1_destruct_r} = {6 {(\lizzieLet34_4Lcall_main_map'_Int_Int3_1sc_0_12_1isZacL_2_1gacM_2_1q1acP_1_1q2acQ_1_1Lcall_main_map'_Int_Int2_r  && \lizzieLet34_4Lcall_main_map'_Int_Int3_1sc_0_12_1isZacL_2_1gacM_2_1q1acP_1_1q2acQ_1_1Lcall_main_map'_Int_Int2_d [0])}};
  
  /* buf (Ty CTmain_map'_Int_Int) : (lizzieLet34_4Lcall_main_map'_Int_Int3_1sc_0_12_1isZacL_2_1gacM_2_1q1acP_1_1q2acQ_1_1Lcall_main_map'_Int_Int2,CTmain_map'_Int_Int) > (lizzieLet35_1_argbuf,CTmain_map'_Int_Int) */
  \CTmain_map'_Int_Int_t  \lizzieLet34_4Lcall_main_map'_Int_Int3_1sc_0_12_1isZacL_2_1gacM_2_1q1acP_1_1q2acQ_1_1Lcall_main_map'_Int_Int2_bufchan_d ;
  logic \lizzieLet34_4Lcall_main_map'_Int_Int3_1sc_0_12_1isZacL_2_1gacM_2_1q1acP_1_1q2acQ_1_1Lcall_main_map'_Int_Int2_bufchan_r ;
  assign \lizzieLet34_4Lcall_main_map'_Int_Int3_1sc_0_12_1isZacL_2_1gacM_2_1q1acP_1_1q2acQ_1_1Lcall_main_map'_Int_Int2_r  = ((! \lizzieLet34_4Lcall_main_map'_Int_Int3_1sc_0_12_1isZacL_2_1gacM_2_1q1acP_1_1q2acQ_1_1Lcall_main_map'_Int_Int2_bufchan_d [0]) || \lizzieLet34_4Lcall_main_map'_Int_Int3_1sc_0_12_1isZacL_2_1gacM_2_1q1acP_1_1q2acQ_1_1Lcall_main_map'_Int_Int2_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet34_4Lcall_main_map'_Int_Int3_1sc_0_12_1isZacL_2_1gacM_2_1q1acP_1_1q2acQ_1_1Lcall_main_map'_Int_Int2_bufchan_d  <= {67'd0,
                                                                                                                                   1'd0};
    else
      if (\lizzieLet34_4Lcall_main_map'_Int_Int3_1sc_0_12_1isZacL_2_1gacM_2_1q1acP_1_1q2acQ_1_1Lcall_main_map'_Int_Int2_r )
        \lizzieLet34_4Lcall_main_map'_Int_Int3_1sc_0_12_1isZacL_2_1gacM_2_1q1acP_1_1q2acQ_1_1Lcall_main_map'_Int_Int2_bufchan_d  <= \lizzieLet34_4Lcall_main_map'_Int_Int3_1sc_0_12_1isZacL_2_1gacM_2_1q1acP_1_1q2acQ_1_1Lcall_main_map'_Int_Int2_d ;
  \CTmain_map'_Int_Int_t  \lizzieLet34_4Lcall_main_map'_Int_Int3_1sc_0_12_1isZacL_2_1gacM_2_1q1acP_1_1q2acQ_1_1Lcall_main_map'_Int_Int2_bufchan_buf ;
  assign \lizzieLet34_4Lcall_main_map'_Int_Int3_1sc_0_12_1isZacL_2_1gacM_2_1q1acP_1_1q2acQ_1_1Lcall_main_map'_Int_Int2_bufchan_r  = (! \lizzieLet34_4Lcall_main_map'_Int_Int3_1sc_0_12_1isZacL_2_1gacM_2_1q1acP_1_1q2acQ_1_1Lcall_main_map'_Int_Int2_bufchan_buf [0]);
  assign lizzieLet35_1_argbuf_d = (\lizzieLet34_4Lcall_main_map'_Int_Int3_1sc_0_12_1isZacL_2_1gacM_2_1q1acP_1_1q2acQ_1_1Lcall_main_map'_Int_Int2_bufchan_buf [0] ? \lizzieLet34_4Lcall_main_map'_Int_Int3_1sc_0_12_1isZacL_2_1gacM_2_1q1acP_1_1q2acQ_1_1Lcall_main_map'_Int_Int2_bufchan_buf  :
                                   \lizzieLet34_4Lcall_main_map'_Int_Int3_1sc_0_12_1isZacL_2_1gacM_2_1q1acP_1_1q2acQ_1_1Lcall_main_map'_Int_Int2_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet34_4Lcall_main_map'_Int_Int3_1sc_0_12_1isZacL_2_1gacM_2_1q1acP_1_1q2acQ_1_1Lcall_main_map'_Int_Int2_bufchan_buf  <= {67'd0,
                                                                                                                                     1'd0};
    else
      if ((lizzieLet35_1_argbuf_r && \lizzieLet34_4Lcall_main_map'_Int_Int3_1sc_0_12_1isZacL_2_1gacM_2_1q1acP_1_1q2acQ_1_1Lcall_main_map'_Int_Int2_bufchan_buf [0]))
        \lizzieLet34_4Lcall_main_map'_Int_Int3_1sc_0_12_1isZacL_2_1gacM_2_1q1acP_1_1q2acQ_1_1Lcall_main_map'_Int_Int2_bufchan_buf  <= {67'd0,
                                                                                                                                       1'd0};
      else if (((! lizzieLet35_1_argbuf_r) && (! \lizzieLet34_4Lcall_main_map'_Int_Int3_1sc_0_12_1isZacL_2_1gacM_2_1q1acP_1_1q2acQ_1_1Lcall_main_map'_Int_Int2_bufchan_buf [0])))
        \lizzieLet34_4Lcall_main_map'_Int_Int3_1sc_0_12_1isZacL_2_1gacM_2_1q1acP_1_1q2acQ_1_1Lcall_main_map'_Int_Int2_bufchan_buf  <= \lizzieLet34_4Lcall_main_map'_Int_Int3_1sc_0_12_1isZacL_2_1gacM_2_1q1acP_1_1q2acQ_1_1Lcall_main_map'_Int_Int2_bufchan_d ;
  
  /* fork (Ty Pointer_QTree_Int) : (lizzieLet34_4Lmain_map'_Int_Intsbos,Pointer_QTree_Int) > [(lizzieLet34_4Lmain_map'_Int_Intsbos_1_merge_merge_fork_1,Pointer_QTree_Int),
                                                                                         (lizzieLet34_4Lmain_map'_Int_Intsbos_1_merge_merge_fork_2,Pointer_QTree_Int)] */
  logic [1:0] \lizzieLet34_4Lmain_map'_Int_Intsbos_emitted ;
  logic [1:0] \lizzieLet34_4Lmain_map'_Int_Intsbos_done ;
  assign \lizzieLet34_4Lmain_map'_Int_Intsbos_1_merge_merge_fork_1_d  = {\lizzieLet34_4Lmain_map'_Int_Intsbos_d [16:1],
                                                                         (\lizzieLet34_4Lmain_map'_Int_Intsbos_d [0] && (! \lizzieLet34_4Lmain_map'_Int_Intsbos_emitted [0]))};
  assign \lizzieLet34_4Lmain_map'_Int_Intsbos_1_merge_merge_fork_2_d  = {\lizzieLet34_4Lmain_map'_Int_Intsbos_d [16:1],
                                                                         (\lizzieLet34_4Lmain_map'_Int_Intsbos_d [0] && (! \lizzieLet34_4Lmain_map'_Int_Intsbos_emitted [1]))};
  assign \lizzieLet34_4Lmain_map'_Int_Intsbos_done  = (\lizzieLet34_4Lmain_map'_Int_Intsbos_emitted  | ({\lizzieLet34_4Lmain_map'_Int_Intsbos_1_merge_merge_fork_2_d [0],
                                                                                                         \lizzieLet34_4Lmain_map'_Int_Intsbos_1_merge_merge_fork_1_d [0]} & {\lizzieLet34_4Lmain_map'_Int_Intsbos_1_merge_merge_fork_2_r ,
                                                                                                                                                                             \lizzieLet34_4Lmain_map'_Int_Intsbos_1_merge_merge_fork_1_r }));
  assign \lizzieLet34_4Lmain_map'_Int_Intsbos_r  = (& \lizzieLet34_4Lmain_map'_Int_Intsbos_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet34_4Lmain_map'_Int_Intsbos_emitted  <= 2'd0;
    else
      \lizzieLet34_4Lmain_map'_Int_Intsbos_emitted  <= (\lizzieLet34_4Lmain_map'_Int_Intsbos_r  ? 2'd0 :
                                                        \lizzieLet34_4Lmain_map'_Int_Intsbos_done );
  
  /* togo (Ty Pointer_QTree_Int) : (lizzieLet34_4Lmain_map'_Int_Intsbos_1_merge_merge_fork_1,Pointer_QTree_Int) > (call_main_map'_Int_Int_goConst,Go) */
  assign \call_main_map'_Int_Int_goConst_d  = \lizzieLet34_4Lmain_map'_Int_Intsbos_1_merge_merge_fork_1_d [0];
  assign \lizzieLet34_4Lmain_map'_Int_Intsbos_1_merge_merge_fork_1_r  = \call_main_map'_Int_Int_goConst_r ;
  
  /* buf (Ty Pointer_QTree_Int) : (lizzieLet34_4Lmain_map'_Int_Intsbos_1_merge_merge_fork_2,Pointer_QTree_Int) > (main_map'_Int_Int_resbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t \lizzieLet34_4Lmain_map'_Int_Intsbos_1_merge_merge_fork_2_bufchan_d ;
  logic \lizzieLet34_4Lmain_map'_Int_Intsbos_1_merge_merge_fork_2_bufchan_r ;
  assign \lizzieLet34_4Lmain_map'_Int_Intsbos_1_merge_merge_fork_2_r  = ((! \lizzieLet34_4Lmain_map'_Int_Intsbos_1_merge_merge_fork_2_bufchan_d [0]) || \lizzieLet34_4Lmain_map'_Int_Intsbos_1_merge_merge_fork_2_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet34_4Lmain_map'_Int_Intsbos_1_merge_merge_fork_2_bufchan_d  <= {16'd0,
                                                                               1'd0};
    else
      if (\lizzieLet34_4Lmain_map'_Int_Intsbos_1_merge_merge_fork_2_r )
        \lizzieLet34_4Lmain_map'_Int_Intsbos_1_merge_merge_fork_2_bufchan_d  <= \lizzieLet34_4Lmain_map'_Int_Intsbos_1_merge_merge_fork_2_d ;
  Pointer_QTree_Int_t \lizzieLet34_4Lmain_map'_Int_Intsbos_1_merge_merge_fork_2_bufchan_buf ;
  assign \lizzieLet34_4Lmain_map'_Int_Intsbos_1_merge_merge_fork_2_bufchan_r  = (! \lizzieLet34_4Lmain_map'_Int_Intsbos_1_merge_merge_fork_2_bufchan_buf [0]);
  assign \main_map'_Int_Int_resbuf_d  = (\lizzieLet34_4Lmain_map'_Int_Intsbos_1_merge_merge_fork_2_bufchan_buf [0] ? \lizzieLet34_4Lmain_map'_Int_Intsbos_1_merge_merge_fork_2_bufchan_buf  :
                                         \lizzieLet34_4Lmain_map'_Int_Intsbos_1_merge_merge_fork_2_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet34_4Lmain_map'_Int_Intsbos_1_merge_merge_fork_2_bufchan_buf  <= {16'd0,
                                                                                 1'd0};
    else
      if ((\main_map'_Int_Int_resbuf_r  && \lizzieLet34_4Lmain_map'_Int_Intsbos_1_merge_merge_fork_2_bufchan_buf [0]))
        \lizzieLet34_4Lmain_map'_Int_Intsbos_1_merge_merge_fork_2_bufchan_buf  <= {16'd0,
                                                                                   1'd0};
      else if (((! \main_map'_Int_Int_resbuf_r ) && (! \lizzieLet34_4Lmain_map'_Int_Intsbos_1_merge_merge_fork_2_bufchan_buf [0])))
        \lizzieLet34_4Lmain_map'_Int_Intsbos_1_merge_merge_fork_2_bufchan_buf  <= \lizzieLet34_4Lmain_map'_Int_Intsbos_1_merge_merge_fork_2_bufchan_d ;
  
  /* destruct (Ty CTmap''_map''_Int_Int_Int,
          Dcon Lcall_map''_map''_Int_Int_Int0) : (lizzieLet39_1Lcall_map''_map''_Int_Int_Int0,CTmap''_map''_Int_Int_Int) > [(es_2_4_destruct,Pointer_QTree_Int),
                                                                                                                            (es_3_7_destruct,Pointer_QTree_Int),
                                                                                                                            (es_4_7_destruct,Pointer_QTree_Int),
                                                                                                                            (sc_0_19_destruct,Pointer_CTmap''_map''_Int_Int_Int)] */
  logic [3:0] \lizzieLet39_1Lcall_map''_map''_Int_Int_Int0_emitted ;
  logic [3:0] \lizzieLet39_1Lcall_map''_map''_Int_Int_Int0_done ;
  assign es_2_4_destruct_d = {\lizzieLet39_1Lcall_map''_map''_Int_Int_Int0_d [19:4],
                              (\lizzieLet39_1Lcall_map''_map''_Int_Int_Int0_d [0] && (! \lizzieLet39_1Lcall_map''_map''_Int_Int_Int0_emitted [0]))};
  assign es_3_7_destruct_d = {\lizzieLet39_1Lcall_map''_map''_Int_Int_Int0_d [35:20],
                              (\lizzieLet39_1Lcall_map''_map''_Int_Int_Int0_d [0] && (! \lizzieLet39_1Lcall_map''_map''_Int_Int_Int0_emitted [1]))};
  assign es_4_7_destruct_d = {\lizzieLet39_1Lcall_map''_map''_Int_Int_Int0_d [51:36],
                              (\lizzieLet39_1Lcall_map''_map''_Int_Int_Int0_d [0] && (! \lizzieLet39_1Lcall_map''_map''_Int_Int_Int0_emitted [2]))};
  assign sc_0_19_destruct_d = {\lizzieLet39_1Lcall_map''_map''_Int_Int_Int0_d [67:52],
                               (\lizzieLet39_1Lcall_map''_map''_Int_Int_Int0_d [0] && (! \lizzieLet39_1Lcall_map''_map''_Int_Int_Int0_emitted [3]))};
  assign \lizzieLet39_1Lcall_map''_map''_Int_Int_Int0_done  = (\lizzieLet39_1Lcall_map''_map''_Int_Int_Int0_emitted  | ({sc_0_19_destruct_d[0],
                                                                                                                         es_4_7_destruct_d[0],
                                                                                                                         es_3_7_destruct_d[0],
                                                                                                                         es_2_4_destruct_d[0]} & {sc_0_19_destruct_r,
                                                                                                                                                  es_4_7_destruct_r,
                                                                                                                                                  es_3_7_destruct_r,
                                                                                                                                                  es_2_4_destruct_r}));
  assign \lizzieLet39_1Lcall_map''_map''_Int_Int_Int0_r  = (& \lizzieLet39_1Lcall_map''_map''_Int_Int_Int0_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet39_1Lcall_map''_map''_Int_Int_Int0_emitted  <= 4'd0;
    else
      \lizzieLet39_1Lcall_map''_map''_Int_Int_Int0_emitted  <= (\lizzieLet39_1Lcall_map''_map''_Int_Int_Int0_r  ? 4'd0 :
                                                                \lizzieLet39_1Lcall_map''_map''_Int_Int_Int0_done );
  
  /* destruct (Ty CTmap''_map''_Int_Int_Int,
          Dcon Lcall_map''_map''_Int_Int_Int1) : (lizzieLet39_1Lcall_map''_map''_Int_Int_Int1,CTmap''_map''_Int_Int_Int) > [(es_3_6_destruct,Pointer_QTree_Int),
                                                                                                                            (es_4_6_destruct,Pointer_QTree_Int),
                                                                                                                            (sc_0_18_destruct,Pointer_CTmap''_map''_Int_Int_Int),
                                                                                                                            (isZacT_4_destruct,MyDTInt_Bool),
                                                                                                                            (gacU_4_destruct,MyDTInt_Int_Int),
                                                                                                                            (v'acV_4_destruct,Int),
                                                                                                                            (q1acY_3_destruct,Pointer_QTree_Int)] */
  logic [6:0] \lizzieLet39_1Lcall_map''_map''_Int_Int_Int1_emitted ;
  logic [6:0] \lizzieLet39_1Lcall_map''_map''_Int_Int_Int1_done ;
  assign es_3_6_destruct_d = {\lizzieLet39_1Lcall_map''_map''_Int_Int_Int1_d [19:4],
                              (\lizzieLet39_1Lcall_map''_map''_Int_Int_Int1_d [0] && (! \lizzieLet39_1Lcall_map''_map''_Int_Int_Int1_emitted [0]))};
  assign es_4_6_destruct_d = {\lizzieLet39_1Lcall_map''_map''_Int_Int_Int1_d [35:20],
                              (\lizzieLet39_1Lcall_map''_map''_Int_Int_Int1_d [0] && (! \lizzieLet39_1Lcall_map''_map''_Int_Int_Int1_emitted [1]))};
  assign sc_0_18_destruct_d = {\lizzieLet39_1Lcall_map''_map''_Int_Int_Int1_d [51:36],
                               (\lizzieLet39_1Lcall_map''_map''_Int_Int_Int1_d [0] && (! \lizzieLet39_1Lcall_map''_map''_Int_Int_Int1_emitted [2]))};
  assign isZacT_4_destruct_d = (\lizzieLet39_1Lcall_map''_map''_Int_Int_Int1_d [0] && (! \lizzieLet39_1Lcall_map''_map''_Int_Int_Int1_emitted [3]));
  assign gacU_4_destruct_d = (\lizzieLet39_1Lcall_map''_map''_Int_Int_Int1_d [0] && (! \lizzieLet39_1Lcall_map''_map''_Int_Int_Int1_emitted [4]));
  assign \v'acV_4_destruct_d  = {\lizzieLet39_1Lcall_map''_map''_Int_Int_Int1_d [83:52],
                                 (\lizzieLet39_1Lcall_map''_map''_Int_Int_Int1_d [0] && (! \lizzieLet39_1Lcall_map''_map''_Int_Int_Int1_emitted [5]))};
  assign q1acY_3_destruct_d = {\lizzieLet39_1Lcall_map''_map''_Int_Int_Int1_d [99:84],
                               (\lizzieLet39_1Lcall_map''_map''_Int_Int_Int1_d [0] && (! \lizzieLet39_1Lcall_map''_map''_Int_Int_Int1_emitted [6]))};
  assign \lizzieLet39_1Lcall_map''_map''_Int_Int_Int1_done  = (\lizzieLet39_1Lcall_map''_map''_Int_Int_Int1_emitted  | ({q1acY_3_destruct_d[0],
                                                                                                                         \v'acV_4_destruct_d [0],
                                                                                                                         gacU_4_destruct_d[0],
                                                                                                                         isZacT_4_destruct_d[0],
                                                                                                                         sc_0_18_destruct_d[0],
                                                                                                                         es_4_6_destruct_d[0],
                                                                                                                         es_3_6_destruct_d[0]} & {q1acY_3_destruct_r,
                                                                                                                                                  \v'acV_4_destruct_r ,
                                                                                                                                                  gacU_4_destruct_r,
                                                                                                                                                  isZacT_4_destruct_r,
                                                                                                                                                  sc_0_18_destruct_r,
                                                                                                                                                  es_4_6_destruct_r,
                                                                                                                                                  es_3_6_destruct_r}));
  assign \lizzieLet39_1Lcall_map''_map''_Int_Int_Int1_r  = (& \lizzieLet39_1Lcall_map''_map''_Int_Int_Int1_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet39_1Lcall_map''_map''_Int_Int_Int1_emitted  <= 7'd0;
    else
      \lizzieLet39_1Lcall_map''_map''_Int_Int_Int1_emitted  <= (\lizzieLet39_1Lcall_map''_map''_Int_Int_Int1_r  ? 7'd0 :
                                                                \lizzieLet39_1Lcall_map''_map''_Int_Int_Int1_done );
  
  /* destruct (Ty CTmap''_map''_Int_Int_Int,
          Dcon Lcall_map''_map''_Int_Int_Int2) : (lizzieLet39_1Lcall_map''_map''_Int_Int_Int2,CTmap''_map''_Int_Int_Int) > [(es_4_5_destruct,Pointer_QTree_Int),
                                                                                                                            (sc_0_17_destruct,Pointer_CTmap''_map''_Int_Int_Int),
                                                                                                                            (isZacT_3_destruct,MyDTInt_Bool),
                                                                                                                            (gacU_3_destruct,MyDTInt_Int_Int),
                                                                                                                            (v'acV_3_destruct,Int),
                                                                                                                            (q1acY_2_destruct,Pointer_QTree_Int),
                                                                                                                            (q2acZ_2_destruct,Pointer_QTree_Int)] */
  logic [6:0] \lizzieLet39_1Lcall_map''_map''_Int_Int_Int2_emitted ;
  logic [6:0] \lizzieLet39_1Lcall_map''_map''_Int_Int_Int2_done ;
  assign es_4_5_destruct_d = {\lizzieLet39_1Lcall_map''_map''_Int_Int_Int2_d [19:4],
                              (\lizzieLet39_1Lcall_map''_map''_Int_Int_Int2_d [0] && (! \lizzieLet39_1Lcall_map''_map''_Int_Int_Int2_emitted [0]))};
  assign sc_0_17_destruct_d = {\lizzieLet39_1Lcall_map''_map''_Int_Int_Int2_d [35:20],
                               (\lizzieLet39_1Lcall_map''_map''_Int_Int_Int2_d [0] && (! \lizzieLet39_1Lcall_map''_map''_Int_Int_Int2_emitted [1]))};
  assign isZacT_3_destruct_d = (\lizzieLet39_1Lcall_map''_map''_Int_Int_Int2_d [0] && (! \lizzieLet39_1Lcall_map''_map''_Int_Int_Int2_emitted [2]));
  assign gacU_3_destruct_d = (\lizzieLet39_1Lcall_map''_map''_Int_Int_Int2_d [0] && (! \lizzieLet39_1Lcall_map''_map''_Int_Int_Int2_emitted [3]));
  assign \v'acV_3_destruct_d  = {\lizzieLet39_1Lcall_map''_map''_Int_Int_Int2_d [67:36],
                                 (\lizzieLet39_1Lcall_map''_map''_Int_Int_Int2_d [0] && (! \lizzieLet39_1Lcall_map''_map''_Int_Int_Int2_emitted [4]))};
  assign q1acY_2_destruct_d = {\lizzieLet39_1Lcall_map''_map''_Int_Int_Int2_d [83:68],
                               (\lizzieLet39_1Lcall_map''_map''_Int_Int_Int2_d [0] && (! \lizzieLet39_1Lcall_map''_map''_Int_Int_Int2_emitted [5]))};
  assign q2acZ_2_destruct_d = {\lizzieLet39_1Lcall_map''_map''_Int_Int_Int2_d [99:84],
                               (\lizzieLet39_1Lcall_map''_map''_Int_Int_Int2_d [0] && (! \lizzieLet39_1Lcall_map''_map''_Int_Int_Int2_emitted [6]))};
  assign \lizzieLet39_1Lcall_map''_map''_Int_Int_Int2_done  = (\lizzieLet39_1Lcall_map''_map''_Int_Int_Int2_emitted  | ({q2acZ_2_destruct_d[0],
                                                                                                                         q1acY_2_destruct_d[0],
                                                                                                                         \v'acV_3_destruct_d [0],
                                                                                                                         gacU_3_destruct_d[0],
                                                                                                                         isZacT_3_destruct_d[0],
                                                                                                                         sc_0_17_destruct_d[0],
                                                                                                                         es_4_5_destruct_d[0]} & {q2acZ_2_destruct_r,
                                                                                                                                                  q1acY_2_destruct_r,
                                                                                                                                                  \v'acV_3_destruct_r ,
                                                                                                                                                  gacU_3_destruct_r,
                                                                                                                                                  isZacT_3_destruct_r,
                                                                                                                                                  sc_0_17_destruct_r,
                                                                                                                                                  es_4_5_destruct_r}));
  assign \lizzieLet39_1Lcall_map''_map''_Int_Int_Int2_r  = (& \lizzieLet39_1Lcall_map''_map''_Int_Int_Int2_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet39_1Lcall_map''_map''_Int_Int_Int2_emitted  <= 7'd0;
    else
      \lizzieLet39_1Lcall_map''_map''_Int_Int_Int2_emitted  <= (\lizzieLet39_1Lcall_map''_map''_Int_Int_Int2_r  ? 7'd0 :
                                                                \lizzieLet39_1Lcall_map''_map''_Int_Int_Int2_done );
  
  /* destruct (Ty CTmap''_map''_Int_Int_Int,
          Dcon Lcall_map''_map''_Int_Int_Int3) : (lizzieLet39_1Lcall_map''_map''_Int_Int_Int3,CTmap''_map''_Int_Int_Int) > [(sc_0_16_destruct,Pointer_CTmap''_map''_Int_Int_Int),
                                                                                                                            (isZacT_2_destruct,MyDTInt_Bool),
                                                                                                                            (gacU_2_destruct,MyDTInt_Int_Int),
                                                                                                                            (v'acV_2_destruct,Int),
                                                                                                                            (q1acY_1_destruct,Pointer_QTree_Int),
                                                                                                                            (q2acZ_1_destruct,Pointer_QTree_Int),
                                                                                                                            (q3ad0_1_destruct,Pointer_QTree_Int)] */
  logic [6:0] \lizzieLet39_1Lcall_map''_map''_Int_Int_Int3_emitted ;
  logic [6:0] \lizzieLet39_1Lcall_map''_map''_Int_Int_Int3_done ;
  assign sc_0_16_destruct_d = {\lizzieLet39_1Lcall_map''_map''_Int_Int_Int3_d [19:4],
                               (\lizzieLet39_1Lcall_map''_map''_Int_Int_Int3_d [0] && (! \lizzieLet39_1Lcall_map''_map''_Int_Int_Int3_emitted [0]))};
  assign isZacT_2_destruct_d = (\lizzieLet39_1Lcall_map''_map''_Int_Int_Int3_d [0] && (! \lizzieLet39_1Lcall_map''_map''_Int_Int_Int3_emitted [1]));
  assign gacU_2_destruct_d = (\lizzieLet39_1Lcall_map''_map''_Int_Int_Int3_d [0] && (! \lizzieLet39_1Lcall_map''_map''_Int_Int_Int3_emitted [2]));
  assign \v'acV_2_destruct_d  = {\lizzieLet39_1Lcall_map''_map''_Int_Int_Int3_d [51:20],
                                 (\lizzieLet39_1Lcall_map''_map''_Int_Int_Int3_d [0] && (! \lizzieLet39_1Lcall_map''_map''_Int_Int_Int3_emitted [3]))};
  assign q1acY_1_destruct_d = {\lizzieLet39_1Lcall_map''_map''_Int_Int_Int3_d [67:52],
                               (\lizzieLet39_1Lcall_map''_map''_Int_Int_Int3_d [0] && (! \lizzieLet39_1Lcall_map''_map''_Int_Int_Int3_emitted [4]))};
  assign q2acZ_1_destruct_d = {\lizzieLet39_1Lcall_map''_map''_Int_Int_Int3_d [83:68],
                               (\lizzieLet39_1Lcall_map''_map''_Int_Int_Int3_d [0] && (! \lizzieLet39_1Lcall_map''_map''_Int_Int_Int3_emitted [5]))};
  assign q3ad0_1_destruct_d = {\lizzieLet39_1Lcall_map''_map''_Int_Int_Int3_d [99:84],
                               (\lizzieLet39_1Lcall_map''_map''_Int_Int_Int3_d [0] && (! \lizzieLet39_1Lcall_map''_map''_Int_Int_Int3_emitted [6]))};
  assign \lizzieLet39_1Lcall_map''_map''_Int_Int_Int3_done  = (\lizzieLet39_1Lcall_map''_map''_Int_Int_Int3_emitted  | ({q3ad0_1_destruct_d[0],
                                                                                                                         q2acZ_1_destruct_d[0],
                                                                                                                         q1acY_1_destruct_d[0],
                                                                                                                         \v'acV_2_destruct_d [0],
                                                                                                                         gacU_2_destruct_d[0],
                                                                                                                         isZacT_2_destruct_d[0],
                                                                                                                         sc_0_16_destruct_d[0]} & {q3ad0_1_destruct_r,
                                                                                                                                                   q2acZ_1_destruct_r,
                                                                                                                                                   q1acY_1_destruct_r,
                                                                                                                                                   \v'acV_2_destruct_r ,
                                                                                                                                                   gacU_2_destruct_r,
                                                                                                                                                   isZacT_2_destruct_r,
                                                                                                                                                   sc_0_16_destruct_r}));
  assign \lizzieLet39_1Lcall_map''_map''_Int_Int_Int3_r  = (& \lizzieLet39_1Lcall_map''_map''_Int_Int_Int3_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet39_1Lcall_map''_map''_Int_Int_Int3_emitted  <= 7'd0;
    else
      \lizzieLet39_1Lcall_map''_map''_Int_Int_Int3_emitted  <= (\lizzieLet39_1Lcall_map''_map''_Int_Int_Int3_r  ? 7'd0 :
                                                                \lizzieLet39_1Lcall_map''_map''_Int_Int_Int3_done );
  
  /* demux (Ty CTmap''_map''_Int_Int_Int,
       Ty CTmap''_map''_Int_Int_Int) : (lizzieLet39_2,CTmap''_map''_Int_Int_Int) (lizzieLet39_1,CTmap''_map''_Int_Int_Int) > [(_12,CTmap''_map''_Int_Int_Int),
                                                                                                                              (lizzieLet39_1Lcall_map''_map''_Int_Int_Int3,CTmap''_map''_Int_Int_Int),
                                                                                                                              (lizzieLet39_1Lcall_map''_map''_Int_Int_Int2,CTmap''_map''_Int_Int_Int),
                                                                                                                              (lizzieLet39_1Lcall_map''_map''_Int_Int_Int1,CTmap''_map''_Int_Int_Int),
                                                                                                                              (lizzieLet39_1Lcall_map''_map''_Int_Int_Int0,CTmap''_map''_Int_Int_Int)] */
  logic [4:0] lizzieLet39_1_onehotd;
  always_comb
    if ((lizzieLet39_2_d[0] && lizzieLet39_1_d[0]))
      unique case (lizzieLet39_2_d[3:1])
        3'd0: lizzieLet39_1_onehotd = 5'd1;
        3'd1: lizzieLet39_1_onehotd = 5'd2;
        3'd2: lizzieLet39_1_onehotd = 5'd4;
        3'd3: lizzieLet39_1_onehotd = 5'd8;
        3'd4: lizzieLet39_1_onehotd = 5'd16;
        default: lizzieLet39_1_onehotd = 5'd0;
      endcase
    else lizzieLet39_1_onehotd = 5'd0;
  assign _12_d = {lizzieLet39_1_d[99:1], lizzieLet39_1_onehotd[0]};
  assign \lizzieLet39_1Lcall_map''_map''_Int_Int_Int3_d  = {lizzieLet39_1_d[99:1],
                                                            lizzieLet39_1_onehotd[1]};
  assign \lizzieLet39_1Lcall_map''_map''_Int_Int_Int2_d  = {lizzieLet39_1_d[99:1],
                                                            lizzieLet39_1_onehotd[2]};
  assign \lizzieLet39_1Lcall_map''_map''_Int_Int_Int1_d  = {lizzieLet39_1_d[99:1],
                                                            lizzieLet39_1_onehotd[3]};
  assign \lizzieLet39_1Lcall_map''_map''_Int_Int_Int0_d  = {lizzieLet39_1_d[99:1],
                                                            lizzieLet39_1_onehotd[4]};
  assign lizzieLet39_1_r = (| (lizzieLet39_1_onehotd & {\lizzieLet39_1Lcall_map''_map''_Int_Int_Int0_r ,
                                                        \lizzieLet39_1Lcall_map''_map''_Int_Int_Int1_r ,
                                                        \lizzieLet39_1Lcall_map''_map''_Int_Int_Int2_r ,
                                                        \lizzieLet39_1Lcall_map''_map''_Int_Int_Int3_r ,
                                                        _12_r}));
  assign lizzieLet39_2_r = lizzieLet39_1_r;
  
  /* demux (Ty CTmap''_map''_Int_Int_Int,
       Ty Go) : (lizzieLet39_3,CTmap''_map''_Int_Int_Int) (go_21_goMux_data,Go) > [(_11,Go),
                                                                                   (lizzieLet39_3Lcall_map''_map''_Int_Int_Int3,Go),
                                                                                   (lizzieLet39_3Lcall_map''_map''_Int_Int_Int2,Go),
                                                                                   (lizzieLet39_3Lcall_map''_map''_Int_Int_Int1,Go),
                                                                                   (lizzieLet39_3Lcall_map''_map''_Int_Int_Int0,Go)] */
  logic [4:0] go_21_goMux_data_onehotd;
  always_comb
    if ((lizzieLet39_3_d[0] && go_21_goMux_data_d[0]))
      unique case (lizzieLet39_3_d[3:1])
        3'd0: go_21_goMux_data_onehotd = 5'd1;
        3'd1: go_21_goMux_data_onehotd = 5'd2;
        3'd2: go_21_goMux_data_onehotd = 5'd4;
        3'd3: go_21_goMux_data_onehotd = 5'd8;
        3'd4: go_21_goMux_data_onehotd = 5'd16;
        default: go_21_goMux_data_onehotd = 5'd0;
      endcase
    else go_21_goMux_data_onehotd = 5'd0;
  assign _11_d = go_21_goMux_data_onehotd[0];
  assign \lizzieLet39_3Lcall_map''_map''_Int_Int_Int3_d  = go_21_goMux_data_onehotd[1];
  assign \lizzieLet39_3Lcall_map''_map''_Int_Int_Int2_d  = go_21_goMux_data_onehotd[2];
  assign \lizzieLet39_3Lcall_map''_map''_Int_Int_Int1_d  = go_21_goMux_data_onehotd[3];
  assign \lizzieLet39_3Lcall_map''_map''_Int_Int_Int0_d  = go_21_goMux_data_onehotd[4];
  assign go_21_goMux_data_r = (| (go_21_goMux_data_onehotd & {\lizzieLet39_3Lcall_map''_map''_Int_Int_Int0_r ,
                                                              \lizzieLet39_3Lcall_map''_map''_Int_Int_Int1_r ,
                                                              \lizzieLet39_3Lcall_map''_map''_Int_Int_Int2_r ,
                                                              \lizzieLet39_3Lcall_map''_map''_Int_Int_Int3_r ,
                                                              _11_r}));
  assign lizzieLet39_3_r = go_21_goMux_data_r;
  
  /* buf (Ty Go) : (lizzieLet39_3Lcall_map''_map''_Int_Int_Int0,Go) > (lizzieLet39_3Lcall_map''_map''_Int_Int_Int0_1_argbuf,Go) */
  Go_t \lizzieLet39_3Lcall_map''_map''_Int_Int_Int0_bufchan_d ;
  logic \lizzieLet39_3Lcall_map''_map''_Int_Int_Int0_bufchan_r ;
  assign \lizzieLet39_3Lcall_map''_map''_Int_Int_Int0_r  = ((! \lizzieLet39_3Lcall_map''_map''_Int_Int_Int0_bufchan_d [0]) || \lizzieLet39_3Lcall_map''_map''_Int_Int_Int0_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet39_3Lcall_map''_map''_Int_Int_Int0_bufchan_d  <= 1'd0;
    else
      if (\lizzieLet39_3Lcall_map''_map''_Int_Int_Int0_r )
        \lizzieLet39_3Lcall_map''_map''_Int_Int_Int0_bufchan_d  <= \lizzieLet39_3Lcall_map''_map''_Int_Int_Int0_d ;
  Go_t \lizzieLet39_3Lcall_map''_map''_Int_Int_Int0_bufchan_buf ;
  assign \lizzieLet39_3Lcall_map''_map''_Int_Int_Int0_bufchan_r  = (! \lizzieLet39_3Lcall_map''_map''_Int_Int_Int0_bufchan_buf [0]);
  assign \lizzieLet39_3Lcall_map''_map''_Int_Int_Int0_1_argbuf_d  = (\lizzieLet39_3Lcall_map''_map''_Int_Int_Int0_bufchan_buf [0] ? \lizzieLet39_3Lcall_map''_map''_Int_Int_Int0_bufchan_buf  :
                                                                     \lizzieLet39_3Lcall_map''_map''_Int_Int_Int0_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet39_3Lcall_map''_map''_Int_Int_Int0_bufchan_buf  <= 1'd0;
    else
      if ((\lizzieLet39_3Lcall_map''_map''_Int_Int_Int0_1_argbuf_r  && \lizzieLet39_3Lcall_map''_map''_Int_Int_Int0_bufchan_buf [0]))
        \lizzieLet39_3Lcall_map''_map''_Int_Int_Int0_bufchan_buf  <= 1'd0;
      else if (((! \lizzieLet39_3Lcall_map''_map''_Int_Int_Int0_1_argbuf_r ) && (! \lizzieLet39_3Lcall_map''_map''_Int_Int_Int0_bufchan_buf [0])))
        \lizzieLet39_3Lcall_map''_map''_Int_Int_Int0_bufchan_buf  <= \lizzieLet39_3Lcall_map''_map''_Int_Int_Int0_bufchan_d ;
  
  /* buf (Ty Go) : (lizzieLet39_3Lcall_map''_map''_Int_Int_Int1,Go) > (lizzieLet39_3Lcall_map''_map''_Int_Int_Int1_1_argbuf,Go) */
  Go_t \lizzieLet39_3Lcall_map''_map''_Int_Int_Int1_bufchan_d ;
  logic \lizzieLet39_3Lcall_map''_map''_Int_Int_Int1_bufchan_r ;
  assign \lizzieLet39_3Lcall_map''_map''_Int_Int_Int1_r  = ((! \lizzieLet39_3Lcall_map''_map''_Int_Int_Int1_bufchan_d [0]) || \lizzieLet39_3Lcall_map''_map''_Int_Int_Int1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet39_3Lcall_map''_map''_Int_Int_Int1_bufchan_d  <= 1'd0;
    else
      if (\lizzieLet39_3Lcall_map''_map''_Int_Int_Int1_r )
        \lizzieLet39_3Lcall_map''_map''_Int_Int_Int1_bufchan_d  <= \lizzieLet39_3Lcall_map''_map''_Int_Int_Int1_d ;
  Go_t \lizzieLet39_3Lcall_map''_map''_Int_Int_Int1_bufchan_buf ;
  assign \lizzieLet39_3Lcall_map''_map''_Int_Int_Int1_bufchan_r  = (! \lizzieLet39_3Lcall_map''_map''_Int_Int_Int1_bufchan_buf [0]);
  assign \lizzieLet39_3Lcall_map''_map''_Int_Int_Int1_1_argbuf_d  = (\lizzieLet39_3Lcall_map''_map''_Int_Int_Int1_bufchan_buf [0] ? \lizzieLet39_3Lcall_map''_map''_Int_Int_Int1_bufchan_buf  :
                                                                     \lizzieLet39_3Lcall_map''_map''_Int_Int_Int1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet39_3Lcall_map''_map''_Int_Int_Int1_bufchan_buf  <= 1'd0;
    else
      if ((\lizzieLet39_3Lcall_map''_map''_Int_Int_Int1_1_argbuf_r  && \lizzieLet39_3Lcall_map''_map''_Int_Int_Int1_bufchan_buf [0]))
        \lizzieLet39_3Lcall_map''_map''_Int_Int_Int1_bufchan_buf  <= 1'd0;
      else if (((! \lizzieLet39_3Lcall_map''_map''_Int_Int_Int1_1_argbuf_r ) && (! \lizzieLet39_3Lcall_map''_map''_Int_Int_Int1_bufchan_buf [0])))
        \lizzieLet39_3Lcall_map''_map''_Int_Int_Int1_bufchan_buf  <= \lizzieLet39_3Lcall_map''_map''_Int_Int_Int1_bufchan_d ;
  
  /* buf (Ty Go) : (lizzieLet39_3Lcall_map''_map''_Int_Int_Int2,Go) > (lizzieLet39_3Lcall_map''_map''_Int_Int_Int2_1_argbuf,Go) */
  Go_t \lizzieLet39_3Lcall_map''_map''_Int_Int_Int2_bufchan_d ;
  logic \lizzieLet39_3Lcall_map''_map''_Int_Int_Int2_bufchan_r ;
  assign \lizzieLet39_3Lcall_map''_map''_Int_Int_Int2_r  = ((! \lizzieLet39_3Lcall_map''_map''_Int_Int_Int2_bufchan_d [0]) || \lizzieLet39_3Lcall_map''_map''_Int_Int_Int2_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet39_3Lcall_map''_map''_Int_Int_Int2_bufchan_d  <= 1'd0;
    else
      if (\lizzieLet39_3Lcall_map''_map''_Int_Int_Int2_r )
        \lizzieLet39_3Lcall_map''_map''_Int_Int_Int2_bufchan_d  <= \lizzieLet39_3Lcall_map''_map''_Int_Int_Int2_d ;
  Go_t \lizzieLet39_3Lcall_map''_map''_Int_Int_Int2_bufchan_buf ;
  assign \lizzieLet39_3Lcall_map''_map''_Int_Int_Int2_bufchan_r  = (! \lizzieLet39_3Lcall_map''_map''_Int_Int_Int2_bufchan_buf [0]);
  assign \lizzieLet39_3Lcall_map''_map''_Int_Int_Int2_1_argbuf_d  = (\lizzieLet39_3Lcall_map''_map''_Int_Int_Int2_bufchan_buf [0] ? \lizzieLet39_3Lcall_map''_map''_Int_Int_Int2_bufchan_buf  :
                                                                     \lizzieLet39_3Lcall_map''_map''_Int_Int_Int2_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet39_3Lcall_map''_map''_Int_Int_Int2_bufchan_buf  <= 1'd0;
    else
      if ((\lizzieLet39_3Lcall_map''_map''_Int_Int_Int2_1_argbuf_r  && \lizzieLet39_3Lcall_map''_map''_Int_Int_Int2_bufchan_buf [0]))
        \lizzieLet39_3Lcall_map''_map''_Int_Int_Int2_bufchan_buf  <= 1'd0;
      else if (((! \lizzieLet39_3Lcall_map''_map''_Int_Int_Int2_1_argbuf_r ) && (! \lizzieLet39_3Lcall_map''_map''_Int_Int_Int2_bufchan_buf [0])))
        \lizzieLet39_3Lcall_map''_map''_Int_Int_Int2_bufchan_buf  <= \lizzieLet39_3Lcall_map''_map''_Int_Int_Int2_bufchan_d ;
  
  /* buf (Ty Go) : (lizzieLet39_3Lcall_map''_map''_Int_Int_Int3,Go) > (lizzieLet39_3Lcall_map''_map''_Int_Int_Int3_1_argbuf,Go) */
  Go_t \lizzieLet39_3Lcall_map''_map''_Int_Int_Int3_bufchan_d ;
  logic \lizzieLet39_3Lcall_map''_map''_Int_Int_Int3_bufchan_r ;
  assign \lizzieLet39_3Lcall_map''_map''_Int_Int_Int3_r  = ((! \lizzieLet39_3Lcall_map''_map''_Int_Int_Int3_bufchan_d [0]) || \lizzieLet39_3Lcall_map''_map''_Int_Int_Int3_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet39_3Lcall_map''_map''_Int_Int_Int3_bufchan_d  <= 1'd0;
    else
      if (\lizzieLet39_3Lcall_map''_map''_Int_Int_Int3_r )
        \lizzieLet39_3Lcall_map''_map''_Int_Int_Int3_bufchan_d  <= \lizzieLet39_3Lcall_map''_map''_Int_Int_Int3_d ;
  Go_t \lizzieLet39_3Lcall_map''_map''_Int_Int_Int3_bufchan_buf ;
  assign \lizzieLet39_3Lcall_map''_map''_Int_Int_Int3_bufchan_r  = (! \lizzieLet39_3Lcall_map''_map''_Int_Int_Int3_bufchan_buf [0]);
  assign \lizzieLet39_3Lcall_map''_map''_Int_Int_Int3_1_argbuf_d  = (\lizzieLet39_3Lcall_map''_map''_Int_Int_Int3_bufchan_buf [0] ? \lizzieLet39_3Lcall_map''_map''_Int_Int_Int3_bufchan_buf  :
                                                                     \lizzieLet39_3Lcall_map''_map''_Int_Int_Int3_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet39_3Lcall_map''_map''_Int_Int_Int3_bufchan_buf  <= 1'd0;
    else
      if ((\lizzieLet39_3Lcall_map''_map''_Int_Int_Int3_1_argbuf_r  && \lizzieLet39_3Lcall_map''_map''_Int_Int_Int3_bufchan_buf [0]))
        \lizzieLet39_3Lcall_map''_map''_Int_Int_Int3_bufchan_buf  <= 1'd0;
      else if (((! \lizzieLet39_3Lcall_map''_map''_Int_Int_Int3_1_argbuf_r ) && (! \lizzieLet39_3Lcall_map''_map''_Int_Int_Int3_bufchan_buf [0])))
        \lizzieLet39_3Lcall_map''_map''_Int_Int_Int3_bufchan_buf  <= \lizzieLet39_3Lcall_map''_map''_Int_Int_Int3_bufchan_d ;
  
  /* demux (Ty CTmap''_map''_Int_Int_Int,
       Ty Pointer_QTree_Int) : (lizzieLet39_4,CTmap''_map''_Int_Int_Int) (srtarg_0_3_goMux_mux,Pointer_QTree_Int) > [(lizzieLet39_4Lmap''_map''_Int_Int_Intsbos,Pointer_QTree_Int),
                                                                                                                     (lizzieLet39_4Lcall_map''_map''_Int_Int_Int3,Pointer_QTree_Int),
                                                                                                                     (lizzieLet39_4Lcall_map''_map''_Int_Int_Int2,Pointer_QTree_Int),
                                                                                                                     (lizzieLet39_4Lcall_map''_map''_Int_Int_Int1,Pointer_QTree_Int),
                                                                                                                     (lizzieLet39_4Lcall_map''_map''_Int_Int_Int0,Pointer_QTree_Int)] */
  logic [4:0] srtarg_0_3_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet39_4_d[0] && srtarg_0_3_goMux_mux_d[0]))
      unique case (lizzieLet39_4_d[3:1])
        3'd0: srtarg_0_3_goMux_mux_onehotd = 5'd1;
        3'd1: srtarg_0_3_goMux_mux_onehotd = 5'd2;
        3'd2: srtarg_0_3_goMux_mux_onehotd = 5'd4;
        3'd3: srtarg_0_3_goMux_mux_onehotd = 5'd8;
        3'd4: srtarg_0_3_goMux_mux_onehotd = 5'd16;
        default: srtarg_0_3_goMux_mux_onehotd = 5'd0;
      endcase
    else srtarg_0_3_goMux_mux_onehotd = 5'd0;
  assign \lizzieLet39_4Lmap''_map''_Int_Int_Intsbos_d  = {srtarg_0_3_goMux_mux_d[16:1],
                                                          srtarg_0_3_goMux_mux_onehotd[0]};
  assign \lizzieLet39_4Lcall_map''_map''_Int_Int_Int3_d  = {srtarg_0_3_goMux_mux_d[16:1],
                                                            srtarg_0_3_goMux_mux_onehotd[1]};
  assign \lizzieLet39_4Lcall_map''_map''_Int_Int_Int2_d  = {srtarg_0_3_goMux_mux_d[16:1],
                                                            srtarg_0_3_goMux_mux_onehotd[2]};
  assign \lizzieLet39_4Lcall_map''_map''_Int_Int_Int1_d  = {srtarg_0_3_goMux_mux_d[16:1],
                                                            srtarg_0_3_goMux_mux_onehotd[3]};
  assign \lizzieLet39_4Lcall_map''_map''_Int_Int_Int0_d  = {srtarg_0_3_goMux_mux_d[16:1],
                                                            srtarg_0_3_goMux_mux_onehotd[4]};
  assign srtarg_0_3_goMux_mux_r = (| (srtarg_0_3_goMux_mux_onehotd & {\lizzieLet39_4Lcall_map''_map''_Int_Int_Int0_r ,
                                                                      \lizzieLet39_4Lcall_map''_map''_Int_Int_Int1_r ,
                                                                      \lizzieLet39_4Lcall_map''_map''_Int_Int_Int2_r ,
                                                                      \lizzieLet39_4Lcall_map''_map''_Int_Int_Int3_r ,
                                                                      \lizzieLet39_4Lmap''_map''_Int_Int_Intsbos_r }));
  assign lizzieLet39_4_r = srtarg_0_3_goMux_mux_r;
  
  /* dcon (Ty QTree_Int,
      Dcon QNode_Int) : [(lizzieLet39_4Lcall_map''_map''_Int_Int_Int0,Pointer_QTree_Int),
                         (es_2_4_destruct,Pointer_QTree_Int),
                         (es_3_7_destruct,Pointer_QTree_Int),
                         (es_4_7_destruct,Pointer_QTree_Int)] > (lizzieLet39_4Lcall_map''_map''_Int_Int_Int0_1es_2_4_1es_3_7_1es_4_7_1QNode_Int,QTree_Int) */
  assign \lizzieLet39_4Lcall_map''_map''_Int_Int_Int0_1es_2_4_1es_3_7_1es_4_7_1QNode_Int_d  = QNode_Int_dc((& {\lizzieLet39_4Lcall_map''_map''_Int_Int_Int0_d [0],
                                                                                                               es_2_4_destruct_d[0],
                                                                                                               es_3_7_destruct_d[0],
                                                                                                               es_4_7_destruct_d[0]}), \lizzieLet39_4Lcall_map''_map''_Int_Int_Int0_d , es_2_4_destruct_d, es_3_7_destruct_d, es_4_7_destruct_d);
  assign {\lizzieLet39_4Lcall_map''_map''_Int_Int_Int0_r ,
          es_2_4_destruct_r,
          es_3_7_destruct_r,
          es_4_7_destruct_r} = {4 {(\lizzieLet39_4Lcall_map''_map''_Int_Int_Int0_1es_2_4_1es_3_7_1es_4_7_1QNode_Int_r  && \lizzieLet39_4Lcall_map''_map''_Int_Int_Int0_1es_2_4_1es_3_7_1es_4_7_1QNode_Int_d [0])}};
  
  /* buf (Ty QTree_Int) : (lizzieLet39_4Lcall_map''_map''_Int_Int_Int0_1es_2_4_1es_3_7_1es_4_7_1QNode_Int,QTree_Int) > (lizzieLet43_1_argbuf,QTree_Int) */
  QTree_Int_t \lizzieLet39_4Lcall_map''_map''_Int_Int_Int0_1es_2_4_1es_3_7_1es_4_7_1QNode_Int_bufchan_d ;
  logic \lizzieLet39_4Lcall_map''_map''_Int_Int_Int0_1es_2_4_1es_3_7_1es_4_7_1QNode_Int_bufchan_r ;
  assign \lizzieLet39_4Lcall_map''_map''_Int_Int_Int0_1es_2_4_1es_3_7_1es_4_7_1QNode_Int_r  = ((! \lizzieLet39_4Lcall_map''_map''_Int_Int_Int0_1es_2_4_1es_3_7_1es_4_7_1QNode_Int_bufchan_d [0]) || \lizzieLet39_4Lcall_map''_map''_Int_Int_Int0_1es_2_4_1es_3_7_1es_4_7_1QNode_Int_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet39_4Lcall_map''_map''_Int_Int_Int0_1es_2_4_1es_3_7_1es_4_7_1QNode_Int_bufchan_d  <= {66'd0,
                                                                                                     1'd0};
    else
      if (\lizzieLet39_4Lcall_map''_map''_Int_Int_Int0_1es_2_4_1es_3_7_1es_4_7_1QNode_Int_r )
        \lizzieLet39_4Lcall_map''_map''_Int_Int_Int0_1es_2_4_1es_3_7_1es_4_7_1QNode_Int_bufchan_d  <= \lizzieLet39_4Lcall_map''_map''_Int_Int_Int0_1es_2_4_1es_3_7_1es_4_7_1QNode_Int_d ;
  QTree_Int_t \lizzieLet39_4Lcall_map''_map''_Int_Int_Int0_1es_2_4_1es_3_7_1es_4_7_1QNode_Int_bufchan_buf ;
  assign \lizzieLet39_4Lcall_map''_map''_Int_Int_Int0_1es_2_4_1es_3_7_1es_4_7_1QNode_Int_bufchan_r  = (! \lizzieLet39_4Lcall_map''_map''_Int_Int_Int0_1es_2_4_1es_3_7_1es_4_7_1QNode_Int_bufchan_buf [0]);
  assign lizzieLet43_1_argbuf_d = (\lizzieLet39_4Lcall_map''_map''_Int_Int_Int0_1es_2_4_1es_3_7_1es_4_7_1QNode_Int_bufchan_buf [0] ? \lizzieLet39_4Lcall_map''_map''_Int_Int_Int0_1es_2_4_1es_3_7_1es_4_7_1QNode_Int_bufchan_buf  :
                                   \lizzieLet39_4Lcall_map''_map''_Int_Int_Int0_1es_2_4_1es_3_7_1es_4_7_1QNode_Int_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet39_4Lcall_map''_map''_Int_Int_Int0_1es_2_4_1es_3_7_1es_4_7_1QNode_Int_bufchan_buf  <= {66'd0,
                                                                                                       1'd0};
    else
      if ((lizzieLet43_1_argbuf_r && \lizzieLet39_4Lcall_map''_map''_Int_Int_Int0_1es_2_4_1es_3_7_1es_4_7_1QNode_Int_bufchan_buf [0]))
        \lizzieLet39_4Lcall_map''_map''_Int_Int_Int0_1es_2_4_1es_3_7_1es_4_7_1QNode_Int_bufchan_buf  <= {66'd0,
                                                                                                         1'd0};
      else if (((! lizzieLet43_1_argbuf_r) && (! \lizzieLet39_4Lcall_map''_map''_Int_Int_Int0_1es_2_4_1es_3_7_1es_4_7_1QNode_Int_bufchan_buf [0])))
        \lizzieLet39_4Lcall_map''_map''_Int_Int_Int0_1es_2_4_1es_3_7_1es_4_7_1QNode_Int_bufchan_buf  <= \lizzieLet39_4Lcall_map''_map''_Int_Int_Int0_1es_2_4_1es_3_7_1es_4_7_1QNode_Int_bufchan_d ;
  
  /* dcon (Ty CTmap''_map''_Int_Int_Int,
      Dcon Lcall_map''_map''_Int_Int_Int0) : [(lizzieLet39_4Lcall_map''_map''_Int_Int_Int1,Pointer_QTree_Int),
                                              (es_3_6_destruct,Pointer_QTree_Int),
                                              (es_4_6_destruct,Pointer_QTree_Int),
                                              (sc_0_18_destruct,Pointer_CTmap''_map''_Int_Int_Int)] > (lizzieLet39_4Lcall_map''_map''_Int_Int_Int1_1es_3_6_1es_4_6_1sc_0_18_1Lcall_map''_map''_Int_Int_Int0,CTmap''_map''_Int_Int_Int) */
  assign \lizzieLet39_4Lcall_map''_map''_Int_Int_Int1_1es_3_6_1es_4_6_1sc_0_18_1Lcall_map''_map''_Int_Int_Int0_d  = \Lcall_map''_map''_Int_Int_Int0_dc ((& {\lizzieLet39_4Lcall_map''_map''_Int_Int_Int1_d [0],
                                                                                                                                                            es_3_6_destruct_d[0],
                                                                                                                                                            es_4_6_destruct_d[0],
                                                                                                                                                            sc_0_18_destruct_d[0]}), \lizzieLet39_4Lcall_map''_map''_Int_Int_Int1_d , es_3_6_destruct_d, es_4_6_destruct_d, sc_0_18_destruct_d);
  assign {\lizzieLet39_4Lcall_map''_map''_Int_Int_Int1_r ,
          es_3_6_destruct_r,
          es_4_6_destruct_r,
          sc_0_18_destruct_r} = {4 {(\lizzieLet39_4Lcall_map''_map''_Int_Int_Int1_1es_3_6_1es_4_6_1sc_0_18_1Lcall_map''_map''_Int_Int_Int0_r  && \lizzieLet39_4Lcall_map''_map''_Int_Int_Int1_1es_3_6_1es_4_6_1sc_0_18_1Lcall_map''_map''_Int_Int_Int0_d [0])}};
  
  /* buf (Ty CTmap''_map''_Int_Int_Int) : (lizzieLet39_4Lcall_map''_map''_Int_Int_Int1_1es_3_6_1es_4_6_1sc_0_18_1Lcall_map''_map''_Int_Int_Int0,CTmap''_map''_Int_Int_Int) > (lizzieLet42_1_argbuf,CTmap''_map''_Int_Int_Int) */
  \CTmap''_map''_Int_Int_Int_t  \lizzieLet39_4Lcall_map''_map''_Int_Int_Int1_1es_3_6_1es_4_6_1sc_0_18_1Lcall_map''_map''_Int_Int_Int0_bufchan_d ;
  logic \lizzieLet39_4Lcall_map''_map''_Int_Int_Int1_1es_3_6_1es_4_6_1sc_0_18_1Lcall_map''_map''_Int_Int_Int0_bufchan_r ;
  assign \lizzieLet39_4Lcall_map''_map''_Int_Int_Int1_1es_3_6_1es_4_6_1sc_0_18_1Lcall_map''_map''_Int_Int_Int0_r  = ((! \lizzieLet39_4Lcall_map''_map''_Int_Int_Int1_1es_3_6_1es_4_6_1sc_0_18_1Lcall_map''_map''_Int_Int_Int0_bufchan_d [0]) || \lizzieLet39_4Lcall_map''_map''_Int_Int_Int1_1es_3_6_1es_4_6_1sc_0_18_1Lcall_map''_map''_Int_Int_Int0_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet39_4Lcall_map''_map''_Int_Int_Int1_1es_3_6_1es_4_6_1sc_0_18_1Lcall_map''_map''_Int_Int_Int0_bufchan_d  <= {99'd0,
                                                                                                                           1'd0};
    else
      if (\lizzieLet39_4Lcall_map''_map''_Int_Int_Int1_1es_3_6_1es_4_6_1sc_0_18_1Lcall_map''_map''_Int_Int_Int0_r )
        \lizzieLet39_4Lcall_map''_map''_Int_Int_Int1_1es_3_6_1es_4_6_1sc_0_18_1Lcall_map''_map''_Int_Int_Int0_bufchan_d  <= \lizzieLet39_4Lcall_map''_map''_Int_Int_Int1_1es_3_6_1es_4_6_1sc_0_18_1Lcall_map''_map''_Int_Int_Int0_d ;
  \CTmap''_map''_Int_Int_Int_t  \lizzieLet39_4Lcall_map''_map''_Int_Int_Int1_1es_3_6_1es_4_6_1sc_0_18_1Lcall_map''_map''_Int_Int_Int0_bufchan_buf ;
  assign \lizzieLet39_4Lcall_map''_map''_Int_Int_Int1_1es_3_6_1es_4_6_1sc_0_18_1Lcall_map''_map''_Int_Int_Int0_bufchan_r  = (! \lizzieLet39_4Lcall_map''_map''_Int_Int_Int1_1es_3_6_1es_4_6_1sc_0_18_1Lcall_map''_map''_Int_Int_Int0_bufchan_buf [0]);
  assign lizzieLet42_1_argbuf_d = (\lizzieLet39_4Lcall_map''_map''_Int_Int_Int1_1es_3_6_1es_4_6_1sc_0_18_1Lcall_map''_map''_Int_Int_Int0_bufchan_buf [0] ? \lizzieLet39_4Lcall_map''_map''_Int_Int_Int1_1es_3_6_1es_4_6_1sc_0_18_1Lcall_map''_map''_Int_Int_Int0_bufchan_buf  :
                                   \lizzieLet39_4Lcall_map''_map''_Int_Int_Int1_1es_3_6_1es_4_6_1sc_0_18_1Lcall_map''_map''_Int_Int_Int0_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet39_4Lcall_map''_map''_Int_Int_Int1_1es_3_6_1es_4_6_1sc_0_18_1Lcall_map''_map''_Int_Int_Int0_bufchan_buf  <= {99'd0,
                                                                                                                             1'd0};
    else
      if ((lizzieLet42_1_argbuf_r && \lizzieLet39_4Lcall_map''_map''_Int_Int_Int1_1es_3_6_1es_4_6_1sc_0_18_1Lcall_map''_map''_Int_Int_Int0_bufchan_buf [0]))
        \lizzieLet39_4Lcall_map''_map''_Int_Int_Int1_1es_3_6_1es_4_6_1sc_0_18_1Lcall_map''_map''_Int_Int_Int0_bufchan_buf  <= {99'd0,
                                                                                                                               1'd0};
      else if (((! lizzieLet42_1_argbuf_r) && (! \lizzieLet39_4Lcall_map''_map''_Int_Int_Int1_1es_3_6_1es_4_6_1sc_0_18_1Lcall_map''_map''_Int_Int_Int0_bufchan_buf [0])))
        \lizzieLet39_4Lcall_map''_map''_Int_Int_Int1_1es_3_6_1es_4_6_1sc_0_18_1Lcall_map''_map''_Int_Int_Int0_bufchan_buf  <= \lizzieLet39_4Lcall_map''_map''_Int_Int_Int1_1es_3_6_1es_4_6_1sc_0_18_1Lcall_map''_map''_Int_Int_Int0_bufchan_d ;
  
  /* dcon (Ty CTmap''_map''_Int_Int_Int,
      Dcon Lcall_map''_map''_Int_Int_Int1) : [(lizzieLet39_4Lcall_map''_map''_Int_Int_Int2,Pointer_QTree_Int),
                                              (es_4_5_destruct,Pointer_QTree_Int),
                                              (sc_0_17_destruct,Pointer_CTmap''_map''_Int_Int_Int),
                                              (isZacT_3_1,MyDTInt_Bool),
                                              (gacU_3_1,MyDTInt_Int_Int),
                                              (v'acV_3_1,Int),
                                              (q1acY_2_destruct,Pointer_QTree_Int)] > (lizzieLet39_4Lcall_map''_map''_Int_Int_Int2_1es_4_5_1sc_0_17_1isZacT_3_1gacU_3_1v'acV_3_1q1acY_2_1Lcall_map''_map''_Int_Int_Int1,CTmap''_map''_Int_Int_Int) */
  assign \lizzieLet39_4Lcall_map''_map''_Int_Int_Int2_1es_4_5_1sc_0_17_1isZacT_3_1gacU_3_1v'acV_3_1q1acY_2_1Lcall_map''_map''_Int_Int_Int1_d  = \Lcall_map''_map''_Int_Int_Int1_dc ((& {\lizzieLet39_4Lcall_map''_map''_Int_Int_Int2_d [0],
                                                                                                                                                                                        es_4_5_destruct_d[0],
                                                                                                                                                                                        sc_0_17_destruct_d[0],
                                                                                                                                                                                        isZacT_3_1_d[0],
                                                                                                                                                                                        gacU_3_1_d[0],
                                                                                                                                                                                        \v'acV_3_1_d [0],
                                                                                                                                                                                        q1acY_2_destruct_d[0]}), \lizzieLet39_4Lcall_map''_map''_Int_Int_Int2_d , es_4_5_destruct_d, sc_0_17_destruct_d, isZacT_3_1_d, gacU_3_1_d, \v'acV_3_1_d , q1acY_2_destruct_d);
  assign {\lizzieLet39_4Lcall_map''_map''_Int_Int_Int2_r ,
          es_4_5_destruct_r,
          sc_0_17_destruct_r,
          isZacT_3_1_r,
          gacU_3_1_r,
          \v'acV_3_1_r ,
          q1acY_2_destruct_r} = {7 {(\lizzieLet39_4Lcall_map''_map''_Int_Int_Int2_1es_4_5_1sc_0_17_1isZacT_3_1gacU_3_1v'acV_3_1q1acY_2_1Lcall_map''_map''_Int_Int_Int1_r  && \lizzieLet39_4Lcall_map''_map''_Int_Int_Int2_1es_4_5_1sc_0_17_1isZacT_3_1gacU_3_1v'acV_3_1q1acY_2_1Lcall_map''_map''_Int_Int_Int1_d [0])}};
  
  /* buf (Ty CTmap''_map''_Int_Int_Int) : (lizzieLet39_4Lcall_map''_map''_Int_Int_Int2_1es_4_5_1sc_0_17_1isZacT_3_1gacU_3_1v'acV_3_1q1acY_2_1Lcall_map''_map''_Int_Int_Int1,CTmap''_map''_Int_Int_Int) > (lizzieLet41_1_argbuf,CTmap''_map''_Int_Int_Int) */
  \CTmap''_map''_Int_Int_Int_t  \lizzieLet39_4Lcall_map''_map''_Int_Int_Int2_1es_4_5_1sc_0_17_1isZacT_3_1gacU_3_1v'acV_3_1q1acY_2_1Lcall_map''_map''_Int_Int_Int1_bufchan_d ;
  logic \lizzieLet39_4Lcall_map''_map''_Int_Int_Int2_1es_4_5_1sc_0_17_1isZacT_3_1gacU_3_1v'acV_3_1q1acY_2_1Lcall_map''_map''_Int_Int_Int1_bufchan_r ;
  assign \lizzieLet39_4Lcall_map''_map''_Int_Int_Int2_1es_4_5_1sc_0_17_1isZacT_3_1gacU_3_1v'acV_3_1q1acY_2_1Lcall_map''_map''_Int_Int_Int1_r  = ((! \lizzieLet39_4Lcall_map''_map''_Int_Int_Int2_1es_4_5_1sc_0_17_1isZacT_3_1gacU_3_1v'acV_3_1q1acY_2_1Lcall_map''_map''_Int_Int_Int1_bufchan_d [0]) || \lizzieLet39_4Lcall_map''_map''_Int_Int_Int2_1es_4_5_1sc_0_17_1isZacT_3_1gacU_3_1v'acV_3_1q1acY_2_1Lcall_map''_map''_Int_Int_Int1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet39_4Lcall_map''_map''_Int_Int_Int2_1es_4_5_1sc_0_17_1isZacT_3_1gacU_3_1v'acV_3_1q1acY_2_1Lcall_map''_map''_Int_Int_Int1_bufchan_d  <= {99'd0,
                                                                                                                                                       1'd0};
    else
      if (\lizzieLet39_4Lcall_map''_map''_Int_Int_Int2_1es_4_5_1sc_0_17_1isZacT_3_1gacU_3_1v'acV_3_1q1acY_2_1Lcall_map''_map''_Int_Int_Int1_r )
        \lizzieLet39_4Lcall_map''_map''_Int_Int_Int2_1es_4_5_1sc_0_17_1isZacT_3_1gacU_3_1v'acV_3_1q1acY_2_1Lcall_map''_map''_Int_Int_Int1_bufchan_d  <= \lizzieLet39_4Lcall_map''_map''_Int_Int_Int2_1es_4_5_1sc_0_17_1isZacT_3_1gacU_3_1v'acV_3_1q1acY_2_1Lcall_map''_map''_Int_Int_Int1_d ;
  \CTmap''_map''_Int_Int_Int_t  \lizzieLet39_4Lcall_map''_map''_Int_Int_Int2_1es_4_5_1sc_0_17_1isZacT_3_1gacU_3_1v'acV_3_1q1acY_2_1Lcall_map''_map''_Int_Int_Int1_bufchan_buf ;
  assign \lizzieLet39_4Lcall_map''_map''_Int_Int_Int2_1es_4_5_1sc_0_17_1isZacT_3_1gacU_3_1v'acV_3_1q1acY_2_1Lcall_map''_map''_Int_Int_Int1_bufchan_r  = (! \lizzieLet39_4Lcall_map''_map''_Int_Int_Int2_1es_4_5_1sc_0_17_1isZacT_3_1gacU_3_1v'acV_3_1q1acY_2_1Lcall_map''_map''_Int_Int_Int1_bufchan_buf [0]);
  assign lizzieLet41_1_argbuf_d = (\lizzieLet39_4Lcall_map''_map''_Int_Int_Int2_1es_4_5_1sc_0_17_1isZacT_3_1gacU_3_1v'acV_3_1q1acY_2_1Lcall_map''_map''_Int_Int_Int1_bufchan_buf [0] ? \lizzieLet39_4Lcall_map''_map''_Int_Int_Int2_1es_4_5_1sc_0_17_1isZacT_3_1gacU_3_1v'acV_3_1q1acY_2_1Lcall_map''_map''_Int_Int_Int1_bufchan_buf  :
                                   \lizzieLet39_4Lcall_map''_map''_Int_Int_Int2_1es_4_5_1sc_0_17_1isZacT_3_1gacU_3_1v'acV_3_1q1acY_2_1Lcall_map''_map''_Int_Int_Int1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet39_4Lcall_map''_map''_Int_Int_Int2_1es_4_5_1sc_0_17_1isZacT_3_1gacU_3_1v'acV_3_1q1acY_2_1Lcall_map''_map''_Int_Int_Int1_bufchan_buf  <= {99'd0,
                                                                                                                                                         1'd0};
    else
      if ((lizzieLet41_1_argbuf_r && \lizzieLet39_4Lcall_map''_map''_Int_Int_Int2_1es_4_5_1sc_0_17_1isZacT_3_1gacU_3_1v'acV_3_1q1acY_2_1Lcall_map''_map''_Int_Int_Int1_bufchan_buf [0]))
        \lizzieLet39_4Lcall_map''_map''_Int_Int_Int2_1es_4_5_1sc_0_17_1isZacT_3_1gacU_3_1v'acV_3_1q1acY_2_1Lcall_map''_map''_Int_Int_Int1_bufchan_buf  <= {99'd0,
                                                                                                                                                           1'd0};
      else if (((! lizzieLet41_1_argbuf_r) && (! \lizzieLet39_4Lcall_map''_map''_Int_Int_Int2_1es_4_5_1sc_0_17_1isZacT_3_1gacU_3_1v'acV_3_1q1acY_2_1Lcall_map''_map''_Int_Int_Int1_bufchan_buf [0])))
        \lizzieLet39_4Lcall_map''_map''_Int_Int_Int2_1es_4_5_1sc_0_17_1isZacT_3_1gacU_3_1v'acV_3_1q1acY_2_1Lcall_map''_map''_Int_Int_Int1_bufchan_buf  <= \lizzieLet39_4Lcall_map''_map''_Int_Int_Int2_1es_4_5_1sc_0_17_1isZacT_3_1gacU_3_1v'acV_3_1q1acY_2_1Lcall_map''_map''_Int_Int_Int1_bufchan_d ;
  
  /* dcon (Ty CTmap''_map''_Int_Int_Int,
      Dcon Lcall_map''_map''_Int_Int_Int2) : [(lizzieLet39_4Lcall_map''_map''_Int_Int_Int3,Pointer_QTree_Int),
                                              (sc_0_16_destruct,Pointer_CTmap''_map''_Int_Int_Int),
                                              (isZacT_2_1,MyDTInt_Bool),
                                              (gacU_2_1,MyDTInt_Int_Int),
                                              (v'acV_2_1,Int),
                                              (q1acY_1_destruct,Pointer_QTree_Int),
                                              (q2acZ_1_destruct,Pointer_QTree_Int)] > (lizzieLet39_4Lcall_map''_map''_Int_Int_Int3_1sc_0_16_1isZacT_2_1gacU_2_1v'acV_2_1q1acY_1_1q2acZ_1_1Lcall_map''_map''_Int_Int_Int2,CTmap''_map''_Int_Int_Int) */
  assign \lizzieLet39_4Lcall_map''_map''_Int_Int_Int3_1sc_0_16_1isZacT_2_1gacU_2_1v'acV_2_1q1acY_1_1q2acZ_1_1Lcall_map''_map''_Int_Int_Int2_d  = \Lcall_map''_map''_Int_Int_Int2_dc ((& {\lizzieLet39_4Lcall_map''_map''_Int_Int_Int3_d [0],
                                                                                                                                                                                         sc_0_16_destruct_d[0],
                                                                                                                                                                                         isZacT_2_1_d[0],
                                                                                                                                                                                         gacU_2_1_d[0],
                                                                                                                                                                                         \v'acV_2_1_d [0],
                                                                                                                                                                                         q1acY_1_destruct_d[0],
                                                                                                                                                                                         q2acZ_1_destruct_d[0]}), \lizzieLet39_4Lcall_map''_map''_Int_Int_Int3_d , sc_0_16_destruct_d, isZacT_2_1_d, gacU_2_1_d, \v'acV_2_1_d , q1acY_1_destruct_d, q2acZ_1_destruct_d);
  assign {\lizzieLet39_4Lcall_map''_map''_Int_Int_Int3_r ,
          sc_0_16_destruct_r,
          isZacT_2_1_r,
          gacU_2_1_r,
          \v'acV_2_1_r ,
          q1acY_1_destruct_r,
          q2acZ_1_destruct_r} = {7 {(\lizzieLet39_4Lcall_map''_map''_Int_Int_Int3_1sc_0_16_1isZacT_2_1gacU_2_1v'acV_2_1q1acY_1_1q2acZ_1_1Lcall_map''_map''_Int_Int_Int2_r  && \lizzieLet39_4Lcall_map''_map''_Int_Int_Int3_1sc_0_16_1isZacT_2_1gacU_2_1v'acV_2_1q1acY_1_1q2acZ_1_1Lcall_map''_map''_Int_Int_Int2_d [0])}};
  
  /* buf (Ty CTmap''_map''_Int_Int_Int) : (lizzieLet39_4Lcall_map''_map''_Int_Int_Int3_1sc_0_16_1isZacT_2_1gacU_2_1v'acV_2_1q1acY_1_1q2acZ_1_1Lcall_map''_map''_Int_Int_Int2,CTmap''_map''_Int_Int_Int) > (lizzieLet40_1_argbuf,CTmap''_map''_Int_Int_Int) */
  \CTmap''_map''_Int_Int_Int_t  \lizzieLet39_4Lcall_map''_map''_Int_Int_Int3_1sc_0_16_1isZacT_2_1gacU_2_1v'acV_2_1q1acY_1_1q2acZ_1_1Lcall_map''_map''_Int_Int_Int2_bufchan_d ;
  logic \lizzieLet39_4Lcall_map''_map''_Int_Int_Int3_1sc_0_16_1isZacT_2_1gacU_2_1v'acV_2_1q1acY_1_1q2acZ_1_1Lcall_map''_map''_Int_Int_Int2_bufchan_r ;
  assign \lizzieLet39_4Lcall_map''_map''_Int_Int_Int3_1sc_0_16_1isZacT_2_1gacU_2_1v'acV_2_1q1acY_1_1q2acZ_1_1Lcall_map''_map''_Int_Int_Int2_r  = ((! \lizzieLet39_4Lcall_map''_map''_Int_Int_Int3_1sc_0_16_1isZacT_2_1gacU_2_1v'acV_2_1q1acY_1_1q2acZ_1_1Lcall_map''_map''_Int_Int_Int2_bufchan_d [0]) || \lizzieLet39_4Lcall_map''_map''_Int_Int_Int3_1sc_0_16_1isZacT_2_1gacU_2_1v'acV_2_1q1acY_1_1q2acZ_1_1Lcall_map''_map''_Int_Int_Int2_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet39_4Lcall_map''_map''_Int_Int_Int3_1sc_0_16_1isZacT_2_1gacU_2_1v'acV_2_1q1acY_1_1q2acZ_1_1Lcall_map''_map''_Int_Int_Int2_bufchan_d  <= {99'd0,
                                                                                                                                                        1'd0};
    else
      if (\lizzieLet39_4Lcall_map''_map''_Int_Int_Int3_1sc_0_16_1isZacT_2_1gacU_2_1v'acV_2_1q1acY_1_1q2acZ_1_1Lcall_map''_map''_Int_Int_Int2_r )
        \lizzieLet39_4Lcall_map''_map''_Int_Int_Int3_1sc_0_16_1isZacT_2_1gacU_2_1v'acV_2_1q1acY_1_1q2acZ_1_1Lcall_map''_map''_Int_Int_Int2_bufchan_d  <= \lizzieLet39_4Lcall_map''_map''_Int_Int_Int3_1sc_0_16_1isZacT_2_1gacU_2_1v'acV_2_1q1acY_1_1q2acZ_1_1Lcall_map''_map''_Int_Int_Int2_d ;
  \CTmap''_map''_Int_Int_Int_t  \lizzieLet39_4Lcall_map''_map''_Int_Int_Int3_1sc_0_16_1isZacT_2_1gacU_2_1v'acV_2_1q1acY_1_1q2acZ_1_1Lcall_map''_map''_Int_Int_Int2_bufchan_buf ;
  assign \lizzieLet39_4Lcall_map''_map''_Int_Int_Int3_1sc_0_16_1isZacT_2_1gacU_2_1v'acV_2_1q1acY_1_1q2acZ_1_1Lcall_map''_map''_Int_Int_Int2_bufchan_r  = (! \lizzieLet39_4Lcall_map''_map''_Int_Int_Int3_1sc_0_16_1isZacT_2_1gacU_2_1v'acV_2_1q1acY_1_1q2acZ_1_1Lcall_map''_map''_Int_Int_Int2_bufchan_buf [0]);
  assign lizzieLet40_1_argbuf_d = (\lizzieLet39_4Lcall_map''_map''_Int_Int_Int3_1sc_0_16_1isZacT_2_1gacU_2_1v'acV_2_1q1acY_1_1q2acZ_1_1Lcall_map''_map''_Int_Int_Int2_bufchan_buf [0] ? \lizzieLet39_4Lcall_map''_map''_Int_Int_Int3_1sc_0_16_1isZacT_2_1gacU_2_1v'acV_2_1q1acY_1_1q2acZ_1_1Lcall_map''_map''_Int_Int_Int2_bufchan_buf  :
                                   \lizzieLet39_4Lcall_map''_map''_Int_Int_Int3_1sc_0_16_1isZacT_2_1gacU_2_1v'acV_2_1q1acY_1_1q2acZ_1_1Lcall_map''_map''_Int_Int_Int2_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet39_4Lcall_map''_map''_Int_Int_Int3_1sc_0_16_1isZacT_2_1gacU_2_1v'acV_2_1q1acY_1_1q2acZ_1_1Lcall_map''_map''_Int_Int_Int2_bufchan_buf  <= {99'd0,
                                                                                                                                                          1'd0};
    else
      if ((lizzieLet40_1_argbuf_r && \lizzieLet39_4Lcall_map''_map''_Int_Int_Int3_1sc_0_16_1isZacT_2_1gacU_2_1v'acV_2_1q1acY_1_1q2acZ_1_1Lcall_map''_map''_Int_Int_Int2_bufchan_buf [0]))
        \lizzieLet39_4Lcall_map''_map''_Int_Int_Int3_1sc_0_16_1isZacT_2_1gacU_2_1v'acV_2_1q1acY_1_1q2acZ_1_1Lcall_map''_map''_Int_Int_Int2_bufchan_buf  <= {99'd0,
                                                                                                                                                            1'd0};
      else if (((! lizzieLet40_1_argbuf_r) && (! \lizzieLet39_4Lcall_map''_map''_Int_Int_Int3_1sc_0_16_1isZacT_2_1gacU_2_1v'acV_2_1q1acY_1_1q2acZ_1_1Lcall_map''_map''_Int_Int_Int2_bufchan_buf [0])))
        \lizzieLet39_4Lcall_map''_map''_Int_Int_Int3_1sc_0_16_1isZacT_2_1gacU_2_1v'acV_2_1q1acY_1_1q2acZ_1_1Lcall_map''_map''_Int_Int_Int2_bufchan_buf  <= \lizzieLet39_4Lcall_map''_map''_Int_Int_Int3_1sc_0_16_1isZacT_2_1gacU_2_1v'acV_2_1q1acY_1_1q2acZ_1_1Lcall_map''_map''_Int_Int_Int2_bufchan_d ;
  
  /* fork (Ty Pointer_QTree_Int) : (lizzieLet39_4Lmap''_map''_Int_Int_Intsbos,Pointer_QTree_Int) > [(lizzieLet39_4Lmap''_map''_Int_Int_Intsbos_1_merge_merge_fork_1,Pointer_QTree_Int),
                                                                                               (lizzieLet39_4Lmap''_map''_Int_Int_Intsbos_1_merge_merge_fork_2,Pointer_QTree_Int)] */
  logic [1:0] \lizzieLet39_4Lmap''_map''_Int_Int_Intsbos_emitted ;
  logic [1:0] \lizzieLet39_4Lmap''_map''_Int_Int_Intsbos_done ;
  assign \lizzieLet39_4Lmap''_map''_Int_Int_Intsbos_1_merge_merge_fork_1_d  = {\lizzieLet39_4Lmap''_map''_Int_Int_Intsbos_d [16:1],
                                                                               (\lizzieLet39_4Lmap''_map''_Int_Int_Intsbos_d [0] && (! \lizzieLet39_4Lmap''_map''_Int_Int_Intsbos_emitted [0]))};
  assign \lizzieLet39_4Lmap''_map''_Int_Int_Intsbos_1_merge_merge_fork_2_d  = {\lizzieLet39_4Lmap''_map''_Int_Int_Intsbos_d [16:1],
                                                                               (\lizzieLet39_4Lmap''_map''_Int_Int_Intsbos_d [0] && (! \lizzieLet39_4Lmap''_map''_Int_Int_Intsbos_emitted [1]))};
  assign \lizzieLet39_4Lmap''_map''_Int_Int_Intsbos_done  = (\lizzieLet39_4Lmap''_map''_Int_Int_Intsbos_emitted  | ({\lizzieLet39_4Lmap''_map''_Int_Int_Intsbos_1_merge_merge_fork_2_d [0],
                                                                                                                     \lizzieLet39_4Lmap''_map''_Int_Int_Intsbos_1_merge_merge_fork_1_d [0]} & {\lizzieLet39_4Lmap''_map''_Int_Int_Intsbos_1_merge_merge_fork_2_r ,
                                                                                                                                                                                               \lizzieLet39_4Lmap''_map''_Int_Int_Intsbos_1_merge_merge_fork_1_r }));
  assign \lizzieLet39_4Lmap''_map''_Int_Int_Intsbos_r  = (& \lizzieLet39_4Lmap''_map''_Int_Int_Intsbos_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet39_4Lmap''_map''_Int_Int_Intsbos_emitted  <= 2'd0;
    else
      \lizzieLet39_4Lmap''_map''_Int_Int_Intsbos_emitted  <= (\lizzieLet39_4Lmap''_map''_Int_Int_Intsbos_r  ? 2'd0 :
                                                              \lizzieLet39_4Lmap''_map''_Int_Int_Intsbos_done );
  
  /* togo (Ty Pointer_QTree_Int) : (lizzieLet39_4Lmap''_map''_Int_Int_Intsbos_1_merge_merge_fork_1,Pointer_QTree_Int) > (call_map''_map''_Int_Int_Int_goConst,Go) */
  assign \call_map''_map''_Int_Int_Int_goConst_d  = \lizzieLet39_4Lmap''_map''_Int_Int_Intsbos_1_merge_merge_fork_1_d [0];
  assign \lizzieLet39_4Lmap''_map''_Int_Int_Intsbos_1_merge_merge_fork_1_r  = \call_map''_map''_Int_Int_Int_goConst_r ;
  
  /* buf (Ty Pointer_QTree_Int) : (lizzieLet39_4Lmap''_map''_Int_Int_Intsbos_1_merge_merge_fork_2,Pointer_QTree_Int) > (map''_map''_Int_Int_Int_resbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t \lizzieLet39_4Lmap''_map''_Int_Int_Intsbos_1_merge_merge_fork_2_bufchan_d ;
  logic \lizzieLet39_4Lmap''_map''_Int_Int_Intsbos_1_merge_merge_fork_2_bufchan_r ;
  assign \lizzieLet39_4Lmap''_map''_Int_Int_Intsbos_1_merge_merge_fork_2_r  = ((! \lizzieLet39_4Lmap''_map''_Int_Int_Intsbos_1_merge_merge_fork_2_bufchan_d [0]) || \lizzieLet39_4Lmap''_map''_Int_Int_Intsbos_1_merge_merge_fork_2_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet39_4Lmap''_map''_Int_Int_Intsbos_1_merge_merge_fork_2_bufchan_d  <= {16'd0,
                                                                                     1'd0};
    else
      if (\lizzieLet39_4Lmap''_map''_Int_Int_Intsbos_1_merge_merge_fork_2_r )
        \lizzieLet39_4Lmap''_map''_Int_Int_Intsbos_1_merge_merge_fork_2_bufchan_d  <= \lizzieLet39_4Lmap''_map''_Int_Int_Intsbos_1_merge_merge_fork_2_d ;
  Pointer_QTree_Int_t \lizzieLet39_4Lmap''_map''_Int_Int_Intsbos_1_merge_merge_fork_2_bufchan_buf ;
  assign \lizzieLet39_4Lmap''_map''_Int_Int_Intsbos_1_merge_merge_fork_2_bufchan_r  = (! \lizzieLet39_4Lmap''_map''_Int_Int_Intsbos_1_merge_merge_fork_2_bufchan_buf [0]);
  assign \map''_map''_Int_Int_Int_resbuf_d  = (\lizzieLet39_4Lmap''_map''_Int_Int_Intsbos_1_merge_merge_fork_2_bufchan_buf [0] ? \lizzieLet39_4Lmap''_map''_Int_Int_Intsbos_1_merge_merge_fork_2_bufchan_buf  :
                                               \lizzieLet39_4Lmap''_map''_Int_Int_Intsbos_1_merge_merge_fork_2_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet39_4Lmap''_map''_Int_Int_Intsbos_1_merge_merge_fork_2_bufchan_buf  <= {16'd0,
                                                                                       1'd0};
    else
      if ((\map''_map''_Int_Int_Int_resbuf_r  && \lizzieLet39_4Lmap''_map''_Int_Int_Intsbos_1_merge_merge_fork_2_bufchan_buf [0]))
        \lizzieLet39_4Lmap''_map''_Int_Int_Intsbos_1_merge_merge_fork_2_bufchan_buf  <= {16'd0,
                                                                                         1'd0};
      else if (((! \map''_map''_Int_Int_Int_resbuf_r ) && (! \lizzieLet39_4Lmap''_map''_Int_Int_Intsbos_1_merge_merge_fork_2_bufchan_buf [0])))
        \lizzieLet39_4Lmap''_map''_Int_Int_Intsbos_1_merge_merge_fork_2_bufchan_buf  <= \lizzieLet39_4Lmap''_map''_Int_Int_Intsbos_1_merge_merge_fork_2_bufchan_d ;
  
  /* demux (Ty MyBool,
       Ty Go) : (lizzieLet3_1,MyBool) (arg0_1Dcon_eqZero_3I#_3,Go) > [(lizzieLet3_1MyFalse,Go),
                                                                      (lizzieLet3_1MyTrue,Go)] */
  logic [1:0] \arg0_1Dcon_eqZero_3I#_3_onehotd ;
  always_comb
    if ((lizzieLet3_1_d[0] && \arg0_1Dcon_eqZero_3I#_3_d [0]))
      unique case (lizzieLet3_1_d[1:1])
        1'd0: \arg0_1Dcon_eqZero_3I#_3_onehotd  = 2'd1;
        1'd1: \arg0_1Dcon_eqZero_3I#_3_onehotd  = 2'd2;
        default: \arg0_1Dcon_eqZero_3I#_3_onehotd  = 2'd0;
      endcase
    else \arg0_1Dcon_eqZero_3I#_3_onehotd  = 2'd0;
  assign lizzieLet3_1MyFalse_d = \arg0_1Dcon_eqZero_3I#_3_onehotd [0];
  assign lizzieLet3_1MyTrue_d = \arg0_1Dcon_eqZero_3I#_3_onehotd [1];
  assign \arg0_1Dcon_eqZero_3I#_3_r  = (| (\arg0_1Dcon_eqZero_3I#_3_onehotd  & {lizzieLet3_1MyTrue_r,
                                                                                lizzieLet3_1MyFalse_r}));
  assign lizzieLet3_1_r = \arg0_1Dcon_eqZero_3I#_3_r ;
  
  /* dcon (Ty MyBool,
      Dcon MyFalse) : [(lizzieLet3_1MyFalse,Go)] > (lizzieLet3_1MyFalse_1MyFalse,MyBool) */
  assign lizzieLet3_1MyFalse_1MyFalse_d = MyFalse_dc((& {lizzieLet3_1MyFalse_d[0]}), lizzieLet3_1MyFalse_d);
  assign {lizzieLet3_1MyFalse_r} = {1 {(lizzieLet3_1MyFalse_1MyFalse_r && lizzieLet3_1MyFalse_1MyFalse_d[0])}};
  
  /* dcon (Ty MyBool,
      Dcon MyTrue) : [(lizzieLet3_1MyTrue,Go)] > (lizzieLet3_1MyTrue_1MyTrue,MyBool) */
  assign lizzieLet3_1MyTrue_1MyTrue_d = MyTrue_dc((& {lizzieLet3_1MyTrue_d[0]}), lizzieLet3_1MyTrue_d);
  assign {lizzieLet3_1MyTrue_r} = {1 {(lizzieLet3_1MyTrue_1MyTrue_r && lizzieLet3_1MyTrue_1MyTrue_d[0])}};
  
  /* mux (Ty MyBool,
     Ty MyBool) : (lizzieLet3_2,MyBool) [(lizzieLet3_1MyFalse_1MyFalse,MyBool),
                                         (lizzieLet3_1MyTrue_1MyTrue,MyBool)] > (lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux,MyBool) */
  logic [1:0] lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux;
  logic [1:0] lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_onehot;
  always_comb
    unique case (lizzieLet3_2_d[1:1])
      1'd0:
        {lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_onehot,
         lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux} = {2'd1,
                                                                            lizzieLet3_1MyFalse_1MyFalse_d};
      1'd1:
        {lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_onehot,
         lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux} = {2'd2,
                                                                            lizzieLet3_1MyTrue_1MyTrue_d};
      default:
        {lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_onehot,
         lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux} = {2'd0,
                                                                            {1'd0, 1'd0}};
    endcase
  assign lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_d = {lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux[1:1],
                                                                         (lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux[0] && lizzieLet3_2_d[0])};
  assign lizzieLet3_2_r = (lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_d[0] && lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_r);
  assign {lizzieLet3_1MyTrue_1MyTrue_r,
          lizzieLet3_1MyFalse_1MyFalse_r} = (lizzieLet3_2_r ? lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_onehot :
                                             2'd0);
  
  /* destruct (Ty QTree_Int,
          Dcon QNode_Int) : (lizzieLet4_1QNode_Int,QTree_Int) > [(q1ac0_destruct,Pointer_QTree_Int),
                                                                 (q2ac1_destruct,Pointer_QTree_Int),
                                                                 (q3ac2_destruct,Pointer_QTree_Int),
                                                                 (q4ac3_destruct,Pointer_QTree_Int)] */
  logic [3:0] lizzieLet4_1QNode_Int_emitted;
  logic [3:0] lizzieLet4_1QNode_Int_done;
  assign q1ac0_destruct_d = {lizzieLet4_1QNode_Int_d[18:3],
                             (lizzieLet4_1QNode_Int_d[0] && (! lizzieLet4_1QNode_Int_emitted[0]))};
  assign q2ac1_destruct_d = {lizzieLet4_1QNode_Int_d[34:19],
                             (lizzieLet4_1QNode_Int_d[0] && (! lizzieLet4_1QNode_Int_emitted[1]))};
  assign q3ac2_destruct_d = {lizzieLet4_1QNode_Int_d[50:35],
                             (lizzieLet4_1QNode_Int_d[0] && (! lizzieLet4_1QNode_Int_emitted[2]))};
  assign q4ac3_destruct_d = {lizzieLet4_1QNode_Int_d[66:51],
                             (lizzieLet4_1QNode_Int_d[0] && (! lizzieLet4_1QNode_Int_emitted[3]))};
  assign lizzieLet4_1QNode_Int_done = (lizzieLet4_1QNode_Int_emitted | ({q4ac3_destruct_d[0],
                                                                         q3ac2_destruct_d[0],
                                                                         q2ac1_destruct_d[0],
                                                                         q1ac0_destruct_d[0]} & {q4ac3_destruct_r,
                                                                                                 q3ac2_destruct_r,
                                                                                                 q2ac1_destruct_r,
                                                                                                 q1ac0_destruct_r}));
  assign lizzieLet4_1QNode_Int_r = (& lizzieLet4_1QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_1QNode_Int_emitted <= 4'd0;
    else
      lizzieLet4_1QNode_Int_emitted <= (lizzieLet4_1QNode_Int_r ? 4'd0 :
                                        lizzieLet4_1QNode_Int_done);
  
  /* demux (Ty QTree_Int,
       Ty QTree_Int) : (lizzieLet4_2,QTree_Int) (lizzieLet4_1,QTree_Int) > [(_10,QTree_Int),
                                                                            (_9,QTree_Int),
                                                                            (lizzieLet4_1QNode_Int,QTree_Int),
                                                                            (_8,QTree_Int)] */
  logic [3:0] lizzieLet4_1_onehotd;
  always_comb
    if ((lizzieLet4_2_d[0] && lizzieLet4_1_d[0]))
      unique case (lizzieLet4_2_d[2:1])
        2'd0: lizzieLet4_1_onehotd = 4'd1;
        2'd1: lizzieLet4_1_onehotd = 4'd2;
        2'd2: lizzieLet4_1_onehotd = 4'd4;
        2'd3: lizzieLet4_1_onehotd = 4'd8;
        default: lizzieLet4_1_onehotd = 4'd0;
      endcase
    else lizzieLet4_1_onehotd = 4'd0;
  assign _10_d = {lizzieLet4_1_d[66:1], lizzieLet4_1_onehotd[0]};
  assign _9_d = {lizzieLet4_1_d[66:1], lizzieLet4_1_onehotd[1]};
  assign lizzieLet4_1QNode_Int_d = {lizzieLet4_1_d[66:1],
                                    lizzieLet4_1_onehotd[2]};
  assign _8_d = {lizzieLet4_1_d[66:1], lizzieLet4_1_onehotd[3]};
  assign lizzieLet4_1_r = (| (lizzieLet4_1_onehotd & {_8_r,
                                                      lizzieLet4_1QNode_Int_r,
                                                      _9_r,
                                                      _10_r}));
  assign lizzieLet4_2_r = lizzieLet4_1_r;
  
  /* demux (Ty QTree_Int,
       Ty Go) : (lizzieLet4_3,QTree_Int) (go_11_goMux_data,Go) > [(lizzieLet4_3QNone_Int,Go),
                                                                  (lizzieLet4_3QVal_Int,Go),
                                                                  (lizzieLet4_3QNode_Int,Go),
                                                                  (lizzieLet4_3QError_Int,Go)] */
  logic [3:0] go_11_goMux_data_onehotd;
  always_comb
    if ((lizzieLet4_3_d[0] && go_11_goMux_data_d[0]))
      unique case (lizzieLet4_3_d[2:1])
        2'd0: go_11_goMux_data_onehotd = 4'd1;
        2'd1: go_11_goMux_data_onehotd = 4'd2;
        2'd2: go_11_goMux_data_onehotd = 4'd4;
        2'd3: go_11_goMux_data_onehotd = 4'd8;
        default: go_11_goMux_data_onehotd = 4'd0;
      endcase
    else go_11_goMux_data_onehotd = 4'd0;
  assign lizzieLet4_3QNone_Int_d = go_11_goMux_data_onehotd[0];
  assign lizzieLet4_3QVal_Int_d = go_11_goMux_data_onehotd[1];
  assign lizzieLet4_3QNode_Int_d = go_11_goMux_data_onehotd[2];
  assign lizzieLet4_3QError_Int_d = go_11_goMux_data_onehotd[3];
  assign go_11_goMux_data_r = (| (go_11_goMux_data_onehotd & {lizzieLet4_3QError_Int_r,
                                                              lizzieLet4_3QNode_Int_r,
                                                              lizzieLet4_3QVal_Int_r,
                                                              lizzieLet4_3QNone_Int_r}));
  assign lizzieLet4_3_r = go_11_goMux_data_r;
  
  /* fork (Ty Go) : (lizzieLet4_3QError_Int,Go) > [(lizzieLet4_3QError_Int_1,Go),
                                              (lizzieLet4_3QError_Int_2,Go)] */
  logic [1:0] lizzieLet4_3QError_Int_emitted;
  logic [1:0] lizzieLet4_3QError_Int_done;
  assign lizzieLet4_3QError_Int_1_d = (lizzieLet4_3QError_Int_d[0] && (! lizzieLet4_3QError_Int_emitted[0]));
  assign lizzieLet4_3QError_Int_2_d = (lizzieLet4_3QError_Int_d[0] && (! lizzieLet4_3QError_Int_emitted[1]));
  assign lizzieLet4_3QError_Int_done = (lizzieLet4_3QError_Int_emitted | ({lizzieLet4_3QError_Int_2_d[0],
                                                                           lizzieLet4_3QError_Int_1_d[0]} & {lizzieLet4_3QError_Int_2_r,
                                                                                                             lizzieLet4_3QError_Int_1_r}));
  assign lizzieLet4_3QError_Int_r = (& lizzieLet4_3QError_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3QError_Int_emitted <= 2'd0;
    else
      lizzieLet4_3QError_Int_emitted <= (lizzieLet4_3QError_Int_r ? 2'd0 :
                                         lizzieLet4_3QError_Int_done);
  
  /* buf (Ty Go) : (lizzieLet4_3QError_Int_1,Go) > (lizzieLet4_3QError_Int_1_argbuf,Go) */
  Go_t lizzieLet4_3QError_Int_1_bufchan_d;
  logic lizzieLet4_3QError_Int_1_bufchan_r;
  assign lizzieLet4_3QError_Int_1_r = ((! lizzieLet4_3QError_Int_1_bufchan_d[0]) || lizzieLet4_3QError_Int_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3QError_Int_1_bufchan_d <= 1'd0;
    else
      if (lizzieLet4_3QError_Int_1_r)
        lizzieLet4_3QError_Int_1_bufchan_d <= lizzieLet4_3QError_Int_1_d;
  Go_t lizzieLet4_3QError_Int_1_bufchan_buf;
  assign lizzieLet4_3QError_Int_1_bufchan_r = (! lizzieLet4_3QError_Int_1_bufchan_buf[0]);
  assign lizzieLet4_3QError_Int_1_argbuf_d = (lizzieLet4_3QError_Int_1_bufchan_buf[0] ? lizzieLet4_3QError_Int_1_bufchan_buf :
                                              lizzieLet4_3QError_Int_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3QError_Int_1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet4_3QError_Int_1_argbuf_r && lizzieLet4_3QError_Int_1_bufchan_buf[0]))
        lizzieLet4_3QError_Int_1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet4_3QError_Int_1_argbuf_r) && (! lizzieLet4_3QError_Int_1_bufchan_buf[0])))
        lizzieLet4_3QError_Int_1_bufchan_buf <= lizzieLet4_3QError_Int_1_bufchan_d;
  
  /* const (Ty Int#,
       Lit 0) : (lizzieLet4_3QError_Int_1_argbuf,Go) > (lizzieLet4_3QError_Int_1_argbuf_0,Int#) */
  assign lizzieLet4_3QError_Int_1_argbuf_0_d = {32'd0,
                                                lizzieLet4_3QError_Int_1_argbuf_d[0]};
  assign lizzieLet4_3QError_Int_1_argbuf_r = lizzieLet4_3QError_Int_1_argbuf_0_r;
  
  /* buf (Ty Int#) : (lizzieLet4_3QError_Int_1_argbuf_0,Int#) > (lizzieLet15_1_1_argbuf,Int#) */
  \Int#_t  lizzieLet4_3QError_Int_1_argbuf_0_bufchan_d;
  logic lizzieLet4_3QError_Int_1_argbuf_0_bufchan_r;
  assign lizzieLet4_3QError_Int_1_argbuf_0_r = ((! lizzieLet4_3QError_Int_1_argbuf_0_bufchan_d[0]) || lizzieLet4_3QError_Int_1_argbuf_0_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_3QError_Int_1_argbuf_0_bufchan_d <= {32'd0, 1'd0};
    else
      if (lizzieLet4_3QError_Int_1_argbuf_0_r)
        lizzieLet4_3QError_Int_1_argbuf_0_bufchan_d <= lizzieLet4_3QError_Int_1_argbuf_0_d;
  \Int#_t  lizzieLet4_3QError_Int_1_argbuf_0_bufchan_buf;
  assign lizzieLet4_3QError_Int_1_argbuf_0_bufchan_r = (! lizzieLet4_3QError_Int_1_argbuf_0_bufchan_buf[0]);
  assign lizzieLet15_1_1_argbuf_d = (lizzieLet4_3QError_Int_1_argbuf_0_bufchan_buf[0] ? lizzieLet4_3QError_Int_1_argbuf_0_bufchan_buf :
                                     lizzieLet4_3QError_Int_1_argbuf_0_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_3QError_Int_1_argbuf_0_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((lizzieLet15_1_1_argbuf_r && lizzieLet4_3QError_Int_1_argbuf_0_bufchan_buf[0]))
        lizzieLet4_3QError_Int_1_argbuf_0_bufchan_buf <= {32'd0, 1'd0};
      else if (((! lizzieLet15_1_1_argbuf_r) && (! lizzieLet4_3QError_Int_1_argbuf_0_bufchan_buf[0])))
        lizzieLet4_3QError_Int_1_argbuf_0_bufchan_buf <= lizzieLet4_3QError_Int_1_argbuf_0_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet4_3QError_Int_2,Go) > (lizzieLet4_3QError_Int_2_argbuf,Go) */
  Go_t lizzieLet4_3QError_Int_2_bufchan_d;
  logic lizzieLet4_3QError_Int_2_bufchan_r;
  assign lizzieLet4_3QError_Int_2_r = ((! lizzieLet4_3QError_Int_2_bufchan_d[0]) || lizzieLet4_3QError_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3QError_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet4_3QError_Int_2_r)
        lizzieLet4_3QError_Int_2_bufchan_d <= lizzieLet4_3QError_Int_2_d;
  Go_t lizzieLet4_3QError_Int_2_bufchan_buf;
  assign lizzieLet4_3QError_Int_2_bufchan_r = (! lizzieLet4_3QError_Int_2_bufchan_buf[0]);
  assign lizzieLet4_3QError_Int_2_argbuf_d = (lizzieLet4_3QError_Int_2_bufchan_buf[0] ? lizzieLet4_3QError_Int_2_bufchan_buf :
                                              lizzieLet4_3QError_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3QError_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet4_3QError_Int_2_argbuf_r && lizzieLet4_3QError_Int_2_bufchan_buf[0]))
        lizzieLet4_3QError_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet4_3QError_Int_2_argbuf_r) && (! lizzieLet4_3QError_Int_2_bufchan_buf[0])))
        lizzieLet4_3QError_Int_2_bufchan_buf <= lizzieLet4_3QError_Int_2_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet4_3QNode_Int,Go) > (lizzieLet4_3QNode_Int_1_argbuf,Go) */
  Go_t lizzieLet4_3QNode_Int_bufchan_d;
  logic lizzieLet4_3QNode_Int_bufchan_r;
  assign lizzieLet4_3QNode_Int_r = ((! lizzieLet4_3QNode_Int_bufchan_d[0]) || lizzieLet4_3QNode_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3QNode_Int_bufchan_d <= 1'd0;
    else
      if (lizzieLet4_3QNode_Int_r)
        lizzieLet4_3QNode_Int_bufchan_d <= lizzieLet4_3QNode_Int_d;
  Go_t lizzieLet4_3QNode_Int_bufchan_buf;
  assign lizzieLet4_3QNode_Int_bufchan_r = (! lizzieLet4_3QNode_Int_bufchan_buf[0]);
  assign lizzieLet4_3QNode_Int_1_argbuf_d = (lizzieLet4_3QNode_Int_bufchan_buf[0] ? lizzieLet4_3QNode_Int_bufchan_buf :
                                             lizzieLet4_3QNode_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3QNode_Int_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet4_3QNode_Int_1_argbuf_r && lizzieLet4_3QNode_Int_bufchan_buf[0]))
        lizzieLet4_3QNode_Int_bufchan_buf <= 1'd0;
      else if (((! lizzieLet4_3QNode_Int_1_argbuf_r) && (! lizzieLet4_3QNode_Int_bufchan_buf[0])))
        lizzieLet4_3QNode_Int_bufchan_buf <= lizzieLet4_3QNode_Int_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet4_3QNone_Int,Go) > [(lizzieLet4_3QNone_Int_1,Go),
                                             (lizzieLet4_3QNone_Int_2,Go)] */
  logic [1:0] lizzieLet4_3QNone_Int_emitted;
  logic [1:0] lizzieLet4_3QNone_Int_done;
  assign lizzieLet4_3QNone_Int_1_d = (lizzieLet4_3QNone_Int_d[0] && (! lizzieLet4_3QNone_Int_emitted[0]));
  assign lizzieLet4_3QNone_Int_2_d = (lizzieLet4_3QNone_Int_d[0] && (! lizzieLet4_3QNone_Int_emitted[1]));
  assign lizzieLet4_3QNone_Int_done = (lizzieLet4_3QNone_Int_emitted | ({lizzieLet4_3QNone_Int_2_d[0],
                                                                         lizzieLet4_3QNone_Int_1_d[0]} & {lizzieLet4_3QNone_Int_2_r,
                                                                                                          lizzieLet4_3QNone_Int_1_r}));
  assign lizzieLet4_3QNone_Int_r = (& lizzieLet4_3QNone_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3QNone_Int_emitted <= 2'd0;
    else
      lizzieLet4_3QNone_Int_emitted <= (lizzieLet4_3QNone_Int_r ? 2'd0 :
                                        lizzieLet4_3QNone_Int_done);
  
  /* buf (Ty Go) : (lizzieLet4_3QNone_Int_1,Go) > (lizzieLet4_3QNone_Int_1_argbuf,Go) */
  Go_t lizzieLet4_3QNone_Int_1_bufchan_d;
  logic lizzieLet4_3QNone_Int_1_bufchan_r;
  assign lizzieLet4_3QNone_Int_1_r = ((! lizzieLet4_3QNone_Int_1_bufchan_d[0]) || lizzieLet4_3QNone_Int_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3QNone_Int_1_bufchan_d <= 1'd0;
    else
      if (lizzieLet4_3QNone_Int_1_r)
        lizzieLet4_3QNone_Int_1_bufchan_d <= lizzieLet4_3QNone_Int_1_d;
  Go_t lizzieLet4_3QNone_Int_1_bufchan_buf;
  assign lizzieLet4_3QNone_Int_1_bufchan_r = (! lizzieLet4_3QNone_Int_1_bufchan_buf[0]);
  assign lizzieLet4_3QNone_Int_1_argbuf_d = (lizzieLet4_3QNone_Int_1_bufchan_buf[0] ? lizzieLet4_3QNone_Int_1_bufchan_buf :
                                             lizzieLet4_3QNone_Int_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3QNone_Int_1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet4_3QNone_Int_1_argbuf_r && lizzieLet4_3QNone_Int_1_bufchan_buf[0]))
        lizzieLet4_3QNone_Int_1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet4_3QNone_Int_1_argbuf_r) && (! lizzieLet4_3QNone_Int_1_bufchan_buf[0])))
        lizzieLet4_3QNone_Int_1_bufchan_buf <= lizzieLet4_3QNone_Int_1_bufchan_d;
  
  /* const (Ty Int#,
       Lit 0) : (lizzieLet4_3QNone_Int_1_argbuf,Go) > (lizzieLet4_3QNone_Int_1_argbuf_0,Int#) */
  assign lizzieLet4_3QNone_Int_1_argbuf_0_d = {32'd0,
                                               lizzieLet4_3QNone_Int_1_argbuf_d[0]};
  assign lizzieLet4_3QNone_Int_1_argbuf_r = lizzieLet4_3QNone_Int_1_argbuf_0_r;
  
  /* buf (Ty Int#) : (lizzieLet4_3QNone_Int_1_argbuf_0,Int#) > (lizzieLet15_1_argbuf,Int#) */
  \Int#_t  lizzieLet4_3QNone_Int_1_argbuf_0_bufchan_d;
  logic lizzieLet4_3QNone_Int_1_argbuf_0_bufchan_r;
  assign lizzieLet4_3QNone_Int_1_argbuf_0_r = ((! lizzieLet4_3QNone_Int_1_argbuf_0_bufchan_d[0]) || lizzieLet4_3QNone_Int_1_argbuf_0_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_3QNone_Int_1_argbuf_0_bufchan_d <= {32'd0, 1'd0};
    else
      if (lizzieLet4_3QNone_Int_1_argbuf_0_r)
        lizzieLet4_3QNone_Int_1_argbuf_0_bufchan_d <= lizzieLet4_3QNone_Int_1_argbuf_0_d;
  \Int#_t  lizzieLet4_3QNone_Int_1_argbuf_0_bufchan_buf;
  assign lizzieLet4_3QNone_Int_1_argbuf_0_bufchan_r = (! lizzieLet4_3QNone_Int_1_argbuf_0_bufchan_buf[0]);
  assign lizzieLet15_1_argbuf_d = (lizzieLet4_3QNone_Int_1_argbuf_0_bufchan_buf[0] ? lizzieLet4_3QNone_Int_1_argbuf_0_bufchan_buf :
                                   lizzieLet4_3QNone_Int_1_argbuf_0_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_3QNone_Int_1_argbuf_0_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((lizzieLet15_1_argbuf_r && lizzieLet4_3QNone_Int_1_argbuf_0_bufchan_buf[0]))
        lizzieLet4_3QNone_Int_1_argbuf_0_bufchan_buf <= {32'd0, 1'd0};
      else if (((! lizzieLet15_1_argbuf_r) && (! lizzieLet4_3QNone_Int_1_argbuf_0_bufchan_buf[0])))
        lizzieLet4_3QNone_Int_1_argbuf_0_bufchan_buf <= lizzieLet4_3QNone_Int_1_argbuf_0_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet4_3QNone_Int_2,Go) > (lizzieLet4_3QNone_Int_2_argbuf,Go) */
  Go_t lizzieLet4_3QNone_Int_2_bufchan_d;
  logic lizzieLet4_3QNone_Int_2_bufchan_r;
  assign lizzieLet4_3QNone_Int_2_r = ((! lizzieLet4_3QNone_Int_2_bufchan_d[0]) || lizzieLet4_3QNone_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3QNone_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet4_3QNone_Int_2_r)
        lizzieLet4_3QNone_Int_2_bufchan_d <= lizzieLet4_3QNone_Int_2_d;
  Go_t lizzieLet4_3QNone_Int_2_bufchan_buf;
  assign lizzieLet4_3QNone_Int_2_bufchan_r = (! lizzieLet4_3QNone_Int_2_bufchan_buf[0]);
  assign lizzieLet4_3QNone_Int_2_argbuf_d = (lizzieLet4_3QNone_Int_2_bufchan_buf[0] ? lizzieLet4_3QNone_Int_2_bufchan_buf :
                                             lizzieLet4_3QNone_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3QNone_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet4_3QNone_Int_2_argbuf_r && lizzieLet4_3QNone_Int_2_bufchan_buf[0]))
        lizzieLet4_3QNone_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet4_3QNone_Int_2_argbuf_r) && (! lizzieLet4_3QNone_Int_2_bufchan_buf[0])))
        lizzieLet4_3QNone_Int_2_bufchan_buf <= lizzieLet4_3QNone_Int_2_bufchan_d;
  
  /* mergectrl (Ty C4,Ty Go) : [(lizzieLet4_3QNone_Int_2_argbuf,Go),
                           (lizzieLet25_3Lcall_$wnnz_Int0_1_argbuf,Go),
                           (lizzieLet4_3QVal_Int_2_argbuf,Go),
                           (lizzieLet4_3QError_Int_2_argbuf,Go)] > (go_18_goMux_choice,C4) (go_18_goMux_data,Go) */
  logic [3:0] lizzieLet4_3QNone_Int_2_argbuf_select_d;
  assign lizzieLet4_3QNone_Int_2_argbuf_select_d = ((| lizzieLet4_3QNone_Int_2_argbuf_select_q) ? lizzieLet4_3QNone_Int_2_argbuf_select_q :
                                                    (lizzieLet4_3QNone_Int_2_argbuf_d[0] ? 4'd1 :
                                                     (lizzieLet25_3Lcall_$wnnz_Int0_1_argbuf_d[0] ? 4'd2 :
                                                      (lizzieLet4_3QVal_Int_2_argbuf_d[0] ? 4'd4 :
                                                       (lizzieLet4_3QError_Int_2_argbuf_d[0] ? 4'd8 :
                                                        4'd0)))));
  logic [3:0] lizzieLet4_3QNone_Int_2_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_3QNone_Int_2_argbuf_select_q <= 4'd0;
    else
      lizzieLet4_3QNone_Int_2_argbuf_select_q <= (lizzieLet4_3QNone_Int_2_argbuf_done ? 4'd0 :
                                                  lizzieLet4_3QNone_Int_2_argbuf_select_d);
  logic [1:0] lizzieLet4_3QNone_Int_2_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3QNone_Int_2_argbuf_emit_q <= 2'd0;
    else
      lizzieLet4_3QNone_Int_2_argbuf_emit_q <= (lizzieLet4_3QNone_Int_2_argbuf_done ? 2'd0 :
                                                lizzieLet4_3QNone_Int_2_argbuf_emit_d);
  logic [1:0] lizzieLet4_3QNone_Int_2_argbuf_emit_d;
  assign lizzieLet4_3QNone_Int_2_argbuf_emit_d = (lizzieLet4_3QNone_Int_2_argbuf_emit_q | ({go_18_goMux_choice_d[0],
                                                                                            go_18_goMux_data_d[0]} & {go_18_goMux_choice_r,
                                                                                                                      go_18_goMux_data_r}));
  logic lizzieLet4_3QNone_Int_2_argbuf_done;
  assign lizzieLet4_3QNone_Int_2_argbuf_done = (& lizzieLet4_3QNone_Int_2_argbuf_emit_d);
  assign {lizzieLet4_3QError_Int_2_argbuf_r,
          lizzieLet4_3QVal_Int_2_argbuf_r,
          lizzieLet25_3Lcall_$wnnz_Int0_1_argbuf_r,
          lizzieLet4_3QNone_Int_2_argbuf_r} = (lizzieLet4_3QNone_Int_2_argbuf_done ? lizzieLet4_3QNone_Int_2_argbuf_select_d :
                                               4'd0);
  assign go_18_goMux_data_d = ((lizzieLet4_3QNone_Int_2_argbuf_select_d[0] && (! lizzieLet4_3QNone_Int_2_argbuf_emit_q[0])) ? lizzieLet4_3QNone_Int_2_argbuf_d :
                               ((lizzieLet4_3QNone_Int_2_argbuf_select_d[1] && (! lizzieLet4_3QNone_Int_2_argbuf_emit_q[0])) ? lizzieLet25_3Lcall_$wnnz_Int0_1_argbuf_d :
                                ((lizzieLet4_3QNone_Int_2_argbuf_select_d[2] && (! lizzieLet4_3QNone_Int_2_argbuf_emit_q[0])) ? lizzieLet4_3QVal_Int_2_argbuf_d :
                                 ((lizzieLet4_3QNone_Int_2_argbuf_select_d[3] && (! lizzieLet4_3QNone_Int_2_argbuf_emit_q[0])) ? lizzieLet4_3QError_Int_2_argbuf_d :
                                  1'd0))));
  assign go_18_goMux_choice_d = ((lizzieLet4_3QNone_Int_2_argbuf_select_d[0] && (! lizzieLet4_3QNone_Int_2_argbuf_emit_q[1])) ? C1_4_dc(1'd1) :
                                 ((lizzieLet4_3QNone_Int_2_argbuf_select_d[1] && (! lizzieLet4_3QNone_Int_2_argbuf_emit_q[1])) ? C2_4_dc(1'd1) :
                                  ((lizzieLet4_3QNone_Int_2_argbuf_select_d[2] && (! lizzieLet4_3QNone_Int_2_argbuf_emit_q[1])) ? C3_4_dc(1'd1) :
                                   ((lizzieLet4_3QNone_Int_2_argbuf_select_d[3] && (! lizzieLet4_3QNone_Int_2_argbuf_emit_q[1])) ? C4_4_dc(1'd1) :
                                    {2'd0, 1'd0}))));
  
  /* fork (Ty Go) : (lizzieLet4_3QVal_Int,Go) > [(lizzieLet4_3QVal_Int_1,Go),
                                            (lizzieLet4_3QVal_Int_2,Go)] */
  logic [1:0] lizzieLet4_3QVal_Int_emitted;
  logic [1:0] lizzieLet4_3QVal_Int_done;
  assign lizzieLet4_3QVal_Int_1_d = (lizzieLet4_3QVal_Int_d[0] && (! lizzieLet4_3QVal_Int_emitted[0]));
  assign lizzieLet4_3QVal_Int_2_d = (lizzieLet4_3QVal_Int_d[0] && (! lizzieLet4_3QVal_Int_emitted[1]));
  assign lizzieLet4_3QVal_Int_done = (lizzieLet4_3QVal_Int_emitted | ({lizzieLet4_3QVal_Int_2_d[0],
                                                                       lizzieLet4_3QVal_Int_1_d[0]} & {lizzieLet4_3QVal_Int_2_r,
                                                                                                       lizzieLet4_3QVal_Int_1_r}));
  assign lizzieLet4_3QVal_Int_r = (& lizzieLet4_3QVal_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3QVal_Int_emitted <= 2'd0;
    else
      lizzieLet4_3QVal_Int_emitted <= (lizzieLet4_3QVal_Int_r ? 2'd0 :
                                       lizzieLet4_3QVal_Int_done);
  
  /* buf (Ty Go) : (lizzieLet4_3QVal_Int_1,Go) > (lizzieLet4_3QVal_Int_1_argbuf,Go) */
  Go_t lizzieLet4_3QVal_Int_1_bufchan_d;
  logic lizzieLet4_3QVal_Int_1_bufchan_r;
  assign lizzieLet4_3QVal_Int_1_r = ((! lizzieLet4_3QVal_Int_1_bufchan_d[0]) || lizzieLet4_3QVal_Int_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3QVal_Int_1_bufchan_d <= 1'd0;
    else
      if (lizzieLet4_3QVal_Int_1_r)
        lizzieLet4_3QVal_Int_1_bufchan_d <= lizzieLet4_3QVal_Int_1_d;
  Go_t lizzieLet4_3QVal_Int_1_bufchan_buf;
  assign lizzieLet4_3QVal_Int_1_bufchan_r = (! lizzieLet4_3QVal_Int_1_bufchan_buf[0]);
  assign lizzieLet4_3QVal_Int_1_argbuf_d = (lizzieLet4_3QVal_Int_1_bufchan_buf[0] ? lizzieLet4_3QVal_Int_1_bufchan_buf :
                                            lizzieLet4_3QVal_Int_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3QVal_Int_1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet4_3QVal_Int_1_argbuf_r && lizzieLet4_3QVal_Int_1_bufchan_buf[0]))
        lizzieLet4_3QVal_Int_1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet4_3QVal_Int_1_argbuf_r) && (! lizzieLet4_3QVal_Int_1_bufchan_buf[0])))
        lizzieLet4_3QVal_Int_1_bufchan_buf <= lizzieLet4_3QVal_Int_1_bufchan_d;
  
  /* const (Ty Int#,
       Lit 1) : (lizzieLet4_3QVal_Int_1_argbuf,Go) > (lizzieLet4_3QVal_Int_1_argbuf_1,Int#) */
  assign lizzieLet4_3QVal_Int_1_argbuf_1_d = {32'd1,
                                              lizzieLet4_3QVal_Int_1_argbuf_d[0]};
  assign lizzieLet4_3QVal_Int_1_argbuf_r = lizzieLet4_3QVal_Int_1_argbuf_1_r;
  
  /* buf (Ty Int#) : (lizzieLet4_3QVal_Int_1_argbuf_1,Int#) > (lizzieLet16_1_argbuf,Int#) */
  \Int#_t  lizzieLet4_3QVal_Int_1_argbuf_1_bufchan_d;
  logic lizzieLet4_3QVal_Int_1_argbuf_1_bufchan_r;
  assign lizzieLet4_3QVal_Int_1_argbuf_1_r = ((! lizzieLet4_3QVal_Int_1_argbuf_1_bufchan_d[0]) || lizzieLet4_3QVal_Int_1_argbuf_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_3QVal_Int_1_argbuf_1_bufchan_d <= {32'd0, 1'd0};
    else
      if (lizzieLet4_3QVal_Int_1_argbuf_1_r)
        lizzieLet4_3QVal_Int_1_argbuf_1_bufchan_d <= lizzieLet4_3QVal_Int_1_argbuf_1_d;
  \Int#_t  lizzieLet4_3QVal_Int_1_argbuf_1_bufchan_buf;
  assign lizzieLet4_3QVal_Int_1_argbuf_1_bufchan_r = (! lizzieLet4_3QVal_Int_1_argbuf_1_bufchan_buf[0]);
  assign lizzieLet16_1_argbuf_d = (lizzieLet4_3QVal_Int_1_argbuf_1_bufchan_buf[0] ? lizzieLet4_3QVal_Int_1_argbuf_1_bufchan_buf :
                                   lizzieLet4_3QVal_Int_1_argbuf_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_3QVal_Int_1_argbuf_1_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((lizzieLet16_1_argbuf_r && lizzieLet4_3QVal_Int_1_argbuf_1_bufchan_buf[0]))
        lizzieLet4_3QVal_Int_1_argbuf_1_bufchan_buf <= {32'd0, 1'd0};
      else if (((! lizzieLet16_1_argbuf_r) && (! lizzieLet4_3QVal_Int_1_argbuf_1_bufchan_buf[0])))
        lizzieLet4_3QVal_Int_1_argbuf_1_bufchan_buf <= lizzieLet4_3QVal_Int_1_argbuf_1_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet4_3QVal_Int_2,Go) > (lizzieLet4_3QVal_Int_2_argbuf,Go) */
  Go_t lizzieLet4_3QVal_Int_2_bufchan_d;
  logic lizzieLet4_3QVal_Int_2_bufchan_r;
  assign lizzieLet4_3QVal_Int_2_r = ((! lizzieLet4_3QVal_Int_2_bufchan_d[0]) || lizzieLet4_3QVal_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3QVal_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet4_3QVal_Int_2_r)
        lizzieLet4_3QVal_Int_2_bufchan_d <= lizzieLet4_3QVal_Int_2_d;
  Go_t lizzieLet4_3QVal_Int_2_bufchan_buf;
  assign lizzieLet4_3QVal_Int_2_bufchan_r = (! lizzieLet4_3QVal_Int_2_bufchan_buf[0]);
  assign lizzieLet4_3QVal_Int_2_argbuf_d = (lizzieLet4_3QVal_Int_2_bufchan_buf[0] ? lizzieLet4_3QVal_Int_2_bufchan_buf :
                                            lizzieLet4_3QVal_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3QVal_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet4_3QVal_Int_2_argbuf_r && lizzieLet4_3QVal_Int_2_bufchan_buf[0]))
        lizzieLet4_3QVal_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet4_3QVal_Int_2_argbuf_r) && (! lizzieLet4_3QVal_Int_2_bufchan_buf[0])))
        lizzieLet4_3QVal_Int_2_bufchan_buf <= lizzieLet4_3QVal_Int_2_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_CT$wnnz_Int) : (lizzieLet4_4,QTree_Int) (sc_0_goMux_mux,Pointer_CT$wnnz_Int) > [(lizzieLet4_4QNone_Int,Pointer_CT$wnnz_Int),
                                                                                                  (lizzieLet4_4QVal_Int,Pointer_CT$wnnz_Int),
                                                                                                  (lizzieLet4_4QNode_Int,Pointer_CT$wnnz_Int),
                                                                                                  (lizzieLet4_4QError_Int,Pointer_CT$wnnz_Int)] */
  logic [3:0] sc_0_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet4_4_d[0] && sc_0_goMux_mux_d[0]))
      unique case (lizzieLet4_4_d[2:1])
        2'd0: sc_0_goMux_mux_onehotd = 4'd1;
        2'd1: sc_0_goMux_mux_onehotd = 4'd2;
        2'd2: sc_0_goMux_mux_onehotd = 4'd4;
        2'd3: sc_0_goMux_mux_onehotd = 4'd8;
        default: sc_0_goMux_mux_onehotd = 4'd0;
      endcase
    else sc_0_goMux_mux_onehotd = 4'd0;
  assign lizzieLet4_4QNone_Int_d = {sc_0_goMux_mux_d[16:1],
                                    sc_0_goMux_mux_onehotd[0]};
  assign lizzieLet4_4QVal_Int_d = {sc_0_goMux_mux_d[16:1],
                                   sc_0_goMux_mux_onehotd[1]};
  assign lizzieLet4_4QNode_Int_d = {sc_0_goMux_mux_d[16:1],
                                    sc_0_goMux_mux_onehotd[2]};
  assign lizzieLet4_4QError_Int_d = {sc_0_goMux_mux_d[16:1],
                                     sc_0_goMux_mux_onehotd[3]};
  assign sc_0_goMux_mux_r = (| (sc_0_goMux_mux_onehotd & {lizzieLet4_4QError_Int_r,
                                                          lizzieLet4_4QNode_Int_r,
                                                          lizzieLet4_4QVal_Int_r,
                                                          lizzieLet4_4QNone_Int_r}));
  assign lizzieLet4_4_r = sc_0_goMux_mux_r;
  
  /* buf (Ty Pointer_CT$wnnz_Int) : (lizzieLet4_4QError_Int,Pointer_CT$wnnz_Int) > (lizzieLet4_4QError_Int_1_argbuf,Pointer_CT$wnnz_Int) */
  Pointer_CT$wnnz_Int_t lizzieLet4_4QError_Int_bufchan_d;
  logic lizzieLet4_4QError_Int_bufchan_r;
  assign lizzieLet4_4QError_Int_r = ((! lizzieLet4_4QError_Int_bufchan_d[0]) || lizzieLet4_4QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_4QError_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet4_4QError_Int_r)
        lizzieLet4_4QError_Int_bufchan_d <= lizzieLet4_4QError_Int_d;
  Pointer_CT$wnnz_Int_t lizzieLet4_4QError_Int_bufchan_buf;
  assign lizzieLet4_4QError_Int_bufchan_r = (! lizzieLet4_4QError_Int_bufchan_buf[0]);
  assign lizzieLet4_4QError_Int_1_argbuf_d = (lizzieLet4_4QError_Int_bufchan_buf[0] ? lizzieLet4_4QError_Int_bufchan_buf :
                                              lizzieLet4_4QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_4QError_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet4_4QError_Int_1_argbuf_r && lizzieLet4_4QError_Int_bufchan_buf[0]))
        lizzieLet4_4QError_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet4_4QError_Int_1_argbuf_r) && (! lizzieLet4_4QError_Int_bufchan_buf[0])))
        lizzieLet4_4QError_Int_bufchan_buf <= lizzieLet4_4QError_Int_bufchan_d;
  
  /* dcon (Ty CT$wnnz_Int,
      Dcon Lcall_$wnnz_Int3) : [(lizzieLet4_4QNode_Int,Pointer_CT$wnnz_Int),
                                (q4ac3_destruct,Pointer_QTree_Int),
                                (q3ac2_destruct,Pointer_QTree_Int),
                                (q2ac1_destruct,Pointer_QTree_Int)] > (lizzieLet4_4QNode_Int_1q4ac3_1q3ac2_1q2ac1_1Lcall_$wnnz_Int3,CT$wnnz_Int) */
  assign lizzieLet4_4QNode_Int_1q4ac3_1q3ac2_1q2ac1_1Lcall_$wnnz_Int3_d = Lcall_$wnnz_Int3_dc((& {lizzieLet4_4QNode_Int_d[0],
                                                                                                  q4ac3_destruct_d[0],
                                                                                                  q3ac2_destruct_d[0],
                                                                                                  q2ac1_destruct_d[0]}), lizzieLet4_4QNode_Int_d, q4ac3_destruct_d, q3ac2_destruct_d, q2ac1_destruct_d);
  assign {lizzieLet4_4QNode_Int_r,
          q4ac3_destruct_r,
          q3ac2_destruct_r,
          q2ac1_destruct_r} = {4 {(lizzieLet4_4QNode_Int_1q4ac3_1q3ac2_1q2ac1_1Lcall_$wnnz_Int3_r && lizzieLet4_4QNode_Int_1q4ac3_1q3ac2_1q2ac1_1Lcall_$wnnz_Int3_d[0])}};
  
  /* buf (Ty CT$wnnz_Int) : (lizzieLet4_4QNode_Int_1q4ac3_1q3ac2_1q2ac1_1Lcall_$wnnz_Int3,CT$wnnz_Int) > (lizzieLet5_1_argbuf,CT$wnnz_Int) */
  CT$wnnz_Int_t lizzieLet4_4QNode_Int_1q4ac3_1q3ac2_1q2ac1_1Lcall_$wnnz_Int3_bufchan_d;
  logic lizzieLet4_4QNode_Int_1q4ac3_1q3ac2_1q2ac1_1Lcall_$wnnz_Int3_bufchan_r;
  assign lizzieLet4_4QNode_Int_1q4ac3_1q3ac2_1q2ac1_1Lcall_$wnnz_Int3_r = ((! lizzieLet4_4QNode_Int_1q4ac3_1q3ac2_1q2ac1_1Lcall_$wnnz_Int3_bufchan_d[0]) || lizzieLet4_4QNode_Int_1q4ac3_1q3ac2_1q2ac1_1Lcall_$wnnz_Int3_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_4QNode_Int_1q4ac3_1q3ac2_1q2ac1_1Lcall_$wnnz_Int3_bufchan_d <= {115'd0,
                                                                                 1'd0};
    else
      if (lizzieLet4_4QNode_Int_1q4ac3_1q3ac2_1q2ac1_1Lcall_$wnnz_Int3_r)
        lizzieLet4_4QNode_Int_1q4ac3_1q3ac2_1q2ac1_1Lcall_$wnnz_Int3_bufchan_d <= lizzieLet4_4QNode_Int_1q4ac3_1q3ac2_1q2ac1_1Lcall_$wnnz_Int3_d;
  CT$wnnz_Int_t lizzieLet4_4QNode_Int_1q4ac3_1q3ac2_1q2ac1_1Lcall_$wnnz_Int3_bufchan_buf;
  assign lizzieLet4_4QNode_Int_1q4ac3_1q3ac2_1q2ac1_1Lcall_$wnnz_Int3_bufchan_r = (! lizzieLet4_4QNode_Int_1q4ac3_1q3ac2_1q2ac1_1Lcall_$wnnz_Int3_bufchan_buf[0]);
  assign lizzieLet5_1_argbuf_d = (lizzieLet4_4QNode_Int_1q4ac3_1q3ac2_1q2ac1_1Lcall_$wnnz_Int3_bufchan_buf[0] ? lizzieLet4_4QNode_Int_1q4ac3_1q3ac2_1q2ac1_1Lcall_$wnnz_Int3_bufchan_buf :
                                  lizzieLet4_4QNode_Int_1q4ac3_1q3ac2_1q2ac1_1Lcall_$wnnz_Int3_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_4QNode_Int_1q4ac3_1q3ac2_1q2ac1_1Lcall_$wnnz_Int3_bufchan_buf <= {115'd0,
                                                                                   1'd0};
    else
      if ((lizzieLet5_1_argbuf_r && lizzieLet4_4QNode_Int_1q4ac3_1q3ac2_1q2ac1_1Lcall_$wnnz_Int3_bufchan_buf[0]))
        lizzieLet4_4QNode_Int_1q4ac3_1q3ac2_1q2ac1_1Lcall_$wnnz_Int3_bufchan_buf <= {115'd0,
                                                                                     1'd0};
      else if (((! lizzieLet5_1_argbuf_r) && (! lizzieLet4_4QNode_Int_1q4ac3_1q3ac2_1q2ac1_1Lcall_$wnnz_Int3_bufchan_buf[0])))
        lizzieLet4_4QNode_Int_1q4ac3_1q3ac2_1q2ac1_1Lcall_$wnnz_Int3_bufchan_buf <= lizzieLet4_4QNode_Int_1q4ac3_1q3ac2_1q2ac1_1Lcall_$wnnz_Int3_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz_Int) : (lizzieLet4_4QNone_Int,Pointer_CT$wnnz_Int) > (lizzieLet4_4QNone_Int_1_argbuf,Pointer_CT$wnnz_Int) */
  Pointer_CT$wnnz_Int_t lizzieLet4_4QNone_Int_bufchan_d;
  logic lizzieLet4_4QNone_Int_bufchan_r;
  assign lizzieLet4_4QNone_Int_r = ((! lizzieLet4_4QNone_Int_bufchan_d[0]) || lizzieLet4_4QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_4QNone_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet4_4QNone_Int_r)
        lizzieLet4_4QNone_Int_bufchan_d <= lizzieLet4_4QNone_Int_d;
  Pointer_CT$wnnz_Int_t lizzieLet4_4QNone_Int_bufchan_buf;
  assign lizzieLet4_4QNone_Int_bufchan_r = (! lizzieLet4_4QNone_Int_bufchan_buf[0]);
  assign lizzieLet4_4QNone_Int_1_argbuf_d = (lizzieLet4_4QNone_Int_bufchan_buf[0] ? lizzieLet4_4QNone_Int_bufchan_buf :
                                             lizzieLet4_4QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_4QNone_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet4_4QNone_Int_1_argbuf_r && lizzieLet4_4QNone_Int_bufchan_buf[0]))
        lizzieLet4_4QNone_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet4_4QNone_Int_1_argbuf_r) && (! lizzieLet4_4QNone_Int_bufchan_buf[0])))
        lizzieLet4_4QNone_Int_bufchan_buf <= lizzieLet4_4QNone_Int_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz_Int) : (lizzieLet4_4QVal_Int,Pointer_CT$wnnz_Int) > (lizzieLet4_4QVal_Int_1_argbuf,Pointer_CT$wnnz_Int) */
  Pointer_CT$wnnz_Int_t lizzieLet4_4QVal_Int_bufchan_d;
  logic lizzieLet4_4QVal_Int_bufchan_r;
  assign lizzieLet4_4QVal_Int_r = ((! lizzieLet4_4QVal_Int_bufchan_d[0]) || lizzieLet4_4QVal_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_4QVal_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet4_4QVal_Int_r)
        lizzieLet4_4QVal_Int_bufchan_d <= lizzieLet4_4QVal_Int_d;
  Pointer_CT$wnnz_Int_t lizzieLet4_4QVal_Int_bufchan_buf;
  assign lizzieLet4_4QVal_Int_bufchan_r = (! lizzieLet4_4QVal_Int_bufchan_buf[0]);
  assign lizzieLet4_4QVal_Int_1_argbuf_d = (lizzieLet4_4QVal_Int_bufchan_buf[0] ? lizzieLet4_4QVal_Int_bufchan_buf :
                                            lizzieLet4_4QVal_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_4QVal_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet4_4QVal_Int_1_argbuf_r && lizzieLet4_4QVal_Int_bufchan_buf[0]))
        lizzieLet4_4QVal_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet4_4QVal_Int_1_argbuf_r) && (! lizzieLet4_4QVal_Int_bufchan_buf[0])))
        lizzieLet4_4QVal_Int_bufchan_buf <= lizzieLet4_4QVal_Int_bufchan_d;
  
  /* destruct (Ty QTree_Int,
          Dcon QNode_Int) : (lizzieLet6_1QNode_Int,QTree_Int) > [(q1ad7_destruct,Pointer_QTree_Int),
                                                                 (q2ad8_destruct,Pointer_QTree_Int),
                                                                 (q3ad9_destruct,Pointer_QTree_Int),
                                                                 (q4ada_destruct,Pointer_QTree_Int)] */
  logic [3:0] lizzieLet6_1QNode_Int_emitted;
  logic [3:0] lizzieLet6_1QNode_Int_done;
  assign q1ad7_destruct_d = {lizzieLet6_1QNode_Int_d[18:3],
                             (lizzieLet6_1QNode_Int_d[0] && (! lizzieLet6_1QNode_Int_emitted[0]))};
  assign q2ad8_destruct_d = {lizzieLet6_1QNode_Int_d[34:19],
                             (lizzieLet6_1QNode_Int_d[0] && (! lizzieLet6_1QNode_Int_emitted[1]))};
  assign q3ad9_destruct_d = {lizzieLet6_1QNode_Int_d[50:35],
                             (lizzieLet6_1QNode_Int_d[0] && (! lizzieLet6_1QNode_Int_emitted[2]))};
  assign q4ada_destruct_d = {lizzieLet6_1QNode_Int_d[66:51],
                             (lizzieLet6_1QNode_Int_d[0] && (! lizzieLet6_1QNode_Int_emitted[3]))};
  assign lizzieLet6_1QNode_Int_done = (lizzieLet6_1QNode_Int_emitted | ({q4ada_destruct_d[0],
                                                                         q3ad9_destruct_d[0],
                                                                         q2ad8_destruct_d[0],
                                                                         q1ad7_destruct_d[0]} & {q4ada_destruct_r,
                                                                                                 q3ad9_destruct_r,
                                                                                                 q2ad8_destruct_r,
                                                                                                 q1ad7_destruct_r}));
  assign lizzieLet6_1QNode_Int_r = (& lizzieLet6_1QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_1QNode_Int_emitted <= 4'd0;
    else
      lizzieLet6_1QNode_Int_emitted <= (lizzieLet6_1QNode_Int_r ? 4'd0 :
                                        lizzieLet6_1QNode_Int_done);
  
  /* destruct (Ty QTree_Int,
          Dcon QVal_Int) : (lizzieLet6_1QVal_Int,QTree_Int) > [(vad6_destruct,Int)] */
  assign vad6_destruct_d = {lizzieLet6_1QVal_Int_d[34:3],
                            lizzieLet6_1QVal_Int_d[0]};
  assign lizzieLet6_1QVal_Int_r = vad6_destruct_r;
  
  /* demux (Ty QTree_Int,
       Ty QTree_Int) : (lizzieLet6_2,QTree_Int) (lizzieLet6_1,QTree_Int) > [(_7,QTree_Int),
                                                                            (lizzieLet6_1QVal_Int,QTree_Int),
                                                                            (lizzieLet6_1QNode_Int,QTree_Int),
                                                                            (_6,QTree_Int)] */
  logic [3:0] lizzieLet6_1_onehotd;
  always_comb
    if ((lizzieLet6_2_d[0] && lizzieLet6_1_d[0]))
      unique case (lizzieLet6_2_d[2:1])
        2'd0: lizzieLet6_1_onehotd = 4'd1;
        2'd1: lizzieLet6_1_onehotd = 4'd2;
        2'd2: lizzieLet6_1_onehotd = 4'd4;
        2'd3: lizzieLet6_1_onehotd = 4'd8;
        default: lizzieLet6_1_onehotd = 4'd0;
      endcase
    else lizzieLet6_1_onehotd = 4'd0;
  assign _7_d = {lizzieLet6_1_d[66:1], lizzieLet6_1_onehotd[0]};
  assign lizzieLet6_1QVal_Int_d = {lizzieLet6_1_d[66:1],
                                   lizzieLet6_1_onehotd[1]};
  assign lizzieLet6_1QNode_Int_d = {lizzieLet6_1_d[66:1],
                                    lizzieLet6_1_onehotd[2]};
  assign _6_d = {lizzieLet6_1_d[66:1], lizzieLet6_1_onehotd[3]};
  assign lizzieLet6_1_r = (| (lizzieLet6_1_onehotd & {_6_r,
                                                      lizzieLet6_1QNode_Int_r,
                                                      lizzieLet6_1QVal_Int_r,
                                                      _7_r}));
  assign lizzieLet6_2_r = lizzieLet6_1_r;
  
  /* demux (Ty QTree_Int,
       Ty MyDTInt_Int_Int) : (lizzieLet6_3,QTree_Int) (gad3_goMux_mux,MyDTInt_Int_Int) > [(_5,MyDTInt_Int_Int),
                                                                                          (lizzieLet6_3QVal_Int,MyDTInt_Int_Int),
                                                                                          (lizzieLet6_3QNode_Int,MyDTInt_Int_Int),
                                                                                          (_4,MyDTInt_Int_Int)] */
  logic [3:0] gad3_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet6_3_d[0] && gad3_goMux_mux_d[0]))
      unique case (lizzieLet6_3_d[2:1])
        2'd0: gad3_goMux_mux_onehotd = 4'd1;
        2'd1: gad3_goMux_mux_onehotd = 4'd2;
        2'd2: gad3_goMux_mux_onehotd = 4'd4;
        2'd3: gad3_goMux_mux_onehotd = 4'd8;
        default: gad3_goMux_mux_onehotd = 4'd0;
      endcase
    else gad3_goMux_mux_onehotd = 4'd0;
  assign _5_d = gad3_goMux_mux_onehotd[0];
  assign lizzieLet6_3QVal_Int_d = gad3_goMux_mux_onehotd[1];
  assign lizzieLet6_3QNode_Int_d = gad3_goMux_mux_onehotd[2];
  assign _4_d = gad3_goMux_mux_onehotd[3];
  assign gad3_goMux_mux_r = (| (gad3_goMux_mux_onehotd & {_4_r,
                                                          lizzieLet6_3QNode_Int_r,
                                                          lizzieLet6_3QVal_Int_r,
                                                          _5_r}));
  assign lizzieLet6_3_r = gad3_goMux_mux_r;
  
  /* fork (Ty MyDTInt_Int_Int) : (lizzieLet6_3QNode_Int,MyDTInt_Int_Int) > [(lizzieLet6_3QNode_Int_1,MyDTInt_Int_Int),
                                                                       (lizzieLet6_3QNode_Int_2,MyDTInt_Int_Int)] */
  logic [1:0] lizzieLet6_3QNode_Int_emitted;
  logic [1:0] lizzieLet6_3QNode_Int_done;
  assign lizzieLet6_3QNode_Int_1_d = (lizzieLet6_3QNode_Int_d[0] && (! lizzieLet6_3QNode_Int_emitted[0]));
  assign lizzieLet6_3QNode_Int_2_d = (lizzieLet6_3QNode_Int_d[0] && (! lizzieLet6_3QNode_Int_emitted[1]));
  assign lizzieLet6_3QNode_Int_done = (lizzieLet6_3QNode_Int_emitted | ({lizzieLet6_3QNode_Int_2_d[0],
                                                                         lizzieLet6_3QNode_Int_1_d[0]} & {lizzieLet6_3QNode_Int_2_r,
                                                                                                          lizzieLet6_3QNode_Int_1_r}));
  assign lizzieLet6_3QNode_Int_r = (& lizzieLet6_3QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_3QNode_Int_emitted <= 2'd0;
    else
      lizzieLet6_3QNode_Int_emitted <= (lizzieLet6_3QNode_Int_r ? 2'd0 :
                                        lizzieLet6_3QNode_Int_done);
  
  /* buf (Ty MyDTInt_Int_Int) : (lizzieLet6_3QNode_Int_2,MyDTInt_Int_Int) > (lizzieLet6_3QNode_Int_2_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t lizzieLet6_3QNode_Int_2_bufchan_d;
  logic lizzieLet6_3QNode_Int_2_bufchan_r;
  assign lizzieLet6_3QNode_Int_2_r = ((! lizzieLet6_3QNode_Int_2_bufchan_d[0]) || lizzieLet6_3QNode_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_3QNode_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet6_3QNode_Int_2_r)
        lizzieLet6_3QNode_Int_2_bufchan_d <= lizzieLet6_3QNode_Int_2_d;
  MyDTInt_Int_Int_t lizzieLet6_3QNode_Int_2_bufchan_buf;
  assign lizzieLet6_3QNode_Int_2_bufchan_r = (! lizzieLet6_3QNode_Int_2_bufchan_buf[0]);
  assign lizzieLet6_3QNode_Int_2_argbuf_d = (lizzieLet6_3QNode_Int_2_bufchan_buf[0] ? lizzieLet6_3QNode_Int_2_bufchan_buf :
                                             lizzieLet6_3QNode_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_3QNode_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet6_3QNode_Int_2_argbuf_r && lizzieLet6_3QNode_Int_2_bufchan_buf[0]))
        lizzieLet6_3QNode_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet6_3QNode_Int_2_argbuf_r) && (! lizzieLet6_3QNode_Int_2_bufchan_buf[0])))
        lizzieLet6_3QNode_Int_2_bufchan_buf <= lizzieLet6_3QNode_Int_2_bufchan_d;
  
  /* buf (Ty MyDTInt_Int_Int) : (lizzieLet6_3QVal_Int,MyDTInt_Int_Int) > (lizzieLet6_3QVal_Int_1_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t lizzieLet6_3QVal_Int_bufchan_d;
  logic lizzieLet6_3QVal_Int_bufchan_r;
  assign lizzieLet6_3QVal_Int_r = ((! lizzieLet6_3QVal_Int_bufchan_d[0]) || lizzieLet6_3QVal_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_3QVal_Int_bufchan_d <= 1'd0;
    else
      if (lizzieLet6_3QVal_Int_r)
        lizzieLet6_3QVal_Int_bufchan_d <= lizzieLet6_3QVal_Int_d;
  MyDTInt_Int_Int_t lizzieLet6_3QVal_Int_bufchan_buf;
  assign lizzieLet6_3QVal_Int_bufchan_r = (! lizzieLet6_3QVal_Int_bufchan_buf[0]);
  assign lizzieLet6_3QVal_Int_1_argbuf_d = (lizzieLet6_3QVal_Int_bufchan_buf[0] ? lizzieLet6_3QVal_Int_bufchan_buf :
                                            lizzieLet6_3QVal_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_3QVal_Int_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet6_3QVal_Int_1_argbuf_r && lizzieLet6_3QVal_Int_bufchan_buf[0]))
        lizzieLet6_3QVal_Int_bufchan_buf <= 1'd0;
      else if (((! lizzieLet6_3QVal_Int_1_argbuf_r) && (! lizzieLet6_3QVal_Int_bufchan_buf[0])))
        lizzieLet6_3QVal_Int_bufchan_buf <= lizzieLet6_3QVal_Int_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Go) : (lizzieLet6_4,QTree_Int) (go_12_goMux_data,Go) > [(lizzieLet6_4QNone_Int,Go),
                                                                  (lizzieLet6_4QVal_Int,Go),
                                                                  (lizzieLet6_4QNode_Int,Go),
                                                                  (lizzieLet6_4QError_Int,Go)] */
  logic [3:0] go_12_goMux_data_onehotd;
  always_comb
    if ((lizzieLet6_4_d[0] && go_12_goMux_data_d[0]))
      unique case (lizzieLet6_4_d[2:1])
        2'd0: go_12_goMux_data_onehotd = 4'd1;
        2'd1: go_12_goMux_data_onehotd = 4'd2;
        2'd2: go_12_goMux_data_onehotd = 4'd4;
        2'd3: go_12_goMux_data_onehotd = 4'd8;
        default: go_12_goMux_data_onehotd = 4'd0;
      endcase
    else go_12_goMux_data_onehotd = 4'd0;
  assign lizzieLet6_4QNone_Int_d = go_12_goMux_data_onehotd[0];
  assign lizzieLet6_4QVal_Int_d = go_12_goMux_data_onehotd[1];
  assign lizzieLet6_4QNode_Int_d = go_12_goMux_data_onehotd[2];
  assign lizzieLet6_4QError_Int_d = go_12_goMux_data_onehotd[3];
  assign go_12_goMux_data_r = (| (go_12_goMux_data_onehotd & {lizzieLet6_4QError_Int_r,
                                                              lizzieLet6_4QNode_Int_r,
                                                              lizzieLet6_4QVal_Int_r,
                                                              lizzieLet6_4QNone_Int_r}));
  assign lizzieLet6_4_r = go_12_goMux_data_r;
  
  /* fork (Ty Go) : (lizzieLet6_4QError_Int,Go) > [(lizzieLet6_4QError_Int_1,Go),
                                              (lizzieLet6_4QError_Int_2,Go)] */
  logic [1:0] lizzieLet6_4QError_Int_emitted;
  logic [1:0] lizzieLet6_4QError_Int_done;
  assign lizzieLet6_4QError_Int_1_d = (lizzieLet6_4QError_Int_d[0] && (! lizzieLet6_4QError_Int_emitted[0]));
  assign lizzieLet6_4QError_Int_2_d = (lizzieLet6_4QError_Int_d[0] && (! lizzieLet6_4QError_Int_emitted[1]));
  assign lizzieLet6_4QError_Int_done = (lizzieLet6_4QError_Int_emitted | ({lizzieLet6_4QError_Int_2_d[0],
                                                                           lizzieLet6_4QError_Int_1_d[0]} & {lizzieLet6_4QError_Int_2_r,
                                                                                                             lizzieLet6_4QError_Int_1_r}));
  assign lizzieLet6_4QError_Int_r = (& lizzieLet6_4QError_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_4QError_Int_emitted <= 2'd0;
    else
      lizzieLet6_4QError_Int_emitted <= (lizzieLet6_4QError_Int_r ? 2'd0 :
                                         lizzieLet6_4QError_Int_done);
  
  /* dcon (Ty QTree_Int,
      Dcon QError_Int) : [(lizzieLet6_4QError_Int_1,Go)] > (lizzieLet6_4QError_Int_1QError_Int,QTree_Int) */
  assign lizzieLet6_4QError_Int_1QError_Int_d = QError_Int_dc((& {lizzieLet6_4QError_Int_1_d[0]}), lizzieLet6_4QError_Int_1_d);
  assign {lizzieLet6_4QError_Int_1_r} = {1 {(lizzieLet6_4QError_Int_1QError_Int_r && lizzieLet6_4QError_Int_1QError_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (lizzieLet6_4QError_Int_1QError_Int,QTree_Int) > (lizzieLet9_1_argbuf,QTree_Int) */
  QTree_Int_t lizzieLet6_4QError_Int_1QError_Int_bufchan_d;
  logic lizzieLet6_4QError_Int_1QError_Int_bufchan_r;
  assign lizzieLet6_4QError_Int_1QError_Int_r = ((! lizzieLet6_4QError_Int_1QError_Int_bufchan_d[0]) || lizzieLet6_4QError_Int_1QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_4QError_Int_1QError_Int_bufchan_d <= {66'd0, 1'd0};
    else
      if (lizzieLet6_4QError_Int_1QError_Int_r)
        lizzieLet6_4QError_Int_1QError_Int_bufchan_d <= lizzieLet6_4QError_Int_1QError_Int_d;
  QTree_Int_t lizzieLet6_4QError_Int_1QError_Int_bufchan_buf;
  assign lizzieLet6_4QError_Int_1QError_Int_bufchan_r = (! lizzieLet6_4QError_Int_1QError_Int_bufchan_buf[0]);
  assign lizzieLet9_1_argbuf_d = (lizzieLet6_4QError_Int_1QError_Int_bufchan_buf[0] ? lizzieLet6_4QError_Int_1QError_Int_bufchan_buf :
                                  lizzieLet6_4QError_Int_1QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_4QError_Int_1QError_Int_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((lizzieLet9_1_argbuf_r && lizzieLet6_4QError_Int_1QError_Int_bufchan_buf[0]))
        lizzieLet6_4QError_Int_1QError_Int_bufchan_buf <= {66'd0, 1'd0};
      else if (((! lizzieLet9_1_argbuf_r) && (! lizzieLet6_4QError_Int_1QError_Int_bufchan_buf[0])))
        lizzieLet6_4QError_Int_1QError_Int_bufchan_buf <= lizzieLet6_4QError_Int_1QError_Int_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet6_4QError_Int_2,Go) > (lizzieLet6_4QError_Int_2_argbuf,Go) */
  Go_t lizzieLet6_4QError_Int_2_bufchan_d;
  logic lizzieLet6_4QError_Int_2_bufchan_r;
  assign lizzieLet6_4QError_Int_2_r = ((! lizzieLet6_4QError_Int_2_bufchan_d[0]) || lizzieLet6_4QError_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_4QError_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet6_4QError_Int_2_r)
        lizzieLet6_4QError_Int_2_bufchan_d <= lizzieLet6_4QError_Int_2_d;
  Go_t lizzieLet6_4QError_Int_2_bufchan_buf;
  assign lizzieLet6_4QError_Int_2_bufchan_r = (! lizzieLet6_4QError_Int_2_bufchan_buf[0]);
  assign lizzieLet6_4QError_Int_2_argbuf_d = (lizzieLet6_4QError_Int_2_bufchan_buf[0] ? lizzieLet6_4QError_Int_2_bufchan_buf :
                                              lizzieLet6_4QError_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_4QError_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet6_4QError_Int_2_argbuf_r && lizzieLet6_4QError_Int_2_bufchan_buf[0]))
        lizzieLet6_4QError_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet6_4QError_Int_2_argbuf_r) && (! lizzieLet6_4QError_Int_2_bufchan_buf[0])))
        lizzieLet6_4QError_Int_2_bufchan_buf <= lizzieLet6_4QError_Int_2_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet6_4QNode_Int,Go) > (lizzieLet6_4QNode_Int_1_argbuf,Go) */
  Go_t lizzieLet6_4QNode_Int_bufchan_d;
  logic lizzieLet6_4QNode_Int_bufchan_r;
  assign lizzieLet6_4QNode_Int_r = ((! lizzieLet6_4QNode_Int_bufchan_d[0]) || lizzieLet6_4QNode_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_4QNode_Int_bufchan_d <= 1'd0;
    else
      if (lizzieLet6_4QNode_Int_r)
        lizzieLet6_4QNode_Int_bufchan_d <= lizzieLet6_4QNode_Int_d;
  Go_t lizzieLet6_4QNode_Int_bufchan_buf;
  assign lizzieLet6_4QNode_Int_bufchan_r = (! lizzieLet6_4QNode_Int_bufchan_buf[0]);
  assign lizzieLet6_4QNode_Int_1_argbuf_d = (lizzieLet6_4QNode_Int_bufchan_buf[0] ? lizzieLet6_4QNode_Int_bufchan_buf :
                                             lizzieLet6_4QNode_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_4QNode_Int_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet6_4QNode_Int_1_argbuf_r && lizzieLet6_4QNode_Int_bufchan_buf[0]))
        lizzieLet6_4QNode_Int_bufchan_buf <= 1'd0;
      else if (((! lizzieLet6_4QNode_Int_1_argbuf_r) && (! lizzieLet6_4QNode_Int_bufchan_buf[0])))
        lizzieLet6_4QNode_Int_bufchan_buf <= lizzieLet6_4QNode_Int_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet6_4QNone_Int,Go) > [(lizzieLet6_4QNone_Int_1,Go),
                                             (lizzieLet6_4QNone_Int_2,Go)] */
  logic [1:0] lizzieLet6_4QNone_Int_emitted;
  logic [1:0] lizzieLet6_4QNone_Int_done;
  assign lizzieLet6_4QNone_Int_1_d = (lizzieLet6_4QNone_Int_d[0] && (! lizzieLet6_4QNone_Int_emitted[0]));
  assign lizzieLet6_4QNone_Int_2_d = (lizzieLet6_4QNone_Int_d[0] && (! lizzieLet6_4QNone_Int_emitted[1]));
  assign lizzieLet6_4QNone_Int_done = (lizzieLet6_4QNone_Int_emitted | ({lizzieLet6_4QNone_Int_2_d[0],
                                                                         lizzieLet6_4QNone_Int_1_d[0]} & {lizzieLet6_4QNone_Int_2_r,
                                                                                                          lizzieLet6_4QNone_Int_1_r}));
  assign lizzieLet6_4QNone_Int_r = (& lizzieLet6_4QNone_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_4QNone_Int_emitted <= 2'd0;
    else
      lizzieLet6_4QNone_Int_emitted <= (lizzieLet6_4QNone_Int_r ? 2'd0 :
                                        lizzieLet6_4QNone_Int_done);
  
  /* dcon (Ty QTree_Int,
      Dcon QNone_Int) : [(lizzieLet6_4QNone_Int_1,Go)] > (lizzieLet6_4QNone_Int_1QNone_Int,QTree_Int) */
  assign lizzieLet6_4QNone_Int_1QNone_Int_d = QNone_Int_dc((& {lizzieLet6_4QNone_Int_1_d[0]}), lizzieLet6_4QNone_Int_1_d);
  assign {lizzieLet6_4QNone_Int_1_r} = {1 {(lizzieLet6_4QNone_Int_1QNone_Int_r && lizzieLet6_4QNone_Int_1QNone_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (lizzieLet6_4QNone_Int_1QNone_Int,QTree_Int) > (lizzieLet7_1_argbuf,QTree_Int) */
  QTree_Int_t lizzieLet6_4QNone_Int_1QNone_Int_bufchan_d;
  logic lizzieLet6_4QNone_Int_1QNone_Int_bufchan_r;
  assign lizzieLet6_4QNone_Int_1QNone_Int_r = ((! lizzieLet6_4QNone_Int_1QNone_Int_bufchan_d[0]) || lizzieLet6_4QNone_Int_1QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_4QNone_Int_1QNone_Int_bufchan_d <= {66'd0, 1'd0};
    else
      if (lizzieLet6_4QNone_Int_1QNone_Int_r)
        lizzieLet6_4QNone_Int_1QNone_Int_bufchan_d <= lizzieLet6_4QNone_Int_1QNone_Int_d;
  QTree_Int_t lizzieLet6_4QNone_Int_1QNone_Int_bufchan_buf;
  assign lizzieLet6_4QNone_Int_1QNone_Int_bufchan_r = (! lizzieLet6_4QNone_Int_1QNone_Int_bufchan_buf[0]);
  assign lizzieLet7_1_argbuf_d = (lizzieLet6_4QNone_Int_1QNone_Int_bufchan_buf[0] ? lizzieLet6_4QNone_Int_1QNone_Int_bufchan_buf :
                                  lizzieLet6_4QNone_Int_1QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_4QNone_Int_1QNone_Int_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((lizzieLet7_1_argbuf_r && lizzieLet6_4QNone_Int_1QNone_Int_bufchan_buf[0]))
        lizzieLet6_4QNone_Int_1QNone_Int_bufchan_buf <= {66'd0, 1'd0};
      else if (((! lizzieLet7_1_argbuf_r) && (! lizzieLet6_4QNone_Int_1QNone_Int_bufchan_buf[0])))
        lizzieLet6_4QNone_Int_1QNone_Int_bufchan_buf <= lizzieLet6_4QNone_Int_1QNone_Int_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet6_4QNone_Int_2,Go) > (lizzieLet6_4QNone_Int_2_argbuf,Go) */
  Go_t lizzieLet6_4QNone_Int_2_bufchan_d;
  logic lizzieLet6_4QNone_Int_2_bufchan_r;
  assign lizzieLet6_4QNone_Int_2_r = ((! lizzieLet6_4QNone_Int_2_bufchan_d[0]) || lizzieLet6_4QNone_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_4QNone_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet6_4QNone_Int_2_r)
        lizzieLet6_4QNone_Int_2_bufchan_d <= lizzieLet6_4QNone_Int_2_d;
  Go_t lizzieLet6_4QNone_Int_2_bufchan_buf;
  assign lizzieLet6_4QNone_Int_2_bufchan_r = (! lizzieLet6_4QNone_Int_2_bufchan_buf[0]);
  assign lizzieLet6_4QNone_Int_2_argbuf_d = (lizzieLet6_4QNone_Int_2_bufchan_buf[0] ? lizzieLet6_4QNone_Int_2_bufchan_buf :
                                             lizzieLet6_4QNone_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_4QNone_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet6_4QNone_Int_2_argbuf_r && lizzieLet6_4QNone_Int_2_bufchan_buf[0]))
        lizzieLet6_4QNone_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet6_4QNone_Int_2_argbuf_r) && (! lizzieLet6_4QNone_Int_2_bufchan_buf[0])))
        lizzieLet6_4QNone_Int_2_bufchan_buf <= lizzieLet6_4QNone_Int_2_bufchan_d;
  
  /* mergectrl (Ty C4,Ty Go) : [(lizzieLet6_4QNone_Int_2_argbuf,Go),
                           (lizzieLet29_3Lcall_kron_kron_Int_Int_Int0_1_argbuf,Go),
                           (lizzieLet6_4QVal_Int_2_argbuf,Go),
                           (lizzieLet6_4QError_Int_2_argbuf,Go)] > (go_19_goMux_choice,C4) (go_19_goMux_data,Go) */
  logic [3:0] lizzieLet6_4QNone_Int_2_argbuf_select_d;
  assign lizzieLet6_4QNone_Int_2_argbuf_select_d = ((| lizzieLet6_4QNone_Int_2_argbuf_select_q) ? lizzieLet6_4QNone_Int_2_argbuf_select_q :
                                                    (lizzieLet6_4QNone_Int_2_argbuf_d[0] ? 4'd1 :
                                                     (lizzieLet29_3Lcall_kron_kron_Int_Int_Int0_1_argbuf_d[0] ? 4'd2 :
                                                      (lizzieLet6_4QVal_Int_2_argbuf_d[0] ? 4'd4 :
                                                       (lizzieLet6_4QError_Int_2_argbuf_d[0] ? 4'd8 :
                                                        4'd0)))));
  logic [3:0] lizzieLet6_4QNone_Int_2_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_4QNone_Int_2_argbuf_select_q <= 4'd0;
    else
      lizzieLet6_4QNone_Int_2_argbuf_select_q <= (lizzieLet6_4QNone_Int_2_argbuf_done ? 4'd0 :
                                                  lizzieLet6_4QNone_Int_2_argbuf_select_d);
  logic [1:0] lizzieLet6_4QNone_Int_2_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_4QNone_Int_2_argbuf_emit_q <= 2'd0;
    else
      lizzieLet6_4QNone_Int_2_argbuf_emit_q <= (lizzieLet6_4QNone_Int_2_argbuf_done ? 2'd0 :
                                                lizzieLet6_4QNone_Int_2_argbuf_emit_d);
  logic [1:0] lizzieLet6_4QNone_Int_2_argbuf_emit_d;
  assign lizzieLet6_4QNone_Int_2_argbuf_emit_d = (lizzieLet6_4QNone_Int_2_argbuf_emit_q | ({go_19_goMux_choice_d[0],
                                                                                            go_19_goMux_data_d[0]} & {go_19_goMux_choice_r,
                                                                                                                      go_19_goMux_data_r}));
  logic lizzieLet6_4QNone_Int_2_argbuf_done;
  assign lizzieLet6_4QNone_Int_2_argbuf_done = (& lizzieLet6_4QNone_Int_2_argbuf_emit_d);
  assign {lizzieLet6_4QError_Int_2_argbuf_r,
          lizzieLet6_4QVal_Int_2_argbuf_r,
          lizzieLet29_3Lcall_kron_kron_Int_Int_Int0_1_argbuf_r,
          lizzieLet6_4QNone_Int_2_argbuf_r} = (lizzieLet6_4QNone_Int_2_argbuf_done ? lizzieLet6_4QNone_Int_2_argbuf_select_d :
                                               4'd0);
  assign go_19_goMux_data_d = ((lizzieLet6_4QNone_Int_2_argbuf_select_d[0] && (! lizzieLet6_4QNone_Int_2_argbuf_emit_q[0])) ? lizzieLet6_4QNone_Int_2_argbuf_d :
                               ((lizzieLet6_4QNone_Int_2_argbuf_select_d[1] && (! lizzieLet6_4QNone_Int_2_argbuf_emit_q[0])) ? lizzieLet29_3Lcall_kron_kron_Int_Int_Int0_1_argbuf_d :
                                ((lizzieLet6_4QNone_Int_2_argbuf_select_d[2] && (! lizzieLet6_4QNone_Int_2_argbuf_emit_q[0])) ? lizzieLet6_4QVal_Int_2_argbuf_d :
                                 ((lizzieLet6_4QNone_Int_2_argbuf_select_d[3] && (! lizzieLet6_4QNone_Int_2_argbuf_emit_q[0])) ? lizzieLet6_4QError_Int_2_argbuf_d :
                                  1'd0))));
  assign go_19_goMux_choice_d = ((lizzieLet6_4QNone_Int_2_argbuf_select_d[0] && (! lizzieLet6_4QNone_Int_2_argbuf_emit_q[1])) ? C1_4_dc(1'd1) :
                                 ((lizzieLet6_4QNone_Int_2_argbuf_select_d[1] && (! lizzieLet6_4QNone_Int_2_argbuf_emit_q[1])) ? C2_4_dc(1'd1) :
                                  ((lizzieLet6_4QNone_Int_2_argbuf_select_d[2] && (! lizzieLet6_4QNone_Int_2_argbuf_emit_q[1])) ? C3_4_dc(1'd1) :
                                   ((lizzieLet6_4QNone_Int_2_argbuf_select_d[3] && (! lizzieLet6_4QNone_Int_2_argbuf_emit_q[1])) ? C4_4_dc(1'd1) :
                                    {2'd0, 1'd0}))));
  
  /* fork (Ty Go) : (lizzieLet6_4QVal_Int,Go) > [(lizzieLet6_4QVal_Int_1,Go),
                                            (lizzieLet6_4QVal_Int_2,Go)] */
  logic [1:0] lizzieLet6_4QVal_Int_emitted;
  logic [1:0] lizzieLet6_4QVal_Int_done;
  assign lizzieLet6_4QVal_Int_1_d = (lizzieLet6_4QVal_Int_d[0] && (! lizzieLet6_4QVal_Int_emitted[0]));
  assign lizzieLet6_4QVal_Int_2_d = (lizzieLet6_4QVal_Int_d[0] && (! lizzieLet6_4QVal_Int_emitted[1]));
  assign lizzieLet6_4QVal_Int_done = (lizzieLet6_4QVal_Int_emitted | ({lizzieLet6_4QVal_Int_2_d[0],
                                                                       lizzieLet6_4QVal_Int_1_d[0]} & {lizzieLet6_4QVal_Int_2_r,
                                                                                                       lizzieLet6_4QVal_Int_1_r}));
  assign lizzieLet6_4QVal_Int_r = (& lizzieLet6_4QVal_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_4QVal_Int_emitted <= 2'd0;
    else
      lizzieLet6_4QVal_Int_emitted <= (lizzieLet6_4QVal_Int_r ? 2'd0 :
                                       lizzieLet6_4QVal_Int_done);
  
  /* buf (Ty Go) : (lizzieLet6_4QVal_Int_1,Go) > (lizzieLet6_4QVal_Int_1_argbuf,Go) */
  Go_t lizzieLet6_4QVal_Int_1_bufchan_d;
  logic lizzieLet6_4QVal_Int_1_bufchan_r;
  assign lizzieLet6_4QVal_Int_1_r = ((! lizzieLet6_4QVal_Int_1_bufchan_d[0]) || lizzieLet6_4QVal_Int_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_4QVal_Int_1_bufchan_d <= 1'd0;
    else
      if (lizzieLet6_4QVal_Int_1_r)
        lizzieLet6_4QVal_Int_1_bufchan_d <= lizzieLet6_4QVal_Int_1_d;
  Go_t lizzieLet6_4QVal_Int_1_bufchan_buf;
  assign lizzieLet6_4QVal_Int_1_bufchan_r = (! lizzieLet6_4QVal_Int_1_bufchan_buf[0]);
  assign lizzieLet6_4QVal_Int_1_argbuf_d = (lizzieLet6_4QVal_Int_1_bufchan_buf[0] ? lizzieLet6_4QVal_Int_1_bufchan_buf :
                                            lizzieLet6_4QVal_Int_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_4QVal_Int_1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet6_4QVal_Int_1_argbuf_r && lizzieLet6_4QVal_Int_1_bufchan_buf[0]))
        lizzieLet6_4QVal_Int_1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet6_4QVal_Int_1_argbuf_r) && (! lizzieLet6_4QVal_Int_1_bufchan_buf[0])))
        lizzieLet6_4QVal_Int_1_bufchan_buf <= lizzieLet6_4QVal_Int_1_bufchan_d;
  
  /* dcon (Ty TupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int,
      Dcon TupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int) : [(lizzieLet6_4QVal_Int_1_argbuf,Go),
                                                                                (lizzieLet6_5QVal_Int_1_argbuf,MyDTInt_Bool),
                                                                                (lizzieLet6_3QVal_Int_1_argbuf,MyDTInt_Int_Int),
                                                                                (vad6_1_argbuf,Int),
                                                                                (lizzieLet6_6QVal_Int_1_argbuf,Pointer_QTree_Int)] > (map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int_1,TupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int) */
  assign \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int_1_d  = TupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int_dc((& {lizzieLet6_4QVal_Int_1_argbuf_d[0],
                                                                                                                                                                                 lizzieLet6_5QVal_Int_1_argbuf_d[0],
                                                                                                                                                                                 lizzieLet6_3QVal_Int_1_argbuf_d[0],
                                                                                                                                                                                 vad6_1_argbuf_d[0],
                                                                                                                                                                                 lizzieLet6_6QVal_Int_1_argbuf_d[0]}), lizzieLet6_4QVal_Int_1_argbuf_d, lizzieLet6_5QVal_Int_1_argbuf_d, lizzieLet6_3QVal_Int_1_argbuf_d, vad6_1_argbuf_d, lizzieLet6_6QVal_Int_1_argbuf_d);
  assign {lizzieLet6_4QVal_Int_1_argbuf_r,
          lizzieLet6_5QVal_Int_1_argbuf_r,
          lizzieLet6_3QVal_Int_1_argbuf_r,
          vad6_1_argbuf_r,
          lizzieLet6_6QVal_Int_1_argbuf_r} = {5 {(\map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int_1_r  && \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int_1_d [0])}};
  
  /* buf (Ty Go) : (lizzieLet6_4QVal_Int_2,Go) > (lizzieLet6_4QVal_Int_2_argbuf,Go) */
  Go_t lizzieLet6_4QVal_Int_2_bufchan_d;
  logic lizzieLet6_4QVal_Int_2_bufchan_r;
  assign lizzieLet6_4QVal_Int_2_r = ((! lizzieLet6_4QVal_Int_2_bufchan_d[0]) || lizzieLet6_4QVal_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_4QVal_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet6_4QVal_Int_2_r)
        lizzieLet6_4QVal_Int_2_bufchan_d <= lizzieLet6_4QVal_Int_2_d;
  Go_t lizzieLet6_4QVal_Int_2_bufchan_buf;
  assign lizzieLet6_4QVal_Int_2_bufchan_r = (! lizzieLet6_4QVal_Int_2_bufchan_buf[0]);
  assign lizzieLet6_4QVal_Int_2_argbuf_d = (lizzieLet6_4QVal_Int_2_bufchan_buf[0] ? lizzieLet6_4QVal_Int_2_bufchan_buf :
                                            lizzieLet6_4QVal_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_4QVal_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet6_4QVal_Int_2_argbuf_r && lizzieLet6_4QVal_Int_2_bufchan_buf[0]))
        lizzieLet6_4QVal_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet6_4QVal_Int_2_argbuf_r) && (! lizzieLet6_4QVal_Int_2_bufchan_buf[0])))
        lizzieLet6_4QVal_Int_2_bufchan_buf <= lizzieLet6_4QVal_Int_2_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty MyDTInt_Bool) : (lizzieLet6_5,QTree_Int) (isZad2_goMux_mux,MyDTInt_Bool) > [(_3,MyDTInt_Bool),
                                                                                      (lizzieLet6_5QVal_Int,MyDTInt_Bool),
                                                                                      (lizzieLet6_5QNode_Int,MyDTInt_Bool),
                                                                                      (_2,MyDTInt_Bool)] */
  logic [3:0] isZad2_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet6_5_d[0] && isZad2_goMux_mux_d[0]))
      unique case (lizzieLet6_5_d[2:1])
        2'd0: isZad2_goMux_mux_onehotd = 4'd1;
        2'd1: isZad2_goMux_mux_onehotd = 4'd2;
        2'd2: isZad2_goMux_mux_onehotd = 4'd4;
        2'd3: isZad2_goMux_mux_onehotd = 4'd8;
        default: isZad2_goMux_mux_onehotd = 4'd0;
      endcase
    else isZad2_goMux_mux_onehotd = 4'd0;
  assign _3_d = isZad2_goMux_mux_onehotd[0];
  assign lizzieLet6_5QVal_Int_d = isZad2_goMux_mux_onehotd[1];
  assign lizzieLet6_5QNode_Int_d = isZad2_goMux_mux_onehotd[2];
  assign _2_d = isZad2_goMux_mux_onehotd[3];
  assign isZad2_goMux_mux_r = (| (isZad2_goMux_mux_onehotd & {_2_r,
                                                              lizzieLet6_5QNode_Int_r,
                                                              lizzieLet6_5QVal_Int_r,
                                                              _3_r}));
  assign lizzieLet6_5_r = isZad2_goMux_mux_r;
  
  /* fork (Ty MyDTInt_Bool) : (lizzieLet6_5QNode_Int,MyDTInt_Bool) > [(lizzieLet6_5QNode_Int_1,MyDTInt_Bool),
                                                                 (lizzieLet6_5QNode_Int_2,MyDTInt_Bool)] */
  logic [1:0] lizzieLet6_5QNode_Int_emitted;
  logic [1:0] lizzieLet6_5QNode_Int_done;
  assign lizzieLet6_5QNode_Int_1_d = (lizzieLet6_5QNode_Int_d[0] && (! lizzieLet6_5QNode_Int_emitted[0]));
  assign lizzieLet6_5QNode_Int_2_d = (lizzieLet6_5QNode_Int_d[0] && (! lizzieLet6_5QNode_Int_emitted[1]));
  assign lizzieLet6_5QNode_Int_done = (lizzieLet6_5QNode_Int_emitted | ({lizzieLet6_5QNode_Int_2_d[0],
                                                                         lizzieLet6_5QNode_Int_1_d[0]} & {lizzieLet6_5QNode_Int_2_r,
                                                                                                          lizzieLet6_5QNode_Int_1_r}));
  assign lizzieLet6_5QNode_Int_r = (& lizzieLet6_5QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_5QNode_Int_emitted <= 2'd0;
    else
      lizzieLet6_5QNode_Int_emitted <= (lizzieLet6_5QNode_Int_r ? 2'd0 :
                                        lizzieLet6_5QNode_Int_done);
  
  /* buf (Ty MyDTInt_Bool) : (lizzieLet6_5QNode_Int_2,MyDTInt_Bool) > (lizzieLet6_5QNode_Int_2_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t lizzieLet6_5QNode_Int_2_bufchan_d;
  logic lizzieLet6_5QNode_Int_2_bufchan_r;
  assign lizzieLet6_5QNode_Int_2_r = ((! lizzieLet6_5QNode_Int_2_bufchan_d[0]) || lizzieLet6_5QNode_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_5QNode_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet6_5QNode_Int_2_r)
        lizzieLet6_5QNode_Int_2_bufchan_d <= lizzieLet6_5QNode_Int_2_d;
  MyDTInt_Bool_t lizzieLet6_5QNode_Int_2_bufchan_buf;
  assign lizzieLet6_5QNode_Int_2_bufchan_r = (! lizzieLet6_5QNode_Int_2_bufchan_buf[0]);
  assign lizzieLet6_5QNode_Int_2_argbuf_d = (lizzieLet6_5QNode_Int_2_bufchan_buf[0] ? lizzieLet6_5QNode_Int_2_bufchan_buf :
                                             lizzieLet6_5QNode_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_5QNode_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet6_5QNode_Int_2_argbuf_r && lizzieLet6_5QNode_Int_2_bufchan_buf[0]))
        lizzieLet6_5QNode_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet6_5QNode_Int_2_argbuf_r) && (! lizzieLet6_5QNode_Int_2_bufchan_buf[0])))
        lizzieLet6_5QNode_Int_2_bufchan_buf <= lizzieLet6_5QNode_Int_2_bufchan_d;
  
  /* buf (Ty MyDTInt_Bool) : (lizzieLet6_5QVal_Int,MyDTInt_Bool) > (lizzieLet6_5QVal_Int_1_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t lizzieLet6_5QVal_Int_bufchan_d;
  logic lizzieLet6_5QVal_Int_bufchan_r;
  assign lizzieLet6_5QVal_Int_r = ((! lizzieLet6_5QVal_Int_bufchan_d[0]) || lizzieLet6_5QVal_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_5QVal_Int_bufchan_d <= 1'd0;
    else
      if (lizzieLet6_5QVal_Int_r)
        lizzieLet6_5QVal_Int_bufchan_d <= lizzieLet6_5QVal_Int_d;
  MyDTInt_Bool_t lizzieLet6_5QVal_Int_bufchan_buf;
  assign lizzieLet6_5QVal_Int_bufchan_r = (! lizzieLet6_5QVal_Int_bufchan_buf[0]);
  assign lizzieLet6_5QVal_Int_1_argbuf_d = (lizzieLet6_5QVal_Int_bufchan_buf[0] ? lizzieLet6_5QVal_Int_bufchan_buf :
                                            lizzieLet6_5QVal_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_5QVal_Int_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet6_5QVal_Int_1_argbuf_r && lizzieLet6_5QVal_Int_bufchan_buf[0]))
        lizzieLet6_5QVal_Int_bufchan_buf <= 1'd0;
      else if (((! lizzieLet6_5QVal_Int_1_argbuf_r) && (! lizzieLet6_5QVal_Int_bufchan_buf[0])))
        lizzieLet6_5QVal_Int_bufchan_buf <= lizzieLet6_5QVal_Int_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_QTree_Int) : (lizzieLet6_6,QTree_Int) (m2ad5_goMux_mux,Pointer_QTree_Int) > [(_1,Pointer_QTree_Int),
                                                                                               (lizzieLet6_6QVal_Int,Pointer_QTree_Int),
                                                                                               (lizzieLet6_6QNode_Int,Pointer_QTree_Int),
                                                                                               (_0,Pointer_QTree_Int)] */
  logic [3:0] m2ad5_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet6_6_d[0] && m2ad5_goMux_mux_d[0]))
      unique case (lizzieLet6_6_d[2:1])
        2'd0: m2ad5_goMux_mux_onehotd = 4'd1;
        2'd1: m2ad5_goMux_mux_onehotd = 4'd2;
        2'd2: m2ad5_goMux_mux_onehotd = 4'd4;
        2'd3: m2ad5_goMux_mux_onehotd = 4'd8;
        default: m2ad5_goMux_mux_onehotd = 4'd0;
      endcase
    else m2ad5_goMux_mux_onehotd = 4'd0;
  assign _1_d = {m2ad5_goMux_mux_d[16:1],
                 m2ad5_goMux_mux_onehotd[0]};
  assign lizzieLet6_6QVal_Int_d = {m2ad5_goMux_mux_d[16:1],
                                   m2ad5_goMux_mux_onehotd[1]};
  assign lizzieLet6_6QNode_Int_d = {m2ad5_goMux_mux_d[16:1],
                                    m2ad5_goMux_mux_onehotd[2]};
  assign _0_d = {m2ad5_goMux_mux_d[16:1],
                 m2ad5_goMux_mux_onehotd[3]};
  assign m2ad5_goMux_mux_r = (| (m2ad5_goMux_mux_onehotd & {_0_r,
                                                            lizzieLet6_6QNode_Int_r,
                                                            lizzieLet6_6QVal_Int_r,
                                                            _1_r}));
  assign lizzieLet6_6_r = m2ad5_goMux_mux_r;
  
  /* fork (Ty Pointer_QTree_Int) : (lizzieLet6_6QNode_Int,Pointer_QTree_Int) > [(lizzieLet6_6QNode_Int_1,Pointer_QTree_Int),
                                                                           (lizzieLet6_6QNode_Int_2,Pointer_QTree_Int)] */
  logic [1:0] lizzieLet6_6QNode_Int_emitted;
  logic [1:0] lizzieLet6_6QNode_Int_done;
  assign lizzieLet6_6QNode_Int_1_d = {lizzieLet6_6QNode_Int_d[16:1],
                                      (lizzieLet6_6QNode_Int_d[0] && (! lizzieLet6_6QNode_Int_emitted[0]))};
  assign lizzieLet6_6QNode_Int_2_d = {lizzieLet6_6QNode_Int_d[16:1],
                                      (lizzieLet6_6QNode_Int_d[0] && (! lizzieLet6_6QNode_Int_emitted[1]))};
  assign lizzieLet6_6QNode_Int_done = (lizzieLet6_6QNode_Int_emitted | ({lizzieLet6_6QNode_Int_2_d[0],
                                                                         lizzieLet6_6QNode_Int_1_d[0]} & {lizzieLet6_6QNode_Int_2_r,
                                                                                                          lizzieLet6_6QNode_Int_1_r}));
  assign lizzieLet6_6QNode_Int_r = (& lizzieLet6_6QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_6QNode_Int_emitted <= 2'd0;
    else
      lizzieLet6_6QNode_Int_emitted <= (lizzieLet6_6QNode_Int_r ? 2'd0 :
                                        lizzieLet6_6QNode_Int_done);
  
  /* buf (Ty Pointer_QTree_Int) : (lizzieLet6_6QNode_Int_2,Pointer_QTree_Int) > (lizzieLet6_6QNode_Int_2_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t lizzieLet6_6QNode_Int_2_bufchan_d;
  logic lizzieLet6_6QNode_Int_2_bufchan_r;
  assign lizzieLet6_6QNode_Int_2_r = ((! lizzieLet6_6QNode_Int_2_bufchan_d[0]) || lizzieLet6_6QNode_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_6QNode_Int_2_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet6_6QNode_Int_2_r)
        lizzieLet6_6QNode_Int_2_bufchan_d <= lizzieLet6_6QNode_Int_2_d;
  Pointer_QTree_Int_t lizzieLet6_6QNode_Int_2_bufchan_buf;
  assign lizzieLet6_6QNode_Int_2_bufchan_r = (! lizzieLet6_6QNode_Int_2_bufchan_buf[0]);
  assign lizzieLet6_6QNode_Int_2_argbuf_d = (lizzieLet6_6QNode_Int_2_bufchan_buf[0] ? lizzieLet6_6QNode_Int_2_bufchan_buf :
                                             lizzieLet6_6QNode_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_6QNode_Int_2_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet6_6QNode_Int_2_argbuf_r && lizzieLet6_6QNode_Int_2_bufchan_buf[0]))
        lizzieLet6_6QNode_Int_2_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet6_6QNode_Int_2_argbuf_r) && (! lizzieLet6_6QNode_Int_2_bufchan_buf[0])))
        lizzieLet6_6QNode_Int_2_bufchan_buf <= lizzieLet6_6QNode_Int_2_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (lizzieLet6_6QVal_Int,Pointer_QTree_Int) > (lizzieLet6_6QVal_Int_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t lizzieLet6_6QVal_Int_bufchan_d;
  logic lizzieLet6_6QVal_Int_bufchan_r;
  assign lizzieLet6_6QVal_Int_r = ((! lizzieLet6_6QVal_Int_bufchan_d[0]) || lizzieLet6_6QVal_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_6QVal_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet6_6QVal_Int_r)
        lizzieLet6_6QVal_Int_bufchan_d <= lizzieLet6_6QVal_Int_d;
  Pointer_QTree_Int_t lizzieLet6_6QVal_Int_bufchan_buf;
  assign lizzieLet6_6QVal_Int_bufchan_r = (! lizzieLet6_6QVal_Int_bufchan_buf[0]);
  assign lizzieLet6_6QVal_Int_1_argbuf_d = (lizzieLet6_6QVal_Int_bufchan_buf[0] ? lizzieLet6_6QVal_Int_bufchan_buf :
                                            lizzieLet6_6QVal_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_6QVal_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet6_6QVal_Int_1_argbuf_r && lizzieLet6_6QVal_Int_bufchan_buf[0]))
        lizzieLet6_6QVal_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet6_6QVal_Int_1_argbuf_r) && (! lizzieLet6_6QVal_Int_bufchan_buf[0])))
        lizzieLet6_6QVal_Int_bufchan_buf <= lizzieLet6_6QVal_Int_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_CTkron_kron_Int_Int_Int) : (lizzieLet6_7,QTree_Int) (sc_0_1_goMux_mux,Pointer_CTkron_kron_Int_Int_Int) > [(lizzieLet6_7QNone_Int,Pointer_CTkron_kron_Int_Int_Int),
                                                                                                                            (lizzieLet6_7QVal_Int,Pointer_CTkron_kron_Int_Int_Int),
                                                                                                                            (lizzieLet6_7QNode_Int,Pointer_CTkron_kron_Int_Int_Int),
                                                                                                                            (lizzieLet6_7QError_Int,Pointer_CTkron_kron_Int_Int_Int)] */
  logic [3:0] sc_0_1_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet6_7_d[0] && sc_0_1_goMux_mux_d[0]))
      unique case (lizzieLet6_7_d[2:1])
        2'd0: sc_0_1_goMux_mux_onehotd = 4'd1;
        2'd1: sc_0_1_goMux_mux_onehotd = 4'd2;
        2'd2: sc_0_1_goMux_mux_onehotd = 4'd4;
        2'd3: sc_0_1_goMux_mux_onehotd = 4'd8;
        default: sc_0_1_goMux_mux_onehotd = 4'd0;
      endcase
    else sc_0_1_goMux_mux_onehotd = 4'd0;
  assign lizzieLet6_7QNone_Int_d = {sc_0_1_goMux_mux_d[16:1],
                                    sc_0_1_goMux_mux_onehotd[0]};
  assign lizzieLet6_7QVal_Int_d = {sc_0_1_goMux_mux_d[16:1],
                                   sc_0_1_goMux_mux_onehotd[1]};
  assign lizzieLet6_7QNode_Int_d = {sc_0_1_goMux_mux_d[16:1],
                                    sc_0_1_goMux_mux_onehotd[2]};
  assign lizzieLet6_7QError_Int_d = {sc_0_1_goMux_mux_d[16:1],
                                     sc_0_1_goMux_mux_onehotd[3]};
  assign sc_0_1_goMux_mux_r = (| (sc_0_1_goMux_mux_onehotd & {lizzieLet6_7QError_Int_r,
                                                              lizzieLet6_7QNode_Int_r,
                                                              lizzieLet6_7QVal_Int_r,
                                                              lizzieLet6_7QNone_Int_r}));
  assign lizzieLet6_7_r = sc_0_1_goMux_mux_r;
  
  /* buf (Ty Pointer_CTkron_kron_Int_Int_Int) : (lizzieLet6_7QError_Int,Pointer_CTkron_kron_Int_Int_Int) > (lizzieLet6_7QError_Int_1_argbuf,Pointer_CTkron_kron_Int_Int_Int) */
  Pointer_CTkron_kron_Int_Int_Int_t lizzieLet6_7QError_Int_bufchan_d;
  logic lizzieLet6_7QError_Int_bufchan_r;
  assign lizzieLet6_7QError_Int_r = ((! lizzieLet6_7QError_Int_bufchan_d[0]) || lizzieLet6_7QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_7QError_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet6_7QError_Int_r)
        lizzieLet6_7QError_Int_bufchan_d <= lizzieLet6_7QError_Int_d;
  Pointer_CTkron_kron_Int_Int_Int_t lizzieLet6_7QError_Int_bufchan_buf;
  assign lizzieLet6_7QError_Int_bufchan_r = (! lizzieLet6_7QError_Int_bufchan_buf[0]);
  assign lizzieLet6_7QError_Int_1_argbuf_d = (lizzieLet6_7QError_Int_bufchan_buf[0] ? lizzieLet6_7QError_Int_bufchan_buf :
                                              lizzieLet6_7QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_7QError_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet6_7QError_Int_1_argbuf_r && lizzieLet6_7QError_Int_bufchan_buf[0]))
        lizzieLet6_7QError_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet6_7QError_Int_1_argbuf_r) && (! lizzieLet6_7QError_Int_bufchan_buf[0])))
        lizzieLet6_7QError_Int_bufchan_buf <= lizzieLet6_7QError_Int_bufchan_d;
  
  /* dcon (Ty CTkron_kron_Int_Int_Int,
      Dcon Lcall_kron_kron_Int_Int_Int3) : [(lizzieLet6_7QNode_Int,Pointer_CTkron_kron_Int_Int_Int),
                                            (lizzieLet6_5QNode_Int_1,MyDTInt_Bool),
                                            (lizzieLet6_3QNode_Int_1,MyDTInt_Int_Int),
                                            (q1ad7_destruct,Pointer_QTree_Int),
                                            (lizzieLet6_6QNode_Int_1,Pointer_QTree_Int),
                                            (q2ad8_destruct,Pointer_QTree_Int),
                                            (q3ad9_destruct,Pointer_QTree_Int)] > (lizzieLet6_7QNode_Int_1lizzieLet6_5QNode_Int_1lizzieLet6_3QNode_Int_1q1ad7_1lizzieLet6_6QNode_Int_1q2ad8_1q3ad9_1Lcall_kron_kron_Int_Int_Int3,CTkron_kron_Int_Int_Int) */
  assign lizzieLet6_7QNode_Int_1lizzieLet6_5QNode_Int_1lizzieLet6_3QNode_Int_1q1ad7_1lizzieLet6_6QNode_Int_1q2ad8_1q3ad9_1Lcall_kron_kron_Int_Int_Int3_d = Lcall_kron_kron_Int_Int_Int3_dc((& {lizzieLet6_7QNode_Int_d[0],
                                                                                                                                                                                               lizzieLet6_5QNode_Int_1_d[0],
                                                                                                                                                                                               lizzieLet6_3QNode_Int_1_d[0],
                                                                                                                                                                                               q1ad7_destruct_d[0],
                                                                                                                                                                                               lizzieLet6_6QNode_Int_1_d[0],
                                                                                                                                                                                               q2ad8_destruct_d[0],
                                                                                                                                                                                               q3ad9_destruct_d[0]}), lizzieLet6_7QNode_Int_d, lizzieLet6_5QNode_Int_1_d, lizzieLet6_3QNode_Int_1_d, q1ad7_destruct_d, lizzieLet6_6QNode_Int_1_d, q2ad8_destruct_d, q3ad9_destruct_d);
  assign {lizzieLet6_7QNode_Int_r,
          lizzieLet6_5QNode_Int_1_r,
          lizzieLet6_3QNode_Int_1_r,
          q1ad7_destruct_r,
          lizzieLet6_6QNode_Int_1_r,
          q2ad8_destruct_r,
          q3ad9_destruct_r} = {7 {(lizzieLet6_7QNode_Int_1lizzieLet6_5QNode_Int_1lizzieLet6_3QNode_Int_1q1ad7_1lizzieLet6_6QNode_Int_1q2ad8_1q3ad9_1Lcall_kron_kron_Int_Int_Int3_r && lizzieLet6_7QNode_Int_1lizzieLet6_5QNode_Int_1lizzieLet6_3QNode_Int_1q1ad7_1lizzieLet6_6QNode_Int_1q2ad8_1q3ad9_1Lcall_kron_kron_Int_Int_Int3_d[0])}};
  
  /* buf (Ty CTkron_kron_Int_Int_Int) : (lizzieLet6_7QNode_Int_1lizzieLet6_5QNode_Int_1lizzieLet6_3QNode_Int_1q1ad7_1lizzieLet6_6QNode_Int_1q2ad8_1q3ad9_1Lcall_kron_kron_Int_Int_Int3,CTkron_kron_Int_Int_Int) > (lizzieLet8_1_argbuf,CTkron_kron_Int_Int_Int) */
  CTkron_kron_Int_Int_Int_t lizzieLet6_7QNode_Int_1lizzieLet6_5QNode_Int_1lizzieLet6_3QNode_Int_1q1ad7_1lizzieLet6_6QNode_Int_1q2ad8_1q3ad9_1Lcall_kron_kron_Int_Int_Int3_bufchan_d;
  logic lizzieLet6_7QNode_Int_1lizzieLet6_5QNode_Int_1lizzieLet6_3QNode_Int_1q1ad7_1lizzieLet6_6QNode_Int_1q2ad8_1q3ad9_1Lcall_kron_kron_Int_Int_Int3_bufchan_r;
  assign lizzieLet6_7QNode_Int_1lizzieLet6_5QNode_Int_1lizzieLet6_3QNode_Int_1q1ad7_1lizzieLet6_6QNode_Int_1q2ad8_1q3ad9_1Lcall_kron_kron_Int_Int_Int3_r = ((! lizzieLet6_7QNode_Int_1lizzieLet6_5QNode_Int_1lizzieLet6_3QNode_Int_1q1ad7_1lizzieLet6_6QNode_Int_1q2ad8_1q3ad9_1Lcall_kron_kron_Int_Int_Int3_bufchan_d[0]) || lizzieLet6_7QNode_Int_1lizzieLet6_5QNode_Int_1lizzieLet6_3QNode_Int_1q1ad7_1lizzieLet6_6QNode_Int_1q2ad8_1q3ad9_1Lcall_kron_kron_Int_Int_Int3_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_7QNode_Int_1lizzieLet6_5QNode_Int_1lizzieLet6_3QNode_Int_1q1ad7_1lizzieLet6_6QNode_Int_1q2ad8_1q3ad9_1Lcall_kron_kron_Int_Int_Int3_bufchan_d <= {83'd0,
                                                                                                                                                                  1'd0};
    else
      if (lizzieLet6_7QNode_Int_1lizzieLet6_5QNode_Int_1lizzieLet6_3QNode_Int_1q1ad7_1lizzieLet6_6QNode_Int_1q2ad8_1q3ad9_1Lcall_kron_kron_Int_Int_Int3_r)
        lizzieLet6_7QNode_Int_1lizzieLet6_5QNode_Int_1lizzieLet6_3QNode_Int_1q1ad7_1lizzieLet6_6QNode_Int_1q2ad8_1q3ad9_1Lcall_kron_kron_Int_Int_Int3_bufchan_d <= lizzieLet6_7QNode_Int_1lizzieLet6_5QNode_Int_1lizzieLet6_3QNode_Int_1q1ad7_1lizzieLet6_6QNode_Int_1q2ad8_1q3ad9_1Lcall_kron_kron_Int_Int_Int3_d;
  CTkron_kron_Int_Int_Int_t lizzieLet6_7QNode_Int_1lizzieLet6_5QNode_Int_1lizzieLet6_3QNode_Int_1q1ad7_1lizzieLet6_6QNode_Int_1q2ad8_1q3ad9_1Lcall_kron_kron_Int_Int_Int3_bufchan_buf;
  assign lizzieLet6_7QNode_Int_1lizzieLet6_5QNode_Int_1lizzieLet6_3QNode_Int_1q1ad7_1lizzieLet6_6QNode_Int_1q2ad8_1q3ad9_1Lcall_kron_kron_Int_Int_Int3_bufchan_r = (! lizzieLet6_7QNode_Int_1lizzieLet6_5QNode_Int_1lizzieLet6_3QNode_Int_1q1ad7_1lizzieLet6_6QNode_Int_1q2ad8_1q3ad9_1Lcall_kron_kron_Int_Int_Int3_bufchan_buf[0]);
  assign lizzieLet8_1_argbuf_d = (lizzieLet6_7QNode_Int_1lizzieLet6_5QNode_Int_1lizzieLet6_3QNode_Int_1q1ad7_1lizzieLet6_6QNode_Int_1q2ad8_1q3ad9_1Lcall_kron_kron_Int_Int_Int3_bufchan_buf[0] ? lizzieLet6_7QNode_Int_1lizzieLet6_5QNode_Int_1lizzieLet6_3QNode_Int_1q1ad7_1lizzieLet6_6QNode_Int_1q2ad8_1q3ad9_1Lcall_kron_kron_Int_Int_Int3_bufchan_buf :
                                  lizzieLet6_7QNode_Int_1lizzieLet6_5QNode_Int_1lizzieLet6_3QNode_Int_1q1ad7_1lizzieLet6_6QNode_Int_1q2ad8_1q3ad9_1Lcall_kron_kron_Int_Int_Int3_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_7QNode_Int_1lizzieLet6_5QNode_Int_1lizzieLet6_3QNode_Int_1q1ad7_1lizzieLet6_6QNode_Int_1q2ad8_1q3ad9_1Lcall_kron_kron_Int_Int_Int3_bufchan_buf <= {83'd0,
                                                                                                                                                                    1'd0};
    else
      if ((lizzieLet8_1_argbuf_r && lizzieLet6_7QNode_Int_1lizzieLet6_5QNode_Int_1lizzieLet6_3QNode_Int_1q1ad7_1lizzieLet6_6QNode_Int_1q2ad8_1q3ad9_1Lcall_kron_kron_Int_Int_Int3_bufchan_buf[0]))
        lizzieLet6_7QNode_Int_1lizzieLet6_5QNode_Int_1lizzieLet6_3QNode_Int_1q1ad7_1lizzieLet6_6QNode_Int_1q2ad8_1q3ad9_1Lcall_kron_kron_Int_Int_Int3_bufchan_buf <= {83'd0,
                                                                                                                                                                      1'd0};
      else if (((! lizzieLet8_1_argbuf_r) && (! lizzieLet6_7QNode_Int_1lizzieLet6_5QNode_Int_1lizzieLet6_3QNode_Int_1q1ad7_1lizzieLet6_6QNode_Int_1q2ad8_1q3ad9_1Lcall_kron_kron_Int_Int_Int3_bufchan_buf[0])))
        lizzieLet6_7QNode_Int_1lizzieLet6_5QNode_Int_1lizzieLet6_3QNode_Int_1q1ad7_1lizzieLet6_6QNode_Int_1q2ad8_1q3ad9_1Lcall_kron_kron_Int_Int_Int3_bufchan_buf <= lizzieLet6_7QNode_Int_1lizzieLet6_5QNode_Int_1lizzieLet6_3QNode_Int_1q1ad7_1lizzieLet6_6QNode_Int_1q2ad8_1q3ad9_1Lcall_kron_kron_Int_Int_Int3_bufchan_d;
  
  /* buf (Ty Pointer_CTkron_kron_Int_Int_Int) : (lizzieLet6_7QNone_Int,Pointer_CTkron_kron_Int_Int_Int) > (lizzieLet6_7QNone_Int_1_argbuf,Pointer_CTkron_kron_Int_Int_Int) */
  Pointer_CTkron_kron_Int_Int_Int_t lizzieLet6_7QNone_Int_bufchan_d;
  logic lizzieLet6_7QNone_Int_bufchan_r;
  assign lizzieLet6_7QNone_Int_r = ((! lizzieLet6_7QNone_Int_bufchan_d[0]) || lizzieLet6_7QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_7QNone_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet6_7QNone_Int_r)
        lizzieLet6_7QNone_Int_bufchan_d <= lizzieLet6_7QNone_Int_d;
  Pointer_CTkron_kron_Int_Int_Int_t lizzieLet6_7QNone_Int_bufchan_buf;
  assign lizzieLet6_7QNone_Int_bufchan_r = (! lizzieLet6_7QNone_Int_bufchan_buf[0]);
  assign lizzieLet6_7QNone_Int_1_argbuf_d = (lizzieLet6_7QNone_Int_bufchan_buf[0] ? lizzieLet6_7QNone_Int_bufchan_buf :
                                             lizzieLet6_7QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_7QNone_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet6_7QNone_Int_1_argbuf_r && lizzieLet6_7QNone_Int_bufchan_buf[0]))
        lizzieLet6_7QNone_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet6_7QNone_Int_1_argbuf_r) && (! lizzieLet6_7QNone_Int_bufchan_buf[0])))
        lizzieLet6_7QNone_Int_bufchan_buf <= lizzieLet6_7QNone_Int_bufchan_d;
  
  /* buf (Ty Pointer_CTkron_kron_Int_Int_Int) : (lizzieLet6_7QVal_Int,Pointer_CTkron_kron_Int_Int_Int) > (lizzieLet6_7QVal_Int_1_argbuf,Pointer_CTkron_kron_Int_Int_Int) */
  Pointer_CTkron_kron_Int_Int_Int_t lizzieLet6_7QVal_Int_bufchan_d;
  logic lizzieLet6_7QVal_Int_bufchan_r;
  assign lizzieLet6_7QVal_Int_r = ((! lizzieLet6_7QVal_Int_bufchan_d[0]) || lizzieLet6_7QVal_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_7QVal_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet6_7QVal_Int_r)
        lizzieLet6_7QVal_Int_bufchan_d <= lizzieLet6_7QVal_Int_d;
  Pointer_CTkron_kron_Int_Int_Int_t lizzieLet6_7QVal_Int_bufchan_buf;
  assign lizzieLet6_7QVal_Int_bufchan_r = (! lizzieLet6_7QVal_Int_bufchan_buf[0]);
  assign lizzieLet6_7QVal_Int_1_argbuf_d = (lizzieLet6_7QVal_Int_bufchan_buf[0] ? lizzieLet6_7QVal_Int_bufchan_buf :
                                            lizzieLet6_7QVal_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_7QVal_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet6_7QVal_Int_1_argbuf_r && lizzieLet6_7QVal_Int_bufchan_buf[0]))
        lizzieLet6_7QVal_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet6_7QVal_Int_1_argbuf_r) && (! lizzieLet6_7QVal_Int_bufchan_buf[0])))
        lizzieLet6_7QVal_Int_bufchan_buf <= lizzieLet6_7QVal_Int_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (m1ad4_goMux_mux,Pointer_QTree_Int) > (m1ad4_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t m1ad4_goMux_mux_bufchan_d;
  logic m1ad4_goMux_mux_bufchan_r;
  assign m1ad4_goMux_mux_r = ((! m1ad4_goMux_mux_bufchan_d[0]) || m1ad4_goMux_mux_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m1ad4_goMux_mux_bufchan_d <= {16'd0, 1'd0};
    else
      if (m1ad4_goMux_mux_r)
        m1ad4_goMux_mux_bufchan_d <= m1ad4_goMux_mux_d;
  Pointer_QTree_Int_t m1ad4_goMux_mux_bufchan_buf;
  assign m1ad4_goMux_mux_bufchan_r = (! m1ad4_goMux_mux_bufchan_buf[0]);
  assign m1ad4_1_argbuf_d = (m1ad4_goMux_mux_bufchan_buf[0] ? m1ad4_goMux_mux_bufchan_buf :
                             m1ad4_goMux_mux_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m1ad4_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((m1ad4_1_argbuf_r && m1ad4_goMux_mux_bufchan_buf[0]))
        m1ad4_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
      else if (((! m1ad4_1_argbuf_r) && (! m1ad4_goMux_mux_bufchan_buf[0])))
        m1ad4_goMux_mux_bufchan_buf <= m1ad4_goMux_mux_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (m2ad5_2_2,Pointer_QTree_Int) > (m2ad5_2_2_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t m2ad5_2_2_bufchan_d;
  logic m2ad5_2_2_bufchan_r;
  assign m2ad5_2_2_r = ((! m2ad5_2_2_bufchan_d[0]) || m2ad5_2_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m2ad5_2_2_bufchan_d <= {16'd0, 1'd0};
    else if (m2ad5_2_2_r) m2ad5_2_2_bufchan_d <= m2ad5_2_2_d;
  Pointer_QTree_Int_t m2ad5_2_2_bufchan_buf;
  assign m2ad5_2_2_bufchan_r = (! m2ad5_2_2_bufchan_buf[0]);
  assign m2ad5_2_2_argbuf_d = (m2ad5_2_2_bufchan_buf[0] ? m2ad5_2_2_bufchan_buf :
                               m2ad5_2_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m2ad5_2_2_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((m2ad5_2_2_argbuf_r && m2ad5_2_2_bufchan_buf[0]))
        m2ad5_2_2_bufchan_buf <= {16'd0, 1'd0};
      else if (((! m2ad5_2_2_argbuf_r) && (! m2ad5_2_2_bufchan_buf[0])))
        m2ad5_2_2_bufchan_buf <= m2ad5_2_2_bufchan_d;
  
  /* fork (Ty Pointer_QTree_Int) : (m2ad5_2_destruct,Pointer_QTree_Int) > [(m2ad5_2_1,Pointer_QTree_Int),
                                                                      (m2ad5_2_2,Pointer_QTree_Int)] */
  logic [1:0] m2ad5_2_destruct_emitted;
  logic [1:0] m2ad5_2_destruct_done;
  assign m2ad5_2_1_d = {m2ad5_2_destruct_d[16:1],
                        (m2ad5_2_destruct_d[0] && (! m2ad5_2_destruct_emitted[0]))};
  assign m2ad5_2_2_d = {m2ad5_2_destruct_d[16:1],
                        (m2ad5_2_destruct_d[0] && (! m2ad5_2_destruct_emitted[1]))};
  assign m2ad5_2_destruct_done = (m2ad5_2_destruct_emitted | ({m2ad5_2_2_d[0],
                                                               m2ad5_2_1_d[0]} & {m2ad5_2_2_r,
                                                                                  m2ad5_2_1_r}));
  assign m2ad5_2_destruct_r = (& m2ad5_2_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m2ad5_2_destruct_emitted <= 2'd0;
    else
      m2ad5_2_destruct_emitted <= (m2ad5_2_destruct_r ? 2'd0 :
                                   m2ad5_2_destruct_done);
  
  /* buf (Ty Pointer_QTree_Int) : (m2ad5_3_2,Pointer_QTree_Int) > (m2ad5_3_2_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t m2ad5_3_2_bufchan_d;
  logic m2ad5_3_2_bufchan_r;
  assign m2ad5_3_2_r = ((! m2ad5_3_2_bufchan_d[0]) || m2ad5_3_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m2ad5_3_2_bufchan_d <= {16'd0, 1'd0};
    else if (m2ad5_3_2_r) m2ad5_3_2_bufchan_d <= m2ad5_3_2_d;
  Pointer_QTree_Int_t m2ad5_3_2_bufchan_buf;
  assign m2ad5_3_2_bufchan_r = (! m2ad5_3_2_bufchan_buf[0]);
  assign m2ad5_3_2_argbuf_d = (m2ad5_3_2_bufchan_buf[0] ? m2ad5_3_2_bufchan_buf :
                               m2ad5_3_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m2ad5_3_2_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((m2ad5_3_2_argbuf_r && m2ad5_3_2_bufchan_buf[0]))
        m2ad5_3_2_bufchan_buf <= {16'd0, 1'd0};
      else if (((! m2ad5_3_2_argbuf_r) && (! m2ad5_3_2_bufchan_buf[0])))
        m2ad5_3_2_bufchan_buf <= m2ad5_3_2_bufchan_d;
  
  /* fork (Ty Pointer_QTree_Int) : (m2ad5_3_destruct,Pointer_QTree_Int) > [(m2ad5_3_1,Pointer_QTree_Int),
                                                                      (m2ad5_3_2,Pointer_QTree_Int)] */
  logic [1:0] m2ad5_3_destruct_emitted;
  logic [1:0] m2ad5_3_destruct_done;
  assign m2ad5_3_1_d = {m2ad5_3_destruct_d[16:1],
                        (m2ad5_3_destruct_d[0] && (! m2ad5_3_destruct_emitted[0]))};
  assign m2ad5_3_2_d = {m2ad5_3_destruct_d[16:1],
                        (m2ad5_3_destruct_d[0] && (! m2ad5_3_destruct_emitted[1]))};
  assign m2ad5_3_destruct_done = (m2ad5_3_destruct_emitted | ({m2ad5_3_2_d[0],
                                                               m2ad5_3_1_d[0]} & {m2ad5_3_2_r,
                                                                                  m2ad5_3_1_r}));
  assign m2ad5_3_destruct_r = (& m2ad5_3_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m2ad5_3_destruct_emitted <= 2'd0;
    else
      m2ad5_3_destruct_emitted <= (m2ad5_3_destruct_r ? 2'd0 :
                                   m2ad5_3_destruct_done);
  
  /* buf (Ty Pointer_QTree_Int) : (m2ad5_4_destruct,Pointer_QTree_Int) > (m2ad5_4_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t m2ad5_4_destruct_bufchan_d;
  logic m2ad5_4_destruct_bufchan_r;
  assign m2ad5_4_destruct_r = ((! m2ad5_4_destruct_bufchan_d[0]) || m2ad5_4_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m2ad5_4_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (m2ad5_4_destruct_r)
        m2ad5_4_destruct_bufchan_d <= m2ad5_4_destruct_d;
  Pointer_QTree_Int_t m2ad5_4_destruct_bufchan_buf;
  assign m2ad5_4_destruct_bufchan_r = (! m2ad5_4_destruct_bufchan_buf[0]);
  assign m2ad5_4_1_argbuf_d = (m2ad5_4_destruct_bufchan_buf[0] ? m2ad5_4_destruct_bufchan_buf :
                               m2ad5_4_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m2ad5_4_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((m2ad5_4_1_argbuf_r && m2ad5_4_destruct_bufchan_buf[0]))
        m2ad5_4_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! m2ad5_4_1_argbuf_r) && (! m2ad5_4_destruct_bufchan_buf[0])))
        m2ad5_4_destruct_bufchan_buf <= m2ad5_4_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (macN_goMux_mux,Pointer_QTree_Int) > (macN_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t macN_goMux_mux_bufchan_d;
  logic macN_goMux_mux_bufchan_r;
  assign macN_goMux_mux_r = ((! macN_goMux_mux_bufchan_d[0]) || macN_goMux_mux_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) macN_goMux_mux_bufchan_d <= {16'd0, 1'd0};
    else
      if (macN_goMux_mux_r) macN_goMux_mux_bufchan_d <= macN_goMux_mux_d;
  Pointer_QTree_Int_t macN_goMux_mux_bufchan_buf;
  assign macN_goMux_mux_bufchan_r = (! macN_goMux_mux_bufchan_buf[0]);
  assign macN_1_argbuf_d = (macN_goMux_mux_bufchan_buf[0] ? macN_goMux_mux_bufchan_buf :
                            macN_goMux_mux_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) macN_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((macN_1_argbuf_r && macN_goMux_mux_bufchan_buf[0]))
        macN_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
      else if (((! macN_1_argbuf_r) && (! macN_goMux_mux_bufchan_buf[0])))
        macN_goMux_mux_bufchan_buf <= macN_goMux_mux_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (macW_goMux_mux,Pointer_QTree_Int) > (macW_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t macW_goMux_mux_bufchan_d;
  logic macW_goMux_mux_bufchan_r;
  assign macW_goMux_mux_r = ((! macW_goMux_mux_bufchan_d[0]) || macW_goMux_mux_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) macW_goMux_mux_bufchan_d <= {16'd0, 1'd0};
    else
      if (macW_goMux_mux_r) macW_goMux_mux_bufchan_d <= macW_goMux_mux_d;
  Pointer_QTree_Int_t macW_goMux_mux_bufchan_buf;
  assign macW_goMux_mux_bufchan_r = (! macW_goMux_mux_bufchan_buf[0]);
  assign macW_1_argbuf_d = (macW_goMux_mux_bufchan_buf[0] ? macW_goMux_mux_bufchan_buf :
                            macW_goMux_mux_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) macW_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((macW_1_argbuf_r && macW_goMux_mux_bufchan_buf[0]))
        macW_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
      else if (((! macW_1_argbuf_r) && (! macW_goMux_mux_bufchan_buf[0])))
        macW_goMux_mux_bufchan_buf <= macW_goMux_mux_bufchan_d;
  
  /* destruct (Ty TupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int,
          Dcon TupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int) : (main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int_1,TupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int) > [(main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Intgo_16,Go),
                                                                                                                                                                                                               (main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_IntisZacL_1,MyDTInt_Bool),
                                                                                                                                                                                                               (main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_IntgacM_1,MyDTInt_Int),
                                                                                                                                                                                                               (main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_IntmacN_1,Pointer_QTree_Int)] */
  logic [3:0] \main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int_1_emitted ;
  logic [3:0] \main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int_1_done ;
  assign \main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Intgo_16_d  = (\main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int_1_d [0] && (! \main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int_1_emitted [0]));
  assign \main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_IntisZacL_1_d  = (\main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int_1_d [0] && (! \main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int_1_emitted [1]));
  assign \main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_IntgacM_1_d  = (\main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int_1_d [0] && (! \main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int_1_emitted [2]));
  assign \main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_IntmacN_1_d  = {\main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int_1_d [16:1],
                                                                                              (\main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int_1_d [0] && (! \main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int_1_emitted [3]))};
  assign \main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int_1_done  = (\main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int_1_emitted  | ({\main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_IntmacN_1_d [0],
                                                                                                                                                                                     \main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_IntgacM_1_d [0],
                                                                                                                                                                                     \main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_IntisZacL_1_d [0],
                                                                                                                                                                                     \main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Intgo_16_d [0]} & {\main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_IntmacN_1_r ,
                                                                                                                                                                                                                                                                             \main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_IntgacM_1_r ,
                                                                                                                                                                                                                                                                             \main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_IntisZacL_1_r ,
                                                                                                                                                                                                                                                                             \main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Intgo_16_r }));
  assign \main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int_1_r  = (& \main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int_1_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int_1_emitted  <= 4'd0;
    else
      \main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int_1_emitted  <= (\main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int_1_r  ? 4'd0 :
                                                                                              \main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Int_1_done );
  
  /* buf (Ty MyDTInt_Int) : (main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_IntgacM_1,MyDTInt_Int) > (gacM_1_1_argbuf,MyDTInt_Int) */
  MyDTInt_Int_t \main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_IntgacM_1_bufchan_d ;
  logic \main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_IntgacM_1_bufchan_r ;
  assign \main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_IntgacM_1_r  = ((! \main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_IntgacM_1_bufchan_d [0]) || \main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_IntgacM_1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_IntgacM_1_bufchan_d  <= 1'd0;
    else
      if (\main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_IntgacM_1_r )
        \main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_IntgacM_1_bufchan_d  <= \main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_IntgacM_1_d ;
  MyDTInt_Int_t \main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_IntgacM_1_bufchan_buf ;
  assign \main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_IntgacM_1_bufchan_r  = (! \main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_IntgacM_1_bufchan_buf [0]);
  assign gacM_1_1_argbuf_d = (\main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_IntgacM_1_bufchan_buf [0] ? \main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_IntgacM_1_bufchan_buf  :
                              \main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_IntgacM_1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_IntgacM_1_bufchan_buf  <= 1'd0;
    else
      if ((gacM_1_1_argbuf_r && \main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_IntgacM_1_bufchan_buf [0]))
        \main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_IntgacM_1_bufchan_buf  <= 1'd0;
      else if (((! gacM_1_1_argbuf_r) && (! \main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_IntgacM_1_bufchan_buf [0])))
        \main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_IntgacM_1_bufchan_buf  <= \main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_IntgacM_1_bufchan_d ;
  
  /* fork (Ty Go) : (main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Intgo_16,Go) > [(go_16_1,Go),
                                                                                                    (go_16_2,Go)] */
  logic [1:0] \main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Intgo_16_emitted ;
  logic [1:0] \main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Intgo_16_done ;
  assign go_16_1_d = (\main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Intgo_16_d [0] && (! \main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Intgo_16_emitted [0]));
  assign go_16_2_d = (\main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Intgo_16_d [0] && (! \main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Intgo_16_emitted [1]));
  assign \main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Intgo_16_done  = (\main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Intgo_16_emitted  | ({go_16_2_d[0],
                                                                                                                                                                                           go_16_1_d[0]} & {go_16_2_r,
                                                                                                                                                                                                            go_16_1_r}));
  assign \main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Intgo_16_r  = (& \main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Intgo_16_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Intgo_16_emitted  <= 2'd0;
    else
      \main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Intgo_16_emitted  <= (\main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Intgo_16_r  ? 2'd0 :
                                                                                                 \main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_Intgo_16_done );
  
  /* buf (Ty MyDTInt_Bool) : (main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_IntisZacL_1,MyDTInt_Bool) > (isZacL_1_1_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t \main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_IntisZacL_1_bufchan_d ;
  logic \main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_IntisZacL_1_bufchan_r ;
  assign \main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_IntisZacL_1_r  = ((! \main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_IntisZacL_1_bufchan_d [0]) || \main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_IntisZacL_1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_IntisZacL_1_bufchan_d  <= 1'd0;
    else
      if (\main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_IntisZacL_1_r )
        \main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_IntisZacL_1_bufchan_d  <= \main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_IntisZacL_1_d ;
  MyDTInt_Bool_t \main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_IntisZacL_1_bufchan_buf ;
  assign \main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_IntisZacL_1_bufchan_r  = (! \main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_IntisZacL_1_bufchan_buf [0]);
  assign isZacL_1_1_argbuf_d = (\main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_IntisZacL_1_bufchan_buf [0] ? \main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_IntisZacL_1_bufchan_buf  :
                                \main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_IntisZacL_1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_IntisZacL_1_bufchan_buf  <= 1'd0;
    else
      if ((isZacL_1_1_argbuf_r && \main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_IntisZacL_1_bufchan_buf [0]))
        \main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_IntisZacL_1_bufchan_buf  <= 1'd0;
      else if (((! isZacL_1_1_argbuf_r) && (! \main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_IntisZacL_1_bufchan_buf [0])))
        \main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_IntisZacL_1_bufchan_buf  <= \main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_IntisZacL_1_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Int) : (main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_IntmacN_1,Pointer_QTree_Int) > (macN_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t \main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_IntmacN_1_bufchan_d ;
  logic \main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_IntmacN_1_bufchan_r ;
  assign \main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_IntmacN_1_r  = ((! \main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_IntmacN_1_bufchan_d [0]) || \main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_IntmacN_1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_IntmacN_1_bufchan_d  <= {16'd0,
                                                                                                    1'd0};
    else
      if (\main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_IntmacN_1_r )
        \main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_IntmacN_1_bufchan_d  <= \main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_IntmacN_1_d ;
  Pointer_QTree_Int_t \main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_IntmacN_1_bufchan_buf ;
  assign \main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_IntmacN_1_bufchan_r  = (! \main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_IntmacN_1_bufchan_buf [0]);
  assign macN_1_1_argbuf_d = (\main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_IntmacN_1_bufchan_buf [0] ? \main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_IntmacN_1_bufchan_buf  :
                              \main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_IntmacN_1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_IntmacN_1_bufchan_buf  <= {16'd0,
                                                                                                      1'd0};
    else
      if ((macN_1_1_argbuf_r && \main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_IntmacN_1_bufchan_buf [0]))
        \main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_IntmacN_1_bufchan_buf  <= {16'd0,
                                                                                                        1'd0};
      else if (((! macN_1_1_argbuf_r) && (! \main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_IntmacN_1_bufchan_buf [0])))
        \main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_IntmacN_1_bufchan_buf  <= \main_map'_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int___Pointer_QTree_IntmacN_1_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Int) : (main_map'_Int_Int_resbuf,Pointer_QTree_Int) > (es_0_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t \main_map'_Int_Int_resbuf_bufchan_d ;
  logic \main_map'_Int_Int_resbuf_bufchan_r ;
  assign \main_map'_Int_Int_resbuf_r  = ((! \main_map'_Int_Int_resbuf_bufchan_d [0]) || \main_map'_Int_Int_resbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \main_map'_Int_Int_resbuf_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\main_map'_Int_Int_resbuf_r )
        \main_map'_Int_Int_resbuf_bufchan_d  <= \main_map'_Int_Int_resbuf_d ;
  Pointer_QTree_Int_t \main_map'_Int_Int_resbuf_bufchan_buf ;
  assign \main_map'_Int_Int_resbuf_bufchan_r  = (! \main_map'_Int_Int_resbuf_bufchan_buf [0]);
  assign es_0_1_1_argbuf_d = (\main_map'_Int_Int_resbuf_bufchan_buf [0] ? \main_map'_Int_Int_resbuf_bufchan_buf  :
                              \main_map'_Int_Int_resbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \main_map'_Int_Int_resbuf_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((es_0_1_1_argbuf_r && \main_map'_Int_Int_resbuf_bufchan_buf [0]))
        \main_map'_Int_Int_resbuf_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! es_0_1_1_argbuf_r) && (! \main_map'_Int_Int_resbuf_bufchan_buf [0])))
        \main_map'_Int_Int_resbuf_bufchan_buf  <= \main_map'_Int_Int_resbuf_bufchan_d ;
  
  /* destruct (Ty TupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int,
          Dcon TupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int) : (map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int_1,TupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int) > [(map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Intgo_17,Go),
                                                                                                                                                                                                                                                   (map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntisZacT_1,MyDTInt_Bool),
                                                                                                                                                                                                                                                   (map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntgacU_1,MyDTInt_Int_Int),
                                                                                                                                                                                                                                                   (map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Intv'acV_1,Int),
                                                                                                                                                                                                                                                   (map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntmacW_1,Pointer_QTree_Int)] */
  logic [4:0] \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int_1_emitted ;
  logic [4:0] \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int_1_done ;
  assign \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Intgo_17_d  = (\map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int_1_d [0] && (! \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int_1_emitted [0]));
  assign \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntisZacT_1_d  = (\map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int_1_d [0] && (! \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int_1_emitted [1]));
  assign \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntgacU_1_d  = (\map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int_1_d [0] && (! \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int_1_emitted [2]));
  assign \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Intv'acV_1_d  = {\map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int_1_d [32:1],
                                                                                                               (\map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int_1_d [0] && (! \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int_1_emitted [3]))};
  assign \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntmacW_1_d  = {\map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int_1_d [48:33],
                                                                                                              (\map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int_1_d [0] && (! \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int_1_emitted [4]))};
  assign \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int_1_done  = (\map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int_1_emitted  | ({\map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntmacW_1_d [0],
                                                                                                                                                                                                                     \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Intv'acV_1_d [0],
                                                                                                                                                                                                                     \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntgacU_1_d [0],
                                                                                                                                                                                                                     \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntisZacT_1_d [0],
                                                                                                                                                                                                                     \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Intgo_17_d [0]} & {\map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntmacW_1_r ,
                                                                                                                                                                                                                                                                                                                             \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Intv'acV_1_r ,
                                                                                                                                                                                                                                                                                                                             \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntgacU_1_r ,
                                                                                                                                                                                                                                                                                                                             \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntisZacT_1_r ,
                                                                                                                                                                                                                                                                                                                             \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Intgo_17_r }));
  assign \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int_1_r  = (& \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int_1_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int_1_emitted  <= 5'd0;
    else
      \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int_1_emitted  <= (\map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int_1_r  ? 5'd0 :
                                                                                                              \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int_1_done );
  
  /* buf (Ty MyDTInt_Int_Int) : (map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntgacU_1,MyDTInt_Int_Int) > (gacU_1_1_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntgacU_1_bufchan_d ;
  logic \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntgacU_1_bufchan_r ;
  assign \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntgacU_1_r  = ((! \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntgacU_1_bufchan_d [0]) || \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntgacU_1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntgacU_1_bufchan_d  <= 1'd0;
    else
      if (\map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntgacU_1_r )
        \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntgacU_1_bufchan_d  <= \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntgacU_1_d ;
  MyDTInt_Int_Int_t \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntgacU_1_bufchan_buf ;
  assign \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntgacU_1_bufchan_r  = (! \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntgacU_1_bufchan_buf [0]);
  assign gacU_1_1_argbuf_d = (\map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntgacU_1_bufchan_buf [0] ? \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntgacU_1_bufchan_buf  :
                              \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntgacU_1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntgacU_1_bufchan_buf  <= 1'd0;
    else
      if ((gacU_1_1_argbuf_r && \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntgacU_1_bufchan_buf [0]))
        \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntgacU_1_bufchan_buf  <= 1'd0;
      else if (((! gacU_1_1_argbuf_r) && (! \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntgacU_1_bufchan_buf [0])))
        \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntgacU_1_bufchan_buf  <= \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntgacU_1_bufchan_d ;
  
  /* fork (Ty Go) : (map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Intgo_17,Go) > [(go_17_1,Go),
                                                                                                                    (go_17_2,Go)] */
  logic [1:0] \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Intgo_17_emitted ;
  logic [1:0] \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Intgo_17_done ;
  assign go_17_1_d = (\map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Intgo_17_d [0] && (! \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Intgo_17_emitted [0]));
  assign go_17_2_d = (\map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Intgo_17_d [0] && (! \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Intgo_17_emitted [1]));
  assign \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Intgo_17_done  = (\map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Intgo_17_emitted  | ({go_17_2_d[0],
                                                                                                                                                                                                                           go_17_1_d[0]} & {go_17_2_r,
                                                                                                                                                                                                                                            go_17_1_r}));
  assign \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Intgo_17_r  = (& \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Intgo_17_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Intgo_17_emitted  <= 2'd0;
    else
      \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Intgo_17_emitted  <= (\map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Intgo_17_r  ? 2'd0 :
                                                                                                                 \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Intgo_17_done );
  
  /* buf (Ty MyDTInt_Bool) : (map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntisZacT_1,MyDTInt_Bool) > (isZacT_1_1_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntisZacT_1_bufchan_d ;
  logic \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntisZacT_1_bufchan_r ;
  assign \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntisZacT_1_r  = ((! \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntisZacT_1_bufchan_d [0]) || \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntisZacT_1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntisZacT_1_bufchan_d  <= 1'd0;
    else
      if (\map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntisZacT_1_r )
        \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntisZacT_1_bufchan_d  <= \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntisZacT_1_d ;
  MyDTInt_Bool_t \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntisZacT_1_bufchan_buf ;
  assign \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntisZacT_1_bufchan_r  = (! \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntisZacT_1_bufchan_buf [0]);
  assign isZacT_1_1_argbuf_d = (\map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntisZacT_1_bufchan_buf [0] ? \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntisZacT_1_bufchan_buf  :
                                \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntisZacT_1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntisZacT_1_bufchan_buf  <= 1'd0;
    else
      if ((isZacT_1_1_argbuf_r && \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntisZacT_1_bufchan_buf [0]))
        \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntisZacT_1_bufchan_buf  <= 1'd0;
      else if (((! isZacT_1_1_argbuf_r) && (! \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntisZacT_1_bufchan_buf [0])))
        \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntisZacT_1_bufchan_buf  <= \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntisZacT_1_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Int) : (map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntmacW_1,Pointer_QTree_Int) > (macW_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntmacW_1_bufchan_d ;
  logic \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntmacW_1_bufchan_r ;
  assign \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntmacW_1_r  = ((! \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntmacW_1_bufchan_d [0]) || \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntmacW_1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntmacW_1_bufchan_d  <= {16'd0,
                                                                                                                    1'd0};
    else
      if (\map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntmacW_1_r )
        \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntmacW_1_bufchan_d  <= \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntmacW_1_d ;
  Pointer_QTree_Int_t \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntmacW_1_bufchan_buf ;
  assign \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntmacW_1_bufchan_r  = (! \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntmacW_1_bufchan_buf [0]);
  assign macW_1_1_argbuf_d = (\map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntmacW_1_bufchan_buf [0] ? \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntmacW_1_bufchan_buf  :
                              \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntmacW_1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntmacW_1_bufchan_buf  <= {16'd0,
                                                                                                                      1'd0};
    else
      if ((macW_1_1_argbuf_r && \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntmacW_1_bufchan_buf [0]))
        \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntmacW_1_bufchan_buf  <= {16'd0,
                                                                                                                        1'd0};
      else if (((! macW_1_1_argbuf_r) && (! \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntmacW_1_bufchan_buf [0])))
        \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntmacW_1_bufchan_buf  <= \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntmacW_1_bufchan_d ;
  
  /* buf (Ty Int) : (map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Intv'acV_1,Int) > (v'acV_1_1_argbuf,Int) */
  Int_t \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Intv'acV_1_bufchan_d ;
  logic \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Intv'acV_1_bufchan_r ;
  assign \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Intv'acV_1_r  = ((! \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Intv'acV_1_bufchan_d [0]) || \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Intv'acV_1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Intv'acV_1_bufchan_d  <= {32'd0,
                                                                                                                     1'd0};
    else
      if (\map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Intv'acV_1_r )
        \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Intv'acV_1_bufchan_d  <= \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Intv'acV_1_d ;
  Int_t \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Intv'acV_1_bufchan_buf ;
  assign \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Intv'acV_1_bufchan_r  = (! \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Intv'acV_1_bufchan_buf [0]);
  assign \v'acV_1_1_argbuf_d  = (\map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Intv'acV_1_bufchan_buf [0] ? \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Intv'acV_1_bufchan_buf  :
                                 \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Intv'acV_1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Intv'acV_1_bufchan_buf  <= {32'd0,
                                                                                                                       1'd0};
    else
      if ((\v'acV_1_1_argbuf_r  && \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Intv'acV_1_bufchan_buf [0]))
        \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Intv'acV_1_bufchan_buf  <= {32'd0,
                                                                                                                         1'd0};
      else if (((! \v'acV_1_1_argbuf_r ) && (! \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Intv'acV_1_bufchan_buf [0])))
        \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Intv'acV_1_bufchan_buf  <= \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Intv'acV_1_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Int) : (map''_map''_Int_Int_Int_resbuf,Pointer_QTree_Int) > (lizzieLet12_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t \map''_map''_Int_Int_Int_resbuf_bufchan_d ;
  logic \map''_map''_Int_Int_Int_resbuf_bufchan_r ;
  assign \map''_map''_Int_Int_Int_resbuf_r  = ((! \map''_map''_Int_Int_Int_resbuf_bufchan_d [0]) || \map''_map''_Int_Int_Int_resbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \map''_map''_Int_Int_Int_resbuf_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\map''_map''_Int_Int_Int_resbuf_r )
        \map''_map''_Int_Int_Int_resbuf_bufchan_d  <= \map''_map''_Int_Int_Int_resbuf_d ;
  Pointer_QTree_Int_t \map''_map''_Int_Int_Int_resbuf_bufchan_buf ;
  assign \map''_map''_Int_Int_Int_resbuf_bufchan_r  = (! \map''_map''_Int_Int_Int_resbuf_bufchan_buf [0]);
  assign lizzieLet12_1_argbuf_d = (\map''_map''_Int_Int_Int_resbuf_bufchan_buf [0] ? \map''_map''_Int_Int_Int_resbuf_bufchan_buf  :
                                   \map''_map''_Int_Int_Int_resbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \map''_map''_Int_Int_Int_resbuf_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((lizzieLet12_1_argbuf_r && \map''_map''_Int_Int_Int_resbuf_bufchan_buf [0]))
        \map''_map''_Int_Int_Int_resbuf_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! lizzieLet12_1_argbuf_r) && (! \map''_map''_Int_Int_Int_resbuf_bufchan_buf [0])))
        \map''_map''_Int_Int_Int_resbuf_bufchan_buf  <= \map''_map''_Int_Int_Int_resbuf_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Int) : (q1ac0_destruct,Pointer_QTree_Int) > (q1ac0_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t q1ac0_destruct_bufchan_d;
  logic q1ac0_destruct_bufchan_r;
  assign q1ac0_destruct_r = ((! q1ac0_destruct_bufchan_d[0]) || q1ac0_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q1ac0_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q1ac0_destruct_r) q1ac0_destruct_bufchan_d <= q1ac0_destruct_d;
  Pointer_QTree_Int_t q1ac0_destruct_bufchan_buf;
  assign q1ac0_destruct_bufchan_r = (! q1ac0_destruct_bufchan_buf[0]);
  assign q1ac0_1_argbuf_d = (q1ac0_destruct_bufchan_buf[0] ? q1ac0_destruct_bufchan_buf :
                             q1ac0_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q1ac0_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q1ac0_1_argbuf_r && q1ac0_destruct_bufchan_buf[0]))
        q1ac0_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q1ac0_1_argbuf_r) && (! q1ac0_destruct_bufchan_buf[0])))
        q1ac0_destruct_bufchan_buf <= q1ac0_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (q1acP_3_destruct,Pointer_QTree_Int) > (q1acP_3_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t q1acP_3_destruct_bufchan_d;
  logic q1acP_3_destruct_bufchan_r;
  assign q1acP_3_destruct_r = ((! q1acP_3_destruct_bufchan_d[0]) || q1acP_3_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q1acP_3_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q1acP_3_destruct_r)
        q1acP_3_destruct_bufchan_d <= q1acP_3_destruct_d;
  Pointer_QTree_Int_t q1acP_3_destruct_bufchan_buf;
  assign q1acP_3_destruct_bufchan_r = (! q1acP_3_destruct_bufchan_buf[0]);
  assign q1acP_3_1_argbuf_d = (q1acP_3_destruct_bufchan_buf[0] ? q1acP_3_destruct_bufchan_buf :
                               q1acP_3_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q1acP_3_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q1acP_3_1_argbuf_r && q1acP_3_destruct_bufchan_buf[0]))
        q1acP_3_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q1acP_3_1_argbuf_r) && (! q1acP_3_destruct_bufchan_buf[0])))
        q1acP_3_destruct_bufchan_buf <= q1acP_3_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (q1acY_3_destruct,Pointer_QTree_Int) > (q1acY_3_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t q1acY_3_destruct_bufchan_d;
  logic q1acY_3_destruct_bufchan_r;
  assign q1acY_3_destruct_r = ((! q1acY_3_destruct_bufchan_d[0]) || q1acY_3_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q1acY_3_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q1acY_3_destruct_r)
        q1acY_3_destruct_bufchan_d <= q1acY_3_destruct_d;
  Pointer_QTree_Int_t q1acY_3_destruct_bufchan_buf;
  assign q1acY_3_destruct_bufchan_r = (! q1acY_3_destruct_bufchan_buf[0]);
  assign q1acY_3_1_argbuf_d = (q1acY_3_destruct_bufchan_buf[0] ? q1acY_3_destruct_bufchan_buf :
                               q1acY_3_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q1acY_3_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q1acY_3_1_argbuf_r && q1acY_3_destruct_bufchan_buf[0]))
        q1acY_3_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q1acY_3_1_argbuf_r) && (! q1acY_3_destruct_bufchan_buf[0])))
        q1acY_3_destruct_bufchan_buf <= q1acY_3_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (q1ad7_3_destruct,Pointer_QTree_Int) > (q1ad7_3_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t q1ad7_3_destruct_bufchan_d;
  logic q1ad7_3_destruct_bufchan_r;
  assign q1ad7_3_destruct_r = ((! q1ad7_3_destruct_bufchan_d[0]) || q1ad7_3_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q1ad7_3_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q1ad7_3_destruct_r)
        q1ad7_3_destruct_bufchan_d <= q1ad7_3_destruct_d;
  Pointer_QTree_Int_t q1ad7_3_destruct_bufchan_buf;
  assign q1ad7_3_destruct_bufchan_r = (! q1ad7_3_destruct_bufchan_buf[0]);
  assign q1ad7_3_1_argbuf_d = (q1ad7_3_destruct_bufchan_buf[0] ? q1ad7_3_destruct_bufchan_buf :
                               q1ad7_3_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q1ad7_3_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q1ad7_3_1_argbuf_r && q1ad7_3_destruct_bufchan_buf[0]))
        q1ad7_3_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q1ad7_3_1_argbuf_r) && (! q1ad7_3_destruct_bufchan_buf[0])))
        q1ad7_3_destruct_bufchan_buf <= q1ad7_3_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (q2ac1_1_destruct,Pointer_QTree_Int) > (q2ac1_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t q2ac1_1_destruct_bufchan_d;
  logic q2ac1_1_destruct_bufchan_r;
  assign q2ac1_1_destruct_r = ((! q2ac1_1_destruct_bufchan_d[0]) || q2ac1_1_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q2ac1_1_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q2ac1_1_destruct_r)
        q2ac1_1_destruct_bufchan_d <= q2ac1_1_destruct_d;
  Pointer_QTree_Int_t q2ac1_1_destruct_bufchan_buf;
  assign q2ac1_1_destruct_bufchan_r = (! q2ac1_1_destruct_bufchan_buf[0]);
  assign q2ac1_1_1_argbuf_d = (q2ac1_1_destruct_bufchan_buf[0] ? q2ac1_1_destruct_bufchan_buf :
                               q2ac1_1_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q2ac1_1_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q2ac1_1_1_argbuf_r && q2ac1_1_destruct_bufchan_buf[0]))
        q2ac1_1_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q2ac1_1_1_argbuf_r) && (! q2ac1_1_destruct_bufchan_buf[0])))
        q2ac1_1_destruct_bufchan_buf <= q2ac1_1_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (q2acQ_2_destruct,Pointer_QTree_Int) > (q2acQ_2_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t q2acQ_2_destruct_bufchan_d;
  logic q2acQ_2_destruct_bufchan_r;
  assign q2acQ_2_destruct_r = ((! q2acQ_2_destruct_bufchan_d[0]) || q2acQ_2_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q2acQ_2_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q2acQ_2_destruct_r)
        q2acQ_2_destruct_bufchan_d <= q2acQ_2_destruct_d;
  Pointer_QTree_Int_t q2acQ_2_destruct_bufchan_buf;
  assign q2acQ_2_destruct_bufchan_r = (! q2acQ_2_destruct_bufchan_buf[0]);
  assign q2acQ_2_1_argbuf_d = (q2acQ_2_destruct_bufchan_buf[0] ? q2acQ_2_destruct_bufchan_buf :
                               q2acQ_2_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q2acQ_2_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q2acQ_2_1_argbuf_r && q2acQ_2_destruct_bufchan_buf[0]))
        q2acQ_2_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q2acQ_2_1_argbuf_r) && (! q2acQ_2_destruct_bufchan_buf[0])))
        q2acQ_2_destruct_bufchan_buf <= q2acQ_2_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (q2acZ_2_destruct,Pointer_QTree_Int) > (q2acZ_2_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t q2acZ_2_destruct_bufchan_d;
  logic q2acZ_2_destruct_bufchan_r;
  assign q2acZ_2_destruct_r = ((! q2acZ_2_destruct_bufchan_d[0]) || q2acZ_2_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q2acZ_2_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q2acZ_2_destruct_r)
        q2acZ_2_destruct_bufchan_d <= q2acZ_2_destruct_d;
  Pointer_QTree_Int_t q2acZ_2_destruct_bufchan_buf;
  assign q2acZ_2_destruct_bufchan_r = (! q2acZ_2_destruct_bufchan_buf[0]);
  assign q2acZ_2_1_argbuf_d = (q2acZ_2_destruct_bufchan_buf[0] ? q2acZ_2_destruct_bufchan_buf :
                               q2acZ_2_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q2acZ_2_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q2acZ_2_1_argbuf_r && q2acZ_2_destruct_bufchan_buf[0]))
        q2acZ_2_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q2acZ_2_1_argbuf_r) && (! q2acZ_2_destruct_bufchan_buf[0])))
        q2acZ_2_destruct_bufchan_buf <= q2acZ_2_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (q2ad8_2_destruct,Pointer_QTree_Int) > (q2ad8_2_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t q2ad8_2_destruct_bufchan_d;
  logic q2ad8_2_destruct_bufchan_r;
  assign q2ad8_2_destruct_r = ((! q2ad8_2_destruct_bufchan_d[0]) || q2ad8_2_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q2ad8_2_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q2ad8_2_destruct_r)
        q2ad8_2_destruct_bufchan_d <= q2ad8_2_destruct_d;
  Pointer_QTree_Int_t q2ad8_2_destruct_bufchan_buf;
  assign q2ad8_2_destruct_bufchan_r = (! q2ad8_2_destruct_bufchan_buf[0]);
  assign q2ad8_2_1_argbuf_d = (q2ad8_2_destruct_bufchan_buf[0] ? q2ad8_2_destruct_bufchan_buf :
                               q2ad8_2_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q2ad8_2_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q2ad8_2_1_argbuf_r && q2ad8_2_destruct_bufchan_buf[0]))
        q2ad8_2_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q2ad8_2_1_argbuf_r) && (! q2ad8_2_destruct_bufchan_buf[0])))
        q2ad8_2_destruct_bufchan_buf <= q2ad8_2_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (q3ac2_2_destruct,Pointer_QTree_Int) > (q3ac2_2_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t q3ac2_2_destruct_bufchan_d;
  logic q3ac2_2_destruct_bufchan_r;
  assign q3ac2_2_destruct_r = ((! q3ac2_2_destruct_bufchan_d[0]) || q3ac2_2_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q3ac2_2_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q3ac2_2_destruct_r)
        q3ac2_2_destruct_bufchan_d <= q3ac2_2_destruct_d;
  Pointer_QTree_Int_t q3ac2_2_destruct_bufchan_buf;
  assign q3ac2_2_destruct_bufchan_r = (! q3ac2_2_destruct_bufchan_buf[0]);
  assign q3ac2_2_1_argbuf_d = (q3ac2_2_destruct_bufchan_buf[0] ? q3ac2_2_destruct_bufchan_buf :
                               q3ac2_2_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q3ac2_2_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q3ac2_2_1_argbuf_r && q3ac2_2_destruct_bufchan_buf[0]))
        q3ac2_2_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q3ac2_2_1_argbuf_r) && (! q3ac2_2_destruct_bufchan_buf[0])))
        q3ac2_2_destruct_bufchan_buf <= q3ac2_2_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (q3acR_1_destruct,Pointer_QTree_Int) > (q3acR_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t q3acR_1_destruct_bufchan_d;
  logic q3acR_1_destruct_bufchan_r;
  assign q3acR_1_destruct_r = ((! q3acR_1_destruct_bufchan_d[0]) || q3acR_1_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q3acR_1_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q3acR_1_destruct_r)
        q3acR_1_destruct_bufchan_d <= q3acR_1_destruct_d;
  Pointer_QTree_Int_t q3acR_1_destruct_bufchan_buf;
  assign q3acR_1_destruct_bufchan_r = (! q3acR_1_destruct_bufchan_buf[0]);
  assign q3acR_1_1_argbuf_d = (q3acR_1_destruct_bufchan_buf[0] ? q3acR_1_destruct_bufchan_buf :
                               q3acR_1_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q3acR_1_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q3acR_1_1_argbuf_r && q3acR_1_destruct_bufchan_buf[0]))
        q3acR_1_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q3acR_1_1_argbuf_r) && (! q3acR_1_destruct_bufchan_buf[0])))
        q3acR_1_destruct_bufchan_buf <= q3acR_1_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (q3ad0_1_destruct,Pointer_QTree_Int) > (q3ad0_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t q3ad0_1_destruct_bufchan_d;
  logic q3ad0_1_destruct_bufchan_r;
  assign q3ad0_1_destruct_r = ((! q3ad0_1_destruct_bufchan_d[0]) || q3ad0_1_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q3ad0_1_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q3ad0_1_destruct_r)
        q3ad0_1_destruct_bufchan_d <= q3ad0_1_destruct_d;
  Pointer_QTree_Int_t q3ad0_1_destruct_bufchan_buf;
  assign q3ad0_1_destruct_bufchan_r = (! q3ad0_1_destruct_bufchan_buf[0]);
  assign q3ad0_1_1_argbuf_d = (q3ad0_1_destruct_bufchan_buf[0] ? q3ad0_1_destruct_bufchan_buf :
                               q3ad0_1_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q3ad0_1_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q3ad0_1_1_argbuf_r && q3ad0_1_destruct_bufchan_buf[0]))
        q3ad0_1_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q3ad0_1_1_argbuf_r) && (! q3ad0_1_destruct_bufchan_buf[0])))
        q3ad0_1_destruct_bufchan_buf <= q3ad0_1_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (q3ad9_1_destruct,Pointer_QTree_Int) > (q3ad9_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t q3ad9_1_destruct_bufchan_d;
  logic q3ad9_1_destruct_bufchan_r;
  assign q3ad9_1_destruct_r = ((! q3ad9_1_destruct_bufchan_d[0]) || q3ad9_1_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q3ad9_1_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q3ad9_1_destruct_r)
        q3ad9_1_destruct_bufchan_d <= q3ad9_1_destruct_d;
  Pointer_QTree_Int_t q3ad9_1_destruct_bufchan_buf;
  assign q3ad9_1_destruct_bufchan_r = (! q3ad9_1_destruct_bufchan_buf[0]);
  assign q3ad9_1_1_argbuf_d = (q3ad9_1_destruct_bufchan_buf[0] ? q3ad9_1_destruct_bufchan_buf :
                               q3ad9_1_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q3ad9_1_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q3ad9_1_1_argbuf_r && q3ad9_1_destruct_bufchan_buf[0]))
        q3ad9_1_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q3ad9_1_1_argbuf_r) && (! q3ad9_1_destruct_bufchan_buf[0])))
        q3ad9_1_destruct_bufchan_buf <= q3ad9_1_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (q4ac3_3_destruct,Pointer_QTree_Int) > (q4ac3_3_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t q4ac3_3_destruct_bufchan_d;
  logic q4ac3_3_destruct_bufchan_r;
  assign q4ac3_3_destruct_r = ((! q4ac3_3_destruct_bufchan_d[0]) || q4ac3_3_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q4ac3_3_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q4ac3_3_destruct_r)
        q4ac3_3_destruct_bufchan_d <= q4ac3_3_destruct_d;
  Pointer_QTree_Int_t q4ac3_3_destruct_bufchan_buf;
  assign q4ac3_3_destruct_bufchan_r = (! q4ac3_3_destruct_bufchan_buf[0]);
  assign q4ac3_3_1_argbuf_d = (q4ac3_3_destruct_bufchan_buf[0] ? q4ac3_3_destruct_bufchan_buf :
                               q4ac3_3_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q4ac3_3_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q4ac3_3_1_argbuf_r && q4ac3_3_destruct_bufchan_buf[0]))
        q4ac3_3_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q4ac3_3_1_argbuf_r) && (! q4ac3_3_destruct_bufchan_buf[0])))
        q4ac3_3_destruct_bufchan_buf <= q4ac3_3_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (q4acS_destruct,Pointer_QTree_Int) > (q4acS_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t q4acS_destruct_bufchan_d;
  logic q4acS_destruct_bufchan_r;
  assign q4acS_destruct_r = ((! q4acS_destruct_bufchan_d[0]) || q4acS_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q4acS_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q4acS_destruct_r) q4acS_destruct_bufchan_d <= q4acS_destruct_d;
  Pointer_QTree_Int_t q4acS_destruct_bufchan_buf;
  assign q4acS_destruct_bufchan_r = (! q4acS_destruct_bufchan_buf[0]);
  assign q4acS_1_argbuf_d = (q4acS_destruct_bufchan_buf[0] ? q4acS_destruct_bufchan_buf :
                             q4acS_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q4acS_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q4acS_1_argbuf_r && q4acS_destruct_bufchan_buf[0]))
        q4acS_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q4acS_1_argbuf_r) && (! q4acS_destruct_bufchan_buf[0])))
        q4acS_destruct_bufchan_buf <= q4acS_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (q4ad1_destruct,Pointer_QTree_Int) > (q4ad1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t q4ad1_destruct_bufchan_d;
  logic q4ad1_destruct_bufchan_r;
  assign q4ad1_destruct_r = ((! q4ad1_destruct_bufchan_d[0]) || q4ad1_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q4ad1_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q4ad1_destruct_r) q4ad1_destruct_bufchan_d <= q4ad1_destruct_d;
  Pointer_QTree_Int_t q4ad1_destruct_bufchan_buf;
  assign q4ad1_destruct_bufchan_r = (! q4ad1_destruct_bufchan_buf[0]);
  assign q4ad1_1_argbuf_d = (q4ad1_destruct_bufchan_buf[0] ? q4ad1_destruct_bufchan_buf :
                             q4ad1_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q4ad1_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q4ad1_1_argbuf_r && q4ad1_destruct_bufchan_buf[0]))
        q4ad1_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q4ad1_1_argbuf_r) && (! q4ad1_destruct_bufchan_buf[0])))
        q4ad1_destruct_bufchan_buf <= q4ad1_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (q4ada_destruct,Pointer_QTree_Int) > (q4ada_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t q4ada_destruct_bufchan_d;
  logic q4ada_destruct_bufchan_r;
  assign q4ada_destruct_r = ((! q4ada_destruct_bufchan_d[0]) || q4ada_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q4ada_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q4ada_destruct_r) q4ada_destruct_bufchan_d <= q4ada_destruct_d;
  Pointer_QTree_Int_t q4ada_destruct_bufchan_buf;
  assign q4ada_destruct_bufchan_r = (! q4ada_destruct_bufchan_buf[0]);
  assign q4ada_1_argbuf_d = (q4ada_destruct_bufchan_buf[0] ? q4ada_destruct_bufchan_buf :
                             q4ada_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q4ada_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q4ada_1_argbuf_r && q4ada_destruct_bufchan_buf[0]))
        q4ada_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q4ada_1_argbuf_r) && (! q4ada_destruct_bufchan_buf[0])))
        q4ada_destruct_bufchan_buf <= q4ada_destruct_bufchan_d;
  
  /* buf (Ty CT$wnnz_Int) : (readPointer_CT$wnnz_Intscfarg_0_1_argbuf,CT$wnnz_Int) > (readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb,CT$wnnz_Int) */
  CT$wnnz_Int_t readPointer_CT$wnnz_Intscfarg_0_1_argbuf_bufchan_d;
  logic readPointer_CT$wnnz_Intscfarg_0_1_argbuf_bufchan_r;
  assign readPointer_CT$wnnz_Intscfarg_0_1_argbuf_r = ((! readPointer_CT$wnnz_Intscfarg_0_1_argbuf_bufchan_d[0]) || readPointer_CT$wnnz_Intscfarg_0_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_CT$wnnz_Intscfarg_0_1_argbuf_bufchan_d <= {115'd0,
                                                             1'd0};
    else
      if (readPointer_CT$wnnz_Intscfarg_0_1_argbuf_r)
        readPointer_CT$wnnz_Intscfarg_0_1_argbuf_bufchan_d <= readPointer_CT$wnnz_Intscfarg_0_1_argbuf_d;
  CT$wnnz_Int_t readPointer_CT$wnnz_Intscfarg_0_1_argbuf_bufchan_buf;
  assign readPointer_CT$wnnz_Intscfarg_0_1_argbuf_bufchan_r = (! readPointer_CT$wnnz_Intscfarg_0_1_argbuf_bufchan_buf[0]);
  assign readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb_d = (readPointer_CT$wnnz_Intscfarg_0_1_argbuf_bufchan_buf[0] ? readPointer_CT$wnnz_Intscfarg_0_1_argbuf_bufchan_buf :
                                                           readPointer_CT$wnnz_Intscfarg_0_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_CT$wnnz_Intscfarg_0_1_argbuf_bufchan_buf <= {115'd0,
                                                               1'd0};
    else
      if ((readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb_r && readPointer_CT$wnnz_Intscfarg_0_1_argbuf_bufchan_buf[0]))
        readPointer_CT$wnnz_Intscfarg_0_1_argbuf_bufchan_buf <= {115'd0,
                                                                 1'd0};
      else if (((! readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb_r) && (! readPointer_CT$wnnz_Intscfarg_0_1_argbuf_bufchan_buf[0])))
        readPointer_CT$wnnz_Intscfarg_0_1_argbuf_bufchan_buf <= readPointer_CT$wnnz_Intscfarg_0_1_argbuf_bufchan_d;
  
  /* fork (Ty CT$wnnz_Int) : (readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb,CT$wnnz_Int) > [(lizzieLet25_1,CT$wnnz_Int),
                                                                                      (lizzieLet25_2,CT$wnnz_Int),
                                                                                      (lizzieLet25_3,CT$wnnz_Int),
                                                                                      (lizzieLet25_4,CT$wnnz_Int)] */
  logic [3:0] readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb_emitted;
  logic [3:0] readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb_done;
  assign lizzieLet25_1_d = {readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb_d[115:1],
                            (readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb_d[0] && (! readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb_emitted[0]))};
  assign lizzieLet25_2_d = {readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb_d[115:1],
                            (readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb_d[0] && (! readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb_emitted[1]))};
  assign lizzieLet25_3_d = {readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb_d[115:1],
                            (readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb_d[0] && (! readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb_emitted[2]))};
  assign lizzieLet25_4_d = {readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb_d[115:1],
                            (readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb_d[0] && (! readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb_emitted[3]))};
  assign readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb_done = (readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb_emitted | ({lizzieLet25_4_d[0],
                                                                                                                       lizzieLet25_3_d[0],
                                                                                                                       lizzieLet25_2_d[0],
                                                                                                                       lizzieLet25_1_d[0]} & {lizzieLet25_4_r,
                                                                                                                                              lizzieLet25_3_r,
                                                                                                                                              lizzieLet25_2_r,
                                                                                                                                              lizzieLet25_1_r}));
  assign readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb_r = (& readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb_emitted <= 4'd0;
    else
      readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb_emitted <= (readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb_r ? 4'd0 :
                                                               readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb_done);
  
  /* buf (Ty CTkron_kron_Int_Int_Int) : (readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf,CTkron_kron_Int_Int_Int) > (readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf_rwb,CTkron_kron_Int_Int_Int) */
  CTkron_kron_Int_Int_Int_t readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf_bufchan_d;
  logic readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf_bufchan_r;
  assign readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf_r = ((! readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf_bufchan_d[0]) || readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf_bufchan_d <= {83'd0,
                                                                           1'd0};
    else
      if (readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf_r)
        readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf_bufchan_d <= readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf_d;
  CTkron_kron_Int_Int_Int_t readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf_bufchan_buf;
  assign readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf_bufchan_r = (! readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf_bufchan_buf[0]);
  assign readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf_rwb_d = (readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf_bufchan_buf[0] ? readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf_bufchan_buf :
                                                                         readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf_bufchan_buf <= {83'd0,
                                                                             1'd0};
    else
      if ((readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf_rwb_r && readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf_bufchan_buf[0]))
        readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf_bufchan_buf <= {83'd0,
                                                                               1'd0};
      else if (((! readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf_rwb_r) && (! readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf_bufchan_buf[0])))
        readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf_bufchan_buf <= readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf_bufchan_d;
  
  /* fork (Ty CTkron_kron_Int_Int_Int) : (readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf_rwb,CTkron_kron_Int_Int_Int) > [(lizzieLet29_1,CTkron_kron_Int_Int_Int),
                                                                                                                            (lizzieLet29_2,CTkron_kron_Int_Int_Int),
                                                                                                                            (lizzieLet29_3,CTkron_kron_Int_Int_Int),
                                                                                                                            (lizzieLet29_4,CTkron_kron_Int_Int_Int)] */
  logic [3:0] readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf_rwb_emitted;
  logic [3:0] readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf_rwb_done;
  assign lizzieLet29_1_d = {readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf_rwb_d[83:1],
                            (readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf_rwb_d[0] && (! readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf_rwb_emitted[0]))};
  assign lizzieLet29_2_d = {readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf_rwb_d[83:1],
                            (readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf_rwb_d[0] && (! readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf_rwb_emitted[1]))};
  assign lizzieLet29_3_d = {readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf_rwb_d[83:1],
                            (readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf_rwb_d[0] && (! readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf_rwb_emitted[2]))};
  assign lizzieLet29_4_d = {readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf_rwb_d[83:1],
                            (readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf_rwb_d[0] && (! readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf_rwb_emitted[3]))};
  assign readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf_rwb_done = (readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf_rwb_emitted | ({lizzieLet29_4_d[0],
                                                                                                                                                   lizzieLet29_3_d[0],
                                                                                                                                                   lizzieLet29_2_d[0],
                                                                                                                                                   lizzieLet29_1_d[0]} & {lizzieLet29_4_r,
                                                                                                                                                                          lizzieLet29_3_r,
                                                                                                                                                                          lizzieLet29_2_r,
                                                                                                                                                                          lizzieLet29_1_r}));
  assign readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf_rwb_r = (& readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf_rwb_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf_rwb_emitted <= 4'd0;
    else
      readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf_rwb_emitted <= (readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf_rwb_r ? 4'd0 :
                                                                             readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf_rwb_done);
  
  /* buf (Ty CTmain_map'_Int_Int) : (readPointer_CTmain_map'_Int_Intscfarg_0_2_1_argbuf,CTmain_map'_Int_Int) > (readPointer_CTmain_map'_Int_Intscfarg_0_2_1_argbuf_rwb,CTmain_map'_Int_Int) */
  \CTmain_map'_Int_Int_t  \readPointer_CTmain_map'_Int_Intscfarg_0_2_1_argbuf_bufchan_d ;
  logic \readPointer_CTmain_map'_Int_Intscfarg_0_2_1_argbuf_bufchan_r ;
  assign \readPointer_CTmain_map'_Int_Intscfarg_0_2_1_argbuf_r  = ((! \readPointer_CTmain_map'_Int_Intscfarg_0_2_1_argbuf_bufchan_d [0]) || \readPointer_CTmain_map'_Int_Intscfarg_0_2_1_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \readPointer_CTmain_map'_Int_Intscfarg_0_2_1_argbuf_bufchan_d  <= {67'd0,
                                                                         1'd0};
    else
      if (\readPointer_CTmain_map'_Int_Intscfarg_0_2_1_argbuf_r )
        \readPointer_CTmain_map'_Int_Intscfarg_0_2_1_argbuf_bufchan_d  <= \readPointer_CTmain_map'_Int_Intscfarg_0_2_1_argbuf_d ;
  \CTmain_map'_Int_Int_t  \readPointer_CTmain_map'_Int_Intscfarg_0_2_1_argbuf_bufchan_buf ;
  assign \readPointer_CTmain_map'_Int_Intscfarg_0_2_1_argbuf_bufchan_r  = (! \readPointer_CTmain_map'_Int_Intscfarg_0_2_1_argbuf_bufchan_buf [0]);
  assign \readPointer_CTmain_map'_Int_Intscfarg_0_2_1_argbuf_rwb_d  = (\readPointer_CTmain_map'_Int_Intscfarg_0_2_1_argbuf_bufchan_buf [0] ? \readPointer_CTmain_map'_Int_Intscfarg_0_2_1_argbuf_bufchan_buf  :
                                                                       \readPointer_CTmain_map'_Int_Intscfarg_0_2_1_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \readPointer_CTmain_map'_Int_Intscfarg_0_2_1_argbuf_bufchan_buf  <= {67'd0,
                                                                           1'd0};
    else
      if ((\readPointer_CTmain_map'_Int_Intscfarg_0_2_1_argbuf_rwb_r  && \readPointer_CTmain_map'_Int_Intscfarg_0_2_1_argbuf_bufchan_buf [0]))
        \readPointer_CTmain_map'_Int_Intscfarg_0_2_1_argbuf_bufchan_buf  <= {67'd0,
                                                                             1'd0};
      else if (((! \readPointer_CTmain_map'_Int_Intscfarg_0_2_1_argbuf_rwb_r ) && (! \readPointer_CTmain_map'_Int_Intscfarg_0_2_1_argbuf_bufchan_buf [0])))
        \readPointer_CTmain_map'_Int_Intscfarg_0_2_1_argbuf_bufchan_buf  <= \readPointer_CTmain_map'_Int_Intscfarg_0_2_1_argbuf_bufchan_d ;
  
  /* fork (Ty CTmain_map'_Int_Int) : (readPointer_CTmain_map'_Int_Intscfarg_0_2_1_argbuf_rwb,CTmain_map'_Int_Int) > [(lizzieLet34_1,CTmain_map'_Int_Int),
                                                                                                                (lizzieLet34_2,CTmain_map'_Int_Int),
                                                                                                                (lizzieLet34_3,CTmain_map'_Int_Int),
                                                                                                                (lizzieLet34_4,CTmain_map'_Int_Int)] */
  logic [3:0] \readPointer_CTmain_map'_Int_Intscfarg_0_2_1_argbuf_rwb_emitted ;
  logic [3:0] \readPointer_CTmain_map'_Int_Intscfarg_0_2_1_argbuf_rwb_done ;
  assign lizzieLet34_1_d = {\readPointer_CTmain_map'_Int_Intscfarg_0_2_1_argbuf_rwb_d [67:1],
                            (\readPointer_CTmain_map'_Int_Intscfarg_0_2_1_argbuf_rwb_d [0] && (! \readPointer_CTmain_map'_Int_Intscfarg_0_2_1_argbuf_rwb_emitted [0]))};
  assign lizzieLet34_2_d = {\readPointer_CTmain_map'_Int_Intscfarg_0_2_1_argbuf_rwb_d [67:1],
                            (\readPointer_CTmain_map'_Int_Intscfarg_0_2_1_argbuf_rwb_d [0] && (! \readPointer_CTmain_map'_Int_Intscfarg_0_2_1_argbuf_rwb_emitted [1]))};
  assign lizzieLet34_3_d = {\readPointer_CTmain_map'_Int_Intscfarg_0_2_1_argbuf_rwb_d [67:1],
                            (\readPointer_CTmain_map'_Int_Intscfarg_0_2_1_argbuf_rwb_d [0] && (! \readPointer_CTmain_map'_Int_Intscfarg_0_2_1_argbuf_rwb_emitted [2]))};
  assign lizzieLet34_4_d = {\readPointer_CTmain_map'_Int_Intscfarg_0_2_1_argbuf_rwb_d [67:1],
                            (\readPointer_CTmain_map'_Int_Intscfarg_0_2_1_argbuf_rwb_d [0] && (! \readPointer_CTmain_map'_Int_Intscfarg_0_2_1_argbuf_rwb_emitted [3]))};
  assign \readPointer_CTmain_map'_Int_Intscfarg_0_2_1_argbuf_rwb_done  = (\readPointer_CTmain_map'_Int_Intscfarg_0_2_1_argbuf_rwb_emitted  | ({lizzieLet34_4_d[0],
                                                                                                                                               lizzieLet34_3_d[0],
                                                                                                                                               lizzieLet34_2_d[0],
                                                                                                                                               lizzieLet34_1_d[0]} & {lizzieLet34_4_r,
                                                                                                                                                                      lizzieLet34_3_r,
                                                                                                                                                                      lizzieLet34_2_r,
                                                                                                                                                                      lizzieLet34_1_r}));
  assign \readPointer_CTmain_map'_Int_Intscfarg_0_2_1_argbuf_rwb_r  = (& \readPointer_CTmain_map'_Int_Intscfarg_0_2_1_argbuf_rwb_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \readPointer_CTmain_map'_Int_Intscfarg_0_2_1_argbuf_rwb_emitted  <= 4'd0;
    else
      \readPointer_CTmain_map'_Int_Intscfarg_0_2_1_argbuf_rwb_emitted  <= (\readPointer_CTmain_map'_Int_Intscfarg_0_2_1_argbuf_rwb_r  ? 4'd0 :
                                                                           \readPointer_CTmain_map'_Int_Intscfarg_0_2_1_argbuf_rwb_done );
  
  /* buf (Ty CTmap''_map''_Int_Int_Int) : (readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf,CTmap''_map''_Int_Int_Int) > (readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf_rwb,CTmap''_map''_Int_Int_Int) */
  \CTmap''_map''_Int_Int_Int_t  \readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf_bufchan_d ;
  logic \readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf_bufchan_r ;
  assign \readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf_r  = ((! \readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf_bufchan_d [0]) || \readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf_bufchan_d  <= {99'd0,
                                                                               1'd0};
    else
      if (\readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf_r )
        \readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf_bufchan_d  <= \readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf_d ;
  \CTmap''_map''_Int_Int_Int_t  \readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf_bufchan_buf ;
  assign \readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf_bufchan_r  = (! \readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf_bufchan_buf [0]);
  assign \readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf_rwb_d  = (\readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf_bufchan_buf [0] ? \readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf_bufchan_buf  :
                                                                             \readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf_bufchan_buf  <= {99'd0,
                                                                                 1'd0};
    else
      if ((\readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf_rwb_r  && \readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf_bufchan_buf [0]))
        \readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf_bufchan_buf  <= {99'd0,
                                                                                   1'd0};
      else if (((! \readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf_rwb_r ) && (! \readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf_bufchan_buf [0])))
        \readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf_bufchan_buf  <= \readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf_bufchan_d ;
  
  /* fork (Ty CTmap''_map''_Int_Int_Int) : (readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf_rwb,CTmap''_map''_Int_Int_Int) > [(lizzieLet39_1,CTmap''_map''_Int_Int_Int),
                                                                                                                                  (lizzieLet39_2,CTmap''_map''_Int_Int_Int),
                                                                                                                                  (lizzieLet39_3,CTmap''_map''_Int_Int_Int),
                                                                                                                                  (lizzieLet39_4,CTmap''_map''_Int_Int_Int)] */
  logic [3:0] \readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf_rwb_emitted ;
  logic [3:0] \readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf_rwb_done ;
  assign lizzieLet39_1_d = {\readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf_rwb_d [99:1],
                            (\readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf_rwb_d [0] && (! \readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf_rwb_emitted [0]))};
  assign lizzieLet39_2_d = {\readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf_rwb_d [99:1],
                            (\readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf_rwb_d [0] && (! \readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf_rwb_emitted [1]))};
  assign lizzieLet39_3_d = {\readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf_rwb_d [99:1],
                            (\readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf_rwb_d [0] && (! \readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf_rwb_emitted [2]))};
  assign lizzieLet39_4_d = {\readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf_rwb_d [99:1],
                            (\readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf_rwb_d [0] && (! \readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf_rwb_emitted [3]))};
  assign \readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf_rwb_done  = (\readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf_rwb_emitted  | ({lizzieLet39_4_d[0],
                                                                                                                                                           lizzieLet39_3_d[0],
                                                                                                                                                           lizzieLet39_2_d[0],
                                                                                                                                                           lizzieLet39_1_d[0]} & {lizzieLet39_4_r,
                                                                                                                                                                                  lizzieLet39_3_r,
                                                                                                                                                                                  lizzieLet39_2_r,
                                                                                                                                                                                  lizzieLet39_1_r}));
  assign \readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf_rwb_r  = (& \readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf_rwb_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf_rwb_emitted  <= 4'd0;
    else
      \readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf_rwb_emitted  <= (\readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf_rwb_r  ? 4'd0 :
                                                                                 \readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf_rwb_done );
  
  /* buf (Ty QTree_Int) : (readPointer_QTree_Intm1ad4_1_argbuf,QTree_Int) > (readPointer_QTree_Intm1ad4_1_argbuf_rwb,QTree_Int) */
  QTree_Int_t readPointer_QTree_Intm1ad4_1_argbuf_bufchan_d;
  logic readPointer_QTree_Intm1ad4_1_argbuf_bufchan_r;
  assign readPointer_QTree_Intm1ad4_1_argbuf_r = ((! readPointer_QTree_Intm1ad4_1_argbuf_bufchan_d[0]) || readPointer_QTree_Intm1ad4_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Intm1ad4_1_argbuf_bufchan_d <= {66'd0, 1'd0};
    else
      if (readPointer_QTree_Intm1ad4_1_argbuf_r)
        readPointer_QTree_Intm1ad4_1_argbuf_bufchan_d <= readPointer_QTree_Intm1ad4_1_argbuf_d;
  QTree_Int_t readPointer_QTree_Intm1ad4_1_argbuf_bufchan_buf;
  assign readPointer_QTree_Intm1ad4_1_argbuf_bufchan_r = (! readPointer_QTree_Intm1ad4_1_argbuf_bufchan_buf[0]);
  assign readPointer_QTree_Intm1ad4_1_argbuf_rwb_d = (readPointer_QTree_Intm1ad4_1_argbuf_bufchan_buf[0] ? readPointer_QTree_Intm1ad4_1_argbuf_bufchan_buf :
                                                      readPointer_QTree_Intm1ad4_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Intm1ad4_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((readPointer_QTree_Intm1ad4_1_argbuf_rwb_r && readPointer_QTree_Intm1ad4_1_argbuf_bufchan_buf[0]))
        readPointer_QTree_Intm1ad4_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
      else if (((! readPointer_QTree_Intm1ad4_1_argbuf_rwb_r) && (! readPointer_QTree_Intm1ad4_1_argbuf_bufchan_buf[0])))
        readPointer_QTree_Intm1ad4_1_argbuf_bufchan_buf <= readPointer_QTree_Intm1ad4_1_argbuf_bufchan_d;
  
  /* fork (Ty QTree_Int) : (readPointer_QTree_Intm1ad4_1_argbuf_rwb,QTree_Int) > [(lizzieLet6_1,QTree_Int),
                                                                             (lizzieLet6_2,QTree_Int),
                                                                             (lizzieLet6_3,QTree_Int),
                                                                             (lizzieLet6_4,QTree_Int),
                                                                             (lizzieLet6_5,QTree_Int),
                                                                             (lizzieLet6_6,QTree_Int),
                                                                             (lizzieLet6_7,QTree_Int)] */
  logic [6:0] readPointer_QTree_Intm1ad4_1_argbuf_rwb_emitted;
  logic [6:0] readPointer_QTree_Intm1ad4_1_argbuf_rwb_done;
  assign lizzieLet6_1_d = {readPointer_QTree_Intm1ad4_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_Intm1ad4_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intm1ad4_1_argbuf_rwb_emitted[0]))};
  assign lizzieLet6_2_d = {readPointer_QTree_Intm1ad4_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_Intm1ad4_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intm1ad4_1_argbuf_rwb_emitted[1]))};
  assign lizzieLet6_3_d = {readPointer_QTree_Intm1ad4_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_Intm1ad4_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intm1ad4_1_argbuf_rwb_emitted[2]))};
  assign lizzieLet6_4_d = {readPointer_QTree_Intm1ad4_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_Intm1ad4_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intm1ad4_1_argbuf_rwb_emitted[3]))};
  assign lizzieLet6_5_d = {readPointer_QTree_Intm1ad4_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_Intm1ad4_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intm1ad4_1_argbuf_rwb_emitted[4]))};
  assign lizzieLet6_6_d = {readPointer_QTree_Intm1ad4_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_Intm1ad4_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intm1ad4_1_argbuf_rwb_emitted[5]))};
  assign lizzieLet6_7_d = {readPointer_QTree_Intm1ad4_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_Intm1ad4_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intm1ad4_1_argbuf_rwb_emitted[6]))};
  assign readPointer_QTree_Intm1ad4_1_argbuf_rwb_done = (readPointer_QTree_Intm1ad4_1_argbuf_rwb_emitted | ({lizzieLet6_7_d[0],
                                                                                                             lizzieLet6_6_d[0],
                                                                                                             lizzieLet6_5_d[0],
                                                                                                             lizzieLet6_4_d[0],
                                                                                                             lizzieLet6_3_d[0],
                                                                                                             lizzieLet6_2_d[0],
                                                                                                             lizzieLet6_1_d[0]} & {lizzieLet6_7_r,
                                                                                                                                   lizzieLet6_6_r,
                                                                                                                                   lizzieLet6_5_r,
                                                                                                                                   lizzieLet6_4_r,
                                                                                                                                   lizzieLet6_3_r,
                                                                                                                                   lizzieLet6_2_r,
                                                                                                                                   lizzieLet6_1_r}));
  assign readPointer_QTree_Intm1ad4_1_argbuf_rwb_r = (& readPointer_QTree_Intm1ad4_1_argbuf_rwb_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Intm1ad4_1_argbuf_rwb_emitted <= 7'd0;
    else
      readPointer_QTree_Intm1ad4_1_argbuf_rwb_emitted <= (readPointer_QTree_Intm1ad4_1_argbuf_rwb_r ? 7'd0 :
                                                          readPointer_QTree_Intm1ad4_1_argbuf_rwb_done);
  
  /* buf (Ty QTree_Int) : (readPointer_QTree_IntmacN_1_argbuf,QTree_Int) > (readPointer_QTree_IntmacN_1_argbuf_rwb,QTree_Int) */
  QTree_Int_t readPointer_QTree_IntmacN_1_argbuf_bufchan_d;
  logic readPointer_QTree_IntmacN_1_argbuf_bufchan_r;
  assign readPointer_QTree_IntmacN_1_argbuf_r = ((! readPointer_QTree_IntmacN_1_argbuf_bufchan_d[0]) || readPointer_QTree_IntmacN_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_IntmacN_1_argbuf_bufchan_d <= {66'd0, 1'd0};
    else
      if (readPointer_QTree_IntmacN_1_argbuf_r)
        readPointer_QTree_IntmacN_1_argbuf_bufchan_d <= readPointer_QTree_IntmacN_1_argbuf_d;
  QTree_Int_t readPointer_QTree_IntmacN_1_argbuf_bufchan_buf;
  assign readPointer_QTree_IntmacN_1_argbuf_bufchan_r = (! readPointer_QTree_IntmacN_1_argbuf_bufchan_buf[0]);
  assign readPointer_QTree_IntmacN_1_argbuf_rwb_d = (readPointer_QTree_IntmacN_1_argbuf_bufchan_buf[0] ? readPointer_QTree_IntmacN_1_argbuf_bufchan_buf :
                                                     readPointer_QTree_IntmacN_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_IntmacN_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((readPointer_QTree_IntmacN_1_argbuf_rwb_r && readPointer_QTree_IntmacN_1_argbuf_bufchan_buf[0]))
        readPointer_QTree_IntmacN_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
      else if (((! readPointer_QTree_IntmacN_1_argbuf_rwb_r) && (! readPointer_QTree_IntmacN_1_argbuf_bufchan_buf[0])))
        readPointer_QTree_IntmacN_1_argbuf_bufchan_buf <= readPointer_QTree_IntmacN_1_argbuf_bufchan_d;
  
  /* fork (Ty QTree_Int) : (readPointer_QTree_IntmacN_1_argbuf_rwb,QTree_Int) > [(lizzieLet10_1,QTree_Int),
                                                                            (lizzieLet10_2,QTree_Int),
                                                                            (lizzieLet10_3,QTree_Int),
                                                                            (lizzieLet10_4,QTree_Int),
                                                                            (lizzieLet10_5,QTree_Int),
                                                                            (lizzieLet10_6,QTree_Int)] */
  logic [5:0] readPointer_QTree_IntmacN_1_argbuf_rwb_emitted;
  logic [5:0] readPointer_QTree_IntmacN_1_argbuf_rwb_done;
  assign lizzieLet10_1_d = {readPointer_QTree_IntmacN_1_argbuf_rwb_d[66:1],
                            (readPointer_QTree_IntmacN_1_argbuf_rwb_d[0] && (! readPointer_QTree_IntmacN_1_argbuf_rwb_emitted[0]))};
  assign lizzieLet10_2_d = {readPointer_QTree_IntmacN_1_argbuf_rwb_d[66:1],
                            (readPointer_QTree_IntmacN_1_argbuf_rwb_d[0] && (! readPointer_QTree_IntmacN_1_argbuf_rwb_emitted[1]))};
  assign lizzieLet10_3_d = {readPointer_QTree_IntmacN_1_argbuf_rwb_d[66:1],
                            (readPointer_QTree_IntmacN_1_argbuf_rwb_d[0] && (! readPointer_QTree_IntmacN_1_argbuf_rwb_emitted[2]))};
  assign lizzieLet10_4_d = {readPointer_QTree_IntmacN_1_argbuf_rwb_d[66:1],
                            (readPointer_QTree_IntmacN_1_argbuf_rwb_d[0] && (! readPointer_QTree_IntmacN_1_argbuf_rwb_emitted[3]))};
  assign lizzieLet10_5_d = {readPointer_QTree_IntmacN_1_argbuf_rwb_d[66:1],
                            (readPointer_QTree_IntmacN_1_argbuf_rwb_d[0] && (! readPointer_QTree_IntmacN_1_argbuf_rwb_emitted[4]))};
  assign lizzieLet10_6_d = {readPointer_QTree_IntmacN_1_argbuf_rwb_d[66:1],
                            (readPointer_QTree_IntmacN_1_argbuf_rwb_d[0] && (! readPointer_QTree_IntmacN_1_argbuf_rwb_emitted[5]))};
  assign readPointer_QTree_IntmacN_1_argbuf_rwb_done = (readPointer_QTree_IntmacN_1_argbuf_rwb_emitted | ({lizzieLet10_6_d[0],
                                                                                                           lizzieLet10_5_d[0],
                                                                                                           lizzieLet10_4_d[0],
                                                                                                           lizzieLet10_3_d[0],
                                                                                                           lizzieLet10_2_d[0],
                                                                                                           lizzieLet10_1_d[0]} & {lizzieLet10_6_r,
                                                                                                                                  lizzieLet10_5_r,
                                                                                                                                  lizzieLet10_4_r,
                                                                                                                                  lizzieLet10_3_r,
                                                                                                                                  lizzieLet10_2_r,
                                                                                                                                  lizzieLet10_1_r}));
  assign readPointer_QTree_IntmacN_1_argbuf_rwb_r = (& readPointer_QTree_IntmacN_1_argbuf_rwb_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_IntmacN_1_argbuf_rwb_emitted <= 6'd0;
    else
      readPointer_QTree_IntmacN_1_argbuf_rwb_emitted <= (readPointer_QTree_IntmacN_1_argbuf_rwb_r ? 6'd0 :
                                                         readPointer_QTree_IntmacN_1_argbuf_rwb_done);
  
  /* buf (Ty QTree_Int) : (readPointer_QTree_IntmacW_1_argbuf,QTree_Int) > (readPointer_QTree_IntmacW_1_argbuf_rwb,QTree_Int) */
  QTree_Int_t readPointer_QTree_IntmacW_1_argbuf_bufchan_d;
  logic readPointer_QTree_IntmacW_1_argbuf_bufchan_r;
  assign readPointer_QTree_IntmacW_1_argbuf_r = ((! readPointer_QTree_IntmacW_1_argbuf_bufchan_d[0]) || readPointer_QTree_IntmacW_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_IntmacW_1_argbuf_bufchan_d <= {66'd0, 1'd0};
    else
      if (readPointer_QTree_IntmacW_1_argbuf_r)
        readPointer_QTree_IntmacW_1_argbuf_bufchan_d <= readPointer_QTree_IntmacW_1_argbuf_d;
  QTree_Int_t readPointer_QTree_IntmacW_1_argbuf_bufchan_buf;
  assign readPointer_QTree_IntmacW_1_argbuf_bufchan_r = (! readPointer_QTree_IntmacW_1_argbuf_bufchan_buf[0]);
  assign readPointer_QTree_IntmacW_1_argbuf_rwb_d = (readPointer_QTree_IntmacW_1_argbuf_bufchan_buf[0] ? readPointer_QTree_IntmacW_1_argbuf_bufchan_buf :
                                                     readPointer_QTree_IntmacW_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_IntmacW_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((readPointer_QTree_IntmacW_1_argbuf_rwb_r && readPointer_QTree_IntmacW_1_argbuf_bufchan_buf[0]))
        readPointer_QTree_IntmacW_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
      else if (((! readPointer_QTree_IntmacW_1_argbuf_rwb_r) && (! readPointer_QTree_IntmacW_1_argbuf_bufchan_buf[0])))
        readPointer_QTree_IntmacW_1_argbuf_bufchan_buf <= readPointer_QTree_IntmacW_1_argbuf_bufchan_d;
  
  /* fork (Ty QTree_Int) : (readPointer_QTree_IntmacW_1_argbuf_rwb,QTree_Int) > [(lizzieLet16_1_1,QTree_Int),
                                                                            (lizzieLet16_1_2,QTree_Int),
                                                                            (lizzieLet16_1_3,QTree_Int),
                                                                            (lizzieLet16_1_4,QTree_Int),
                                                                            (lizzieLet16_1_5,QTree_Int),
                                                                            (lizzieLet16_1_6,QTree_Int),
                                                                            (lizzieLet16_1_7,QTree_Int)] */
  logic [6:0] readPointer_QTree_IntmacW_1_argbuf_rwb_emitted;
  logic [6:0] readPointer_QTree_IntmacW_1_argbuf_rwb_done;
  assign lizzieLet16_1_1_d = {readPointer_QTree_IntmacW_1_argbuf_rwb_d[66:1],
                              (readPointer_QTree_IntmacW_1_argbuf_rwb_d[0] && (! readPointer_QTree_IntmacW_1_argbuf_rwb_emitted[0]))};
  assign lizzieLet16_1_2_d = {readPointer_QTree_IntmacW_1_argbuf_rwb_d[66:1],
                              (readPointer_QTree_IntmacW_1_argbuf_rwb_d[0] && (! readPointer_QTree_IntmacW_1_argbuf_rwb_emitted[1]))};
  assign lizzieLet16_1_3_d = {readPointer_QTree_IntmacW_1_argbuf_rwb_d[66:1],
                              (readPointer_QTree_IntmacW_1_argbuf_rwb_d[0] && (! readPointer_QTree_IntmacW_1_argbuf_rwb_emitted[2]))};
  assign lizzieLet16_1_4_d = {readPointer_QTree_IntmacW_1_argbuf_rwb_d[66:1],
                              (readPointer_QTree_IntmacW_1_argbuf_rwb_d[0] && (! readPointer_QTree_IntmacW_1_argbuf_rwb_emitted[3]))};
  assign lizzieLet16_1_5_d = {readPointer_QTree_IntmacW_1_argbuf_rwb_d[66:1],
                              (readPointer_QTree_IntmacW_1_argbuf_rwb_d[0] && (! readPointer_QTree_IntmacW_1_argbuf_rwb_emitted[4]))};
  assign lizzieLet16_1_6_d = {readPointer_QTree_IntmacW_1_argbuf_rwb_d[66:1],
                              (readPointer_QTree_IntmacW_1_argbuf_rwb_d[0] && (! readPointer_QTree_IntmacW_1_argbuf_rwb_emitted[5]))};
  assign lizzieLet16_1_7_d = {readPointer_QTree_IntmacW_1_argbuf_rwb_d[66:1],
                              (readPointer_QTree_IntmacW_1_argbuf_rwb_d[0] && (! readPointer_QTree_IntmacW_1_argbuf_rwb_emitted[6]))};
  assign readPointer_QTree_IntmacW_1_argbuf_rwb_done = (readPointer_QTree_IntmacW_1_argbuf_rwb_emitted | ({lizzieLet16_1_7_d[0],
                                                                                                           lizzieLet16_1_6_d[0],
                                                                                                           lizzieLet16_1_5_d[0],
                                                                                                           lizzieLet16_1_4_d[0],
                                                                                                           lizzieLet16_1_3_d[0],
                                                                                                           lizzieLet16_1_2_d[0],
                                                                                                           lizzieLet16_1_1_d[0]} & {lizzieLet16_1_7_r,
                                                                                                                                    lizzieLet16_1_6_r,
                                                                                                                                    lizzieLet16_1_5_r,
                                                                                                                                    lizzieLet16_1_4_r,
                                                                                                                                    lizzieLet16_1_3_r,
                                                                                                                                    lizzieLet16_1_2_r,
                                                                                                                                    lizzieLet16_1_1_r}));
  assign readPointer_QTree_IntmacW_1_argbuf_rwb_r = (& readPointer_QTree_IntmacW_1_argbuf_rwb_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_IntmacW_1_argbuf_rwb_emitted <= 7'd0;
    else
      readPointer_QTree_IntmacW_1_argbuf_rwb_emitted <= (readPointer_QTree_IntmacW_1_argbuf_rwb_r ? 7'd0 :
                                                         readPointer_QTree_IntmacW_1_argbuf_rwb_done);
  
  /* buf (Ty QTree_Int) : (readPointer_QTree_Intwsvt_1_1_argbuf,QTree_Int) > (readPointer_QTree_Intwsvt_1_1_argbuf_rwb,QTree_Int) */
  QTree_Int_t readPointer_QTree_Intwsvt_1_1_argbuf_bufchan_d;
  logic readPointer_QTree_Intwsvt_1_1_argbuf_bufchan_r;
  assign readPointer_QTree_Intwsvt_1_1_argbuf_r = ((! readPointer_QTree_Intwsvt_1_1_argbuf_bufchan_d[0]) || readPointer_QTree_Intwsvt_1_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Intwsvt_1_1_argbuf_bufchan_d <= {66'd0, 1'd0};
    else
      if (readPointer_QTree_Intwsvt_1_1_argbuf_r)
        readPointer_QTree_Intwsvt_1_1_argbuf_bufchan_d <= readPointer_QTree_Intwsvt_1_1_argbuf_d;
  QTree_Int_t readPointer_QTree_Intwsvt_1_1_argbuf_bufchan_buf;
  assign readPointer_QTree_Intwsvt_1_1_argbuf_bufchan_r = (! readPointer_QTree_Intwsvt_1_1_argbuf_bufchan_buf[0]);
  assign readPointer_QTree_Intwsvt_1_1_argbuf_rwb_d = (readPointer_QTree_Intwsvt_1_1_argbuf_bufchan_buf[0] ? readPointer_QTree_Intwsvt_1_1_argbuf_bufchan_buf :
                                                       readPointer_QTree_Intwsvt_1_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Intwsvt_1_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((readPointer_QTree_Intwsvt_1_1_argbuf_rwb_r && readPointer_QTree_Intwsvt_1_1_argbuf_bufchan_buf[0]))
        readPointer_QTree_Intwsvt_1_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
      else if (((! readPointer_QTree_Intwsvt_1_1_argbuf_rwb_r) && (! readPointer_QTree_Intwsvt_1_1_argbuf_bufchan_buf[0])))
        readPointer_QTree_Intwsvt_1_1_argbuf_bufchan_buf <= readPointer_QTree_Intwsvt_1_1_argbuf_bufchan_d;
  
  /* fork (Ty QTree_Int) : (readPointer_QTree_Intwsvt_1_1_argbuf_rwb,QTree_Int) > [(lizzieLet4_1,QTree_Int),
                                                                              (lizzieLet4_2,QTree_Int),
                                                                              (lizzieLet4_3,QTree_Int),
                                                                              (lizzieLet4_4,QTree_Int)] */
  logic [3:0] readPointer_QTree_Intwsvt_1_1_argbuf_rwb_emitted;
  logic [3:0] readPointer_QTree_Intwsvt_1_1_argbuf_rwb_done;
  assign lizzieLet4_1_d = {readPointer_QTree_Intwsvt_1_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_Intwsvt_1_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intwsvt_1_1_argbuf_rwb_emitted[0]))};
  assign lizzieLet4_2_d = {readPointer_QTree_Intwsvt_1_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_Intwsvt_1_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intwsvt_1_1_argbuf_rwb_emitted[1]))};
  assign lizzieLet4_3_d = {readPointer_QTree_Intwsvt_1_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_Intwsvt_1_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intwsvt_1_1_argbuf_rwb_emitted[2]))};
  assign lizzieLet4_4_d = {readPointer_QTree_Intwsvt_1_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_Intwsvt_1_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intwsvt_1_1_argbuf_rwb_emitted[3]))};
  assign readPointer_QTree_Intwsvt_1_1_argbuf_rwb_done = (readPointer_QTree_Intwsvt_1_1_argbuf_rwb_emitted | ({lizzieLet4_4_d[0],
                                                                                                               lizzieLet4_3_d[0],
                                                                                                               lizzieLet4_2_d[0],
                                                                                                               lizzieLet4_1_d[0]} & {lizzieLet4_4_r,
                                                                                                                                     lizzieLet4_3_r,
                                                                                                                                     lizzieLet4_2_r,
                                                                                                                                     lizzieLet4_1_r}));
  assign readPointer_QTree_Intwsvt_1_1_argbuf_rwb_r = (& readPointer_QTree_Intwsvt_1_1_argbuf_rwb_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Intwsvt_1_1_argbuf_rwb_emitted <= 4'd0;
    else
      readPointer_QTree_Intwsvt_1_1_argbuf_rwb_emitted <= (readPointer_QTree_Intwsvt_1_1_argbuf_rwb_r ? 4'd0 :
                                                           readPointer_QTree_Intwsvt_1_1_argbuf_rwb_done);
  
  /* buf (Ty Pointer_CTkron_kron_Int_Int_Int) : (sc_0_11_destruct,Pointer_CTkron_kron_Int_Int_Int) > (sc_0_11_1_argbuf,Pointer_CTkron_kron_Int_Int_Int) */
  Pointer_CTkron_kron_Int_Int_Int_t sc_0_11_destruct_bufchan_d;
  logic sc_0_11_destruct_bufchan_r;
  assign sc_0_11_destruct_r = ((! sc_0_11_destruct_bufchan_d[0]) || sc_0_11_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) sc_0_11_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (sc_0_11_destruct_r)
        sc_0_11_destruct_bufchan_d <= sc_0_11_destruct_d;
  Pointer_CTkron_kron_Int_Int_Int_t sc_0_11_destruct_bufchan_buf;
  assign sc_0_11_destruct_bufchan_r = (! sc_0_11_destruct_bufchan_buf[0]);
  assign sc_0_11_1_argbuf_d = (sc_0_11_destruct_bufchan_buf[0] ? sc_0_11_destruct_bufchan_buf :
                               sc_0_11_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) sc_0_11_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((sc_0_11_1_argbuf_r && sc_0_11_destruct_bufchan_buf[0]))
        sc_0_11_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! sc_0_11_1_argbuf_r) && (! sc_0_11_destruct_bufchan_buf[0])))
        sc_0_11_destruct_bufchan_buf <= sc_0_11_destruct_bufchan_d;
  
  /* buf (Ty Pointer_CTmain_map'_Int_Int) : (sc_0_15_destruct,Pointer_CTmain_map'_Int_Int) > (sc_0_15_1_argbuf,Pointer_CTmain_map'_Int_Int) */
  \Pointer_CTmain_map'_Int_Int_t  sc_0_15_destruct_bufchan_d;
  logic sc_0_15_destruct_bufchan_r;
  assign sc_0_15_destruct_r = ((! sc_0_15_destruct_bufchan_d[0]) || sc_0_15_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) sc_0_15_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (sc_0_15_destruct_r)
        sc_0_15_destruct_bufchan_d <= sc_0_15_destruct_d;
  \Pointer_CTmain_map'_Int_Int_t  sc_0_15_destruct_bufchan_buf;
  assign sc_0_15_destruct_bufchan_r = (! sc_0_15_destruct_bufchan_buf[0]);
  assign sc_0_15_1_argbuf_d = (sc_0_15_destruct_bufchan_buf[0] ? sc_0_15_destruct_bufchan_buf :
                               sc_0_15_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) sc_0_15_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((sc_0_15_1_argbuf_r && sc_0_15_destruct_bufchan_buf[0]))
        sc_0_15_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! sc_0_15_1_argbuf_r) && (! sc_0_15_destruct_bufchan_buf[0])))
        sc_0_15_destruct_bufchan_buf <= sc_0_15_destruct_bufchan_d;
  
  /* buf (Ty Pointer_CTmap''_map''_Int_Int_Int) : (sc_0_19_destruct,Pointer_CTmap''_map''_Int_Int_Int) > (sc_0_19_1_argbuf,Pointer_CTmap''_map''_Int_Int_Int) */
  \Pointer_CTmap''_map''_Int_Int_Int_t  sc_0_19_destruct_bufchan_d;
  logic sc_0_19_destruct_bufchan_r;
  assign sc_0_19_destruct_r = ((! sc_0_19_destruct_bufchan_d[0]) || sc_0_19_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) sc_0_19_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (sc_0_19_destruct_r)
        sc_0_19_destruct_bufchan_d <= sc_0_19_destruct_d;
  \Pointer_CTmap''_map''_Int_Int_Int_t  sc_0_19_destruct_bufchan_buf;
  assign sc_0_19_destruct_bufchan_r = (! sc_0_19_destruct_bufchan_buf[0]);
  assign sc_0_19_1_argbuf_d = (sc_0_19_destruct_bufchan_buf[0] ? sc_0_19_destruct_bufchan_buf :
                               sc_0_19_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) sc_0_19_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((sc_0_19_1_argbuf_r && sc_0_19_destruct_bufchan_buf[0]))
        sc_0_19_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! sc_0_19_1_argbuf_r) && (! sc_0_19_destruct_bufchan_buf[0])))
        sc_0_19_destruct_bufchan_buf <= sc_0_19_destruct_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz_Int) : (sc_0_7_destruct,Pointer_CT$wnnz_Int) > (sc_0_7_1_argbuf,Pointer_CT$wnnz_Int) */
  Pointer_CT$wnnz_Int_t sc_0_7_destruct_bufchan_d;
  logic sc_0_7_destruct_bufchan_r;
  assign sc_0_7_destruct_r = ((! sc_0_7_destruct_bufchan_d[0]) || sc_0_7_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) sc_0_7_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (sc_0_7_destruct_r)
        sc_0_7_destruct_bufchan_d <= sc_0_7_destruct_d;
  Pointer_CT$wnnz_Int_t sc_0_7_destruct_bufchan_buf;
  assign sc_0_7_destruct_bufchan_r = (! sc_0_7_destruct_bufchan_buf[0]);
  assign sc_0_7_1_argbuf_d = (sc_0_7_destruct_bufchan_buf[0] ? sc_0_7_destruct_bufchan_buf :
                              sc_0_7_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) sc_0_7_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((sc_0_7_1_argbuf_r && sc_0_7_destruct_bufchan_buf[0]))
        sc_0_7_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! sc_0_7_1_argbuf_r) && (! sc_0_7_destruct_bufchan_buf[0])))
        sc_0_7_destruct_bufchan_buf <= sc_0_7_destruct_bufchan_d;
  
  /* buf (Ty Pointer_CTkron_kron_Int_Int_Int) : (scfarg_0_1_goMux_mux,Pointer_CTkron_kron_Int_Int_Int) > (scfarg_0_1_1_argbuf,Pointer_CTkron_kron_Int_Int_Int) */
  Pointer_CTkron_kron_Int_Int_Int_t scfarg_0_1_goMux_mux_bufchan_d;
  logic scfarg_0_1_goMux_mux_bufchan_r;
  assign scfarg_0_1_goMux_mux_r = ((! scfarg_0_1_goMux_mux_bufchan_d[0]) || scfarg_0_1_goMux_mux_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      scfarg_0_1_goMux_mux_bufchan_d <= {16'd0, 1'd0};
    else
      if (scfarg_0_1_goMux_mux_r)
        scfarg_0_1_goMux_mux_bufchan_d <= scfarg_0_1_goMux_mux_d;
  Pointer_CTkron_kron_Int_Int_Int_t scfarg_0_1_goMux_mux_bufchan_buf;
  assign scfarg_0_1_goMux_mux_bufchan_r = (! scfarg_0_1_goMux_mux_bufchan_buf[0]);
  assign scfarg_0_1_1_argbuf_d = (scfarg_0_1_goMux_mux_bufchan_buf[0] ? scfarg_0_1_goMux_mux_bufchan_buf :
                                  scfarg_0_1_goMux_mux_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      scfarg_0_1_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((scfarg_0_1_1_argbuf_r && scfarg_0_1_goMux_mux_bufchan_buf[0]))
        scfarg_0_1_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
      else if (((! scfarg_0_1_1_argbuf_r) && (! scfarg_0_1_goMux_mux_bufchan_buf[0])))
        scfarg_0_1_goMux_mux_bufchan_buf <= scfarg_0_1_goMux_mux_bufchan_d;
  
  /* buf (Ty Pointer_CTmain_map'_Int_Int) : (scfarg_0_2_goMux_mux,Pointer_CTmain_map'_Int_Int) > (scfarg_0_2_1_argbuf,Pointer_CTmain_map'_Int_Int) */
  \Pointer_CTmain_map'_Int_Int_t  scfarg_0_2_goMux_mux_bufchan_d;
  logic scfarg_0_2_goMux_mux_bufchan_r;
  assign scfarg_0_2_goMux_mux_r = ((! scfarg_0_2_goMux_mux_bufchan_d[0]) || scfarg_0_2_goMux_mux_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      scfarg_0_2_goMux_mux_bufchan_d <= {16'd0, 1'd0};
    else
      if (scfarg_0_2_goMux_mux_r)
        scfarg_0_2_goMux_mux_bufchan_d <= scfarg_0_2_goMux_mux_d;
  \Pointer_CTmain_map'_Int_Int_t  scfarg_0_2_goMux_mux_bufchan_buf;
  assign scfarg_0_2_goMux_mux_bufchan_r = (! scfarg_0_2_goMux_mux_bufchan_buf[0]);
  assign scfarg_0_2_1_argbuf_d = (scfarg_0_2_goMux_mux_bufchan_buf[0] ? scfarg_0_2_goMux_mux_bufchan_buf :
                                  scfarg_0_2_goMux_mux_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      scfarg_0_2_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((scfarg_0_2_1_argbuf_r && scfarg_0_2_goMux_mux_bufchan_buf[0]))
        scfarg_0_2_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
      else if (((! scfarg_0_2_1_argbuf_r) && (! scfarg_0_2_goMux_mux_bufchan_buf[0])))
        scfarg_0_2_goMux_mux_bufchan_buf <= scfarg_0_2_goMux_mux_bufchan_d;
  
  /* buf (Ty Pointer_CTmap''_map''_Int_Int_Int) : (scfarg_0_3_goMux_mux,Pointer_CTmap''_map''_Int_Int_Int) > (scfarg_0_3_1_argbuf,Pointer_CTmap''_map''_Int_Int_Int) */
  \Pointer_CTmap''_map''_Int_Int_Int_t  scfarg_0_3_goMux_mux_bufchan_d;
  logic scfarg_0_3_goMux_mux_bufchan_r;
  assign scfarg_0_3_goMux_mux_r = ((! scfarg_0_3_goMux_mux_bufchan_d[0]) || scfarg_0_3_goMux_mux_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      scfarg_0_3_goMux_mux_bufchan_d <= {16'd0, 1'd0};
    else
      if (scfarg_0_3_goMux_mux_r)
        scfarg_0_3_goMux_mux_bufchan_d <= scfarg_0_3_goMux_mux_d;
  \Pointer_CTmap''_map''_Int_Int_Int_t  scfarg_0_3_goMux_mux_bufchan_buf;
  assign scfarg_0_3_goMux_mux_bufchan_r = (! scfarg_0_3_goMux_mux_bufchan_buf[0]);
  assign scfarg_0_3_1_argbuf_d = (scfarg_0_3_goMux_mux_bufchan_buf[0] ? scfarg_0_3_goMux_mux_bufchan_buf :
                                  scfarg_0_3_goMux_mux_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      scfarg_0_3_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((scfarg_0_3_1_argbuf_r && scfarg_0_3_goMux_mux_bufchan_buf[0]))
        scfarg_0_3_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
      else if (((! scfarg_0_3_1_argbuf_r) && (! scfarg_0_3_goMux_mux_bufchan_buf[0])))
        scfarg_0_3_goMux_mux_bufchan_buf <= scfarg_0_3_goMux_mux_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz_Int) : (scfarg_0_goMux_mux,Pointer_CT$wnnz_Int) > (scfarg_0_1_argbuf,Pointer_CT$wnnz_Int) */
  Pointer_CT$wnnz_Int_t scfarg_0_goMux_mux_bufchan_d;
  logic scfarg_0_goMux_mux_bufchan_r;
  assign scfarg_0_goMux_mux_r = ((! scfarg_0_goMux_mux_bufchan_d[0]) || scfarg_0_goMux_mux_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) scfarg_0_goMux_mux_bufchan_d <= {16'd0, 1'd0};
    else
      if (scfarg_0_goMux_mux_r)
        scfarg_0_goMux_mux_bufchan_d <= scfarg_0_goMux_mux_d;
  Pointer_CT$wnnz_Int_t scfarg_0_goMux_mux_bufchan_buf;
  assign scfarg_0_goMux_mux_bufchan_r = (! scfarg_0_goMux_mux_bufchan_buf[0]);
  assign scfarg_0_1_argbuf_d = (scfarg_0_goMux_mux_bufchan_buf[0] ? scfarg_0_goMux_mux_bufchan_buf :
                                scfarg_0_goMux_mux_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      scfarg_0_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((scfarg_0_1_argbuf_r && scfarg_0_goMux_mux_bufchan_buf[0]))
        scfarg_0_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
      else if (((! scfarg_0_1_argbuf_r) && (! scfarg_0_goMux_mux_bufchan_buf[0])))
        scfarg_0_goMux_mux_bufchan_buf <= scfarg_0_goMux_mux_bufchan_d;
  
  /* buf (Ty Int) : (v'acV_2_2,Int) > (v'acV_2_2_argbuf,Int) */
  Int_t \v'acV_2_2_bufchan_d ;
  logic \v'acV_2_2_bufchan_r ;
  assign \v'acV_2_2_r  = ((! \v'acV_2_2_bufchan_d [0]) || \v'acV_2_2_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \v'acV_2_2_bufchan_d  <= {32'd0, 1'd0};
    else if (\v'acV_2_2_r ) \v'acV_2_2_bufchan_d  <= \v'acV_2_2_d ;
  Int_t \v'acV_2_2_bufchan_buf ;
  assign \v'acV_2_2_bufchan_r  = (! \v'acV_2_2_bufchan_buf [0]);
  assign \v'acV_2_2_argbuf_d  = (\v'acV_2_2_bufchan_buf [0] ? \v'acV_2_2_bufchan_buf  :
                                 \v'acV_2_2_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \v'acV_2_2_bufchan_buf  <= {32'd0, 1'd0};
    else
      if ((\v'acV_2_2_argbuf_r  && \v'acV_2_2_bufchan_buf [0]))
        \v'acV_2_2_bufchan_buf  <= {32'd0, 1'd0};
      else if (((! \v'acV_2_2_argbuf_r ) && (! \v'acV_2_2_bufchan_buf [0])))
        \v'acV_2_2_bufchan_buf  <= \v'acV_2_2_bufchan_d ;
  
  /* fork (Ty Int) : (v'acV_2_destruct,Int) > [(v'acV_2_1,Int),
                                          (v'acV_2_2,Int)] */
  logic [1:0] \v'acV_2_destruct_emitted ;
  logic [1:0] \v'acV_2_destruct_done ;
  assign \v'acV_2_1_d  = {\v'acV_2_destruct_d [32:1],
                          (\v'acV_2_destruct_d [0] && (! \v'acV_2_destruct_emitted [0]))};
  assign \v'acV_2_2_d  = {\v'acV_2_destruct_d [32:1],
                          (\v'acV_2_destruct_d [0] && (! \v'acV_2_destruct_emitted [1]))};
  assign \v'acV_2_destruct_done  = (\v'acV_2_destruct_emitted  | ({\v'acV_2_2_d [0],
                                                                   \v'acV_2_1_d [0]} & {\v'acV_2_2_r ,
                                                                                        \v'acV_2_1_r }));
  assign \v'acV_2_destruct_r  = (& \v'acV_2_destruct_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \v'acV_2_destruct_emitted  <= 2'd0;
    else
      \v'acV_2_destruct_emitted  <= (\v'acV_2_destruct_r  ? 2'd0 :
                                     \v'acV_2_destruct_done );
  
  /* buf (Ty Int) : (v'acV_3_2,Int) > (v'acV_3_2_argbuf,Int) */
  Int_t \v'acV_3_2_bufchan_d ;
  logic \v'acV_3_2_bufchan_r ;
  assign \v'acV_3_2_r  = ((! \v'acV_3_2_bufchan_d [0]) || \v'acV_3_2_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \v'acV_3_2_bufchan_d  <= {32'd0, 1'd0};
    else if (\v'acV_3_2_r ) \v'acV_3_2_bufchan_d  <= \v'acV_3_2_d ;
  Int_t \v'acV_3_2_bufchan_buf ;
  assign \v'acV_3_2_bufchan_r  = (! \v'acV_3_2_bufchan_buf [0]);
  assign \v'acV_3_2_argbuf_d  = (\v'acV_3_2_bufchan_buf [0] ? \v'acV_3_2_bufchan_buf  :
                                 \v'acV_3_2_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \v'acV_3_2_bufchan_buf  <= {32'd0, 1'd0};
    else
      if ((\v'acV_3_2_argbuf_r  && \v'acV_3_2_bufchan_buf [0]))
        \v'acV_3_2_bufchan_buf  <= {32'd0, 1'd0};
      else if (((! \v'acV_3_2_argbuf_r ) && (! \v'acV_3_2_bufchan_buf [0])))
        \v'acV_3_2_bufchan_buf  <= \v'acV_3_2_bufchan_d ;
  
  /* fork (Ty Int) : (v'acV_3_destruct,Int) > [(v'acV_3_1,Int),
                                          (v'acV_3_2,Int)] */
  logic [1:0] \v'acV_3_destruct_emitted ;
  logic [1:0] \v'acV_3_destruct_done ;
  assign \v'acV_3_1_d  = {\v'acV_3_destruct_d [32:1],
                          (\v'acV_3_destruct_d [0] && (! \v'acV_3_destruct_emitted [0]))};
  assign \v'acV_3_2_d  = {\v'acV_3_destruct_d [32:1],
                          (\v'acV_3_destruct_d [0] && (! \v'acV_3_destruct_emitted [1]))};
  assign \v'acV_3_destruct_done  = (\v'acV_3_destruct_emitted  | ({\v'acV_3_2_d [0],
                                                                   \v'acV_3_1_d [0]} & {\v'acV_3_2_r ,
                                                                                        \v'acV_3_1_r }));
  assign \v'acV_3_destruct_r  = (& \v'acV_3_destruct_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \v'acV_3_destruct_emitted  <= 2'd0;
    else
      \v'acV_3_destruct_emitted  <= (\v'acV_3_destruct_r  ? 2'd0 :
                                     \v'acV_3_destruct_done );
  
  /* buf (Ty Int) : (v'acV_4_destruct,Int) > (v'acV_4_1_argbuf,Int) */
  Int_t \v'acV_4_destruct_bufchan_d ;
  logic \v'acV_4_destruct_bufchan_r ;
  assign \v'acV_4_destruct_r  = ((! \v'acV_4_destruct_bufchan_d [0]) || \v'acV_4_destruct_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \v'acV_4_destruct_bufchan_d  <= {32'd0, 1'd0};
    else
      if (\v'acV_4_destruct_r )
        \v'acV_4_destruct_bufchan_d  <= \v'acV_4_destruct_d ;
  Int_t \v'acV_4_destruct_bufchan_buf ;
  assign \v'acV_4_destruct_bufchan_r  = (! \v'acV_4_destruct_bufchan_buf [0]);
  assign \v'acV_4_1_argbuf_d  = (\v'acV_4_destruct_bufchan_buf [0] ? \v'acV_4_destruct_bufchan_buf  :
                                 \v'acV_4_destruct_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \v'acV_4_destruct_bufchan_buf  <= {32'd0, 1'd0};
    else
      if ((\v'acV_4_1_argbuf_r  && \v'acV_4_destruct_bufchan_buf [0]))
        \v'acV_4_destruct_bufchan_buf  <= {32'd0, 1'd0};
      else if (((! \v'acV_4_1_argbuf_r ) && (! \v'acV_4_destruct_bufchan_buf [0])))
        \v'acV_4_destruct_bufchan_buf  <= \v'acV_4_destruct_bufchan_d ;
  
  /* buf (Ty Int) : (vacO_destruct,Int) > (vacO_1_argbuf,Int) */
  Int_t vacO_destruct_bufchan_d;
  logic vacO_destruct_bufchan_r;
  assign vacO_destruct_r = ((! vacO_destruct_bufchan_d[0]) || vacO_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) vacO_destruct_bufchan_d <= {32'd0, 1'd0};
    else
      if (vacO_destruct_r) vacO_destruct_bufchan_d <= vacO_destruct_d;
  Int_t vacO_destruct_bufchan_buf;
  assign vacO_destruct_bufchan_r = (! vacO_destruct_bufchan_buf[0]);
  assign vacO_1_argbuf_d = (vacO_destruct_bufchan_buf[0] ? vacO_destruct_bufchan_buf :
                            vacO_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) vacO_destruct_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((vacO_1_argbuf_r && vacO_destruct_bufchan_buf[0]))
        vacO_destruct_bufchan_buf <= {32'd0, 1'd0};
      else if (((! vacO_1_argbuf_r) && (! vacO_destruct_bufchan_buf[0])))
        vacO_destruct_bufchan_buf <= vacO_destruct_bufchan_d;
  
  /* buf (Ty Int) : (vacX_destruct,Int) > (vacX_1_argbuf,Int) */
  Int_t vacX_destruct_bufchan_d;
  logic vacX_destruct_bufchan_r;
  assign vacX_destruct_r = ((! vacX_destruct_bufchan_d[0]) || vacX_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) vacX_destruct_bufchan_d <= {32'd0, 1'd0};
    else
      if (vacX_destruct_r) vacX_destruct_bufchan_d <= vacX_destruct_d;
  Int_t vacX_destruct_bufchan_buf;
  assign vacX_destruct_bufchan_r = (! vacX_destruct_bufchan_buf[0]);
  assign vacX_1_argbuf_d = (vacX_destruct_bufchan_buf[0] ? vacX_destruct_bufchan_buf :
                            vacX_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) vacX_destruct_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((vacX_1_argbuf_r && vacX_destruct_bufchan_buf[0]))
        vacX_destruct_bufchan_buf <= {32'd0, 1'd0};
      else if (((! vacX_1_argbuf_r) && (! vacX_destruct_bufchan_buf[0])))
        vacX_destruct_bufchan_buf <= vacX_destruct_bufchan_d;
  
  /* buf (Ty Int) : (vad6_destruct,Int) > (vad6_1_argbuf,Int) */
  Int_t vad6_destruct_bufchan_d;
  logic vad6_destruct_bufchan_r;
  assign vad6_destruct_r = ((! vad6_destruct_bufchan_d[0]) || vad6_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) vad6_destruct_bufchan_d <= {32'd0, 1'd0};
    else
      if (vad6_destruct_r) vad6_destruct_bufchan_d <= vad6_destruct_d;
  Int_t vad6_destruct_bufchan_buf;
  assign vad6_destruct_bufchan_r = (! vad6_destruct_bufchan_buf[0]);
  assign vad6_1_argbuf_d = (vad6_destruct_bufchan_buf[0] ? vad6_destruct_bufchan_buf :
                            vad6_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) vad6_destruct_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((vad6_1_argbuf_r && vad6_destruct_bufchan_buf[0]))
        vad6_destruct_bufchan_buf <= {32'd0, 1'd0};
      else if (((! vad6_1_argbuf_r) && (! vad6_destruct_bufchan_buf[0])))
        vad6_destruct_bufchan_buf <= vad6_destruct_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz_Int) : (writeCT$wnnz_IntlizzieLet0_1_argbuf,Pointer_CT$wnnz_Int) > (writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb,Pointer_CT$wnnz_Int) */
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet0_1_argbuf_bufchan_d;
  logic writeCT$wnnz_IntlizzieLet0_1_argbuf_bufchan_r;
  assign writeCT$wnnz_IntlizzieLet0_1_argbuf_r = ((! writeCT$wnnz_IntlizzieLet0_1_argbuf_bufchan_d[0]) || writeCT$wnnz_IntlizzieLet0_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnz_IntlizzieLet0_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCT$wnnz_IntlizzieLet0_1_argbuf_r)
        writeCT$wnnz_IntlizzieLet0_1_argbuf_bufchan_d <= writeCT$wnnz_IntlizzieLet0_1_argbuf_d;
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet0_1_argbuf_bufchan_buf;
  assign writeCT$wnnz_IntlizzieLet0_1_argbuf_bufchan_r = (! writeCT$wnnz_IntlizzieLet0_1_argbuf_bufchan_buf[0]);
  assign writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb_d = (writeCT$wnnz_IntlizzieLet0_1_argbuf_bufchan_buf[0] ? writeCT$wnnz_IntlizzieLet0_1_argbuf_bufchan_buf :
                                                      writeCT$wnnz_IntlizzieLet0_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnz_IntlizzieLet0_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb_r && writeCT$wnnz_IntlizzieLet0_1_argbuf_bufchan_buf[0]))
        writeCT$wnnz_IntlizzieLet0_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb_r) && (! writeCT$wnnz_IntlizzieLet0_1_argbuf_bufchan_buf[0])))
        writeCT$wnnz_IntlizzieLet0_1_argbuf_bufchan_buf <= writeCT$wnnz_IntlizzieLet0_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz_Int) : (writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb,Pointer_CT$wnnz_Int) > (lizzieLet17_1_argbuf,Pointer_CT$wnnz_Int) */
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb_bufchan_d;
  logic writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb_bufchan_r;
  assign writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb_r = ((! writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb_bufchan_d[0]) || writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb_r)
        writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb_bufchan_d <= writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb_d;
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb_bufchan_buf;
  assign writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb_bufchan_r = (! writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet17_1_argbuf_d = (writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb_bufchan_buf[0] ? writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb_bufchan_buf :
                                   writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                              1'd0};
    else
      if ((lizzieLet17_1_argbuf_r && writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb_bufchan_buf[0]))
        writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
      else if (((! lizzieLet17_1_argbuf_r) && (! writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb_bufchan_buf[0])))
        writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb_bufchan_buf <= writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz_Int) : (writeCT$wnnz_IntlizzieLet26_1_argbuf,Pointer_CT$wnnz_Int) > (writeCT$wnnz_IntlizzieLet26_1_argbuf_rwb,Pointer_CT$wnnz_Int) */
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet26_1_argbuf_bufchan_d;
  logic writeCT$wnnz_IntlizzieLet26_1_argbuf_bufchan_r;
  assign writeCT$wnnz_IntlizzieLet26_1_argbuf_r = ((! writeCT$wnnz_IntlizzieLet26_1_argbuf_bufchan_d[0]) || writeCT$wnnz_IntlizzieLet26_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnz_IntlizzieLet26_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCT$wnnz_IntlizzieLet26_1_argbuf_r)
        writeCT$wnnz_IntlizzieLet26_1_argbuf_bufchan_d <= writeCT$wnnz_IntlizzieLet26_1_argbuf_d;
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet26_1_argbuf_bufchan_buf;
  assign writeCT$wnnz_IntlizzieLet26_1_argbuf_bufchan_r = (! writeCT$wnnz_IntlizzieLet26_1_argbuf_bufchan_buf[0]);
  assign writeCT$wnnz_IntlizzieLet26_1_argbuf_rwb_d = (writeCT$wnnz_IntlizzieLet26_1_argbuf_bufchan_buf[0] ? writeCT$wnnz_IntlizzieLet26_1_argbuf_bufchan_buf :
                                                       writeCT$wnnz_IntlizzieLet26_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnz_IntlizzieLet26_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeCT$wnnz_IntlizzieLet26_1_argbuf_rwb_r && writeCT$wnnz_IntlizzieLet26_1_argbuf_bufchan_buf[0]))
        writeCT$wnnz_IntlizzieLet26_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeCT$wnnz_IntlizzieLet26_1_argbuf_rwb_r) && (! writeCT$wnnz_IntlizzieLet26_1_argbuf_bufchan_buf[0])))
        writeCT$wnnz_IntlizzieLet26_1_argbuf_bufchan_buf <= writeCT$wnnz_IntlizzieLet26_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz_Int) : (writeCT$wnnz_IntlizzieLet26_1_argbuf_rwb,Pointer_CT$wnnz_Int) > (sca2_1_argbuf,Pointer_CT$wnnz_Int) */
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet26_1_argbuf_rwb_bufchan_d;
  logic writeCT$wnnz_IntlizzieLet26_1_argbuf_rwb_bufchan_r;
  assign writeCT$wnnz_IntlizzieLet26_1_argbuf_rwb_r = ((! writeCT$wnnz_IntlizzieLet26_1_argbuf_rwb_bufchan_d[0]) || writeCT$wnnz_IntlizzieLet26_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnz_IntlizzieLet26_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                             1'd0};
    else
      if (writeCT$wnnz_IntlizzieLet26_1_argbuf_rwb_r)
        writeCT$wnnz_IntlizzieLet26_1_argbuf_rwb_bufchan_d <= writeCT$wnnz_IntlizzieLet26_1_argbuf_rwb_d;
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet26_1_argbuf_rwb_bufchan_buf;
  assign writeCT$wnnz_IntlizzieLet26_1_argbuf_rwb_bufchan_r = (! writeCT$wnnz_IntlizzieLet26_1_argbuf_rwb_bufchan_buf[0]);
  assign sca2_1_argbuf_d = (writeCT$wnnz_IntlizzieLet26_1_argbuf_rwb_bufchan_buf[0] ? writeCT$wnnz_IntlizzieLet26_1_argbuf_rwb_bufchan_buf :
                            writeCT$wnnz_IntlizzieLet26_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnz_IntlizzieLet26_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
    else
      if ((sca2_1_argbuf_r && writeCT$wnnz_IntlizzieLet26_1_argbuf_rwb_bufchan_buf[0]))
        writeCT$wnnz_IntlizzieLet26_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                 1'd0};
      else if (((! sca2_1_argbuf_r) && (! writeCT$wnnz_IntlizzieLet26_1_argbuf_rwb_bufchan_buf[0])))
        writeCT$wnnz_IntlizzieLet26_1_argbuf_rwb_bufchan_buf <= writeCT$wnnz_IntlizzieLet26_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz_Int) : (writeCT$wnnz_IntlizzieLet27_1_argbuf,Pointer_CT$wnnz_Int) > (writeCT$wnnz_IntlizzieLet27_1_argbuf_rwb,Pointer_CT$wnnz_Int) */
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet27_1_argbuf_bufchan_d;
  logic writeCT$wnnz_IntlizzieLet27_1_argbuf_bufchan_r;
  assign writeCT$wnnz_IntlizzieLet27_1_argbuf_r = ((! writeCT$wnnz_IntlizzieLet27_1_argbuf_bufchan_d[0]) || writeCT$wnnz_IntlizzieLet27_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnz_IntlizzieLet27_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCT$wnnz_IntlizzieLet27_1_argbuf_r)
        writeCT$wnnz_IntlizzieLet27_1_argbuf_bufchan_d <= writeCT$wnnz_IntlizzieLet27_1_argbuf_d;
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet27_1_argbuf_bufchan_buf;
  assign writeCT$wnnz_IntlizzieLet27_1_argbuf_bufchan_r = (! writeCT$wnnz_IntlizzieLet27_1_argbuf_bufchan_buf[0]);
  assign writeCT$wnnz_IntlizzieLet27_1_argbuf_rwb_d = (writeCT$wnnz_IntlizzieLet27_1_argbuf_bufchan_buf[0] ? writeCT$wnnz_IntlizzieLet27_1_argbuf_bufchan_buf :
                                                       writeCT$wnnz_IntlizzieLet27_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnz_IntlizzieLet27_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeCT$wnnz_IntlizzieLet27_1_argbuf_rwb_r && writeCT$wnnz_IntlizzieLet27_1_argbuf_bufchan_buf[0]))
        writeCT$wnnz_IntlizzieLet27_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeCT$wnnz_IntlizzieLet27_1_argbuf_rwb_r) && (! writeCT$wnnz_IntlizzieLet27_1_argbuf_bufchan_buf[0])))
        writeCT$wnnz_IntlizzieLet27_1_argbuf_bufchan_buf <= writeCT$wnnz_IntlizzieLet27_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz_Int) : (writeCT$wnnz_IntlizzieLet27_1_argbuf_rwb,Pointer_CT$wnnz_Int) > (sca1_1_argbuf,Pointer_CT$wnnz_Int) */
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet27_1_argbuf_rwb_bufchan_d;
  logic writeCT$wnnz_IntlizzieLet27_1_argbuf_rwb_bufchan_r;
  assign writeCT$wnnz_IntlizzieLet27_1_argbuf_rwb_r = ((! writeCT$wnnz_IntlizzieLet27_1_argbuf_rwb_bufchan_d[0]) || writeCT$wnnz_IntlizzieLet27_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnz_IntlizzieLet27_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                             1'd0};
    else
      if (writeCT$wnnz_IntlizzieLet27_1_argbuf_rwb_r)
        writeCT$wnnz_IntlizzieLet27_1_argbuf_rwb_bufchan_d <= writeCT$wnnz_IntlizzieLet27_1_argbuf_rwb_d;
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet27_1_argbuf_rwb_bufchan_buf;
  assign writeCT$wnnz_IntlizzieLet27_1_argbuf_rwb_bufchan_r = (! writeCT$wnnz_IntlizzieLet27_1_argbuf_rwb_bufchan_buf[0]);
  assign sca1_1_argbuf_d = (writeCT$wnnz_IntlizzieLet27_1_argbuf_rwb_bufchan_buf[0] ? writeCT$wnnz_IntlizzieLet27_1_argbuf_rwb_bufchan_buf :
                            writeCT$wnnz_IntlizzieLet27_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnz_IntlizzieLet27_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
    else
      if ((sca1_1_argbuf_r && writeCT$wnnz_IntlizzieLet27_1_argbuf_rwb_bufchan_buf[0]))
        writeCT$wnnz_IntlizzieLet27_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                 1'd0};
      else if (((! sca1_1_argbuf_r) && (! writeCT$wnnz_IntlizzieLet27_1_argbuf_rwb_bufchan_buf[0])))
        writeCT$wnnz_IntlizzieLet27_1_argbuf_rwb_bufchan_buf <= writeCT$wnnz_IntlizzieLet27_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz_Int) : (writeCT$wnnz_IntlizzieLet28_1_argbuf,Pointer_CT$wnnz_Int) > (writeCT$wnnz_IntlizzieLet28_1_argbuf_rwb,Pointer_CT$wnnz_Int) */
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet28_1_argbuf_bufchan_d;
  logic writeCT$wnnz_IntlizzieLet28_1_argbuf_bufchan_r;
  assign writeCT$wnnz_IntlizzieLet28_1_argbuf_r = ((! writeCT$wnnz_IntlizzieLet28_1_argbuf_bufchan_d[0]) || writeCT$wnnz_IntlizzieLet28_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnz_IntlizzieLet28_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCT$wnnz_IntlizzieLet28_1_argbuf_r)
        writeCT$wnnz_IntlizzieLet28_1_argbuf_bufchan_d <= writeCT$wnnz_IntlizzieLet28_1_argbuf_d;
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet28_1_argbuf_bufchan_buf;
  assign writeCT$wnnz_IntlizzieLet28_1_argbuf_bufchan_r = (! writeCT$wnnz_IntlizzieLet28_1_argbuf_bufchan_buf[0]);
  assign writeCT$wnnz_IntlizzieLet28_1_argbuf_rwb_d = (writeCT$wnnz_IntlizzieLet28_1_argbuf_bufchan_buf[0] ? writeCT$wnnz_IntlizzieLet28_1_argbuf_bufchan_buf :
                                                       writeCT$wnnz_IntlizzieLet28_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnz_IntlizzieLet28_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeCT$wnnz_IntlizzieLet28_1_argbuf_rwb_r && writeCT$wnnz_IntlizzieLet28_1_argbuf_bufchan_buf[0]))
        writeCT$wnnz_IntlizzieLet28_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeCT$wnnz_IntlizzieLet28_1_argbuf_rwb_r) && (! writeCT$wnnz_IntlizzieLet28_1_argbuf_bufchan_buf[0])))
        writeCT$wnnz_IntlizzieLet28_1_argbuf_bufchan_buf <= writeCT$wnnz_IntlizzieLet28_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz_Int) : (writeCT$wnnz_IntlizzieLet28_1_argbuf_rwb,Pointer_CT$wnnz_Int) > (sca0_1_argbuf,Pointer_CT$wnnz_Int) */
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet28_1_argbuf_rwb_bufchan_d;
  logic writeCT$wnnz_IntlizzieLet28_1_argbuf_rwb_bufchan_r;
  assign writeCT$wnnz_IntlizzieLet28_1_argbuf_rwb_r = ((! writeCT$wnnz_IntlizzieLet28_1_argbuf_rwb_bufchan_d[0]) || writeCT$wnnz_IntlizzieLet28_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnz_IntlizzieLet28_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                             1'd0};
    else
      if (writeCT$wnnz_IntlizzieLet28_1_argbuf_rwb_r)
        writeCT$wnnz_IntlizzieLet28_1_argbuf_rwb_bufchan_d <= writeCT$wnnz_IntlizzieLet28_1_argbuf_rwb_d;
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet28_1_argbuf_rwb_bufchan_buf;
  assign writeCT$wnnz_IntlizzieLet28_1_argbuf_rwb_bufchan_r = (! writeCT$wnnz_IntlizzieLet28_1_argbuf_rwb_bufchan_buf[0]);
  assign sca0_1_argbuf_d = (writeCT$wnnz_IntlizzieLet28_1_argbuf_rwb_bufchan_buf[0] ? writeCT$wnnz_IntlizzieLet28_1_argbuf_rwb_bufchan_buf :
                            writeCT$wnnz_IntlizzieLet28_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnz_IntlizzieLet28_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
    else
      if ((sca0_1_argbuf_r && writeCT$wnnz_IntlizzieLet28_1_argbuf_rwb_bufchan_buf[0]))
        writeCT$wnnz_IntlizzieLet28_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                 1'd0};
      else if (((! sca0_1_argbuf_r) && (! writeCT$wnnz_IntlizzieLet28_1_argbuf_rwb_bufchan_buf[0])))
        writeCT$wnnz_IntlizzieLet28_1_argbuf_rwb_bufchan_buf <= writeCT$wnnz_IntlizzieLet28_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz_Int) : (writeCT$wnnz_IntlizzieLet5_1_argbuf,Pointer_CT$wnnz_Int) > (writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb,Pointer_CT$wnnz_Int) */
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet5_1_argbuf_bufchan_d;
  logic writeCT$wnnz_IntlizzieLet5_1_argbuf_bufchan_r;
  assign writeCT$wnnz_IntlizzieLet5_1_argbuf_r = ((! writeCT$wnnz_IntlizzieLet5_1_argbuf_bufchan_d[0]) || writeCT$wnnz_IntlizzieLet5_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnz_IntlizzieLet5_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCT$wnnz_IntlizzieLet5_1_argbuf_r)
        writeCT$wnnz_IntlizzieLet5_1_argbuf_bufchan_d <= writeCT$wnnz_IntlizzieLet5_1_argbuf_d;
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet5_1_argbuf_bufchan_buf;
  assign writeCT$wnnz_IntlizzieLet5_1_argbuf_bufchan_r = (! writeCT$wnnz_IntlizzieLet5_1_argbuf_bufchan_buf[0]);
  assign writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb_d = (writeCT$wnnz_IntlizzieLet5_1_argbuf_bufchan_buf[0] ? writeCT$wnnz_IntlizzieLet5_1_argbuf_bufchan_buf :
                                                      writeCT$wnnz_IntlizzieLet5_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnz_IntlizzieLet5_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb_r && writeCT$wnnz_IntlizzieLet5_1_argbuf_bufchan_buf[0]))
        writeCT$wnnz_IntlizzieLet5_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb_r) && (! writeCT$wnnz_IntlizzieLet5_1_argbuf_bufchan_buf[0])))
        writeCT$wnnz_IntlizzieLet5_1_argbuf_bufchan_buf <= writeCT$wnnz_IntlizzieLet5_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz_Int) : (writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb,Pointer_CT$wnnz_Int) > (sca3_1_argbuf,Pointer_CT$wnnz_Int) */
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb_bufchan_d;
  logic writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb_bufchan_r;
  assign writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb_r = ((! writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb_bufchan_d[0]) || writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb_r)
        writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb_bufchan_d <= writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb_d;
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb_bufchan_buf;
  assign writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb_bufchan_r = (! writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb_bufchan_buf[0]);
  assign sca3_1_argbuf_d = (writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb_bufchan_buf[0] ? writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb_bufchan_buf :
                            writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                              1'd0};
    else
      if ((sca3_1_argbuf_r && writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb_bufchan_buf[0]))
        writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
      else if (((! sca3_1_argbuf_r) && (! writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb_bufchan_buf[0])))
        writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb_bufchan_buf <= writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CTkron_kron_Int_Int_Int) : (writeCTkron_kron_Int_Int_IntlizzieLet22_1_argbuf,Pointer_CTkron_kron_Int_Int_Int) > (writeCTkron_kron_Int_Int_IntlizzieLet22_1_argbuf_rwb,Pointer_CTkron_kron_Int_Int_Int) */
  Pointer_CTkron_kron_Int_Int_Int_t writeCTkron_kron_Int_Int_IntlizzieLet22_1_argbuf_bufchan_d;
  logic writeCTkron_kron_Int_Int_IntlizzieLet22_1_argbuf_bufchan_r;
  assign writeCTkron_kron_Int_Int_IntlizzieLet22_1_argbuf_r = ((! writeCTkron_kron_Int_Int_IntlizzieLet22_1_argbuf_bufchan_d[0]) || writeCTkron_kron_Int_Int_IntlizzieLet22_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTkron_kron_Int_Int_IntlizzieLet22_1_argbuf_bufchan_d <= {16'd0,
                                                                     1'd0};
    else
      if (writeCTkron_kron_Int_Int_IntlizzieLet22_1_argbuf_r)
        writeCTkron_kron_Int_Int_IntlizzieLet22_1_argbuf_bufchan_d <= writeCTkron_kron_Int_Int_IntlizzieLet22_1_argbuf_d;
  Pointer_CTkron_kron_Int_Int_Int_t writeCTkron_kron_Int_Int_IntlizzieLet22_1_argbuf_bufchan_buf;
  assign writeCTkron_kron_Int_Int_IntlizzieLet22_1_argbuf_bufchan_r = (! writeCTkron_kron_Int_Int_IntlizzieLet22_1_argbuf_bufchan_buf[0]);
  assign writeCTkron_kron_Int_Int_IntlizzieLet22_1_argbuf_rwb_d = (writeCTkron_kron_Int_Int_IntlizzieLet22_1_argbuf_bufchan_buf[0] ? writeCTkron_kron_Int_Int_IntlizzieLet22_1_argbuf_bufchan_buf :
                                                                   writeCTkron_kron_Int_Int_IntlizzieLet22_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTkron_kron_Int_Int_IntlizzieLet22_1_argbuf_bufchan_buf <= {16'd0,
                                                                       1'd0};
    else
      if ((writeCTkron_kron_Int_Int_IntlizzieLet22_1_argbuf_rwb_r && writeCTkron_kron_Int_Int_IntlizzieLet22_1_argbuf_bufchan_buf[0]))
        writeCTkron_kron_Int_Int_IntlizzieLet22_1_argbuf_bufchan_buf <= {16'd0,
                                                                         1'd0};
      else if (((! writeCTkron_kron_Int_Int_IntlizzieLet22_1_argbuf_rwb_r) && (! writeCTkron_kron_Int_Int_IntlizzieLet22_1_argbuf_bufchan_buf[0])))
        writeCTkron_kron_Int_Int_IntlizzieLet22_1_argbuf_bufchan_buf <= writeCTkron_kron_Int_Int_IntlizzieLet22_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CTkron_kron_Int_Int_Int) : (writeCTkron_kron_Int_Int_IntlizzieLet22_1_argbuf_rwb,Pointer_CTkron_kron_Int_Int_Int) > (lizzieLet14_1_1_argbuf,Pointer_CTkron_kron_Int_Int_Int) */
  Pointer_CTkron_kron_Int_Int_Int_t writeCTkron_kron_Int_Int_IntlizzieLet22_1_argbuf_rwb_bufchan_d;
  logic writeCTkron_kron_Int_Int_IntlizzieLet22_1_argbuf_rwb_bufchan_r;
  assign writeCTkron_kron_Int_Int_IntlizzieLet22_1_argbuf_rwb_r = ((! writeCTkron_kron_Int_Int_IntlizzieLet22_1_argbuf_rwb_bufchan_d[0]) || writeCTkron_kron_Int_Int_IntlizzieLet22_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTkron_kron_Int_Int_IntlizzieLet22_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                                         1'd0};
    else
      if (writeCTkron_kron_Int_Int_IntlizzieLet22_1_argbuf_rwb_r)
        writeCTkron_kron_Int_Int_IntlizzieLet22_1_argbuf_rwb_bufchan_d <= writeCTkron_kron_Int_Int_IntlizzieLet22_1_argbuf_rwb_d;
  Pointer_CTkron_kron_Int_Int_Int_t writeCTkron_kron_Int_Int_IntlizzieLet22_1_argbuf_rwb_bufchan_buf;
  assign writeCTkron_kron_Int_Int_IntlizzieLet22_1_argbuf_rwb_bufchan_r = (! writeCTkron_kron_Int_Int_IntlizzieLet22_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet14_1_1_argbuf_d = (writeCTkron_kron_Int_Int_IntlizzieLet22_1_argbuf_rwb_bufchan_buf[0] ? writeCTkron_kron_Int_Int_IntlizzieLet22_1_argbuf_rwb_bufchan_buf :
                                     writeCTkron_kron_Int_Int_IntlizzieLet22_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTkron_kron_Int_Int_IntlizzieLet22_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                           1'd0};
    else
      if ((lizzieLet14_1_1_argbuf_r && writeCTkron_kron_Int_Int_IntlizzieLet22_1_argbuf_rwb_bufchan_buf[0]))
        writeCTkron_kron_Int_Int_IntlizzieLet22_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                             1'd0};
      else if (((! lizzieLet14_1_1_argbuf_r) && (! writeCTkron_kron_Int_Int_IntlizzieLet22_1_argbuf_rwb_bufchan_buf[0])))
        writeCTkron_kron_Int_Int_IntlizzieLet22_1_argbuf_rwb_bufchan_buf <= writeCTkron_kron_Int_Int_IntlizzieLet22_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CTkron_kron_Int_Int_Int) : (writeCTkron_kron_Int_Int_IntlizzieLet30_1_argbuf,Pointer_CTkron_kron_Int_Int_Int) > (writeCTkron_kron_Int_Int_IntlizzieLet30_1_argbuf_rwb,Pointer_CTkron_kron_Int_Int_Int) */
  Pointer_CTkron_kron_Int_Int_Int_t writeCTkron_kron_Int_Int_IntlizzieLet30_1_argbuf_bufchan_d;
  logic writeCTkron_kron_Int_Int_IntlizzieLet30_1_argbuf_bufchan_r;
  assign writeCTkron_kron_Int_Int_IntlizzieLet30_1_argbuf_r = ((! writeCTkron_kron_Int_Int_IntlizzieLet30_1_argbuf_bufchan_d[0]) || writeCTkron_kron_Int_Int_IntlizzieLet30_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTkron_kron_Int_Int_IntlizzieLet30_1_argbuf_bufchan_d <= {16'd0,
                                                                     1'd0};
    else
      if (writeCTkron_kron_Int_Int_IntlizzieLet30_1_argbuf_r)
        writeCTkron_kron_Int_Int_IntlizzieLet30_1_argbuf_bufchan_d <= writeCTkron_kron_Int_Int_IntlizzieLet30_1_argbuf_d;
  Pointer_CTkron_kron_Int_Int_Int_t writeCTkron_kron_Int_Int_IntlizzieLet30_1_argbuf_bufchan_buf;
  assign writeCTkron_kron_Int_Int_IntlizzieLet30_1_argbuf_bufchan_r = (! writeCTkron_kron_Int_Int_IntlizzieLet30_1_argbuf_bufchan_buf[0]);
  assign writeCTkron_kron_Int_Int_IntlizzieLet30_1_argbuf_rwb_d = (writeCTkron_kron_Int_Int_IntlizzieLet30_1_argbuf_bufchan_buf[0] ? writeCTkron_kron_Int_Int_IntlizzieLet30_1_argbuf_bufchan_buf :
                                                                   writeCTkron_kron_Int_Int_IntlizzieLet30_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTkron_kron_Int_Int_IntlizzieLet30_1_argbuf_bufchan_buf <= {16'd0,
                                                                       1'd0};
    else
      if ((writeCTkron_kron_Int_Int_IntlizzieLet30_1_argbuf_rwb_r && writeCTkron_kron_Int_Int_IntlizzieLet30_1_argbuf_bufchan_buf[0]))
        writeCTkron_kron_Int_Int_IntlizzieLet30_1_argbuf_bufchan_buf <= {16'd0,
                                                                         1'd0};
      else if (((! writeCTkron_kron_Int_Int_IntlizzieLet30_1_argbuf_rwb_r) && (! writeCTkron_kron_Int_Int_IntlizzieLet30_1_argbuf_bufchan_buf[0])))
        writeCTkron_kron_Int_Int_IntlizzieLet30_1_argbuf_bufchan_buf <= writeCTkron_kron_Int_Int_IntlizzieLet30_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CTkron_kron_Int_Int_Int) : (writeCTkron_kron_Int_Int_IntlizzieLet30_1_argbuf_rwb,Pointer_CTkron_kron_Int_Int_Int) > (sca2_1_1_argbuf,Pointer_CTkron_kron_Int_Int_Int) */
  Pointer_CTkron_kron_Int_Int_Int_t writeCTkron_kron_Int_Int_IntlizzieLet30_1_argbuf_rwb_bufchan_d;
  logic writeCTkron_kron_Int_Int_IntlizzieLet30_1_argbuf_rwb_bufchan_r;
  assign writeCTkron_kron_Int_Int_IntlizzieLet30_1_argbuf_rwb_r = ((! writeCTkron_kron_Int_Int_IntlizzieLet30_1_argbuf_rwb_bufchan_d[0]) || writeCTkron_kron_Int_Int_IntlizzieLet30_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTkron_kron_Int_Int_IntlizzieLet30_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                                         1'd0};
    else
      if (writeCTkron_kron_Int_Int_IntlizzieLet30_1_argbuf_rwb_r)
        writeCTkron_kron_Int_Int_IntlizzieLet30_1_argbuf_rwb_bufchan_d <= writeCTkron_kron_Int_Int_IntlizzieLet30_1_argbuf_rwb_d;
  Pointer_CTkron_kron_Int_Int_Int_t writeCTkron_kron_Int_Int_IntlizzieLet30_1_argbuf_rwb_bufchan_buf;
  assign writeCTkron_kron_Int_Int_IntlizzieLet30_1_argbuf_rwb_bufchan_r = (! writeCTkron_kron_Int_Int_IntlizzieLet30_1_argbuf_rwb_bufchan_buf[0]);
  assign sca2_1_1_argbuf_d = (writeCTkron_kron_Int_Int_IntlizzieLet30_1_argbuf_rwb_bufchan_buf[0] ? writeCTkron_kron_Int_Int_IntlizzieLet30_1_argbuf_rwb_bufchan_buf :
                              writeCTkron_kron_Int_Int_IntlizzieLet30_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTkron_kron_Int_Int_IntlizzieLet30_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                           1'd0};
    else
      if ((sca2_1_1_argbuf_r && writeCTkron_kron_Int_Int_IntlizzieLet30_1_argbuf_rwb_bufchan_buf[0]))
        writeCTkron_kron_Int_Int_IntlizzieLet30_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                             1'd0};
      else if (((! sca2_1_1_argbuf_r) && (! writeCTkron_kron_Int_Int_IntlizzieLet30_1_argbuf_rwb_bufchan_buf[0])))
        writeCTkron_kron_Int_Int_IntlizzieLet30_1_argbuf_rwb_bufchan_buf <= writeCTkron_kron_Int_Int_IntlizzieLet30_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CTkron_kron_Int_Int_Int) : (writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf,Pointer_CTkron_kron_Int_Int_Int) > (writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf_rwb,Pointer_CTkron_kron_Int_Int_Int) */
  Pointer_CTkron_kron_Int_Int_Int_t writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf_bufchan_d;
  logic writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf_bufchan_r;
  assign writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf_r = ((! writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf_bufchan_d[0]) || writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf_bufchan_d <= {16'd0,
                                                                     1'd0};
    else
      if (writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf_r)
        writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf_bufchan_d <= writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf_d;
  Pointer_CTkron_kron_Int_Int_Int_t writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf_bufchan_buf;
  assign writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf_bufchan_r = (! writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf_bufchan_buf[0]);
  assign writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf_rwb_d = (writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf_bufchan_buf[0] ? writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf_bufchan_buf :
                                                                   writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf_bufchan_buf <= {16'd0,
                                                                       1'd0};
    else
      if ((writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf_rwb_r && writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf_bufchan_buf[0]))
        writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf_bufchan_buf <= {16'd0,
                                                                         1'd0};
      else if (((! writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf_rwb_r) && (! writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf_bufchan_buf[0])))
        writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf_bufchan_buf <= writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CTkron_kron_Int_Int_Int) : (writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf_rwb,Pointer_CTkron_kron_Int_Int_Int) > (sca1_1_1_argbuf,Pointer_CTkron_kron_Int_Int_Int) */
  Pointer_CTkron_kron_Int_Int_Int_t writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf_rwb_bufchan_d;
  logic writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf_rwb_bufchan_r;
  assign writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf_rwb_r = ((! writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf_rwb_bufchan_d[0]) || writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                                         1'd0};
    else
      if (writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf_rwb_r)
        writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf_rwb_bufchan_d <= writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf_rwb_d;
  Pointer_CTkron_kron_Int_Int_Int_t writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf_rwb_bufchan_buf;
  assign writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf_rwb_bufchan_r = (! writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf_rwb_bufchan_buf[0]);
  assign sca1_1_1_argbuf_d = (writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf_rwb_bufchan_buf[0] ? writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf_rwb_bufchan_buf :
                              writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                           1'd0};
    else
      if ((sca1_1_1_argbuf_r && writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf_rwb_bufchan_buf[0]))
        writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                             1'd0};
      else if (((! sca1_1_1_argbuf_r) && (! writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf_rwb_bufchan_buf[0])))
        writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf_rwb_bufchan_buf <= writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CTkron_kron_Int_Int_Int) : (writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf,Pointer_CTkron_kron_Int_Int_Int) > (writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf_rwb,Pointer_CTkron_kron_Int_Int_Int) */
  Pointer_CTkron_kron_Int_Int_Int_t writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf_bufchan_d;
  logic writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf_bufchan_r;
  assign writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf_r = ((! writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf_bufchan_d[0]) || writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf_bufchan_d <= {16'd0,
                                                                     1'd0};
    else
      if (writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf_r)
        writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf_bufchan_d <= writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf_d;
  Pointer_CTkron_kron_Int_Int_Int_t writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf_bufchan_buf;
  assign writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf_bufchan_r = (! writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf_bufchan_buf[0]);
  assign writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf_rwb_d = (writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf_bufchan_buf[0] ? writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf_bufchan_buf :
                                                                   writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf_bufchan_buf <= {16'd0,
                                                                       1'd0};
    else
      if ((writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf_rwb_r && writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf_bufchan_buf[0]))
        writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf_bufchan_buf <= {16'd0,
                                                                         1'd0};
      else if (((! writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf_rwb_r) && (! writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf_bufchan_buf[0])))
        writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf_bufchan_buf <= writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CTkron_kron_Int_Int_Int) : (writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf_rwb,Pointer_CTkron_kron_Int_Int_Int) > (sca0_1_1_argbuf,Pointer_CTkron_kron_Int_Int_Int) */
  Pointer_CTkron_kron_Int_Int_Int_t writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf_rwb_bufchan_d;
  logic writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf_rwb_bufchan_r;
  assign writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf_rwb_r = ((! writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf_rwb_bufchan_d[0]) || writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                                         1'd0};
    else
      if (writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf_rwb_r)
        writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf_rwb_bufchan_d <= writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf_rwb_d;
  Pointer_CTkron_kron_Int_Int_Int_t writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf_rwb_bufchan_buf;
  assign writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf_rwb_bufchan_r = (! writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf_rwb_bufchan_buf[0]);
  assign sca0_1_1_argbuf_d = (writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf_rwb_bufchan_buf[0] ? writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf_rwb_bufchan_buf :
                              writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                           1'd0};
    else
      if ((sca0_1_1_argbuf_r && writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf_rwb_bufchan_buf[0]))
        writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                             1'd0};
      else if (((! sca0_1_1_argbuf_r) && (! writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf_rwb_bufchan_buf[0])))
        writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf_rwb_bufchan_buf <= writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CTkron_kron_Int_Int_Int) : (writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf,Pointer_CTkron_kron_Int_Int_Int) > (writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf_rwb,Pointer_CTkron_kron_Int_Int_Int) */
  Pointer_CTkron_kron_Int_Int_Int_t writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf_bufchan_d;
  logic writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf_bufchan_r;
  assign writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf_r = ((! writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf_bufchan_d[0]) || writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf_bufchan_d <= {16'd0,
                                                                    1'd0};
    else
      if (writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf_r)
        writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf_bufchan_d <= writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf_d;
  Pointer_CTkron_kron_Int_Int_Int_t writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf_bufchan_buf;
  assign writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf_bufchan_r = (! writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf_bufchan_buf[0]);
  assign writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf_rwb_d = (writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf_bufchan_buf[0] ? writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf_bufchan_buf :
                                                                  writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf_bufchan_buf <= {16'd0,
                                                                      1'd0};
    else
      if ((writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf_rwb_r && writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf_bufchan_buf[0]))
        writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf_bufchan_buf <= {16'd0,
                                                                        1'd0};
      else if (((! writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf_rwb_r) && (! writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf_bufchan_buf[0])))
        writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf_bufchan_buf <= writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CTkron_kron_Int_Int_Int) : (writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf_rwb,Pointer_CTkron_kron_Int_Int_Int) > (sca3_1_1_argbuf,Pointer_CTkron_kron_Int_Int_Int) */
  Pointer_CTkron_kron_Int_Int_Int_t writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf_rwb_bufchan_d;
  logic writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf_rwb_bufchan_r;
  assign writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf_rwb_r = ((! writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf_rwb_bufchan_d[0]) || writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                                        1'd0};
    else
      if (writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf_rwb_r)
        writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf_rwb_bufchan_d <= writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf_rwb_d;
  Pointer_CTkron_kron_Int_Int_Int_t writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf_rwb_bufchan_buf;
  assign writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf_rwb_bufchan_r = (! writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf_rwb_bufchan_buf[0]);
  assign sca3_1_1_argbuf_d = (writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf_rwb_bufchan_buf[0] ? writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf_rwb_bufchan_buf :
                              writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                          1'd0};
    else
      if ((sca3_1_1_argbuf_r && writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf_rwb_bufchan_buf[0]))
        writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                            1'd0};
      else if (((! sca3_1_1_argbuf_r) && (! writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf_rwb_bufchan_buf[0])))
        writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf_rwb_bufchan_buf <= writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CTmain_map'_Int_Int) : (writeCTmain_map'_Int_IntlizzieLet14_1_argbuf,Pointer_CTmain_map'_Int_Int) > (writeCTmain_map'_Int_IntlizzieLet14_1_argbuf_rwb,Pointer_CTmain_map'_Int_Int) */
  \Pointer_CTmain_map'_Int_Int_t  \writeCTmain_map'_Int_IntlizzieLet14_1_argbuf_bufchan_d ;
  logic \writeCTmain_map'_Int_IntlizzieLet14_1_argbuf_bufchan_r ;
  assign \writeCTmain_map'_Int_IntlizzieLet14_1_argbuf_r  = ((! \writeCTmain_map'_Int_IntlizzieLet14_1_argbuf_bufchan_d [0]) || \writeCTmain_map'_Int_IntlizzieLet14_1_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmain_map'_Int_IntlizzieLet14_1_argbuf_bufchan_d  <= {16'd0,
                                                                   1'd0};
    else
      if (\writeCTmain_map'_Int_IntlizzieLet14_1_argbuf_r )
        \writeCTmain_map'_Int_IntlizzieLet14_1_argbuf_bufchan_d  <= \writeCTmain_map'_Int_IntlizzieLet14_1_argbuf_d ;
  \Pointer_CTmain_map'_Int_Int_t  \writeCTmain_map'_Int_IntlizzieLet14_1_argbuf_bufchan_buf ;
  assign \writeCTmain_map'_Int_IntlizzieLet14_1_argbuf_bufchan_r  = (! \writeCTmain_map'_Int_IntlizzieLet14_1_argbuf_bufchan_buf [0]);
  assign \writeCTmain_map'_Int_IntlizzieLet14_1_argbuf_rwb_d  = (\writeCTmain_map'_Int_IntlizzieLet14_1_argbuf_bufchan_buf [0] ? \writeCTmain_map'_Int_IntlizzieLet14_1_argbuf_bufchan_buf  :
                                                                 \writeCTmain_map'_Int_IntlizzieLet14_1_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmain_map'_Int_IntlizzieLet14_1_argbuf_bufchan_buf  <= {16'd0,
                                                                     1'd0};
    else
      if ((\writeCTmain_map'_Int_IntlizzieLet14_1_argbuf_rwb_r  && \writeCTmain_map'_Int_IntlizzieLet14_1_argbuf_bufchan_buf [0]))
        \writeCTmain_map'_Int_IntlizzieLet14_1_argbuf_bufchan_buf  <= {16'd0,
                                                                       1'd0};
      else if (((! \writeCTmain_map'_Int_IntlizzieLet14_1_argbuf_rwb_r ) && (! \writeCTmain_map'_Int_IntlizzieLet14_1_argbuf_bufchan_buf [0])))
        \writeCTmain_map'_Int_IntlizzieLet14_1_argbuf_bufchan_buf  <= \writeCTmain_map'_Int_IntlizzieLet14_1_argbuf_bufchan_d ;
  
  /* buf (Ty Pointer_CTmain_map'_Int_Int) : (writeCTmain_map'_Int_IntlizzieLet14_1_argbuf_rwb,Pointer_CTmain_map'_Int_Int) > (sca3_2_1_argbuf,Pointer_CTmain_map'_Int_Int) */
  \Pointer_CTmain_map'_Int_Int_t  \writeCTmain_map'_Int_IntlizzieLet14_1_argbuf_rwb_bufchan_d ;
  logic \writeCTmain_map'_Int_IntlizzieLet14_1_argbuf_rwb_bufchan_r ;
  assign \writeCTmain_map'_Int_IntlizzieLet14_1_argbuf_rwb_r  = ((! \writeCTmain_map'_Int_IntlizzieLet14_1_argbuf_rwb_bufchan_d [0]) || \writeCTmain_map'_Int_IntlizzieLet14_1_argbuf_rwb_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmain_map'_Int_IntlizzieLet14_1_argbuf_rwb_bufchan_d  <= {16'd0,
                                                                       1'd0};
    else
      if (\writeCTmain_map'_Int_IntlizzieLet14_1_argbuf_rwb_r )
        \writeCTmain_map'_Int_IntlizzieLet14_1_argbuf_rwb_bufchan_d  <= \writeCTmain_map'_Int_IntlizzieLet14_1_argbuf_rwb_d ;
  \Pointer_CTmain_map'_Int_Int_t  \writeCTmain_map'_Int_IntlizzieLet14_1_argbuf_rwb_bufchan_buf ;
  assign \writeCTmain_map'_Int_IntlizzieLet14_1_argbuf_rwb_bufchan_r  = (! \writeCTmain_map'_Int_IntlizzieLet14_1_argbuf_rwb_bufchan_buf [0]);
  assign sca3_2_1_argbuf_d = (\writeCTmain_map'_Int_IntlizzieLet14_1_argbuf_rwb_bufchan_buf [0] ? \writeCTmain_map'_Int_IntlizzieLet14_1_argbuf_rwb_bufchan_buf  :
                              \writeCTmain_map'_Int_IntlizzieLet14_1_argbuf_rwb_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmain_map'_Int_IntlizzieLet14_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                         1'd0};
    else
      if ((sca3_2_1_argbuf_r && \writeCTmain_map'_Int_IntlizzieLet14_1_argbuf_rwb_bufchan_buf [0]))
        \writeCTmain_map'_Int_IntlizzieLet14_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                           1'd0};
      else if (((! sca3_2_1_argbuf_r) && (! \writeCTmain_map'_Int_IntlizzieLet14_1_argbuf_rwb_bufchan_buf [0])))
        \writeCTmain_map'_Int_IntlizzieLet14_1_argbuf_rwb_bufchan_buf  <= \writeCTmain_map'_Int_IntlizzieLet14_1_argbuf_rwb_bufchan_d ;
  
  /* buf (Ty Pointer_CTmain_map'_Int_Int) : (writeCTmain_map'_Int_IntlizzieLet23_1_argbuf,Pointer_CTmain_map'_Int_Int) > (writeCTmain_map'_Int_IntlizzieLet23_1_argbuf_rwb,Pointer_CTmain_map'_Int_Int) */
  \Pointer_CTmain_map'_Int_Int_t  \writeCTmain_map'_Int_IntlizzieLet23_1_argbuf_bufchan_d ;
  logic \writeCTmain_map'_Int_IntlizzieLet23_1_argbuf_bufchan_r ;
  assign \writeCTmain_map'_Int_IntlizzieLet23_1_argbuf_r  = ((! \writeCTmain_map'_Int_IntlizzieLet23_1_argbuf_bufchan_d [0]) || \writeCTmain_map'_Int_IntlizzieLet23_1_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmain_map'_Int_IntlizzieLet23_1_argbuf_bufchan_d  <= {16'd0,
                                                                   1'd0};
    else
      if (\writeCTmain_map'_Int_IntlizzieLet23_1_argbuf_r )
        \writeCTmain_map'_Int_IntlizzieLet23_1_argbuf_bufchan_d  <= \writeCTmain_map'_Int_IntlizzieLet23_1_argbuf_d ;
  \Pointer_CTmain_map'_Int_Int_t  \writeCTmain_map'_Int_IntlizzieLet23_1_argbuf_bufchan_buf ;
  assign \writeCTmain_map'_Int_IntlizzieLet23_1_argbuf_bufchan_r  = (! \writeCTmain_map'_Int_IntlizzieLet23_1_argbuf_bufchan_buf [0]);
  assign \writeCTmain_map'_Int_IntlizzieLet23_1_argbuf_rwb_d  = (\writeCTmain_map'_Int_IntlizzieLet23_1_argbuf_bufchan_buf [0] ? \writeCTmain_map'_Int_IntlizzieLet23_1_argbuf_bufchan_buf  :
                                                                 \writeCTmain_map'_Int_IntlizzieLet23_1_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmain_map'_Int_IntlizzieLet23_1_argbuf_bufchan_buf  <= {16'd0,
                                                                     1'd0};
    else
      if ((\writeCTmain_map'_Int_IntlizzieLet23_1_argbuf_rwb_r  && \writeCTmain_map'_Int_IntlizzieLet23_1_argbuf_bufchan_buf [0]))
        \writeCTmain_map'_Int_IntlizzieLet23_1_argbuf_bufchan_buf  <= {16'd0,
                                                                       1'd0};
      else if (((! \writeCTmain_map'_Int_IntlizzieLet23_1_argbuf_rwb_r ) && (! \writeCTmain_map'_Int_IntlizzieLet23_1_argbuf_bufchan_buf [0])))
        \writeCTmain_map'_Int_IntlizzieLet23_1_argbuf_bufchan_buf  <= \writeCTmain_map'_Int_IntlizzieLet23_1_argbuf_bufchan_d ;
  
  /* buf (Ty Pointer_CTmain_map'_Int_Int) : (writeCTmain_map'_Int_IntlizzieLet23_1_argbuf_rwb,Pointer_CTmain_map'_Int_Int) > (lizzieLet5_1_1_argbuf,Pointer_CTmain_map'_Int_Int) */
  \Pointer_CTmain_map'_Int_Int_t  \writeCTmain_map'_Int_IntlizzieLet23_1_argbuf_rwb_bufchan_d ;
  logic \writeCTmain_map'_Int_IntlizzieLet23_1_argbuf_rwb_bufchan_r ;
  assign \writeCTmain_map'_Int_IntlizzieLet23_1_argbuf_rwb_r  = ((! \writeCTmain_map'_Int_IntlizzieLet23_1_argbuf_rwb_bufchan_d [0]) || \writeCTmain_map'_Int_IntlizzieLet23_1_argbuf_rwb_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmain_map'_Int_IntlizzieLet23_1_argbuf_rwb_bufchan_d  <= {16'd0,
                                                                       1'd0};
    else
      if (\writeCTmain_map'_Int_IntlizzieLet23_1_argbuf_rwb_r )
        \writeCTmain_map'_Int_IntlizzieLet23_1_argbuf_rwb_bufchan_d  <= \writeCTmain_map'_Int_IntlizzieLet23_1_argbuf_rwb_d ;
  \Pointer_CTmain_map'_Int_Int_t  \writeCTmain_map'_Int_IntlizzieLet23_1_argbuf_rwb_bufchan_buf ;
  assign \writeCTmain_map'_Int_IntlizzieLet23_1_argbuf_rwb_bufchan_r  = (! \writeCTmain_map'_Int_IntlizzieLet23_1_argbuf_rwb_bufchan_buf [0]);
  assign lizzieLet5_1_1_argbuf_d = (\writeCTmain_map'_Int_IntlizzieLet23_1_argbuf_rwb_bufchan_buf [0] ? \writeCTmain_map'_Int_IntlizzieLet23_1_argbuf_rwb_bufchan_buf  :
                                    \writeCTmain_map'_Int_IntlizzieLet23_1_argbuf_rwb_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmain_map'_Int_IntlizzieLet23_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                         1'd0};
    else
      if ((lizzieLet5_1_1_argbuf_r && \writeCTmain_map'_Int_IntlizzieLet23_1_argbuf_rwb_bufchan_buf [0]))
        \writeCTmain_map'_Int_IntlizzieLet23_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                           1'd0};
      else if (((! lizzieLet5_1_1_argbuf_r) && (! \writeCTmain_map'_Int_IntlizzieLet23_1_argbuf_rwb_bufchan_buf [0])))
        \writeCTmain_map'_Int_IntlizzieLet23_1_argbuf_rwb_bufchan_buf  <= \writeCTmain_map'_Int_IntlizzieLet23_1_argbuf_rwb_bufchan_d ;
  
  /* buf (Ty Pointer_CTmain_map'_Int_Int) : (writeCTmain_map'_Int_IntlizzieLet35_1_argbuf,Pointer_CTmain_map'_Int_Int) > (writeCTmain_map'_Int_IntlizzieLet35_1_argbuf_rwb,Pointer_CTmain_map'_Int_Int) */
  \Pointer_CTmain_map'_Int_Int_t  \writeCTmain_map'_Int_IntlizzieLet35_1_argbuf_bufchan_d ;
  logic \writeCTmain_map'_Int_IntlizzieLet35_1_argbuf_bufchan_r ;
  assign \writeCTmain_map'_Int_IntlizzieLet35_1_argbuf_r  = ((! \writeCTmain_map'_Int_IntlizzieLet35_1_argbuf_bufchan_d [0]) || \writeCTmain_map'_Int_IntlizzieLet35_1_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmain_map'_Int_IntlizzieLet35_1_argbuf_bufchan_d  <= {16'd0,
                                                                   1'd0};
    else
      if (\writeCTmain_map'_Int_IntlizzieLet35_1_argbuf_r )
        \writeCTmain_map'_Int_IntlizzieLet35_1_argbuf_bufchan_d  <= \writeCTmain_map'_Int_IntlizzieLet35_1_argbuf_d ;
  \Pointer_CTmain_map'_Int_Int_t  \writeCTmain_map'_Int_IntlizzieLet35_1_argbuf_bufchan_buf ;
  assign \writeCTmain_map'_Int_IntlizzieLet35_1_argbuf_bufchan_r  = (! \writeCTmain_map'_Int_IntlizzieLet35_1_argbuf_bufchan_buf [0]);
  assign \writeCTmain_map'_Int_IntlizzieLet35_1_argbuf_rwb_d  = (\writeCTmain_map'_Int_IntlizzieLet35_1_argbuf_bufchan_buf [0] ? \writeCTmain_map'_Int_IntlizzieLet35_1_argbuf_bufchan_buf  :
                                                                 \writeCTmain_map'_Int_IntlizzieLet35_1_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmain_map'_Int_IntlizzieLet35_1_argbuf_bufchan_buf  <= {16'd0,
                                                                     1'd0};
    else
      if ((\writeCTmain_map'_Int_IntlizzieLet35_1_argbuf_rwb_r  && \writeCTmain_map'_Int_IntlizzieLet35_1_argbuf_bufchan_buf [0]))
        \writeCTmain_map'_Int_IntlizzieLet35_1_argbuf_bufchan_buf  <= {16'd0,
                                                                       1'd0};
      else if (((! \writeCTmain_map'_Int_IntlizzieLet35_1_argbuf_rwb_r ) && (! \writeCTmain_map'_Int_IntlizzieLet35_1_argbuf_bufchan_buf [0])))
        \writeCTmain_map'_Int_IntlizzieLet35_1_argbuf_bufchan_buf  <= \writeCTmain_map'_Int_IntlizzieLet35_1_argbuf_bufchan_d ;
  
  /* buf (Ty Pointer_CTmain_map'_Int_Int) : (writeCTmain_map'_Int_IntlizzieLet35_1_argbuf_rwb,Pointer_CTmain_map'_Int_Int) > (sca2_2_1_argbuf,Pointer_CTmain_map'_Int_Int) */
  \Pointer_CTmain_map'_Int_Int_t  \writeCTmain_map'_Int_IntlizzieLet35_1_argbuf_rwb_bufchan_d ;
  logic \writeCTmain_map'_Int_IntlizzieLet35_1_argbuf_rwb_bufchan_r ;
  assign \writeCTmain_map'_Int_IntlizzieLet35_1_argbuf_rwb_r  = ((! \writeCTmain_map'_Int_IntlizzieLet35_1_argbuf_rwb_bufchan_d [0]) || \writeCTmain_map'_Int_IntlizzieLet35_1_argbuf_rwb_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmain_map'_Int_IntlizzieLet35_1_argbuf_rwb_bufchan_d  <= {16'd0,
                                                                       1'd0};
    else
      if (\writeCTmain_map'_Int_IntlizzieLet35_1_argbuf_rwb_r )
        \writeCTmain_map'_Int_IntlizzieLet35_1_argbuf_rwb_bufchan_d  <= \writeCTmain_map'_Int_IntlizzieLet35_1_argbuf_rwb_d ;
  \Pointer_CTmain_map'_Int_Int_t  \writeCTmain_map'_Int_IntlizzieLet35_1_argbuf_rwb_bufchan_buf ;
  assign \writeCTmain_map'_Int_IntlizzieLet35_1_argbuf_rwb_bufchan_r  = (! \writeCTmain_map'_Int_IntlizzieLet35_1_argbuf_rwb_bufchan_buf [0]);
  assign sca2_2_1_argbuf_d = (\writeCTmain_map'_Int_IntlizzieLet35_1_argbuf_rwb_bufchan_buf [0] ? \writeCTmain_map'_Int_IntlizzieLet35_1_argbuf_rwb_bufchan_buf  :
                              \writeCTmain_map'_Int_IntlizzieLet35_1_argbuf_rwb_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmain_map'_Int_IntlizzieLet35_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                         1'd0};
    else
      if ((sca2_2_1_argbuf_r && \writeCTmain_map'_Int_IntlizzieLet35_1_argbuf_rwb_bufchan_buf [0]))
        \writeCTmain_map'_Int_IntlizzieLet35_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                           1'd0};
      else if (((! sca2_2_1_argbuf_r) && (! \writeCTmain_map'_Int_IntlizzieLet35_1_argbuf_rwb_bufchan_buf [0])))
        \writeCTmain_map'_Int_IntlizzieLet35_1_argbuf_rwb_bufchan_buf  <= \writeCTmain_map'_Int_IntlizzieLet35_1_argbuf_rwb_bufchan_d ;
  
  /* buf (Ty Pointer_CTmain_map'_Int_Int) : (writeCTmain_map'_Int_IntlizzieLet36_1_argbuf,Pointer_CTmain_map'_Int_Int) > (writeCTmain_map'_Int_IntlizzieLet36_1_argbuf_rwb,Pointer_CTmain_map'_Int_Int) */
  \Pointer_CTmain_map'_Int_Int_t  \writeCTmain_map'_Int_IntlizzieLet36_1_argbuf_bufchan_d ;
  logic \writeCTmain_map'_Int_IntlizzieLet36_1_argbuf_bufchan_r ;
  assign \writeCTmain_map'_Int_IntlizzieLet36_1_argbuf_r  = ((! \writeCTmain_map'_Int_IntlizzieLet36_1_argbuf_bufchan_d [0]) || \writeCTmain_map'_Int_IntlizzieLet36_1_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmain_map'_Int_IntlizzieLet36_1_argbuf_bufchan_d  <= {16'd0,
                                                                   1'd0};
    else
      if (\writeCTmain_map'_Int_IntlizzieLet36_1_argbuf_r )
        \writeCTmain_map'_Int_IntlizzieLet36_1_argbuf_bufchan_d  <= \writeCTmain_map'_Int_IntlizzieLet36_1_argbuf_d ;
  \Pointer_CTmain_map'_Int_Int_t  \writeCTmain_map'_Int_IntlizzieLet36_1_argbuf_bufchan_buf ;
  assign \writeCTmain_map'_Int_IntlizzieLet36_1_argbuf_bufchan_r  = (! \writeCTmain_map'_Int_IntlizzieLet36_1_argbuf_bufchan_buf [0]);
  assign \writeCTmain_map'_Int_IntlizzieLet36_1_argbuf_rwb_d  = (\writeCTmain_map'_Int_IntlizzieLet36_1_argbuf_bufchan_buf [0] ? \writeCTmain_map'_Int_IntlizzieLet36_1_argbuf_bufchan_buf  :
                                                                 \writeCTmain_map'_Int_IntlizzieLet36_1_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmain_map'_Int_IntlizzieLet36_1_argbuf_bufchan_buf  <= {16'd0,
                                                                     1'd0};
    else
      if ((\writeCTmain_map'_Int_IntlizzieLet36_1_argbuf_rwb_r  && \writeCTmain_map'_Int_IntlizzieLet36_1_argbuf_bufchan_buf [0]))
        \writeCTmain_map'_Int_IntlizzieLet36_1_argbuf_bufchan_buf  <= {16'd0,
                                                                       1'd0};
      else if (((! \writeCTmain_map'_Int_IntlizzieLet36_1_argbuf_rwb_r ) && (! \writeCTmain_map'_Int_IntlizzieLet36_1_argbuf_bufchan_buf [0])))
        \writeCTmain_map'_Int_IntlizzieLet36_1_argbuf_bufchan_buf  <= \writeCTmain_map'_Int_IntlizzieLet36_1_argbuf_bufchan_d ;
  
  /* buf (Ty Pointer_CTmain_map'_Int_Int) : (writeCTmain_map'_Int_IntlizzieLet36_1_argbuf_rwb,Pointer_CTmain_map'_Int_Int) > (sca1_2_1_argbuf,Pointer_CTmain_map'_Int_Int) */
  \Pointer_CTmain_map'_Int_Int_t  \writeCTmain_map'_Int_IntlizzieLet36_1_argbuf_rwb_bufchan_d ;
  logic \writeCTmain_map'_Int_IntlizzieLet36_1_argbuf_rwb_bufchan_r ;
  assign \writeCTmain_map'_Int_IntlizzieLet36_1_argbuf_rwb_r  = ((! \writeCTmain_map'_Int_IntlizzieLet36_1_argbuf_rwb_bufchan_d [0]) || \writeCTmain_map'_Int_IntlizzieLet36_1_argbuf_rwb_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmain_map'_Int_IntlizzieLet36_1_argbuf_rwb_bufchan_d  <= {16'd0,
                                                                       1'd0};
    else
      if (\writeCTmain_map'_Int_IntlizzieLet36_1_argbuf_rwb_r )
        \writeCTmain_map'_Int_IntlizzieLet36_1_argbuf_rwb_bufchan_d  <= \writeCTmain_map'_Int_IntlizzieLet36_1_argbuf_rwb_d ;
  \Pointer_CTmain_map'_Int_Int_t  \writeCTmain_map'_Int_IntlizzieLet36_1_argbuf_rwb_bufchan_buf ;
  assign \writeCTmain_map'_Int_IntlizzieLet36_1_argbuf_rwb_bufchan_r  = (! \writeCTmain_map'_Int_IntlizzieLet36_1_argbuf_rwb_bufchan_buf [0]);
  assign sca1_2_1_argbuf_d = (\writeCTmain_map'_Int_IntlizzieLet36_1_argbuf_rwb_bufchan_buf [0] ? \writeCTmain_map'_Int_IntlizzieLet36_1_argbuf_rwb_bufchan_buf  :
                              \writeCTmain_map'_Int_IntlizzieLet36_1_argbuf_rwb_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmain_map'_Int_IntlizzieLet36_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                         1'd0};
    else
      if ((sca1_2_1_argbuf_r && \writeCTmain_map'_Int_IntlizzieLet36_1_argbuf_rwb_bufchan_buf [0]))
        \writeCTmain_map'_Int_IntlizzieLet36_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                           1'd0};
      else if (((! sca1_2_1_argbuf_r) && (! \writeCTmain_map'_Int_IntlizzieLet36_1_argbuf_rwb_bufchan_buf [0])))
        \writeCTmain_map'_Int_IntlizzieLet36_1_argbuf_rwb_bufchan_buf  <= \writeCTmain_map'_Int_IntlizzieLet36_1_argbuf_rwb_bufchan_d ;
  
  /* buf (Ty Pointer_CTmain_map'_Int_Int) : (writeCTmain_map'_Int_IntlizzieLet37_1_argbuf,Pointer_CTmain_map'_Int_Int) > (writeCTmain_map'_Int_IntlizzieLet37_1_argbuf_rwb,Pointer_CTmain_map'_Int_Int) */
  \Pointer_CTmain_map'_Int_Int_t  \writeCTmain_map'_Int_IntlizzieLet37_1_argbuf_bufchan_d ;
  logic \writeCTmain_map'_Int_IntlizzieLet37_1_argbuf_bufchan_r ;
  assign \writeCTmain_map'_Int_IntlizzieLet37_1_argbuf_r  = ((! \writeCTmain_map'_Int_IntlizzieLet37_1_argbuf_bufchan_d [0]) || \writeCTmain_map'_Int_IntlizzieLet37_1_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmain_map'_Int_IntlizzieLet37_1_argbuf_bufchan_d  <= {16'd0,
                                                                   1'd0};
    else
      if (\writeCTmain_map'_Int_IntlizzieLet37_1_argbuf_r )
        \writeCTmain_map'_Int_IntlizzieLet37_1_argbuf_bufchan_d  <= \writeCTmain_map'_Int_IntlizzieLet37_1_argbuf_d ;
  \Pointer_CTmain_map'_Int_Int_t  \writeCTmain_map'_Int_IntlizzieLet37_1_argbuf_bufchan_buf ;
  assign \writeCTmain_map'_Int_IntlizzieLet37_1_argbuf_bufchan_r  = (! \writeCTmain_map'_Int_IntlizzieLet37_1_argbuf_bufchan_buf [0]);
  assign \writeCTmain_map'_Int_IntlizzieLet37_1_argbuf_rwb_d  = (\writeCTmain_map'_Int_IntlizzieLet37_1_argbuf_bufchan_buf [0] ? \writeCTmain_map'_Int_IntlizzieLet37_1_argbuf_bufchan_buf  :
                                                                 \writeCTmain_map'_Int_IntlizzieLet37_1_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmain_map'_Int_IntlizzieLet37_1_argbuf_bufchan_buf  <= {16'd0,
                                                                     1'd0};
    else
      if ((\writeCTmain_map'_Int_IntlizzieLet37_1_argbuf_rwb_r  && \writeCTmain_map'_Int_IntlizzieLet37_1_argbuf_bufchan_buf [0]))
        \writeCTmain_map'_Int_IntlizzieLet37_1_argbuf_bufchan_buf  <= {16'd0,
                                                                       1'd0};
      else if (((! \writeCTmain_map'_Int_IntlizzieLet37_1_argbuf_rwb_r ) && (! \writeCTmain_map'_Int_IntlizzieLet37_1_argbuf_bufchan_buf [0])))
        \writeCTmain_map'_Int_IntlizzieLet37_1_argbuf_bufchan_buf  <= \writeCTmain_map'_Int_IntlizzieLet37_1_argbuf_bufchan_d ;
  
  /* buf (Ty Pointer_CTmain_map'_Int_Int) : (writeCTmain_map'_Int_IntlizzieLet37_1_argbuf_rwb,Pointer_CTmain_map'_Int_Int) > (sca0_2_1_argbuf,Pointer_CTmain_map'_Int_Int) */
  \Pointer_CTmain_map'_Int_Int_t  \writeCTmain_map'_Int_IntlizzieLet37_1_argbuf_rwb_bufchan_d ;
  logic \writeCTmain_map'_Int_IntlizzieLet37_1_argbuf_rwb_bufchan_r ;
  assign \writeCTmain_map'_Int_IntlizzieLet37_1_argbuf_rwb_r  = ((! \writeCTmain_map'_Int_IntlizzieLet37_1_argbuf_rwb_bufchan_d [0]) || \writeCTmain_map'_Int_IntlizzieLet37_1_argbuf_rwb_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmain_map'_Int_IntlizzieLet37_1_argbuf_rwb_bufchan_d  <= {16'd0,
                                                                       1'd0};
    else
      if (\writeCTmain_map'_Int_IntlizzieLet37_1_argbuf_rwb_r )
        \writeCTmain_map'_Int_IntlizzieLet37_1_argbuf_rwb_bufchan_d  <= \writeCTmain_map'_Int_IntlizzieLet37_1_argbuf_rwb_d ;
  \Pointer_CTmain_map'_Int_Int_t  \writeCTmain_map'_Int_IntlizzieLet37_1_argbuf_rwb_bufchan_buf ;
  assign \writeCTmain_map'_Int_IntlizzieLet37_1_argbuf_rwb_bufchan_r  = (! \writeCTmain_map'_Int_IntlizzieLet37_1_argbuf_rwb_bufchan_buf [0]);
  assign sca0_2_1_argbuf_d = (\writeCTmain_map'_Int_IntlizzieLet37_1_argbuf_rwb_bufchan_buf [0] ? \writeCTmain_map'_Int_IntlizzieLet37_1_argbuf_rwb_bufchan_buf  :
                              \writeCTmain_map'_Int_IntlizzieLet37_1_argbuf_rwb_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmain_map'_Int_IntlizzieLet37_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                         1'd0};
    else
      if ((sca0_2_1_argbuf_r && \writeCTmain_map'_Int_IntlizzieLet37_1_argbuf_rwb_bufchan_buf [0]))
        \writeCTmain_map'_Int_IntlizzieLet37_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                           1'd0};
      else if (((! sca0_2_1_argbuf_r) && (! \writeCTmain_map'_Int_IntlizzieLet37_1_argbuf_rwb_bufchan_buf [0])))
        \writeCTmain_map'_Int_IntlizzieLet37_1_argbuf_rwb_bufchan_buf  <= \writeCTmain_map'_Int_IntlizzieLet37_1_argbuf_rwb_bufchan_d ;
  
  /* buf (Ty Pointer_CTmap''_map''_Int_Int_Int) : (writeCTmap''_map''_Int_Int_IntlizzieLet20_1_argbuf,Pointer_CTmap''_map''_Int_Int_Int) > (writeCTmap''_map''_Int_Int_IntlizzieLet20_1_argbuf_rwb,Pointer_CTmap''_map''_Int_Int_Int) */
  \Pointer_CTmap''_map''_Int_Int_Int_t  \writeCTmap''_map''_Int_Int_IntlizzieLet20_1_argbuf_bufchan_d ;
  logic \writeCTmap''_map''_Int_Int_IntlizzieLet20_1_argbuf_bufchan_r ;
  assign \writeCTmap''_map''_Int_Int_IntlizzieLet20_1_argbuf_r  = ((! \writeCTmap''_map''_Int_Int_IntlizzieLet20_1_argbuf_bufchan_d [0]) || \writeCTmap''_map''_Int_Int_IntlizzieLet20_1_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmap''_map''_Int_Int_IntlizzieLet20_1_argbuf_bufchan_d  <= {16'd0,
                                                                         1'd0};
    else
      if (\writeCTmap''_map''_Int_Int_IntlizzieLet20_1_argbuf_r )
        \writeCTmap''_map''_Int_Int_IntlizzieLet20_1_argbuf_bufchan_d  <= \writeCTmap''_map''_Int_Int_IntlizzieLet20_1_argbuf_d ;
  \Pointer_CTmap''_map''_Int_Int_Int_t  \writeCTmap''_map''_Int_Int_IntlizzieLet20_1_argbuf_bufchan_buf ;
  assign \writeCTmap''_map''_Int_Int_IntlizzieLet20_1_argbuf_bufchan_r  = (! \writeCTmap''_map''_Int_Int_IntlizzieLet20_1_argbuf_bufchan_buf [0]);
  assign \writeCTmap''_map''_Int_Int_IntlizzieLet20_1_argbuf_rwb_d  = (\writeCTmap''_map''_Int_Int_IntlizzieLet20_1_argbuf_bufchan_buf [0] ? \writeCTmap''_map''_Int_Int_IntlizzieLet20_1_argbuf_bufchan_buf  :
                                                                       \writeCTmap''_map''_Int_Int_IntlizzieLet20_1_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmap''_map''_Int_Int_IntlizzieLet20_1_argbuf_bufchan_buf  <= {16'd0,
                                                                           1'd0};
    else
      if ((\writeCTmap''_map''_Int_Int_IntlizzieLet20_1_argbuf_rwb_r  && \writeCTmap''_map''_Int_Int_IntlizzieLet20_1_argbuf_bufchan_buf [0]))
        \writeCTmap''_map''_Int_Int_IntlizzieLet20_1_argbuf_bufchan_buf  <= {16'd0,
                                                                             1'd0};
      else if (((! \writeCTmap''_map''_Int_Int_IntlizzieLet20_1_argbuf_rwb_r ) && (! \writeCTmap''_map''_Int_Int_IntlizzieLet20_1_argbuf_bufchan_buf [0])))
        \writeCTmap''_map''_Int_Int_IntlizzieLet20_1_argbuf_bufchan_buf  <= \writeCTmap''_map''_Int_Int_IntlizzieLet20_1_argbuf_bufchan_d ;
  
  /* buf (Ty Pointer_CTmap''_map''_Int_Int_Int) : (writeCTmap''_map''_Int_Int_IntlizzieLet20_1_argbuf_rwb,Pointer_CTmap''_map''_Int_Int_Int) > (sca3_3_1_argbuf,Pointer_CTmap''_map''_Int_Int_Int) */
  \Pointer_CTmap''_map''_Int_Int_Int_t  \writeCTmap''_map''_Int_Int_IntlizzieLet20_1_argbuf_rwb_bufchan_d ;
  logic \writeCTmap''_map''_Int_Int_IntlizzieLet20_1_argbuf_rwb_bufchan_r ;
  assign \writeCTmap''_map''_Int_Int_IntlizzieLet20_1_argbuf_rwb_r  = ((! \writeCTmap''_map''_Int_Int_IntlizzieLet20_1_argbuf_rwb_bufchan_d [0]) || \writeCTmap''_map''_Int_Int_IntlizzieLet20_1_argbuf_rwb_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmap''_map''_Int_Int_IntlizzieLet20_1_argbuf_rwb_bufchan_d  <= {16'd0,
                                                                             1'd0};
    else
      if (\writeCTmap''_map''_Int_Int_IntlizzieLet20_1_argbuf_rwb_r )
        \writeCTmap''_map''_Int_Int_IntlizzieLet20_1_argbuf_rwb_bufchan_d  <= \writeCTmap''_map''_Int_Int_IntlizzieLet20_1_argbuf_rwb_d ;
  \Pointer_CTmap''_map''_Int_Int_Int_t  \writeCTmap''_map''_Int_Int_IntlizzieLet20_1_argbuf_rwb_bufchan_buf ;
  assign \writeCTmap''_map''_Int_Int_IntlizzieLet20_1_argbuf_rwb_bufchan_r  = (! \writeCTmap''_map''_Int_Int_IntlizzieLet20_1_argbuf_rwb_bufchan_buf [0]);
  assign sca3_3_1_argbuf_d = (\writeCTmap''_map''_Int_Int_IntlizzieLet20_1_argbuf_rwb_bufchan_buf [0] ? \writeCTmap''_map''_Int_Int_IntlizzieLet20_1_argbuf_rwb_bufchan_buf  :
                              \writeCTmap''_map''_Int_Int_IntlizzieLet20_1_argbuf_rwb_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmap''_map''_Int_Int_IntlizzieLet20_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                               1'd0};
    else
      if ((sca3_3_1_argbuf_r && \writeCTmap''_map''_Int_Int_IntlizzieLet20_1_argbuf_rwb_bufchan_buf [0]))
        \writeCTmap''_map''_Int_Int_IntlizzieLet20_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                                 1'd0};
      else if (((! sca3_3_1_argbuf_r) && (! \writeCTmap''_map''_Int_Int_IntlizzieLet20_1_argbuf_rwb_bufchan_buf [0])))
        \writeCTmap''_map''_Int_Int_IntlizzieLet20_1_argbuf_rwb_bufchan_buf  <= \writeCTmap''_map''_Int_Int_IntlizzieLet20_1_argbuf_rwb_bufchan_d ;
  
  /* buf (Ty Pointer_CTmap''_map''_Int_Int_Int) : (writeCTmap''_map''_Int_Int_IntlizzieLet24_1_argbuf,Pointer_CTmap''_map''_Int_Int_Int) > (writeCTmap''_map''_Int_Int_IntlizzieLet24_1_argbuf_rwb,Pointer_CTmap''_map''_Int_Int_Int) */
  \Pointer_CTmap''_map''_Int_Int_Int_t  \writeCTmap''_map''_Int_Int_IntlizzieLet24_1_argbuf_bufchan_d ;
  logic \writeCTmap''_map''_Int_Int_IntlizzieLet24_1_argbuf_bufchan_r ;
  assign \writeCTmap''_map''_Int_Int_IntlizzieLet24_1_argbuf_r  = ((! \writeCTmap''_map''_Int_Int_IntlizzieLet24_1_argbuf_bufchan_d [0]) || \writeCTmap''_map''_Int_Int_IntlizzieLet24_1_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmap''_map''_Int_Int_IntlizzieLet24_1_argbuf_bufchan_d  <= {16'd0,
                                                                         1'd0};
    else
      if (\writeCTmap''_map''_Int_Int_IntlizzieLet24_1_argbuf_r )
        \writeCTmap''_map''_Int_Int_IntlizzieLet24_1_argbuf_bufchan_d  <= \writeCTmap''_map''_Int_Int_IntlizzieLet24_1_argbuf_d ;
  \Pointer_CTmap''_map''_Int_Int_Int_t  \writeCTmap''_map''_Int_Int_IntlizzieLet24_1_argbuf_bufchan_buf ;
  assign \writeCTmap''_map''_Int_Int_IntlizzieLet24_1_argbuf_bufchan_r  = (! \writeCTmap''_map''_Int_Int_IntlizzieLet24_1_argbuf_bufchan_buf [0]);
  assign \writeCTmap''_map''_Int_Int_IntlizzieLet24_1_argbuf_rwb_d  = (\writeCTmap''_map''_Int_Int_IntlizzieLet24_1_argbuf_bufchan_buf [0] ? \writeCTmap''_map''_Int_Int_IntlizzieLet24_1_argbuf_bufchan_buf  :
                                                                       \writeCTmap''_map''_Int_Int_IntlizzieLet24_1_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmap''_map''_Int_Int_IntlizzieLet24_1_argbuf_bufchan_buf  <= {16'd0,
                                                                           1'd0};
    else
      if ((\writeCTmap''_map''_Int_Int_IntlizzieLet24_1_argbuf_rwb_r  && \writeCTmap''_map''_Int_Int_IntlizzieLet24_1_argbuf_bufchan_buf [0]))
        \writeCTmap''_map''_Int_Int_IntlizzieLet24_1_argbuf_bufchan_buf  <= {16'd0,
                                                                             1'd0};
      else if (((! \writeCTmap''_map''_Int_Int_IntlizzieLet24_1_argbuf_rwb_r ) && (! \writeCTmap''_map''_Int_Int_IntlizzieLet24_1_argbuf_bufchan_buf [0])))
        \writeCTmap''_map''_Int_Int_IntlizzieLet24_1_argbuf_bufchan_buf  <= \writeCTmap''_map''_Int_Int_IntlizzieLet24_1_argbuf_bufchan_d ;
  
  /* buf (Ty Pointer_CTmap''_map''_Int_Int_Int) : (writeCTmap''_map''_Int_Int_IntlizzieLet24_1_argbuf_rwb,Pointer_CTmap''_map''_Int_Int_Int) > (lizzieLet10_1_1_argbuf,Pointer_CTmap''_map''_Int_Int_Int) */
  \Pointer_CTmap''_map''_Int_Int_Int_t  \writeCTmap''_map''_Int_Int_IntlizzieLet24_1_argbuf_rwb_bufchan_d ;
  logic \writeCTmap''_map''_Int_Int_IntlizzieLet24_1_argbuf_rwb_bufchan_r ;
  assign \writeCTmap''_map''_Int_Int_IntlizzieLet24_1_argbuf_rwb_r  = ((! \writeCTmap''_map''_Int_Int_IntlizzieLet24_1_argbuf_rwb_bufchan_d [0]) || \writeCTmap''_map''_Int_Int_IntlizzieLet24_1_argbuf_rwb_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmap''_map''_Int_Int_IntlizzieLet24_1_argbuf_rwb_bufchan_d  <= {16'd0,
                                                                             1'd0};
    else
      if (\writeCTmap''_map''_Int_Int_IntlizzieLet24_1_argbuf_rwb_r )
        \writeCTmap''_map''_Int_Int_IntlizzieLet24_1_argbuf_rwb_bufchan_d  <= \writeCTmap''_map''_Int_Int_IntlizzieLet24_1_argbuf_rwb_d ;
  \Pointer_CTmap''_map''_Int_Int_Int_t  \writeCTmap''_map''_Int_Int_IntlizzieLet24_1_argbuf_rwb_bufchan_buf ;
  assign \writeCTmap''_map''_Int_Int_IntlizzieLet24_1_argbuf_rwb_bufchan_r  = (! \writeCTmap''_map''_Int_Int_IntlizzieLet24_1_argbuf_rwb_bufchan_buf [0]);
  assign lizzieLet10_1_1_argbuf_d = (\writeCTmap''_map''_Int_Int_IntlizzieLet24_1_argbuf_rwb_bufchan_buf [0] ? \writeCTmap''_map''_Int_Int_IntlizzieLet24_1_argbuf_rwb_bufchan_buf  :
                                     \writeCTmap''_map''_Int_Int_IntlizzieLet24_1_argbuf_rwb_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmap''_map''_Int_Int_IntlizzieLet24_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                               1'd0};
    else
      if ((lizzieLet10_1_1_argbuf_r && \writeCTmap''_map''_Int_Int_IntlizzieLet24_1_argbuf_rwb_bufchan_buf [0]))
        \writeCTmap''_map''_Int_Int_IntlizzieLet24_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                                 1'd0};
      else if (((! lizzieLet10_1_1_argbuf_r) && (! \writeCTmap''_map''_Int_Int_IntlizzieLet24_1_argbuf_rwb_bufchan_buf [0])))
        \writeCTmap''_map''_Int_Int_IntlizzieLet24_1_argbuf_rwb_bufchan_buf  <= \writeCTmap''_map''_Int_Int_IntlizzieLet24_1_argbuf_rwb_bufchan_d ;
  
  /* buf (Ty Pointer_CTmap''_map''_Int_Int_Int) : (writeCTmap''_map''_Int_Int_IntlizzieLet40_1_argbuf,Pointer_CTmap''_map''_Int_Int_Int) > (writeCTmap''_map''_Int_Int_IntlizzieLet40_1_argbuf_rwb,Pointer_CTmap''_map''_Int_Int_Int) */
  \Pointer_CTmap''_map''_Int_Int_Int_t  \writeCTmap''_map''_Int_Int_IntlizzieLet40_1_argbuf_bufchan_d ;
  logic \writeCTmap''_map''_Int_Int_IntlizzieLet40_1_argbuf_bufchan_r ;
  assign \writeCTmap''_map''_Int_Int_IntlizzieLet40_1_argbuf_r  = ((! \writeCTmap''_map''_Int_Int_IntlizzieLet40_1_argbuf_bufchan_d [0]) || \writeCTmap''_map''_Int_Int_IntlizzieLet40_1_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmap''_map''_Int_Int_IntlizzieLet40_1_argbuf_bufchan_d  <= {16'd0,
                                                                         1'd0};
    else
      if (\writeCTmap''_map''_Int_Int_IntlizzieLet40_1_argbuf_r )
        \writeCTmap''_map''_Int_Int_IntlizzieLet40_1_argbuf_bufchan_d  <= \writeCTmap''_map''_Int_Int_IntlizzieLet40_1_argbuf_d ;
  \Pointer_CTmap''_map''_Int_Int_Int_t  \writeCTmap''_map''_Int_Int_IntlizzieLet40_1_argbuf_bufchan_buf ;
  assign \writeCTmap''_map''_Int_Int_IntlizzieLet40_1_argbuf_bufchan_r  = (! \writeCTmap''_map''_Int_Int_IntlizzieLet40_1_argbuf_bufchan_buf [0]);
  assign \writeCTmap''_map''_Int_Int_IntlizzieLet40_1_argbuf_rwb_d  = (\writeCTmap''_map''_Int_Int_IntlizzieLet40_1_argbuf_bufchan_buf [0] ? \writeCTmap''_map''_Int_Int_IntlizzieLet40_1_argbuf_bufchan_buf  :
                                                                       \writeCTmap''_map''_Int_Int_IntlizzieLet40_1_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmap''_map''_Int_Int_IntlizzieLet40_1_argbuf_bufchan_buf  <= {16'd0,
                                                                           1'd0};
    else
      if ((\writeCTmap''_map''_Int_Int_IntlizzieLet40_1_argbuf_rwb_r  && \writeCTmap''_map''_Int_Int_IntlizzieLet40_1_argbuf_bufchan_buf [0]))
        \writeCTmap''_map''_Int_Int_IntlizzieLet40_1_argbuf_bufchan_buf  <= {16'd0,
                                                                             1'd0};
      else if (((! \writeCTmap''_map''_Int_Int_IntlizzieLet40_1_argbuf_rwb_r ) && (! \writeCTmap''_map''_Int_Int_IntlizzieLet40_1_argbuf_bufchan_buf [0])))
        \writeCTmap''_map''_Int_Int_IntlizzieLet40_1_argbuf_bufchan_buf  <= \writeCTmap''_map''_Int_Int_IntlizzieLet40_1_argbuf_bufchan_d ;
  
  /* buf (Ty Pointer_CTmap''_map''_Int_Int_Int) : (writeCTmap''_map''_Int_Int_IntlizzieLet40_1_argbuf_rwb,Pointer_CTmap''_map''_Int_Int_Int) > (sca2_3_1_argbuf,Pointer_CTmap''_map''_Int_Int_Int) */
  \Pointer_CTmap''_map''_Int_Int_Int_t  \writeCTmap''_map''_Int_Int_IntlizzieLet40_1_argbuf_rwb_bufchan_d ;
  logic \writeCTmap''_map''_Int_Int_IntlizzieLet40_1_argbuf_rwb_bufchan_r ;
  assign \writeCTmap''_map''_Int_Int_IntlizzieLet40_1_argbuf_rwb_r  = ((! \writeCTmap''_map''_Int_Int_IntlizzieLet40_1_argbuf_rwb_bufchan_d [0]) || \writeCTmap''_map''_Int_Int_IntlizzieLet40_1_argbuf_rwb_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmap''_map''_Int_Int_IntlizzieLet40_1_argbuf_rwb_bufchan_d  <= {16'd0,
                                                                             1'd0};
    else
      if (\writeCTmap''_map''_Int_Int_IntlizzieLet40_1_argbuf_rwb_r )
        \writeCTmap''_map''_Int_Int_IntlizzieLet40_1_argbuf_rwb_bufchan_d  <= \writeCTmap''_map''_Int_Int_IntlizzieLet40_1_argbuf_rwb_d ;
  \Pointer_CTmap''_map''_Int_Int_Int_t  \writeCTmap''_map''_Int_Int_IntlizzieLet40_1_argbuf_rwb_bufchan_buf ;
  assign \writeCTmap''_map''_Int_Int_IntlizzieLet40_1_argbuf_rwb_bufchan_r  = (! \writeCTmap''_map''_Int_Int_IntlizzieLet40_1_argbuf_rwb_bufchan_buf [0]);
  assign sca2_3_1_argbuf_d = (\writeCTmap''_map''_Int_Int_IntlizzieLet40_1_argbuf_rwb_bufchan_buf [0] ? \writeCTmap''_map''_Int_Int_IntlizzieLet40_1_argbuf_rwb_bufchan_buf  :
                              \writeCTmap''_map''_Int_Int_IntlizzieLet40_1_argbuf_rwb_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmap''_map''_Int_Int_IntlizzieLet40_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                               1'd0};
    else
      if ((sca2_3_1_argbuf_r && \writeCTmap''_map''_Int_Int_IntlizzieLet40_1_argbuf_rwb_bufchan_buf [0]))
        \writeCTmap''_map''_Int_Int_IntlizzieLet40_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                                 1'd0};
      else if (((! sca2_3_1_argbuf_r) && (! \writeCTmap''_map''_Int_Int_IntlizzieLet40_1_argbuf_rwb_bufchan_buf [0])))
        \writeCTmap''_map''_Int_Int_IntlizzieLet40_1_argbuf_rwb_bufchan_buf  <= \writeCTmap''_map''_Int_Int_IntlizzieLet40_1_argbuf_rwb_bufchan_d ;
  
  /* buf (Ty Pointer_CTmap''_map''_Int_Int_Int) : (writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf,Pointer_CTmap''_map''_Int_Int_Int) > (writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf_rwb,Pointer_CTmap''_map''_Int_Int_Int) */
  \Pointer_CTmap''_map''_Int_Int_Int_t  \writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf_bufchan_d ;
  logic \writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf_bufchan_r ;
  assign \writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf_r  = ((! \writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf_bufchan_d [0]) || \writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf_bufchan_d  <= {16'd0,
                                                                         1'd0};
    else
      if (\writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf_r )
        \writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf_bufchan_d  <= \writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf_d ;
  \Pointer_CTmap''_map''_Int_Int_Int_t  \writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf_bufchan_buf ;
  assign \writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf_bufchan_r  = (! \writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf_bufchan_buf [0]);
  assign \writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf_rwb_d  = (\writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf_bufchan_buf [0] ? \writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf_bufchan_buf  :
                                                                       \writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf_bufchan_buf  <= {16'd0,
                                                                           1'd0};
    else
      if ((\writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf_rwb_r  && \writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf_bufchan_buf [0]))
        \writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf_bufchan_buf  <= {16'd0,
                                                                             1'd0};
      else if (((! \writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf_rwb_r ) && (! \writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf_bufchan_buf [0])))
        \writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf_bufchan_buf  <= \writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf_bufchan_d ;
  
  /* buf (Ty Pointer_CTmap''_map''_Int_Int_Int) : (writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf_rwb,Pointer_CTmap''_map''_Int_Int_Int) > (sca1_3_1_argbuf,Pointer_CTmap''_map''_Int_Int_Int) */
  \Pointer_CTmap''_map''_Int_Int_Int_t  \writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf_rwb_bufchan_d ;
  logic \writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf_rwb_bufchan_r ;
  assign \writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf_rwb_r  = ((! \writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf_rwb_bufchan_d [0]) || \writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf_rwb_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf_rwb_bufchan_d  <= {16'd0,
                                                                             1'd0};
    else
      if (\writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf_rwb_r )
        \writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf_rwb_bufchan_d  <= \writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf_rwb_d ;
  \Pointer_CTmap''_map''_Int_Int_Int_t  \writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf_rwb_bufchan_buf ;
  assign \writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf_rwb_bufchan_r  = (! \writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf_rwb_bufchan_buf [0]);
  assign sca1_3_1_argbuf_d = (\writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf_rwb_bufchan_buf [0] ? \writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf_rwb_bufchan_buf  :
                              \writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf_rwb_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                               1'd0};
    else
      if ((sca1_3_1_argbuf_r && \writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf_rwb_bufchan_buf [0]))
        \writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                                 1'd0};
      else if (((! sca1_3_1_argbuf_r) && (! \writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf_rwb_bufchan_buf [0])))
        \writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf_rwb_bufchan_buf  <= \writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf_rwb_bufchan_d ;
  
  /* buf (Ty Pointer_CTmap''_map''_Int_Int_Int) : (writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf,Pointer_CTmap''_map''_Int_Int_Int) > (writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf_rwb,Pointer_CTmap''_map''_Int_Int_Int) */
  \Pointer_CTmap''_map''_Int_Int_Int_t  \writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf_bufchan_d ;
  logic \writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf_bufchan_r ;
  assign \writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf_r  = ((! \writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf_bufchan_d [0]) || \writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf_bufchan_d  <= {16'd0,
                                                                         1'd0};
    else
      if (\writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf_r )
        \writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf_bufchan_d  <= \writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf_d ;
  \Pointer_CTmap''_map''_Int_Int_Int_t  \writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf_bufchan_buf ;
  assign \writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf_bufchan_r  = (! \writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf_bufchan_buf [0]);
  assign \writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf_rwb_d  = (\writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf_bufchan_buf [0] ? \writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf_bufchan_buf  :
                                                                       \writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf_bufchan_buf  <= {16'd0,
                                                                           1'd0};
    else
      if ((\writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf_rwb_r  && \writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf_bufchan_buf [0]))
        \writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf_bufchan_buf  <= {16'd0,
                                                                             1'd0};
      else if (((! \writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf_rwb_r ) && (! \writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf_bufchan_buf [0])))
        \writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf_bufchan_buf  <= \writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf_bufchan_d ;
  
  /* buf (Ty Pointer_CTmap''_map''_Int_Int_Int) : (writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf_rwb,Pointer_CTmap''_map''_Int_Int_Int) > (sca0_3_1_argbuf,Pointer_CTmap''_map''_Int_Int_Int) */
  \Pointer_CTmap''_map''_Int_Int_Int_t  \writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf_rwb_bufchan_d ;
  logic \writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf_rwb_bufchan_r ;
  assign \writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf_rwb_r  = ((! \writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf_rwb_bufchan_d [0]) || \writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf_rwb_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf_rwb_bufchan_d  <= {16'd0,
                                                                             1'd0};
    else
      if (\writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf_rwb_r )
        \writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf_rwb_bufchan_d  <= \writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf_rwb_d ;
  \Pointer_CTmap''_map''_Int_Int_Int_t  \writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf_rwb_bufchan_buf ;
  assign \writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf_rwb_bufchan_r  = (! \writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf_rwb_bufchan_buf [0]);
  assign sca0_3_1_argbuf_d = (\writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf_rwb_bufchan_buf [0] ? \writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf_rwb_bufchan_buf  :
                              \writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf_rwb_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                               1'd0};
    else
      if ((sca0_3_1_argbuf_r && \writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf_rwb_bufchan_buf [0]))
        \writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                                 1'd0};
      else if (((! sca0_3_1_argbuf_r) && (! \writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf_rwb_bufchan_buf [0])))
        \writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf_rwb_bufchan_buf  <= \writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf_rwb_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet11_1_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet11_1_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet11_1_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet11_1_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet11_1_1_argbuf_r = ((! writeQTree_IntlizzieLet11_1_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet11_1_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet11_1_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet11_1_1_argbuf_r)
        writeQTree_IntlizzieLet11_1_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet11_1_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet11_1_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet11_1_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet11_1_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet11_1_1_argbuf_rwb_d = (writeQTree_IntlizzieLet11_1_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet11_1_1_argbuf_bufchan_buf :
                                                       writeQTree_IntlizzieLet11_1_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet11_1_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet11_1_1_argbuf_rwb_r && writeQTree_IntlizzieLet11_1_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet11_1_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet11_1_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet11_1_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet11_1_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet11_1_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet11_1_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet1_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet11_1_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet11_1_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet11_1_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet11_1_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet11_1_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet11_1_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                             1'd0};
    else
      if (writeQTree_IntlizzieLet11_1_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet11_1_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet11_1_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet11_1_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet11_1_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet11_1_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet1_1_1_argbuf_d = (writeQTree_IntlizzieLet11_1_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet11_1_1_argbuf_rwb_bufchan_buf :
                                    writeQTree_IntlizzieLet11_1_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet11_1_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
    else
      if ((lizzieLet1_1_1_argbuf_r && writeQTree_IntlizzieLet11_1_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet11_1_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                 1'd0};
      else if (((! lizzieLet1_1_1_argbuf_r) && (! writeQTree_IntlizzieLet11_1_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet11_1_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet11_1_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet12_1_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet12_1_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet12_1_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet12_1_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet12_1_1_argbuf_r = ((! writeQTree_IntlizzieLet12_1_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet12_1_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet12_1_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet12_1_1_argbuf_r)
        writeQTree_IntlizzieLet12_1_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet12_1_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet12_1_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet12_1_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet12_1_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet12_1_1_argbuf_rwb_d = (writeQTree_IntlizzieLet12_1_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet12_1_1_argbuf_bufchan_buf :
                                                       writeQTree_IntlizzieLet12_1_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet12_1_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet12_1_1_argbuf_rwb_r && writeQTree_IntlizzieLet12_1_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet12_1_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet12_1_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet12_1_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet12_1_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet12_1_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet12_1_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet2_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet12_1_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet12_1_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet12_1_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet12_1_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet12_1_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet12_1_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                             1'd0};
    else
      if (writeQTree_IntlizzieLet12_1_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet12_1_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet12_1_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet12_1_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet12_1_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet12_1_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet2_1_1_argbuf_d = (writeQTree_IntlizzieLet12_1_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet12_1_1_argbuf_rwb_bufchan_buf :
                                    writeQTree_IntlizzieLet12_1_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet12_1_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
    else
      if ((lizzieLet2_1_1_argbuf_r && writeQTree_IntlizzieLet12_1_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet12_1_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                 1'd0};
      else if (((! lizzieLet2_1_1_argbuf_r) && (! writeQTree_IntlizzieLet12_1_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet12_1_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet12_1_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet13_1_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet13_1_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet13_1_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet13_1_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet13_1_1_argbuf_r = ((! writeQTree_IntlizzieLet13_1_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet13_1_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet13_1_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet13_1_1_argbuf_r)
        writeQTree_IntlizzieLet13_1_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet13_1_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet13_1_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet13_1_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet13_1_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet13_1_1_argbuf_rwb_d = (writeQTree_IntlizzieLet13_1_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet13_1_1_argbuf_bufchan_buf :
                                                       writeQTree_IntlizzieLet13_1_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet13_1_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet13_1_1_argbuf_rwb_r && writeQTree_IntlizzieLet13_1_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet13_1_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet13_1_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet13_1_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet13_1_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet13_1_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet13_1_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet3_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet13_1_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet13_1_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet13_1_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet13_1_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet13_1_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet13_1_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                             1'd0};
    else
      if (writeQTree_IntlizzieLet13_1_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet13_1_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet13_1_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet13_1_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet13_1_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet13_1_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet3_1_1_argbuf_d = (writeQTree_IntlizzieLet13_1_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet13_1_1_argbuf_rwb_bufchan_buf :
                                    writeQTree_IntlizzieLet13_1_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet13_1_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
    else
      if ((lizzieLet3_1_1_argbuf_r && writeQTree_IntlizzieLet13_1_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet13_1_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                 1'd0};
      else if (((! lizzieLet3_1_1_argbuf_r) && (! writeQTree_IntlizzieLet13_1_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet13_1_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet13_1_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet15_2_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet15_2_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet15_2_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet15_2_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet15_2_1_argbuf_r = ((! writeQTree_IntlizzieLet15_2_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet15_2_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet15_2_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet15_2_1_argbuf_r)
        writeQTree_IntlizzieLet15_2_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet15_2_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet15_2_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet15_2_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet15_2_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet15_2_1_argbuf_rwb_d = (writeQTree_IntlizzieLet15_2_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet15_2_1_argbuf_bufchan_buf :
                                                       writeQTree_IntlizzieLet15_2_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet15_2_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet15_2_1_argbuf_rwb_r && writeQTree_IntlizzieLet15_2_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet15_2_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet15_2_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet15_2_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet15_2_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet15_2_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet15_2_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet4_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet15_2_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet15_2_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet15_2_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet15_2_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet15_2_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet15_2_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                             1'd0};
    else
      if (writeQTree_IntlizzieLet15_2_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet15_2_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet15_2_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet15_2_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet15_2_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet15_2_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet4_1_1_argbuf_d = (writeQTree_IntlizzieLet15_2_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet15_2_1_argbuf_rwb_bufchan_buf :
                                    writeQTree_IntlizzieLet15_2_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet15_2_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
    else
      if ((lizzieLet4_1_1_argbuf_r && writeQTree_IntlizzieLet15_2_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet15_2_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                 1'd0};
      else if (((! lizzieLet4_1_1_argbuf_r) && (! writeQTree_IntlizzieLet15_2_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet15_2_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet15_2_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet17_1_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet17_1_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet17_1_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet17_1_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet17_1_1_argbuf_r = ((! writeQTree_IntlizzieLet17_1_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet17_1_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet17_1_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet17_1_1_argbuf_r)
        writeQTree_IntlizzieLet17_1_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet17_1_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet17_1_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet17_1_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet17_1_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet17_1_1_argbuf_rwb_d = (writeQTree_IntlizzieLet17_1_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet17_1_1_argbuf_bufchan_buf :
                                                       writeQTree_IntlizzieLet17_1_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet17_1_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet17_1_1_argbuf_rwb_r && writeQTree_IntlizzieLet17_1_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet17_1_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet17_1_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet17_1_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet17_1_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet17_1_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet17_1_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet6_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet17_1_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet17_1_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet17_1_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet17_1_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet17_1_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet17_1_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                             1'd0};
    else
      if (writeQTree_IntlizzieLet17_1_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet17_1_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet17_1_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet17_1_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet17_1_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet17_1_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet6_1_1_argbuf_d = (writeQTree_IntlizzieLet17_1_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet17_1_1_argbuf_rwb_bufchan_buf :
                                    writeQTree_IntlizzieLet17_1_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet17_1_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
    else
      if ((lizzieLet6_1_1_argbuf_r && writeQTree_IntlizzieLet17_1_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet17_1_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                 1'd0};
      else if (((! lizzieLet6_1_1_argbuf_r) && (! writeQTree_IntlizzieLet17_1_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet17_1_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet17_1_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet18_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet18_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet18_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet18_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet18_1_argbuf_r = ((! writeQTree_IntlizzieLet18_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet18_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet18_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet18_1_argbuf_r)
        writeQTree_IntlizzieLet18_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet18_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet18_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet18_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet18_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet18_1_argbuf_rwb_d = (writeQTree_IntlizzieLet18_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet18_1_argbuf_bufchan_buf :
                                                     writeQTree_IntlizzieLet18_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet18_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet18_1_argbuf_rwb_r && writeQTree_IntlizzieLet18_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet18_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet18_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet18_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet18_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet18_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet18_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet7_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet18_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet18_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet18_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet18_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet18_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet18_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet18_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet18_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet18_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet18_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet18_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet18_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet7_1_1_argbuf_d = (writeQTree_IntlizzieLet18_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet18_1_argbuf_rwb_bufchan_buf :
                                    writeQTree_IntlizzieLet18_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet18_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((lizzieLet7_1_1_argbuf_r && writeQTree_IntlizzieLet18_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet18_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! lizzieLet7_1_1_argbuf_r) && (! writeQTree_IntlizzieLet18_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet18_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet18_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet19_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet19_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet19_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet19_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet19_1_argbuf_r = ((! writeQTree_IntlizzieLet19_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet19_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet19_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet19_1_argbuf_r)
        writeQTree_IntlizzieLet19_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet19_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet19_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet19_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet19_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet19_1_argbuf_rwb_d = (writeQTree_IntlizzieLet19_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet19_1_argbuf_bufchan_buf :
                                                     writeQTree_IntlizzieLet19_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet19_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet19_1_argbuf_rwb_r && writeQTree_IntlizzieLet19_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet19_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet19_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet19_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet19_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet19_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet19_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet8_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet19_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet19_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet19_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet19_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet19_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet19_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet19_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet19_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet19_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet19_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet19_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet19_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet8_1_1_argbuf_d = (writeQTree_IntlizzieLet19_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet19_1_argbuf_rwb_bufchan_buf :
                                    writeQTree_IntlizzieLet19_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet19_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((lizzieLet8_1_1_argbuf_r && writeQTree_IntlizzieLet19_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet19_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! lizzieLet8_1_1_argbuf_r) && (! writeQTree_IntlizzieLet19_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet19_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet19_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet21_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet21_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet21_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet21_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet21_1_argbuf_r = ((! writeQTree_IntlizzieLet21_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet21_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet21_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet21_1_argbuf_r)
        writeQTree_IntlizzieLet21_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet21_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet21_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet21_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet21_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet21_1_argbuf_rwb_d = (writeQTree_IntlizzieLet21_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet21_1_argbuf_bufchan_buf :
                                                     writeQTree_IntlizzieLet21_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet21_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet21_1_argbuf_rwb_r && writeQTree_IntlizzieLet21_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet21_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet21_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet21_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet21_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet21_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet21_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet9_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet21_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet21_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet21_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet21_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet21_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet21_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet21_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet21_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet21_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet21_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet21_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet21_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet9_1_1_argbuf_d = (writeQTree_IntlizzieLet21_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet21_1_argbuf_rwb_bufchan_buf :
                                    writeQTree_IntlizzieLet21_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet21_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((lizzieLet9_1_1_argbuf_r && writeQTree_IntlizzieLet21_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet21_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! lizzieLet9_1_1_argbuf_r) && (! writeQTree_IntlizzieLet21_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet21_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet21_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet33_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet33_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet33_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet33_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet33_1_argbuf_r = ((! writeQTree_IntlizzieLet33_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet33_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet33_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet33_1_argbuf_r)
        writeQTree_IntlizzieLet33_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet33_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet33_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet33_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet33_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet33_1_argbuf_rwb_d = (writeQTree_IntlizzieLet33_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet33_1_argbuf_bufchan_buf :
                                                     writeQTree_IntlizzieLet33_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet33_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet33_1_argbuf_rwb_r && writeQTree_IntlizzieLet33_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet33_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet33_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet33_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet33_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet33_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet33_1_argbuf_rwb,Pointer_QTree_Int) > (contRet_0_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet33_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet33_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet33_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet33_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet33_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet33_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet33_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet33_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet33_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet33_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet33_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet33_1_argbuf_rwb_bufchan_buf[0]);
  assign contRet_0_1_1_argbuf_d = (writeQTree_IntlizzieLet33_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet33_1_argbuf_rwb_bufchan_buf :
                                   writeQTree_IntlizzieLet33_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet33_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((contRet_0_1_1_argbuf_r && writeQTree_IntlizzieLet33_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet33_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! contRet_0_1_1_argbuf_r) && (! writeQTree_IntlizzieLet33_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet33_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet33_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet38_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet38_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet38_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet38_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet38_1_argbuf_r = ((! writeQTree_IntlizzieLet38_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet38_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet38_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet38_1_argbuf_r)
        writeQTree_IntlizzieLet38_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet38_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet38_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet38_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet38_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet38_1_argbuf_rwb_d = (writeQTree_IntlizzieLet38_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet38_1_argbuf_bufchan_buf :
                                                     writeQTree_IntlizzieLet38_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet38_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet38_1_argbuf_rwb_r && writeQTree_IntlizzieLet38_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet38_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet38_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet38_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet38_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet38_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet38_1_argbuf_rwb,Pointer_QTree_Int) > (contRet_0_2_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet38_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet38_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet38_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet38_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet38_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet38_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet38_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet38_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet38_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet38_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet38_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet38_1_argbuf_rwb_bufchan_buf[0]);
  assign contRet_0_2_1_argbuf_d = (writeQTree_IntlizzieLet38_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet38_1_argbuf_rwb_bufchan_buf :
                                   writeQTree_IntlizzieLet38_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet38_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((contRet_0_2_1_argbuf_r && writeQTree_IntlizzieLet38_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet38_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! contRet_0_2_1_argbuf_r) && (! writeQTree_IntlizzieLet38_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet38_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet38_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet43_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet43_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet43_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet43_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet43_1_argbuf_r = ((! writeQTree_IntlizzieLet43_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet43_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet43_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet43_1_argbuf_r)
        writeQTree_IntlizzieLet43_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet43_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet43_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet43_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet43_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet43_1_argbuf_rwb_d = (writeQTree_IntlizzieLet43_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet43_1_argbuf_bufchan_buf :
                                                     writeQTree_IntlizzieLet43_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet43_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet43_1_argbuf_rwb_r && writeQTree_IntlizzieLet43_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet43_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet43_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet43_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet43_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet43_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet43_1_argbuf_rwb,Pointer_QTree_Int) > (contRet_0_3_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet43_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet43_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet43_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet43_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet43_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet43_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet43_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet43_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet43_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet43_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet43_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet43_1_argbuf_rwb_bufchan_buf[0]);
  assign contRet_0_3_1_argbuf_d = (writeQTree_IntlizzieLet43_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet43_1_argbuf_rwb_bufchan_buf :
                                   writeQTree_IntlizzieLet43_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet43_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((contRet_0_3_1_argbuf_r && writeQTree_IntlizzieLet43_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet43_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! contRet_0_3_1_argbuf_r) && (! writeQTree_IntlizzieLet43_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet43_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet43_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet7_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet7_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet7_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet7_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet7_1_argbuf_r = ((! writeQTree_IntlizzieLet7_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet7_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet7_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet7_1_argbuf_r)
        writeQTree_IntlizzieLet7_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet7_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet7_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet7_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet7_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet7_1_argbuf_rwb_d = (writeQTree_IntlizzieLet7_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet7_1_argbuf_bufchan_buf :
                                                    writeQTree_IntlizzieLet7_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet7_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet7_1_argbuf_rwb_r && writeQTree_IntlizzieLet7_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet7_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet7_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet7_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet7_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet7_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet7_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet11_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet7_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet7_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet7_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet7_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet7_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet7_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet7_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet7_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet7_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet7_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet7_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet7_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet11_1_argbuf_d = (writeQTree_IntlizzieLet7_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet7_1_argbuf_rwb_bufchan_buf :
                                   writeQTree_IntlizzieLet7_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet7_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet11_1_argbuf_r && writeQTree_IntlizzieLet7_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet7_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet11_1_argbuf_r) && (! writeQTree_IntlizzieLet7_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet7_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet7_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet9_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet9_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet9_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet9_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet9_1_argbuf_r = ((! writeQTree_IntlizzieLet9_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet9_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet9_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet9_1_argbuf_r)
        writeQTree_IntlizzieLet9_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet9_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet9_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet9_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet9_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet9_1_argbuf_rwb_d = (writeQTree_IntlizzieLet9_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet9_1_argbuf_bufchan_buf :
                                                    writeQTree_IntlizzieLet9_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet9_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet9_1_argbuf_rwb_r && writeQTree_IntlizzieLet9_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet9_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet9_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet9_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet9_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet9_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet9_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet13_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet9_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet9_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet9_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet9_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet9_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet9_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet9_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet9_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet9_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet9_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet9_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet9_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet13_1_argbuf_d = (writeQTree_IntlizzieLet9_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet9_1_argbuf_rwb_bufchan_buf :
                                   writeQTree_IntlizzieLet9_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet9_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet13_1_argbuf_r && writeQTree_IntlizzieLet9_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet9_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet13_1_argbuf_r) && (! writeQTree_IntlizzieLet9_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet9_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet9_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (wsvt_1_goMux_mux,Pointer_QTree_Int) > (wsvt_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t wsvt_1_goMux_mux_bufchan_d;
  logic wsvt_1_goMux_mux_bufchan_r;
  assign wsvt_1_goMux_mux_r = ((! wsvt_1_goMux_mux_bufchan_d[0]) || wsvt_1_goMux_mux_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) wsvt_1_goMux_mux_bufchan_d <= {16'd0, 1'd0};
    else
      if (wsvt_1_goMux_mux_r)
        wsvt_1_goMux_mux_bufchan_d <= wsvt_1_goMux_mux_d;
  Pointer_QTree_Int_t wsvt_1_goMux_mux_bufchan_buf;
  assign wsvt_1_goMux_mux_bufchan_r = (! wsvt_1_goMux_mux_bufchan_buf[0]);
  assign wsvt_1_1_argbuf_d = (wsvt_1_goMux_mux_bufchan_buf[0] ? wsvt_1_goMux_mux_bufchan_buf :
                              wsvt_1_goMux_mux_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) wsvt_1_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((wsvt_1_1_argbuf_r && wsvt_1_goMux_mux_bufchan_buf[0]))
        wsvt_1_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
      else if (((! wsvt_1_1_argbuf_r) && (! wsvt_1_goMux_mux_bufchan_buf[0])))
        wsvt_1_goMux_mux_bufchan_buf <= wsvt_1_goMux_mux_bufchan_d;
  
  /* buf (Ty CT$wnnz_Int) : (wwsvw_1_1lizzieLet25_4Lcall_$wnnz_Int2_1sc_0_5_1q4ac3_2_1Lcall_$wnnz_Int1,CT$wnnz_Int) > (lizzieLet27_1_argbuf,CT$wnnz_Int) */
  CT$wnnz_Int_t wwsvw_1_1lizzieLet25_4Lcall_$wnnz_Int2_1sc_0_5_1q4ac3_2_1Lcall_$wnnz_Int1_bufchan_d;
  logic wwsvw_1_1lizzieLet25_4Lcall_$wnnz_Int2_1sc_0_5_1q4ac3_2_1Lcall_$wnnz_Int1_bufchan_r;
  assign wwsvw_1_1lizzieLet25_4Lcall_$wnnz_Int2_1sc_0_5_1q4ac3_2_1Lcall_$wnnz_Int1_r = ((! wwsvw_1_1lizzieLet25_4Lcall_$wnnz_Int2_1sc_0_5_1q4ac3_2_1Lcall_$wnnz_Int1_bufchan_d[0]) || wwsvw_1_1lizzieLet25_4Lcall_$wnnz_Int2_1sc_0_5_1q4ac3_2_1Lcall_$wnnz_Int1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      wwsvw_1_1lizzieLet25_4Lcall_$wnnz_Int2_1sc_0_5_1q4ac3_2_1Lcall_$wnnz_Int1_bufchan_d <= {115'd0,
                                                                                              1'd0};
    else
      if (wwsvw_1_1lizzieLet25_4Lcall_$wnnz_Int2_1sc_0_5_1q4ac3_2_1Lcall_$wnnz_Int1_r)
        wwsvw_1_1lizzieLet25_4Lcall_$wnnz_Int2_1sc_0_5_1q4ac3_2_1Lcall_$wnnz_Int1_bufchan_d <= wwsvw_1_1lizzieLet25_4Lcall_$wnnz_Int2_1sc_0_5_1q4ac3_2_1Lcall_$wnnz_Int1_d;
  CT$wnnz_Int_t wwsvw_1_1lizzieLet25_4Lcall_$wnnz_Int2_1sc_0_5_1q4ac3_2_1Lcall_$wnnz_Int1_bufchan_buf;
  assign wwsvw_1_1lizzieLet25_4Lcall_$wnnz_Int2_1sc_0_5_1q4ac3_2_1Lcall_$wnnz_Int1_bufchan_r = (! wwsvw_1_1lizzieLet25_4Lcall_$wnnz_Int2_1sc_0_5_1q4ac3_2_1Lcall_$wnnz_Int1_bufchan_buf[0]);
  assign lizzieLet27_1_argbuf_d = (wwsvw_1_1lizzieLet25_4Lcall_$wnnz_Int2_1sc_0_5_1q4ac3_2_1Lcall_$wnnz_Int1_bufchan_buf[0] ? wwsvw_1_1lizzieLet25_4Lcall_$wnnz_Int2_1sc_0_5_1q4ac3_2_1Lcall_$wnnz_Int1_bufchan_buf :
                                   wwsvw_1_1lizzieLet25_4Lcall_$wnnz_Int2_1sc_0_5_1q4ac3_2_1Lcall_$wnnz_Int1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      wwsvw_1_1lizzieLet25_4Lcall_$wnnz_Int2_1sc_0_5_1q4ac3_2_1Lcall_$wnnz_Int1_bufchan_buf <= {115'd0,
                                                                                                1'd0};
    else
      if ((lizzieLet27_1_argbuf_r && wwsvw_1_1lizzieLet25_4Lcall_$wnnz_Int2_1sc_0_5_1q4ac3_2_1Lcall_$wnnz_Int1_bufchan_buf[0]))
        wwsvw_1_1lizzieLet25_4Lcall_$wnnz_Int2_1sc_0_5_1q4ac3_2_1Lcall_$wnnz_Int1_bufchan_buf <= {115'd0,
                                                                                                  1'd0};
      else if (((! lizzieLet27_1_argbuf_r) && (! wwsvw_1_1lizzieLet25_4Lcall_$wnnz_Int2_1sc_0_5_1q4ac3_2_1Lcall_$wnnz_Int1_bufchan_buf[0])))
        wwsvw_1_1lizzieLet25_4Lcall_$wnnz_Int2_1sc_0_5_1q4ac3_2_1Lcall_$wnnz_Int1_bufchan_buf <= wwsvw_1_1lizzieLet25_4Lcall_$wnnz_Int2_1sc_0_5_1q4ac3_2_1Lcall_$wnnz_Int1_bufchan_d;
  
  /* dcon (Ty CT$wnnz_Int,
      Dcon Lcall_$wnnz_Int1) : [(wwsvw_1_destruct,Int#),
                                (lizzieLet25_4Lcall_$wnnz_Int2,Int#),
                                (sc_0_5_destruct,Pointer_CT$wnnz_Int),
                                (q4ac3_2_destruct,Pointer_QTree_Int)] > (wwsvw_1_1lizzieLet25_4Lcall_$wnnz_Int2_1sc_0_5_1q4ac3_2_1Lcall_$wnnz_Int1,CT$wnnz_Int) */
  assign wwsvw_1_1lizzieLet25_4Lcall_$wnnz_Int2_1sc_0_5_1q4ac3_2_1Lcall_$wnnz_Int1_d = Lcall_$wnnz_Int1_dc((& {wwsvw_1_destruct_d[0],
                                                                                                               lizzieLet25_4Lcall_$wnnz_Int2_d[0],
                                                                                                               sc_0_5_destruct_d[0],
                                                                                                               q4ac3_2_destruct_d[0]}), wwsvw_1_destruct_d, lizzieLet25_4Lcall_$wnnz_Int2_d, sc_0_5_destruct_d, q4ac3_2_destruct_d);
  assign {wwsvw_1_destruct_r,
          lizzieLet25_4Lcall_$wnnz_Int2_r,
          sc_0_5_destruct_r,
          q4ac3_2_destruct_r} = {4 {(wwsvw_1_1lizzieLet25_4Lcall_$wnnz_Int2_1sc_0_5_1q4ac3_2_1Lcall_$wnnz_Int1_r && wwsvw_1_1lizzieLet25_4Lcall_$wnnz_Int2_1sc_0_5_1q4ac3_2_1Lcall_$wnnz_Int1_d[0])}};
  
  /* buf (Ty CT$wnnz_Int) : (wwsvw_2_1ww1XwI_1_1lizzieLet25_4Lcall_$wnnz_Int1_1sc_0_6_1Lcall_$wnnz_Int0,CT$wnnz_Int) > (lizzieLet28_1_argbuf,CT$wnnz_Int) */
  CT$wnnz_Int_t wwsvw_2_1ww1XwI_1_1lizzieLet25_4Lcall_$wnnz_Int1_1sc_0_6_1Lcall_$wnnz_Int0_bufchan_d;
  logic wwsvw_2_1ww1XwI_1_1lizzieLet25_4Lcall_$wnnz_Int1_1sc_0_6_1Lcall_$wnnz_Int0_bufchan_r;
  assign wwsvw_2_1ww1XwI_1_1lizzieLet25_4Lcall_$wnnz_Int1_1sc_0_6_1Lcall_$wnnz_Int0_r = ((! wwsvw_2_1ww1XwI_1_1lizzieLet25_4Lcall_$wnnz_Int1_1sc_0_6_1Lcall_$wnnz_Int0_bufchan_d[0]) || wwsvw_2_1ww1XwI_1_1lizzieLet25_4Lcall_$wnnz_Int1_1sc_0_6_1Lcall_$wnnz_Int0_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      wwsvw_2_1ww1XwI_1_1lizzieLet25_4Lcall_$wnnz_Int1_1sc_0_6_1Lcall_$wnnz_Int0_bufchan_d <= {115'd0,
                                                                                               1'd0};
    else
      if (wwsvw_2_1ww1XwI_1_1lizzieLet25_4Lcall_$wnnz_Int1_1sc_0_6_1Lcall_$wnnz_Int0_r)
        wwsvw_2_1ww1XwI_1_1lizzieLet25_4Lcall_$wnnz_Int1_1sc_0_6_1Lcall_$wnnz_Int0_bufchan_d <= wwsvw_2_1ww1XwI_1_1lizzieLet25_4Lcall_$wnnz_Int1_1sc_0_6_1Lcall_$wnnz_Int0_d;
  CT$wnnz_Int_t wwsvw_2_1ww1XwI_1_1lizzieLet25_4Lcall_$wnnz_Int1_1sc_0_6_1Lcall_$wnnz_Int0_bufchan_buf;
  assign wwsvw_2_1ww1XwI_1_1lizzieLet25_4Lcall_$wnnz_Int1_1sc_0_6_1Lcall_$wnnz_Int0_bufchan_r = (! wwsvw_2_1ww1XwI_1_1lizzieLet25_4Lcall_$wnnz_Int1_1sc_0_6_1Lcall_$wnnz_Int0_bufchan_buf[0]);
  assign lizzieLet28_1_argbuf_d = (wwsvw_2_1ww1XwI_1_1lizzieLet25_4Lcall_$wnnz_Int1_1sc_0_6_1Lcall_$wnnz_Int0_bufchan_buf[0] ? wwsvw_2_1ww1XwI_1_1lizzieLet25_4Lcall_$wnnz_Int1_1sc_0_6_1Lcall_$wnnz_Int0_bufchan_buf :
                                   wwsvw_2_1ww1XwI_1_1lizzieLet25_4Lcall_$wnnz_Int1_1sc_0_6_1Lcall_$wnnz_Int0_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      wwsvw_2_1ww1XwI_1_1lizzieLet25_4Lcall_$wnnz_Int1_1sc_0_6_1Lcall_$wnnz_Int0_bufchan_buf <= {115'd0,
                                                                                                 1'd0};
    else
      if ((lizzieLet28_1_argbuf_r && wwsvw_2_1ww1XwI_1_1lizzieLet25_4Lcall_$wnnz_Int1_1sc_0_6_1Lcall_$wnnz_Int0_bufchan_buf[0]))
        wwsvw_2_1ww1XwI_1_1lizzieLet25_4Lcall_$wnnz_Int1_1sc_0_6_1Lcall_$wnnz_Int0_bufchan_buf <= {115'd0,
                                                                                                   1'd0};
      else if (((! lizzieLet28_1_argbuf_r) && (! wwsvw_2_1ww1XwI_1_1lizzieLet25_4Lcall_$wnnz_Int1_1sc_0_6_1Lcall_$wnnz_Int0_bufchan_buf[0])))
        wwsvw_2_1ww1XwI_1_1lizzieLet25_4Lcall_$wnnz_Int1_1sc_0_6_1Lcall_$wnnz_Int0_bufchan_buf <= wwsvw_2_1ww1XwI_1_1lizzieLet25_4Lcall_$wnnz_Int1_1sc_0_6_1Lcall_$wnnz_Int0_bufchan_d;
  
  /* dcon (Ty CT$wnnz_Int,
      Dcon Lcall_$wnnz_Int0) : [(wwsvw_2_destruct,Int#),
                                (ww1XwI_1_destruct,Int#),
                                (lizzieLet25_4Lcall_$wnnz_Int1,Int#),
                                (sc_0_6_destruct,Pointer_CT$wnnz_Int)] > (wwsvw_2_1ww1XwI_1_1lizzieLet25_4Lcall_$wnnz_Int1_1sc_0_6_1Lcall_$wnnz_Int0,CT$wnnz_Int) */
  assign wwsvw_2_1ww1XwI_1_1lizzieLet25_4Lcall_$wnnz_Int1_1sc_0_6_1Lcall_$wnnz_Int0_d = Lcall_$wnnz_Int0_dc((& {wwsvw_2_destruct_d[0],
                                                                                                                ww1XwI_1_destruct_d[0],
                                                                                                                lizzieLet25_4Lcall_$wnnz_Int1_d[0],
                                                                                                                sc_0_6_destruct_d[0]}), wwsvw_2_destruct_d, ww1XwI_1_destruct_d, lizzieLet25_4Lcall_$wnnz_Int1_d, sc_0_6_destruct_d);
  assign {wwsvw_2_destruct_r,
          ww1XwI_1_destruct_r,
          lizzieLet25_4Lcall_$wnnz_Int1_r,
          sc_0_6_destruct_r} = {4 {(wwsvw_2_1ww1XwI_1_1lizzieLet25_4Lcall_$wnnz_Int1_1sc_0_6_1Lcall_$wnnz_Int0_r && wwsvw_2_1ww1XwI_1_1lizzieLet25_4Lcall_$wnnz_Int1_1sc_0_6_1Lcall_$wnnz_Int0_d[0])}};
  
  /* op_add (Ty Int#) : (wwsvw_3_1ww1XwI_2_1_Add32,Int#) (ww2XwL_1_destruct,Int#) > (es_6_1ww2XwL_1_1_Add32,Int#) */
  assign es_6_1ww2XwL_1_1_Add32_d = {(wwsvw_3_1ww1XwI_2_1_Add32_d[32:1] + ww2XwL_1_destruct_d[32:1]),
                                     (wwsvw_3_1ww1XwI_2_1_Add32_d[0] && ww2XwL_1_destruct_d[0])};
  assign {wwsvw_3_1ww1XwI_2_1_Add32_r,
          ww2XwL_1_destruct_r} = {2 {(es_6_1ww2XwL_1_1_Add32_r && es_6_1ww2XwL_1_1_Add32_d[0])}};
  
  /* op_add (Ty Int#) : (wwsvw_3_destruct,Int#) (ww1XwI_2_destruct,Int#) > (wwsvw_3_1ww1XwI_2_1_Add32,Int#) */
  assign wwsvw_3_1ww1XwI_2_1_Add32_d = {(wwsvw_3_destruct_d[32:1] + ww1XwI_2_destruct_d[32:1]),
                                        (wwsvw_3_destruct_d[0] && ww1XwI_2_destruct_d[0])};
  assign {wwsvw_3_destruct_r,
          ww1XwI_2_destruct_r} = {2 {(wwsvw_3_1ww1XwI_2_1_Add32_r && wwsvw_3_1ww1XwI_2_1_Add32_d[0])}};
  
  /* buf (Ty Int) : (xacr_1,Int) > (xacr_1_argbuf,Int) */
  Int_t xacr_1_bufchan_d;
  logic xacr_1_bufchan_r;
  assign xacr_1_r = ((! xacr_1_bufchan_d[0]) || xacr_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) xacr_1_bufchan_d <= {32'd0, 1'd0};
    else if (xacr_1_r) xacr_1_bufchan_d <= xacr_1_d;
  Int_t xacr_1_bufchan_buf;
  assign xacr_1_bufchan_r = (! xacr_1_bufchan_buf[0]);
  assign xacr_1_argbuf_d = (xacr_1_bufchan_buf[0] ? xacr_1_bufchan_buf :
                            xacr_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) xacr_1_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((xacr_1_argbuf_r && xacr_1_bufchan_buf[0]))
        xacr_1_bufchan_buf <= {32'd0, 1'd0};
      else if (((! xacr_1_argbuf_r) && (! xacr_1_bufchan_buf[0])))
        xacr_1_bufchan_buf <= xacr_1_bufchan_d;
  
  /* buf (Ty Int) : (xacr_1_1,Int) > (xacr_1_1_argbuf,Int) */
  Int_t xacr_1_1_bufchan_d;
  logic xacr_1_1_bufchan_r;
  assign xacr_1_1_r = ((! xacr_1_1_bufchan_d[0]) || xacr_1_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) xacr_1_1_bufchan_d <= {32'd0, 1'd0};
    else if (xacr_1_1_r) xacr_1_1_bufchan_d <= xacr_1_1_d;
  Int_t xacr_1_1_bufchan_buf;
  assign xacr_1_1_bufchan_r = (! xacr_1_1_bufchan_buf[0]);
  assign xacr_1_1_argbuf_d = (xacr_1_1_bufchan_buf[0] ? xacr_1_1_bufchan_buf :
                              xacr_1_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) xacr_1_1_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((xacr_1_1_argbuf_r && xacr_1_1_bufchan_buf[0]))
        xacr_1_1_bufchan_buf <= {32'd0, 1'd0};
      else if (((! xacr_1_1_argbuf_r) && (! xacr_1_1_bufchan_buf[0])))
        xacr_1_1_bufchan_buf <= xacr_1_1_bufchan_d;
  
  /* dcon (Ty Int,
      Dcon I#) : [(xaqa_1lizzieLet0_1_1_Add32,Int#)] > (es_0_2_1I#,Int) */
  assign \es_0_2_1I#_d  = \I#_dc ((& {xaqa_1lizzieLet0_1_1_Add32_d[0]}), xaqa_1lizzieLet0_1_1_Add32_d);
  assign {xaqa_1lizzieLet0_1_1_Add32_r} = {1 {(\es_0_2_1I#_r  && \es_0_2_1I#_d [0])}};
  
  /* op_add (Ty Int#) : (xaqa_destruct,Int#) (arg0_2_1Dcon_main1_3I#_1_argbuf_2,Int#) > (xaqa_1lizzieLet0_1_1_Add32,Int#) */
  assign xaqa_1lizzieLet0_1_1_Add32_d = {(xaqa_destruct_d[32:1] + \arg0_2_1Dcon_main1_3I#_1_argbuf_2_d [32:1]),
                                         (xaqa_destruct_d[0] && \arg0_2_1Dcon_main1_3I#_1_argbuf_2_d [0])};
  assign {xaqa_destruct_r,
          \arg0_2_1Dcon_main1_3I#_1_argbuf_2_r } = {2 {(xaqa_1lizzieLet0_1_1_Add32_r && xaqa_1lizzieLet0_1_1_Add32_d[0])}};
endmodule