`timescale 1ns/1ns
import mMaskAdd_package::*;

module mMaskAdd(
  input logic clk,
  input logic reset,
  input Go_t \\QTree_Bool_src_d ,
  output logic \\QTree_Bool_src_r ,
  input QTree_Bool_t dummy_write_QTree_Bool_d,
  output logic dummy_write_QTree_Bool_r,
  input Go_t \\MaskQTree_src_d ,
  output logic \\MaskQTree_src_r ,
  input MaskQTree_t dummy_write_MaskQTree_d,
  output logic dummy_write_MaskQTree_r,
  input Go_t sourceGo_d,
  output logic sourceGo_r,
  input Pointer_MaskQTree_t m1a82_0_d,
  output logic m1a82_0_r,
  input Pointer_QTree_Bool_t m2a83_1_d,
  output logic m2a83_1_r,
  input Pointer_QTree_Bool_t m3a84_2_d,
  output logic m3a84_2_r,
  output \Word16#_t  forkHP1_QTree_Bool_snk_dout,
  input logic forkHP1_QTree_Bool_snk_rout,
  output Pointer_QTree_Bool_t dummy_write_QTree_Bool_sink_dout,
  input logic dummy_write_QTree_Bool_sink_rout,
  output \Word16#_t  forkHP1_MaskQTree_snk_dout,
  input logic forkHP1_MaskQTree_snk_rout,
  output Pointer_MaskQTree_t dummy_write_MaskQTree_sink_dout,
  input logic dummy_write_MaskQTree_sink_rout,
  output Pointer_QTree_Bool_t f_resbuf_dout,
  input logic f_resbuf_rout
  );
  /* --define=INPUTS=((__05CQTree_Bool_src, 0, 1, Go), (dummy_write_QTree_Bool, 66, 73786976294838206464, QTree_Bool), (__05CMaskQTree_src, 0, 1, Go), (dummy_write_MaskQTree, 66, 73786976294838206464, MaskQTree), (sourceGo, 0, 1, Go), (m1a82_0, 16, 65536, Pointer_MaskQTree), (m2a83_1, 16, 65536, Pointer_QTree_Bool), (m3a84_2, 16, 65536, Pointer_QTree_Bool)) */
  /* --define=TAPS=() */
  /* --define=OUTPUTS=((forkHP1_QTree_Bool_snk, 16, 65536, Word16__023), (dummy_write_QTree_Bool_sink, 16, 65536, Pointer_QTree_Bool), (forkHP1_MaskQTree_snk, 16, 65536, Word16__023), (dummy_write_MaskQTree_sink, 16, 65536, Pointer_MaskQTree), (f_resbuf, 16, 65536, Pointer_QTree_Bool)) */
  /* TYPE_START
QTree_Bool 16 2 (0,[0]) (1,[1]) (2,[16p,16p,16p,16p]) (3,[0])
CTf 16 3 (0,[0]) (1,[16p,16p,16p,16p,16p,16p,16p,16p,16p,16p]) (2,[16p,16p,16p,16p,16p,16p,16p,16p]) (3,[16p,16p,16p,16p,16p,16p]) (4,[16p,16p,16p,16p])
CTf__027 16 3 (0,[0]) (1,[16p,16p,16p,16p,16p,16p,16p]) (2,[16p,16p,16p,16p,16p,16p]) (3,[16p,16p,16p,16p,16p]) (4,[16p,16p,16p,16p])
CTf__027__027__027__027__027__027__027__027__027_f__027__027__027__027__027__027__027__027__027_Bool 16 3 (0,[0]) (1,[16p,16p,16p,16p,16p,16p,16p]) (2,[16p,16p,16p,16p,16p,16p]) (3,[16p,16p,16p,16p,16p]) (4,[16p,16p,16p,16p])
MaskQTree 16 2 (0,[0]) (1,[0]) (2,[16p,16p,16p,16p])
TupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_CTf__027__027__027__027__027__027__027__027__027_f__027__027__027__027__027__027__027__027__027_Bool 16 0 (0,[0,16p,16p,16p])
TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf__027 16 0 (0,[0,16p,16p,16p])
TupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf 16 0 (0,[0,16p,16p,16p,16p])
TupGo___Pointer_MaskQTree___Pointer_QTree_Bool 16 0 (0,[0,16p,16p])
TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool 16 0 (0,[0,16p,16p])
TupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool 16 0 (0,[0,16p,16p,16p])
TYPE_END */
  /*  */
  /*  */
  Go_t goFork_d;
  logic goFork_r;
  Go_t goFor_2_d;
  logic goFor_2_r;
  Go_t goFor_3_d;
  logic goFor_3_r;
  Go_t goFor_4_d;
  logic goFor_4_r;
  Go_t goFor_5_d;
  logic goFor_5_r;
  Go_t goFor_6_d;
  logic goFor_6_r;
  Go_t goFor_7_d;
  logic goFor_7_r;
  \Word16#_t  initHP_QTree_Bool_d;
  logic initHP_QTree_Bool_r;
  \Word16#_t  incrHP_QTree_Bool_d;
  logic incrHP_QTree_Bool_r;
  Go_t incrHP_mergeQTree_Bool_d;
  logic incrHP_mergeQTree_Bool_r;
  Go_t incrHP_QTree_Bool1_d;
  logic incrHP_QTree_Bool1_r;
  Go_t incrHP_QTree_Bool2_d;
  logic incrHP_QTree_Bool2_r;
  \Word16#_t  addHP_QTree_Bool_d;
  logic addHP_QTree_Bool_r;
  \Word16#_t  mergeHP_QTree_Bool_d;
  logic mergeHP_QTree_Bool_r;
  Go_t incrHP_mergeQTree_Bool_buf_d;
  logic incrHP_mergeQTree_Bool_buf_r;
  \Word16#_t  mergeHP_QTree_Bool_buf_d;
  logic mergeHP_QTree_Bool_buf_r;
  Go_t go_1_dummy_write_QTree_Bool_d;
  logic go_1_dummy_write_QTree_Bool_r;
  Go_t go_2_dummy_write_QTree_Bool_d;
  logic go_2_dummy_write_QTree_Bool_r;
  \Word16#_t  forkHP1_QTree_Bool_d;
  logic forkHP1_QTree_Bool_r;
  \Word16#_t  forkHP1_QTree_Bool_snk_d;
  logic forkHP1_QTree_Bool_snk_r;
  \Word16#_t  forkHP1_QTree_Boo3_d;
  logic forkHP1_QTree_Boo3_r;
  \Word16#_t  forkHP1_QTree_Boo4_d;
  logic forkHP1_QTree_Boo4_r;
  C2_t memMergeChoice_QTree_Bool_d;
  logic memMergeChoice_QTree_Bool_r;
  MemIn_QTree_Bool_t memMergeIn_QTree_Bool_d;
  logic memMergeIn_QTree_Bool_r;
  MemOut_QTree_Bool_t memOut_QTree_Bool_d;
  logic memOut_QTree_Bool_r;
  MemOut_QTree_Bool_t memReadOut_QTree_Bool_d;
  logic memReadOut_QTree_Bool_r;
  MemOut_QTree_Bool_t memWriteOut_QTree_Bool_d;
  logic memWriteOut_QTree_Bool_r;
  MemIn_QTree_Bool_t memMergeIn_QTree_Bool_dbuf_d;
  logic memMergeIn_QTree_Bool_dbuf_r;
  MemIn_QTree_Bool_t memMergeIn_QTree_Bool_rbuf_d;
  logic memMergeIn_QTree_Bool_rbuf_r;
  MemOut_QTree_Bool_t memOut_QTree_Bool_dbuf_d;
  logic memOut_QTree_Bool_dbuf_r;
  MemOut_QTree_Bool_t memOut_QTree_Bool_rbuf_d;
  logic memOut_QTree_Bool_rbuf_r;
  C5_t readMerge_choice_QTree_Bool_d;
  logic readMerge_choice_QTree_Bool_r;
  Pointer_QTree_Bool_t readMerge_data_QTree_Bool_d;
  logic readMerge_data_QTree_Bool_r;
  QTree_Bool_t readPointer_QTree_Boolm2a86_1_argbuf_d;
  logic readPointer_QTree_Boolm2a86_1_argbuf_r;
  QTree_Bool_t readPointer_QTree_Boolm2a8H_1_argbuf_d;
  logic readPointer_QTree_Boolm2a8H_1_argbuf_r;
  QTree_Bool_t readPointer_QTree_Boolm3a87_1_argbuf_d;
  logic readPointer_QTree_Boolm3a87_1_argbuf_r;
  QTree_Bool_t readPointer_QTree_Boolm3a8I_1_argbuf_d;
  logic readPointer_QTree_Boolm3a8I_1_argbuf_r;
  QTree_Bool_t \readPointer_QTree_Boolq4'a8x_1_argbuf_d ;
  logic \readPointer_QTree_Boolq4'a8x_1_argbuf_r ;
  \Word16#_t  destructReadIn_QTree_Bool_d;
  logic destructReadIn_QTree_Bool_r;
  MemIn_QTree_Bool_t dconReadIn_QTree_Bool_d;
  logic dconReadIn_QTree_Bool_r;
  QTree_Bool_t destructReadOut_QTree_Bool_d;
  logic destructReadOut_QTree_Bool_r;
  C30_t writeMerge_choice_QTree_Bool_d;
  logic writeMerge_choice_QTree_Bool_r;
  QTree_Bool_t writeMerge_data_QTree_Bool_d;
  logic writeMerge_data_QTree_Bool_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet10_1_argbuf_d;
  logic writeQTree_BoollizzieLet10_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet11_1_argbuf_d;
  logic writeQTree_BoollizzieLet11_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet12_1_argbuf_d;
  logic writeQTree_BoollizzieLet12_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet13_1_1_argbuf_d;
  logic writeQTree_BoollizzieLet13_1_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet15_1_1_argbuf_d;
  logic writeQTree_BoollizzieLet15_1_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet16_1_1_argbuf_d;
  logic writeQTree_BoollizzieLet16_1_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet18_1_1_argbuf_d;
  logic writeQTree_BoollizzieLet18_1_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet19_2_1_argbuf_d;
  logic writeQTree_BoollizzieLet19_2_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet1_1_argbuf_d;
  logic writeQTree_BoollizzieLet1_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet22_1_1_argbuf_d;
  logic writeQTree_BoollizzieLet22_1_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet25_1_1_argbuf_d;
  logic writeQTree_BoollizzieLet25_1_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet26_1_1_argbuf_d;
  logic writeQTree_BoollizzieLet26_1_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet28_1_argbuf_d;
  logic writeQTree_BoollizzieLet28_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet30_1_argbuf_d;
  logic writeQTree_BoollizzieLet30_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet31_1_argbuf_d;
  logic writeQTree_BoollizzieLet31_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet33_1_argbuf_d;
  logic writeQTree_BoollizzieLet33_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet35_1_argbuf_d;
  logic writeQTree_BoollizzieLet35_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet36_1_argbuf_d;
  logic writeQTree_BoollizzieLet36_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet38_1_argbuf_d;
  logic writeQTree_BoollizzieLet38_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet42_1_argbuf_d;
  logic writeQTree_BoollizzieLet42_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet47_1_argbuf_d;
  logic writeQTree_BoollizzieLet47_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet4_1_argbuf_d;
  logic writeQTree_BoollizzieLet4_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet52_1_argbuf_d;
  logic writeQTree_BoollizzieLet52_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet57_1_argbuf_d;
  logic writeQTree_BoollizzieLet57_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet5_1_argbuf_d;
  logic writeQTree_BoollizzieLet5_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet6_1_argbuf_d;
  logic writeQTree_BoollizzieLet6_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet7_1_argbuf_d;
  logic writeQTree_BoollizzieLet7_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet9_1_1_argbuf_d;
  logic writeQTree_BoollizzieLet9_1_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet9_1_argbuf_d;
  logic writeQTree_BoollizzieLet9_1_argbuf_r;
  Pointer_QTree_Bool_t dummy_write_QTree_Bool_sink_d;
  logic dummy_write_QTree_Bool_sink_r;
  MemIn_QTree_Bool_t dconWriteIn_QTree_Bool_d;
  logic dconWriteIn_QTree_Bool_r;
  Pointer_QTree_Bool_t dconPtr_QTree_Bool_d;
  logic dconPtr_QTree_Bool_r;
  Pointer_QTree_Bool_t _130_d;
  logic _130_r;
  assign _130_r = 1'd1;
  Pointer_QTree_Bool_t demuxWriteResult_QTree_Bool_d;
  logic demuxWriteResult_QTree_Bool_r;
  \Word16#_t  initHP_CTf_d;
  logic initHP_CTf_r;
  \Word16#_t  incrHP_CTf_d;
  logic incrHP_CTf_r;
  Go_t incrHP_mergeCTf_d;
  logic incrHP_mergeCTf_r;
  Go_t incrHP_CTf1_d;
  logic incrHP_CTf1_r;
  Go_t incrHP_CTf2_d;
  logic incrHP_CTf2_r;
  \Word16#_t  addHP_CTf_d;
  logic addHP_CTf_r;
  \Word16#_t  mergeHP_CTf_d;
  logic mergeHP_CTf_r;
  Go_t incrHP_mergeCTf_buf_d;
  logic incrHP_mergeCTf_buf_r;
  \Word16#_t  mergeHP_CTf_buf_d;
  logic mergeHP_CTf_buf_r;
  \Word16#_t  forkHP1_CTf_d;
  logic forkHP1_CTf_r;
  \Word16#_t  forkHP1_CT2_d;
  logic forkHP1_CT2_r;
  \Word16#_t  forkHP1_CT3_d;
  logic forkHP1_CT3_r;
  C2_t memMergeChoice_CTf_d;
  logic memMergeChoice_CTf_r;
  MemIn_CTf_t memMergeIn_CTf_d;
  logic memMergeIn_CTf_r;
  MemOut_CTf_t memOut_CTf_d;
  logic memOut_CTf_r;
  MemOut_CTf_t memReadOut_CTf_d;
  logic memReadOut_CTf_r;
  MemOut_CTf_t memWriteOut_CTf_d;
  logic memWriteOut_CTf_r;
  MemIn_CTf_t memMergeIn_CTf_dbuf_d;
  logic memMergeIn_CTf_dbuf_r;
  MemIn_CTf_t memMergeIn_CTf_rbuf_d;
  logic memMergeIn_CTf_rbuf_r;
  MemOut_CTf_t memOut_CTf_dbuf_d;
  logic memOut_CTf_dbuf_r;
  MemOut_CTf_t memOut_CTf_rbuf_d;
  logic memOut_CTf_rbuf_r;
  \Word16#_t  destructReadIn_CTf_d;
  logic destructReadIn_CTf_r;
  MemIn_CTf_t dconReadIn_CTf_d;
  logic dconReadIn_CTf_r;
  CTf_t readPointer_CTfscfarg_0_1_argbuf_d;
  logic readPointer_CTfscfarg_0_1_argbuf_r;
  C5_t writeMerge_choice_CTf_d;
  logic writeMerge_choice_CTf_r;
  CTf_t writeMerge_data_CTf_d;
  logic writeMerge_data_CTf_r;
  Pointer_CTf_t writeCTflizzieLet17_1_1_argbuf_d;
  logic writeCTflizzieLet17_1_1_argbuf_r;
  Pointer_CTf_t writeCTflizzieLet39_1_argbuf_d;
  logic writeCTflizzieLet39_1_argbuf_r;
  Pointer_CTf_t writeCTflizzieLet44_1_argbuf_d;
  logic writeCTflizzieLet44_1_argbuf_r;
  Pointer_CTf_t writeCTflizzieLet45_1_argbuf_d;
  logic writeCTflizzieLet45_1_argbuf_r;
  Pointer_CTf_t writeCTflizzieLet46_1_argbuf_d;
  logic writeCTflizzieLet46_1_argbuf_r;
  MemIn_CTf_t dconWriteIn_CTf_d;
  logic dconWriteIn_CTf_r;
  Pointer_CTf_t dconPtr_CTf_d;
  logic dconPtr_CTf_r;
  Pointer_CTf_t _129_d;
  logic _129_r;
  assign _129_r = 1'd1;
  Pointer_CTf_t demuxWriteResult_CTf_d;
  logic demuxWriteResult_CTf_r;
  \Word16#_t  \initHP_CTf'_d ;
  logic \initHP_CTf'_r ;
  \Word16#_t  \incrHP_CTf'_d ;
  logic \incrHP_CTf'_r ;
  Go_t \incrHP_mergeCTf'_d ;
  logic \incrHP_mergeCTf'_r ;
  Go_t \incrHP_CTf'1_d ;
  logic \incrHP_CTf'1_r ;
  Go_t \incrHP_CTf'2_d ;
  logic \incrHP_CTf'2_r ;
  \Word16#_t  \addHP_CTf'_d ;
  logic \addHP_CTf'_r ;
  \Word16#_t  \mergeHP_CTf'_d ;
  logic \mergeHP_CTf'_r ;
  Go_t \incrHP_mergeCTf'_buf_d ;
  logic \incrHP_mergeCTf'_buf_r ;
  \Word16#_t  \mergeHP_CTf'_buf_d ;
  logic \mergeHP_CTf'_buf_r ;
  \Word16#_t  \forkHP1_CTf'_d ;
  logic \forkHP1_CTf'_r ;
  \Word16#_t  forkHP1_CTf2_d;
  logic forkHP1_CTf2_r;
  \Word16#_t  forkHP1_CTf3_d;
  logic forkHP1_CTf3_r;
  C2_t \memMergeChoice_CTf'_d ;
  logic \memMergeChoice_CTf'_r ;
  \MemIn_CTf'_t  \memMergeIn_CTf'_d ;
  logic \memMergeIn_CTf'_r ;
  \MemOut_CTf'_t  \memOut_CTf'_d ;
  logic \memOut_CTf'_r ;
  \MemOut_CTf'_t  \memReadOut_CTf'_d ;
  logic \memReadOut_CTf'_r ;
  \MemOut_CTf'_t  \memWriteOut_CTf'_d ;
  logic \memWriteOut_CTf'_r ;
  \MemIn_CTf'_t  \memMergeIn_CTf'_dbuf_d ;
  logic \memMergeIn_CTf'_dbuf_r ;
  \MemIn_CTf'_t  \memMergeIn_CTf'_rbuf_d ;
  logic \memMergeIn_CTf'_rbuf_r ;
  \MemOut_CTf'_t  \memOut_CTf'_dbuf_d ;
  logic \memOut_CTf'_dbuf_r ;
  \MemOut_CTf'_t  \memOut_CTf'_rbuf_d ;
  logic \memOut_CTf'_rbuf_r ;
  \Word16#_t  \destructReadIn_CTf'_d ;
  logic \destructReadIn_CTf'_r ;
  \MemIn_CTf'_t  \dconReadIn_CTf'_d ;
  logic \dconReadIn_CTf'_r ;
  \CTf'_t  \readPointer_CTf'scfarg_0_1_1_argbuf_d ;
  logic \readPointer_CTf'scfarg_0_1_1_argbuf_r ;
  C5_t \writeMerge_choice_CTf'_d ;
  logic \writeMerge_choice_CTf'_r ;
  \CTf'_t  \writeMerge_data_CTf'_d ;
  logic \writeMerge_data_CTf'_r ;
  \Pointer_CTf'_t  \writeCTf'lizzieLet29_1_argbuf_d ;
  logic \writeCTf'lizzieLet29_1_argbuf_r ;
  \Pointer_CTf'_t  \writeCTf'lizzieLet40_1_argbuf_d ;
  logic \writeCTf'lizzieLet40_1_argbuf_r ;
  \Pointer_CTf'_t  \writeCTf'lizzieLet49_1_argbuf_d ;
  logic \writeCTf'lizzieLet49_1_argbuf_r ;
  \Pointer_CTf'_t  \writeCTf'lizzieLet50_1_argbuf_d ;
  logic \writeCTf'lizzieLet50_1_argbuf_r ;
  \Pointer_CTf'_t  \writeCTf'lizzieLet51_1_argbuf_d ;
  logic \writeCTf'lizzieLet51_1_argbuf_r ;
  \MemIn_CTf'_t  \dconWriteIn_CTf'_d ;
  logic \dconWriteIn_CTf'_r ;
  \Pointer_CTf'_t  \dconPtr_CTf'_d ;
  logic \dconPtr_CTf'_r ;
  \Pointer_CTf'_t  _128_d;
  logic _128_r;
  assign _128_r = 1'd1;
  \Pointer_CTf'_t  \demuxWriteResult_CTf'_d ;
  logic \demuxWriteResult_CTf'_r ;
  \Word16#_t  \initHP_CTf'''''''''_f'''''''''_Bool_d ;
  logic \initHP_CTf'''''''''_f'''''''''_Bool_r ;
  \Word16#_t  \incrHP_CTf'''''''''_f'''''''''_Bool_d ;
  logic \incrHP_CTf'''''''''_f'''''''''_Bool_r ;
  Go_t \incrHP_mergeCTf'''''''''_f'''''''''_Bool_d ;
  logic \incrHP_mergeCTf'''''''''_f'''''''''_Bool_r ;
  Go_t \incrHP_CTf'''''''''_f'''''''''_Bool1_d ;
  logic \incrHP_CTf'''''''''_f'''''''''_Bool1_r ;
  Go_t \incrHP_CTf'''''''''_f'''''''''_Bool2_d ;
  logic \incrHP_CTf'''''''''_f'''''''''_Bool2_r ;
  \Word16#_t  \addHP_CTf'''''''''_f'''''''''_Bool_d ;
  logic \addHP_CTf'''''''''_f'''''''''_Bool_r ;
  \Word16#_t  \mergeHP_CTf'''''''''_f'''''''''_Bool_d ;
  logic \mergeHP_CTf'''''''''_f'''''''''_Bool_r ;
  Go_t \incrHP_mergeCTf'''''''''_f'''''''''_Bool_buf_d ;
  logic \incrHP_mergeCTf'''''''''_f'''''''''_Bool_buf_r ;
  \Word16#_t  \mergeHP_CTf'''''''''_f'''''''''_Bool_buf_d ;
  logic \mergeHP_CTf'''''''''_f'''''''''_Bool_buf_r ;
  \Word16#_t  \forkHP1_CTf'''''''''_f'''''''''_Bool_d ;
  logic \forkHP1_CTf'''''''''_f'''''''''_Bool_r ;
  \Word16#_t  \forkHP1_CTf'''''''''_f'''''''''_Boo2_d ;
  logic \forkHP1_CTf'''''''''_f'''''''''_Boo2_r ;
  \Word16#_t  \forkHP1_CTf'''''''''_f'''''''''_Boo3_d ;
  logic \forkHP1_CTf'''''''''_f'''''''''_Boo3_r ;
  C2_t \memMergeChoice_CTf'''''''''_f'''''''''_Bool_d ;
  logic \memMergeChoice_CTf'''''''''_f'''''''''_Bool_r ;
  \MemIn_CTf'''''''''_f'''''''''_Bool_t  \memMergeIn_CTf'''''''''_f'''''''''_Bool_d ;
  logic \memMergeIn_CTf'''''''''_f'''''''''_Bool_r ;
  \MemOut_CTf'''''''''_f'''''''''_Bool_t  \memOut_CTf'''''''''_f'''''''''_Bool_d ;
  logic \memOut_CTf'''''''''_f'''''''''_Bool_r ;
  \MemOut_CTf'''''''''_f'''''''''_Bool_t  \memReadOut_CTf'''''''''_f'''''''''_Bool_d ;
  logic \memReadOut_CTf'''''''''_f'''''''''_Bool_r ;
  \MemOut_CTf'''''''''_f'''''''''_Bool_t  \memWriteOut_CTf'''''''''_f'''''''''_Bool_d ;
  logic \memWriteOut_CTf'''''''''_f'''''''''_Bool_r ;
  \MemIn_CTf'''''''''_f'''''''''_Bool_t  \memMergeIn_CTf'''''''''_f'''''''''_Bool_dbuf_d ;
  logic \memMergeIn_CTf'''''''''_f'''''''''_Bool_dbuf_r ;
  \MemIn_CTf'''''''''_f'''''''''_Bool_t  \memMergeIn_CTf'''''''''_f'''''''''_Bool_rbuf_d ;
  logic \memMergeIn_CTf'''''''''_f'''''''''_Bool_rbuf_r ;
  \MemOut_CTf'''''''''_f'''''''''_Bool_t  \memOut_CTf'''''''''_f'''''''''_Bool_dbuf_d ;
  logic \memOut_CTf'''''''''_f'''''''''_Bool_dbuf_r ;
  \MemOut_CTf'''''''''_f'''''''''_Bool_t  \memOut_CTf'''''''''_f'''''''''_Bool_rbuf_d ;
  logic \memOut_CTf'''''''''_f'''''''''_Bool_rbuf_r ;
  \Word16#_t  \destructReadIn_CTf'''''''''_f'''''''''_Bool_d ;
  logic \destructReadIn_CTf'''''''''_f'''''''''_Bool_r ;
  \MemIn_CTf'''''''''_f'''''''''_Bool_t  \dconReadIn_CTf'''''''''_f'''''''''_Bool_d ;
  logic \dconReadIn_CTf'''''''''_f'''''''''_Bool_r ;
  \CTf'''''''''_f'''''''''_Bool_t  \readPointer_CTf'''''''''_f'''''''''_Boolscfarg_0_2_1_argbuf_d ;
  logic \readPointer_CTf'''''''''_f'''''''''_Boolscfarg_0_2_1_argbuf_r ;
  C5_t \writeMerge_choice_CTf'''''''''_f'''''''''_Bool_d ;
  logic \writeMerge_choice_CTf'''''''''_f'''''''''_Bool_r ;
  \CTf'''''''''_f'''''''''_Bool_t  \writeMerge_data_CTf'''''''''_f'''''''''_Bool_d ;
  logic \writeMerge_data_CTf'''''''''_f'''''''''_Bool_r ;
  \Pointer_CTf'''''''''_f'''''''''_Bool_t  \writeCTf'''''''''_f'''''''''_BoollizzieLet37_1_argbuf_d ;
  logic \writeCTf'''''''''_f'''''''''_BoollizzieLet37_1_argbuf_r ;
  \Pointer_CTf'''''''''_f'''''''''_Bool_t  \writeCTf'''''''''_f'''''''''_BoollizzieLet41_1_argbuf_d ;
  logic \writeCTf'''''''''_f'''''''''_BoollizzieLet41_1_argbuf_r ;
  \Pointer_CTf'''''''''_f'''''''''_Bool_t  \writeCTf'''''''''_f'''''''''_BoollizzieLet54_1_argbuf_d ;
  logic \writeCTf'''''''''_f'''''''''_BoollizzieLet54_1_argbuf_r ;
  \Pointer_CTf'''''''''_f'''''''''_Bool_t  \writeCTf'''''''''_f'''''''''_BoollizzieLet55_1_argbuf_d ;
  logic \writeCTf'''''''''_f'''''''''_BoollizzieLet55_1_argbuf_r ;
  \Pointer_CTf'''''''''_f'''''''''_Bool_t  \writeCTf'''''''''_f'''''''''_BoollizzieLet56_1_argbuf_d ;
  logic \writeCTf'''''''''_f'''''''''_BoollizzieLet56_1_argbuf_r ;
  \MemIn_CTf'''''''''_f'''''''''_Bool_t  \dconWriteIn_CTf'''''''''_f'''''''''_Bool_d ;
  logic \dconWriteIn_CTf'''''''''_f'''''''''_Bool_r ;
  \Pointer_CTf'''''''''_f'''''''''_Bool_t  \dconPtr_CTf'''''''''_f'''''''''_Bool_d ;
  logic \dconPtr_CTf'''''''''_f'''''''''_Bool_r ;
  \Pointer_CTf'''''''''_f'''''''''_Bool_t  _127_d;
  logic _127_r;
  assign _127_r = 1'd1;
  \Pointer_CTf'''''''''_f'''''''''_Bool_t  \demuxWriteResult_CTf'''''''''_f'''''''''_Bool_d ;
  logic \demuxWriteResult_CTf'''''''''_f'''''''''_Bool_r ;
  \Word16#_t  initHP_MaskQTree_d;
  logic initHP_MaskQTree_r;
  \Word16#_t  incrHP_MaskQTree_d;
  logic incrHP_MaskQTree_r;
  Go_t incrHP_mergeMaskQTree_d;
  logic incrHP_mergeMaskQTree_r;
  Go_t incrHP_MaskQTree1_d;
  logic incrHP_MaskQTree1_r;
  Go_t incrHP_MaskQTree2_d;
  logic incrHP_MaskQTree2_r;
  \Word16#_t  addHP_MaskQTree_d;
  logic addHP_MaskQTree_r;
  \Word16#_t  mergeHP_MaskQTree_d;
  logic mergeHP_MaskQTree_r;
  Go_t incrHP_mergeMaskQTree_buf_d;
  logic incrHP_mergeMaskQTree_buf_r;
  \Word16#_t  mergeHP_MaskQTree_buf_d;
  logic mergeHP_MaskQTree_buf_r;
  Go_t go_1_dummy_write_MaskQTree_d;
  logic go_1_dummy_write_MaskQTree_r;
  Go_t go_2_dummy_write_MaskQTree_d;
  logic go_2_dummy_write_MaskQTree_r;
  \Word16#_t  forkHP1_MaskQTree_d;
  logic forkHP1_MaskQTree_r;
  \Word16#_t  forkHP1_MaskQTree_snk_d;
  logic forkHP1_MaskQTree_snk_r;
  \Word16#_t  forkHP1_MaskQTre3_d;
  logic forkHP1_MaskQTre3_r;
  \Word16#_t  forkHP1_MaskQTre4_d;
  logic forkHP1_MaskQTre4_r;
  C2_t memMergeChoice_MaskQTree_d;
  logic memMergeChoice_MaskQTree_r;
  MemIn_MaskQTree_t memMergeIn_MaskQTree_d;
  logic memMergeIn_MaskQTree_r;
  MemOut_MaskQTree_t memOut_MaskQTree_d;
  logic memOut_MaskQTree_r;
  MemOut_MaskQTree_t memReadOut_MaskQTree_d;
  logic memReadOut_MaskQTree_r;
  MemOut_MaskQTree_t memWriteOut_MaskQTree_d;
  logic memWriteOut_MaskQTree_r;
  MemIn_MaskQTree_t memMergeIn_MaskQTree_dbuf_d;
  logic memMergeIn_MaskQTree_dbuf_r;
  MemIn_MaskQTree_t memMergeIn_MaskQTree_rbuf_d;
  logic memMergeIn_MaskQTree_rbuf_r;
  MemOut_MaskQTree_t memOut_MaskQTree_dbuf_d;
  logic memOut_MaskQTree_dbuf_r;
  MemOut_MaskQTree_t memOut_MaskQTree_rbuf_d;
  logic memOut_MaskQTree_rbuf_r;
  C2_t readMerge_choice_MaskQTree_d;
  logic readMerge_choice_MaskQTree_r;
  Pointer_MaskQTree_t readMerge_data_MaskQTree_d;
  logic readMerge_data_MaskQTree_r;
  MaskQTree_t readPointer_MaskQTreem1a85_1_argbuf_d;
  logic readPointer_MaskQTreem1a85_1_argbuf_r;
  MaskQTree_t readPointer_MaskQTreeq4a8w_1_argbuf_d;
  logic readPointer_MaskQTreeq4a8w_1_argbuf_r;
  \Word16#_t  destructReadIn_MaskQTree_d;
  logic destructReadIn_MaskQTree_r;
  MemIn_MaskQTree_t dconReadIn_MaskQTree_d;
  logic dconReadIn_MaskQTree_r;
  MaskQTree_t destructReadOut_MaskQTree_d;
  logic destructReadOut_MaskQTree_r;
  MemIn_MaskQTree_t dconWriteIn_MaskQTree_d;
  logic dconWriteIn_MaskQTree_r;
  Pointer_MaskQTree_t dconPtr_MaskQTree_d;
  logic dconPtr_MaskQTree_r;
  Pointer_MaskQTree_t _126_d;
  logic _126_r;
  assign _126_r = 1'd1;
  Pointer_MaskQTree_t dummy_write_MaskQTree_sink_d;
  logic dummy_write_MaskQTree_sink_r;
  Go_t go_1_argbuf_d;
  logic go_1_argbuf_r;
  Go_t \call_f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_CTf'''''''''_f'''''''''_Boolgo_4_d ;
  logic \call_f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_CTf'''''''''_f'''''''''_Boolgo_4_r ;
  Pointer_MaskQTree_t \call_f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_CTf'''''''''_f'''''''''_Boolq4a8w_d ;
  logic \call_f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_CTf'''''''''_f'''''''''_Boolq4a8w_r ;
  Pointer_QTree_Bool_t \call_f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_CTf'''''''''_f'''''''''_Boolq4'a8x_d ;
  logic \call_f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_CTf'''''''''_f'''''''''_Boolq4'a8x_r ;
  \Pointer_CTf'''''''''_f'''''''''_Bool_t  \call_f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_CTf'''''''''_f'''''''''_Boolsc_0_2_d ;
  logic \call_f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_CTf'''''''''_f'''''''''_Boolsc_0_2_r ;
  Go_t \call_f'''''''''_f'''''''''_Bool_initBufi_d ;
  logic \call_f'''''''''_f'''''''''_Bool_initBufi_r ;
  C5_t go_4_goMux_choice_d;
  logic go_4_goMux_choice_r;
  Go_t go_4_goMux_data_d;
  logic go_4_goMux_data_r;
  Go_t \call_f'''''''''_f'''''''''_Bool_unlockFork1_d ;
  logic \call_f'''''''''_f'''''''''_Bool_unlockFork1_r ;
  Go_t \call_f'''''''''_f'''''''''_Bool_unlockFork2_d ;
  logic \call_f'''''''''_f'''''''''_Bool_unlockFork2_r ;
  Go_t \call_f'''''''''_f'''''''''_Bool_unlockFork3_d ;
  logic \call_f'''''''''_f'''''''''_Bool_unlockFork3_r ;
  Go_t \call_f'''''''''_f'''''''''_Bool_unlockFork4_d ;
  logic \call_f'''''''''_f'''''''''_Bool_unlockFork4_r ;
  Go_t \call_f'''''''''_f'''''''''_Bool_initBuf_d ;
  logic \call_f'''''''''_f'''''''''_Bool_initBuf_r ;
  Go_t \call_f'''''''''_f'''''''''_Bool_goMux1_d ;
  logic \call_f'''''''''_f'''''''''_Bool_goMux1_r ;
  Pointer_MaskQTree_t \call_f'''''''''_f'''''''''_Bool_goMux2_d ;
  logic \call_f'''''''''_f'''''''''_Bool_goMux2_r ;
  Pointer_QTree_Bool_t \call_f'''''''''_f'''''''''_Bool_goMux3_d ;
  logic \call_f'''''''''_f'''''''''_Bool_goMux3_r ;
  \Pointer_CTf'''''''''_f'''''''''_Bool_t  \call_f'''''''''_f'''''''''_Bool_goMux4_d ;
  logic \call_f'''''''''_f'''''''''_Bool_goMux4_r ;
  Go_t \call_f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf'go_3_d ;
  logic \call_f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf'go_3_r ;
  Pointer_QTree_Bool_t \call_f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf'm2a8H_d ;
  logic \call_f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf'm2a8H_r ;
  Pointer_QTree_Bool_t \call_f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf'm3a8I_d ;
  logic \call_f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf'm3a8I_r ;
  \Pointer_CTf'_t  \call_f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf'sc_0_1_d ;
  logic \call_f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf'sc_0_1_r ;
  Go_t \call_f'_initBufi_d ;
  logic \call_f'_initBufi_r ;
  C5_t go_3_goMux_choice_d;
  logic go_3_goMux_choice_r;
  Go_t go_3_goMux_data_d;
  logic go_3_goMux_data_r;
  Go_t \call_f'_unlockFork1_d ;
  logic \call_f'_unlockFork1_r ;
  Go_t \call_f'_unlockFork2_d ;
  logic \call_f'_unlockFork2_r ;
  Go_t \call_f'_unlockFork3_d ;
  logic \call_f'_unlockFork3_r ;
  Go_t \call_f'_unlockFork4_d ;
  logic \call_f'_unlockFork4_r ;
  Go_t \call_f'_initBuf_d ;
  logic \call_f'_initBuf_r ;
  Go_t \call_f'_goMux1_d ;
  logic \call_f'_goMux1_r ;
  Pointer_QTree_Bool_t \call_f'_goMux2_d ;
  logic \call_f'_goMux2_r ;
  Pointer_QTree_Bool_t \call_f'_goMux3_d ;
  logic \call_f'_goMux3_r ;
  \Pointer_CTf'_t  \call_f'_goMux4_d ;
  logic \call_f'_goMux4_r ;
  Go_t call_fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfgo_2_d;
  logic call_fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfgo_2_r;
  Pointer_MaskQTree_t call_fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfm1a85_d;
  logic call_fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfm1a85_r;
  Pointer_QTree_Bool_t call_fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfm2a86_d;
  logic call_fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfm2a86_r;
  Pointer_QTree_Bool_t call_fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfm3a87_d;
  logic call_fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfm3a87_r;
  Pointer_CTf_t call_fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfsc_0_d;
  logic call_fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfsc_0_r;
  Go_t call_f_initBufi_d;
  logic call_f_initBufi_r;
  C5_t go_2_goMux_choice_d;
  logic go_2_goMux_choice_r;
  Go_t go_2_goMux_data_d;
  logic go_2_goMux_data_r;
  Go_t call_f_unlockFork1_d;
  logic call_f_unlockFork1_r;
  Go_t call_f_unlockFork2_d;
  logic call_f_unlockFork2_r;
  Go_t call_f_unlockFork3_d;
  logic call_f_unlockFork3_r;
  Go_t call_f_unlockFork4_d;
  logic call_f_unlockFork4_r;
  Go_t call_f_unlockFork5_d;
  logic call_f_unlockFork5_r;
  Go_t call_f_initBuf_d;
  logic call_f_initBuf_r;
  Go_t call_f_goMux1_d;
  logic call_f_goMux1_r;
  Pointer_MaskQTree_t call_f_goMux2_d;
  logic call_f_goMux2_r;
  Pointer_QTree_Bool_t call_f_goMux3_d;
  logic call_f_goMux3_r;
  Pointer_QTree_Bool_t call_f_goMux4_d;
  logic call_f_goMux4_r;
  Pointer_CTf_t call_f_goMux5_d;
  logic call_f_goMux5_r;
  QTree_Bool_t lizzieLet6_1_argbuf_d;
  logic lizzieLet6_1_argbuf_r;
  QTree_Bool_t lizzieLet15_1_1_argbuf_d;
  logic lizzieLet15_1_1_argbuf_r;
  C8_t \f'''''''''_f'''''''''_Bool_choice_d ;
  logic \f'''''''''_f'''''''''_Bool_choice_r ;
  TupGo___Pointer_MaskQTree___Pointer_QTree_Bool_t \f'''''''''_f'''''''''_Bool_data_d ;
  logic \f'''''''''_f'''''''''_Bool_data_r ;
  Go_t go_7_1_d;
  logic go_7_1_r;
  Go_t go_7_2_d;
  logic go_7_2_r;
  Pointer_QTree_Bool_t \q4'a8x_1_1_argbuf_d ;
  logic \q4'a8x_1_1_argbuf_r ;
  Pointer_MaskQTree_t q4a8w_1_1_argbuf_d;
  logic q4a8w_1_1_argbuf_r;
  Pointer_QTree_Bool_t \f'''''''''_f'''''''''_Bool_resbuf_d ;
  logic \f'''''''''_f'''''''''_Bool_resbuf_r ;
  Pointer_QTree_Bool_t \f'''''''''_f'''''''''_Bool_2_argbuf_d ;
  logic \f'''''''''_f'''''''''_Bool_2_argbuf_r ;
  Pointer_QTree_Bool_t \f'''''''''_f'''''''''_Bool_3_argbuf_d ;
  logic \f'''''''''_f'''''''''_Bool_3_argbuf_r ;
  Pointer_QTree_Bool_t \f'''''''''_f'''''''''_Bool_4_argbuf_d ;
  logic \f'''''''''_f'''''''''_Bool_4_argbuf_r ;
  QTree_Bool_t es_0_1es_1_1es_2_1es_3_1QNode_Bool_d;
  logic es_0_1es_1_1es_2_1es_3_1QNode_Bool_r;
  Pointer_QTree_Bool_t \f'''''''''_f'''''''''_Bool_5_argbuf_d ;
  logic \f'''''''''_f'''''''''_Bool_5_argbuf_r ;
  Pointer_QTree_Bool_t \f'''''''''_f'''''''''_Bool_6_argbuf_d ;
  logic \f'''''''''_f'''''''''_Bool_6_argbuf_r ;
  Pointer_QTree_Bool_t \f'''''''''_f'''''''''_Bool_7_argbuf_d ;
  logic \f'''''''''_f'''''''''_Bool_7_argbuf_r ;
  Pointer_QTree_Bool_t \f'''''''''_f'''''''''_Bool_8_argbuf_d ;
  logic \f'''''''''_f'''''''''_Bool_8_argbuf_r ;
  QTree_Bool_t es_4_1es_5_1es_6_1es_7_1QNode_Bool_d;
  logic es_4_1es_5_1es_6_1es_7_1QNode_Bool_r;
  Pointer_QTree_Bool_t \f'''''''''_f'''''''''_Bool_1_d ;
  logic \f'''''''''_f'''''''''_Bool_1_r ;
  Pointer_QTree_Bool_t \f'''''''''_f'''''''''_Bool_2_d ;
  logic \f'''''''''_f'''''''''_Bool_2_r ;
  Pointer_QTree_Bool_t \f'''''''''_f'''''''''_Bool_3_d ;
  logic \f'''''''''_f'''''''''_Bool_3_r ;
  Pointer_QTree_Bool_t \f'''''''''_f'''''''''_Bool_4_d ;
  logic \f'''''''''_f'''''''''_Bool_4_r ;
  Pointer_QTree_Bool_t \f'''''''''_f'''''''''_Bool_5_d ;
  logic \f'''''''''_f'''''''''_Bool_5_r ;
  Pointer_QTree_Bool_t \f'''''''''_f'''''''''_Bool_6_d ;
  logic \f'''''''''_f'''''''''_Bool_6_r ;
  Pointer_QTree_Bool_t \f'''''''''_f'''''''''_Bool_7_d ;
  logic \f'''''''''_f'''''''''_Bool_7_r ;
  Pointer_QTree_Bool_t \f'''''''''_f'''''''''_Bool_8_d ;
  logic \f'''''''''_f'''''''''_Bool_8_r ;
  Go_t \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Boolgo_7_d ;
  logic \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Boolgo_7_r ;
  Pointer_MaskQTree_t \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Boolq4a8w_1_d ;
  logic \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Boolq4a8w_1_r ;
  Pointer_QTree_Bool_t \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Boolq4'a8x_1_d ;
  logic \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Boolq4'a8x_1_r ;
  Go_t \f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolgo_6_d ;
  logic \f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolgo_6_r ;
  Pointer_QTree_Bool_t \f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolm2a8H_1_d ;
  logic \f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolm2a8H_1_r ;
  Pointer_QTree_Bool_t \f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolm3a8I_1_d ;
  logic \f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolm3a8I_1_r ;
  Go_t go_6_1_d;
  logic go_6_1_r;
  Go_t go_6_2_d;
  logic go_6_2_r;
  Pointer_QTree_Bool_t m2a8H_1_1_argbuf_d;
  logic m2a8H_1_1_argbuf_r;
  Pointer_QTree_Bool_t m3a8I_1_1_argbuf_d;
  logic m3a8I_1_1_argbuf_r;
  Pointer_QTree_Bool_t lizzieLet14_1_argbuf_d;
  logic lizzieLet14_1_argbuf_r;
  Go_t fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Boolgo_5_d;
  logic fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Boolgo_5_r;
  Pointer_MaskQTree_t fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Boolm1a85_1_d;
  logic fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Boolm1a85_1_r;
  Pointer_QTree_Bool_t fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Boolm2a86_1_d;
  logic fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Boolm2a86_1_r;
  Pointer_QTree_Bool_t fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Boolm3a87_1_d;
  logic fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Boolm3a87_1_r;
  Go_t go_5_1_d;
  logic go_5_1_r;
  Go_t go_5_2_d;
  logic go_5_2_r;
  Pointer_MaskQTree_t m1a85_1_1_argbuf_d;
  logic m1a85_1_1_argbuf_r;
  Pointer_QTree_Bool_t m2a86_1_1_argbuf_d;
  logic m2a86_1_1_argbuf_r;
  Pointer_QTree_Bool_t m3a87_1_1_argbuf_d;
  logic m3a87_1_1_argbuf_r;
  C12_t go_10_goMux_choice_1_d;
  logic go_10_goMux_choice_1_r;
  C12_t go_10_goMux_choice_2_d;
  logic go_10_goMux_choice_2_r;
  Pointer_QTree_Bool_t srtarg_0_1_goMux_mux_d;
  logic srtarg_0_1_goMux_mux_r;
  \Pointer_CTf'_t  scfarg_0_1_goMux_mux_d;
  logic scfarg_0_1_goMux_mux_r;
  C6_t go_11_goMux_choice_1_d;
  logic go_11_goMux_choice_1_r;
  C6_t go_11_goMux_choice_2_d;
  logic go_11_goMux_choice_2_r;
  Pointer_QTree_Bool_t srtarg_0_2_goMux_mux_d;
  logic srtarg_0_2_goMux_mux_r;
  \Pointer_CTf'''''''''_f'''''''''_Bool_t  scfarg_0_2_goMux_mux_d;
  logic scfarg_0_2_goMux_mux_r;
  TupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool_t fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool_1_d;
  logic fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool_1_r;
  C5_t go_2_goMux_choice_1_d;
  logic go_2_goMux_choice_1_r;
  C5_t go_2_goMux_choice_2_d;
  logic go_2_goMux_choice_2_r;
  C5_t go_2_goMux_choice_3_d;
  logic go_2_goMux_choice_3_r;
  C5_t go_2_goMux_choice_4_d;
  logic go_2_goMux_choice_4_r;
  Pointer_MaskQTree_t m1a85_goMux_mux_d;
  logic m1a85_goMux_mux_r;
  Pointer_QTree_Bool_t m2a86_goMux_mux_d;
  logic m2a86_goMux_mux_r;
  Pointer_QTree_Bool_t m3a87_goMux_mux_d;
  logic m3a87_goMux_mux_r;
  Pointer_CTf_t sc_0_goMux_mux_d;
  logic sc_0_goMux_mux_r;
  C5_t go_3_goMux_choice_1_d;
  logic go_3_goMux_choice_1_r;
  C5_t go_3_goMux_choice_2_d;
  logic go_3_goMux_choice_2_r;
  C5_t go_3_goMux_choice_3_d;
  logic go_3_goMux_choice_3_r;
  Pointer_QTree_Bool_t m2a8H_goMux_mux_d;
  logic m2a8H_goMux_mux_r;
  Pointer_QTree_Bool_t m3a8I_goMux_mux_d;
  logic m3a8I_goMux_mux_r;
  \Pointer_CTf'_t  sc_0_1_goMux_mux_d;
  logic sc_0_1_goMux_mux_r;
  C5_t go_4_goMux_choice_1_d;
  logic go_4_goMux_choice_1_r;
  C5_t go_4_goMux_choice_2_d;
  logic go_4_goMux_choice_2_r;
  C5_t go_4_goMux_choice_3_d;
  logic go_4_goMux_choice_3_r;
  Pointer_MaskQTree_t q4a8w_goMux_mux_d;
  logic q4a8w_goMux_mux_r;
  Pointer_QTree_Bool_t \q4'a8x_goMux_mux_d ;
  logic \q4'a8x_goMux_mux_r ;
  \Pointer_CTf'''''''''_f'''''''''_Bool_t  sc_0_2_goMux_mux_d;
  logic sc_0_2_goMux_mux_r;
  CTf_t go_5_1Lfsbos_d;
  logic go_5_1Lfsbos_r;
  CTf_t lizzieLet39_1_argbuf_d;
  logic lizzieLet39_1_argbuf_r;
  Go_t go_5_2_argbuf_d;
  logic go_5_2_argbuf_r;
  TupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf_t call_fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf_1_d;
  logic call_fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf_1_r;
  \CTf'_t  \go_6_1Lf'sbos_d ;
  logic \go_6_1Lf'sbos_r ;
  \CTf'_t  lizzieLet40_1_argbuf_d;
  logic lizzieLet40_1_argbuf_r;
  Go_t go_6_2_argbuf_d;
  logic go_6_2_argbuf_r;
  \TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf'_t  \call_f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf'_1_d ;
  logic \call_f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf'_1_r ;
  \CTf'''''''''_f'''''''''_Bool_t  \go_7_1Lf'''''''''_f'''''''''_Boolsbos_d ;
  logic \go_7_1Lf'''''''''_f'''''''''_Boolsbos_r ;
  \CTf'''''''''_f'''''''''_Bool_t  lizzieLet41_1_argbuf_d;
  logic lizzieLet41_1_argbuf_r;
  Go_t go_7_2_argbuf_d;
  logic go_7_2_argbuf_r;
  \TupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_CTf'''''''''_f'''''''''_Bool_t  \call_f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_CTf'''''''''_f'''''''''_Bool_1_d ;
  logic \call_f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_CTf'''''''''_f'''''''''_Bool_1_r ;
  QTree_Bool_t lizzieLet0_1_1QVal_Bool_d;
  logic lizzieLet0_1_1QVal_Bool_r;
  C17_t go_9_goMux_choice_1_d;
  logic go_9_goMux_choice_1_r;
  C17_t go_9_goMux_choice_2_d;
  logic go_9_goMux_choice_2_r;
  Pointer_QTree_Bool_t srtarg_0_goMux_mux_d;
  logic srtarg_0_goMux_mux_r;
  Pointer_CTf_t scfarg_0_goMux_mux_d;
  logic scfarg_0_goMux_mux_r;
  Pointer_MaskQTree_t q1a88_destruct_d;
  logic q1a88_destruct_r;
  Pointer_MaskQTree_t q2a89_destruct_d;
  logic q2a89_destruct_r;
  Pointer_MaskQTree_t q3a8a_destruct_d;
  logic q3a8a_destruct_r;
  Pointer_MaskQTree_t q4a8b_destruct_d;
  logic q4a8b_destruct_r;
  QTree_Bool_t lizzieLet42_1_argbuf_d;
  logic lizzieLet42_1_argbuf_r;
  MaskQTree_t _125_d;
  logic _125_r;
  assign _125_r = 1'd1;
  MaskQTree_t _124_d;
  logic _124_r;
  assign _124_r = 1'd1;
  MaskQTree_t lizzieLet0_1MQNode_d;
  logic lizzieLet0_1MQNode_r;
  Go_t lizzieLet0_3MQNone_d;
  logic lizzieLet0_3MQNone_r;
  Go_t lizzieLet0_3MQVal_d;
  logic lizzieLet0_3MQVal_r;
  Go_t lizzieLet0_3MQNode_d;
  logic lizzieLet0_3MQNode_r;
  Go_t lizzieLet0_3MQNone_1_d;
  logic lizzieLet0_3MQNone_1_r;
  Go_t lizzieLet0_3MQNone_2_d;
  logic lizzieLet0_3MQNone_2_r;
  QTree_Bool_t lizzieLet0_3MQNone_1QNone_Bool_d;
  logic lizzieLet0_3MQNone_1QNone_Bool_r;
  QTree_Bool_t lizzieLet1_1_argbuf_d;
  logic lizzieLet1_1_argbuf_r;
  Go_t lizzieLet0_3MQNone_2_argbuf_d;
  logic lizzieLet0_3MQNone_2_argbuf_r;
  C17_t go_9_goMux_choice_d;
  logic go_9_goMux_choice_r;
  Go_t go_9_goMux_data_d;
  logic go_9_goMux_data_r;
  Go_t lizzieLet0_3MQVal_1_d;
  logic lizzieLet0_3MQVal_1_r;
  Go_t lizzieLet0_3MQVal_2_d;
  logic lizzieLet0_3MQVal_2_r;
  Go_t lizzieLet0_3MQVal_1_argbuf_d;
  logic lizzieLet0_3MQVal_1_argbuf_r;
  TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_t \f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_1_d ;
  logic \f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_1_r ;
  Go_t lizzieLet0_3MQVal_2_argbuf_d;
  logic lizzieLet0_3MQVal_2_argbuf_r;
  QTree_Bool_t _123_d;
  logic _123_r;
  assign _123_r = 1'd1;
  QTree_Bool_t _122_d;
  logic _122_r;
  assign _122_r = 1'd1;
  QTree_Bool_t lizzieLet0_4MQNode_d;
  logic lizzieLet0_4MQNode_r;
  QTree_Bool_t lizzieLet0_4MQNode_1_d;
  logic lizzieLet0_4MQNode_1_r;
  QTree_Bool_t lizzieLet0_4MQNode_2_d;
  logic lizzieLet0_4MQNode_2_r;
  QTree_Bool_t lizzieLet0_4MQNode_3_d;
  logic lizzieLet0_4MQNode_3_r;
  QTree_Bool_t lizzieLet0_4MQNode_4_d;
  logic lizzieLet0_4MQNode_4_r;
  QTree_Bool_t lizzieLet0_4MQNode_5_d;
  logic lizzieLet0_4MQNode_5_r;
  QTree_Bool_t lizzieLet0_4MQNode_6_d;
  logic lizzieLet0_4MQNode_6_r;
  QTree_Bool_t lizzieLet0_4MQNode_7_d;
  logic lizzieLet0_4MQNode_7_r;
  QTree_Bool_t lizzieLet0_4MQNode_8_d;
  logic lizzieLet0_4MQNode_8_r;
  QTree_Bool_t lizzieLet0_4MQNode_9_d;
  logic lizzieLet0_4MQNode_9_r;
  Pointer_QTree_Bool_t \q1'a8n_destruct_d ;
  logic \q1'a8n_destruct_r ;
  Pointer_QTree_Bool_t \q2'a8o_destruct_d ;
  logic \q2'a8o_destruct_r ;
  Pointer_QTree_Bool_t \q3'a8p_destruct_d ;
  logic \q3'a8p_destruct_r ;
  Pointer_QTree_Bool_t \q4'a8q_destruct_d ;
  logic \q4'a8q_destruct_r ;
  MyBool_t v1a8h_destruct_d;
  logic v1a8h_destruct_r;
  QTree_Bool_t _121_d;
  logic _121_r;
  assign _121_r = 1'd1;
  QTree_Bool_t lizzieLet0_4MQNode_1QVal_Bool_d;
  logic lizzieLet0_4MQNode_1QVal_Bool_r;
  QTree_Bool_t lizzieLet0_4MQNode_1QNode_Bool_d;
  logic lizzieLet0_4MQNode_1QNode_Bool_r;
  QTree_Bool_t _120_d;
  logic _120_r;
  assign _120_r = 1'd1;
  Go_t lizzieLet0_4MQNode_3QNone_Bool_d;
  logic lizzieLet0_4MQNode_3QNone_Bool_r;
  Go_t lizzieLet0_4MQNode_3QVal_Bool_d;
  logic lizzieLet0_4MQNode_3QVal_Bool_r;
  Go_t lizzieLet0_4MQNode_3QNode_Bool_d;
  logic lizzieLet0_4MQNode_3QNode_Bool_r;
  Go_t lizzieLet0_4MQNode_3QError_Bool_d;
  logic lizzieLet0_4MQNode_3QError_Bool_r;
  Go_t lizzieLet0_4MQNode_3QError_Bool_1_d;
  logic lizzieLet0_4MQNode_3QError_Bool_1_r;
  Go_t lizzieLet0_4MQNode_3QError_Bool_2_d;
  logic lizzieLet0_4MQNode_3QError_Bool_2_r;
  QTree_Bool_t lizzieLet0_4MQNode_3QError_Bool_1QError_Bool_d;
  logic lizzieLet0_4MQNode_3QError_Bool_1QError_Bool_r;
  QTree_Bool_t lizzieLet19_2_1_argbuf_d;
  logic lizzieLet19_2_1_argbuf_r;
  Go_t lizzieLet0_4MQNode_3QError_Bool_2_argbuf_d;
  logic lizzieLet0_4MQNode_3QError_Bool_2_argbuf_r;
  QTree_Bool_t lizzieLet0_4MQNode_4QNone_Bool_d;
  logic lizzieLet0_4MQNode_4QNone_Bool_r;
  QTree_Bool_t lizzieLet0_4MQNode_4QVal_Bool_d;
  logic lizzieLet0_4MQNode_4QVal_Bool_r;
  QTree_Bool_t lizzieLet0_4MQNode_4QNode_Bool_d;
  logic lizzieLet0_4MQNode_4QNode_Bool_r;
  QTree_Bool_t _119_d;
  logic _119_r;
  assign _119_r = 1'd1;
  QTree_Bool_t lizzieLet0_4MQNode_4QNode_Bool_1_d;
  logic lizzieLet0_4MQNode_4QNode_Bool_1_r;
  QTree_Bool_t lizzieLet0_4MQNode_4QNode_Bool_2_d;
  logic lizzieLet0_4MQNode_4QNode_Bool_2_r;
  QTree_Bool_t lizzieLet0_4MQNode_4QNode_Bool_3_d;
  logic lizzieLet0_4MQNode_4QNode_Bool_3_r;
  QTree_Bool_t lizzieLet0_4MQNode_4QNode_Bool_4_d;
  logic lizzieLet0_4MQNode_4QNode_Bool_4_r;
  QTree_Bool_t lizzieLet0_4MQNode_4QNode_Bool_5_d;
  logic lizzieLet0_4MQNode_4QNode_Bool_5_r;
  QTree_Bool_t lizzieLet0_4MQNode_4QNode_Bool_6_d;
  logic lizzieLet0_4MQNode_4QNode_Bool_6_r;
  QTree_Bool_t lizzieLet0_4MQNode_4QNode_Bool_7_d;
  logic lizzieLet0_4MQNode_4QNode_Bool_7_r;
  QTree_Bool_t lizzieLet0_4MQNode_4QNode_Bool_8_d;
  logic lizzieLet0_4MQNode_4QNode_Bool_8_r;
  QTree_Bool_t lizzieLet0_4MQNode_4QNode_Bool_9_d;
  logic lizzieLet0_4MQNode_4QNode_Bool_9_r;
  QTree_Bool_t lizzieLet0_4MQNode_4QNode_Bool_10_d;
  logic lizzieLet0_4MQNode_4QNode_Bool_10_r;
  QTree_Bool_t lizzieLet0_4MQNode_4QNode_Bool_11_d;
  logic lizzieLet0_4MQNode_4QNode_Bool_11_r;
  QTree_Bool_t lizzieLet0_4MQNode_4QNode_Bool_12_d;
  logic lizzieLet0_4MQNode_4QNode_Bool_12_r;
  Pointer_QTree_Bool_t lizzieLet0_4MQNode_4QNode_Bool_10QNone_Bool_d;
  logic lizzieLet0_4MQNode_4QNode_Bool_10QNone_Bool_r;
  Pointer_QTree_Bool_t _118_d;
  logic _118_r;
  assign _118_r = 1'd1;
  Pointer_QTree_Bool_t lizzieLet0_4MQNode_4QNode_Bool_10QNode_Bool_d;
  logic lizzieLet0_4MQNode_4QNode_Bool_10QNode_Bool_r;
  Pointer_QTree_Bool_t _117_d;
  logic _117_r;
  assign _117_r = 1'd1;
  Pointer_QTree_Bool_t lizzieLet0_4MQNode_4QNode_Bool_10QNone_Bool_1_argbuf_d;
  logic lizzieLet0_4MQNode_4QNode_Bool_10QNone_Bool_1_argbuf_r;
  Pointer_QTree_Bool_t lizzieLet0_4MQNode_4QNode_Bool_11QNone_Bool_d;
  logic lizzieLet0_4MQNode_4QNode_Bool_11QNone_Bool_r;
  Pointer_QTree_Bool_t _116_d;
  logic _116_r;
  assign _116_r = 1'd1;
  Pointer_QTree_Bool_t lizzieLet0_4MQNode_4QNode_Bool_11QNode_Bool_d;
  logic lizzieLet0_4MQNode_4QNode_Bool_11QNode_Bool_r;
  Pointer_QTree_Bool_t _115_d;
  logic _115_r;
  assign _115_r = 1'd1;
  Pointer_QTree_Bool_t lizzieLet0_4MQNode_4QNode_Bool_11QNone_Bool_1_argbuf_d;
  logic lizzieLet0_4MQNode_4QNode_Bool_11QNone_Bool_1_argbuf_r;
  Pointer_QTree_Bool_t lizzieLet0_4MQNode_4QNode_Bool_12QNone_Bool_d;
  logic lizzieLet0_4MQNode_4QNode_Bool_12QNone_Bool_r;
  Pointer_QTree_Bool_t _114_d;
  logic _114_r;
  assign _114_r = 1'd1;
  Pointer_QTree_Bool_t lizzieLet0_4MQNode_4QNode_Bool_12QNode_Bool_d;
  logic lizzieLet0_4MQNode_4QNode_Bool_12QNode_Bool_r;
  Pointer_QTree_Bool_t _113_d;
  logic _113_r;
  assign _113_r = 1'd1;
  Pointer_QTree_Bool_t lizzieLet0_4MQNode_4QNode_Bool_12QNode_Bool_1_argbuf_d;
  logic lizzieLet0_4MQNode_4QNode_Bool_12QNode_Bool_1_argbuf_r;
  Pointer_QTree_Bool_t lizzieLet0_4MQNode_4QNode_Bool_12QNone_Bool_1_argbuf_d;
  logic lizzieLet0_4MQNode_4QNode_Bool_12QNone_Bool_1_argbuf_r;
  Pointer_QTree_Bool_t t1a8s_destruct_d;
  logic t1a8s_destruct_r;
  Pointer_QTree_Bool_t t2a8t_destruct_d;
  logic t2a8t_destruct_r;
  Pointer_QTree_Bool_t t3a8u_destruct_d;
  logic t3a8u_destruct_r;
  Pointer_QTree_Bool_t t4a8v_destruct_d;
  logic t4a8v_destruct_r;
  QTree_Bool_t _112_d;
  logic _112_r;
  assign _112_r = 1'd1;
  QTree_Bool_t _111_d;
  logic _111_r;
  assign _111_r = 1'd1;
  QTree_Bool_t lizzieLet0_4MQNode_4QNode_Bool_1QNode_Bool_d;
  logic lizzieLet0_4MQNode_4QNode_Bool_1QNode_Bool_r;
  QTree_Bool_t _110_d;
  logic _110_r;
  assign _110_r = 1'd1;
  Go_t lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_d;
  logic lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_r;
  Go_t lizzieLet0_4MQNode_4QNode_Bool_3QVal_Bool_d;
  logic lizzieLet0_4MQNode_4QNode_Bool_3QVal_Bool_r;
  Go_t lizzieLet0_4MQNode_4QNode_Bool_3QNode_Bool_d;
  logic lizzieLet0_4MQNode_4QNode_Bool_3QNode_Bool_r;
  Go_t lizzieLet0_4MQNode_4QNode_Bool_3QError_Bool_d;
  logic lizzieLet0_4MQNode_4QNode_Bool_3QError_Bool_r;
  Go_t lizzieLet0_4MQNode_4QNode_Bool_3QError_Bool_1_d;
  logic lizzieLet0_4MQNode_4QNode_Bool_3QError_Bool_1_r;
  Go_t lizzieLet0_4MQNode_4QNode_Bool_3QError_Bool_2_d;
  logic lizzieLet0_4MQNode_4QNode_Bool_3QError_Bool_2_r;
  QTree_Bool_t lizzieLet0_4MQNode_4QNode_Bool_3QError_Bool_1QError_Bool_d;
  logic lizzieLet0_4MQNode_4QNode_Bool_3QError_Bool_1QError_Bool_r;
  QTree_Bool_t lizzieLet18_1_1_argbuf_d;
  logic lizzieLet18_1_1_argbuf_r;
  Go_t lizzieLet0_4MQNode_4QNode_Bool_3QError_Bool_2_argbuf_d;
  logic lizzieLet0_4MQNode_4QNode_Bool_3QError_Bool_2_argbuf_r;
  Go_t lizzieLet0_4MQNode_4QNode_Bool_3QNode_Bool_1_argbuf_d;
  logic lizzieLet0_4MQNode_4QNode_Bool_3QNode_Bool_1_argbuf_r;
  Go_t lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_1_d;
  logic lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_1_r;
  Go_t lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_2_d;
  logic lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_2_r;
  Go_t lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_3_d;
  logic lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_3_r;
  Go_t lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_4_d;
  logic lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_4_r;
  Go_t lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_5_d;
  logic lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_5_r;
  Go_t lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_1_argbuf_d;
  logic lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_1_argbuf_r;
  TupGo___Pointer_MaskQTree___Pointer_QTree_Bool_t \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool5_d ;
  logic \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool5_r ;
  Go_t lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_2_argbuf_d;
  logic lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_2_argbuf_r;
  TupGo___Pointer_MaskQTree___Pointer_QTree_Bool_t \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool6_d ;
  logic \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool6_r ;
  Go_t lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_3_argbuf_d;
  logic lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_3_argbuf_r;
  TupGo___Pointer_MaskQTree___Pointer_QTree_Bool_t \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool7_d ;
  logic \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool7_r ;
  Go_t lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_4_argbuf_d;
  logic lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_4_argbuf_r;
  TupGo___Pointer_MaskQTree___Pointer_QTree_Bool_t \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool8_d ;
  logic \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool8_r ;
  Go_t lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_5_argbuf_d;
  logic lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_5_argbuf_r;
  Go_t lizzieLet0_4MQNode_4QNode_Bool_3QVal_Bool_1_d;
  logic lizzieLet0_4MQNode_4QNode_Bool_3QVal_Bool_1_r;
  Go_t lizzieLet0_4MQNode_4QNode_Bool_3QVal_Bool_2_d;
  logic lizzieLet0_4MQNode_4QNode_Bool_3QVal_Bool_2_r;
  QTree_Bool_t lizzieLet0_4MQNode_4QNode_Bool_3QVal_Bool_1QError_Bool_d;
  logic lizzieLet0_4MQNode_4QNode_Bool_3QVal_Bool_1QError_Bool_r;
  QTree_Bool_t lizzieLet16_1_1_argbuf_d;
  logic lizzieLet16_1_1_argbuf_r;
  Go_t lizzieLet0_4MQNode_4QNode_Bool_3QVal_Bool_2_argbuf_d;
  logic lizzieLet0_4MQNode_4QNode_Bool_3QVal_Bool_2_argbuf_r;
  Pointer_CTf_t lizzieLet0_4MQNode_4QNode_Bool_4QNone_Bool_d;
  logic lizzieLet0_4MQNode_4QNode_Bool_4QNone_Bool_r;
  Pointer_CTf_t lizzieLet0_4MQNode_4QNode_Bool_4QVal_Bool_d;
  logic lizzieLet0_4MQNode_4QNode_Bool_4QVal_Bool_r;
  Pointer_CTf_t lizzieLet0_4MQNode_4QNode_Bool_4QNode_Bool_d;
  logic lizzieLet0_4MQNode_4QNode_Bool_4QNode_Bool_r;
  Pointer_CTf_t lizzieLet0_4MQNode_4QNode_Bool_4QError_Bool_d;
  logic lizzieLet0_4MQNode_4QNode_Bool_4QError_Bool_r;
  Pointer_CTf_t lizzieLet0_4MQNode_4QNode_Bool_4QError_Bool_1_argbuf_d;
  logic lizzieLet0_4MQNode_4QNode_Bool_4QError_Bool_1_argbuf_r;
  CTf_t lizzieLet0_4MQNode_4QNode_Bool_4QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_5QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_9QNode_Bool_1t1a8s_1lizzieLet0_4MQNode_4QNode_Bool_6QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_10QNode_Bool_1t2a8t_1lizzieLet0_4MQNode_4QNode_Bool_7QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_11QNode_Bool_1t3a8u_1Lcall_f3_d;
  logic lizzieLet0_4MQNode_4QNode_Bool_4QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_5QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_9QNode_Bool_1t1a8s_1lizzieLet0_4MQNode_4QNode_Bool_6QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_10QNode_Bool_1t2a8t_1lizzieLet0_4MQNode_4QNode_Bool_7QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_11QNode_Bool_1t3a8u_1Lcall_f3_r;
  CTf_t lizzieLet17_1_1_argbuf_d;
  logic lizzieLet17_1_1_argbuf_r;
  Pointer_CTf_t lizzieLet0_4MQNode_4QNode_Bool_4QNone_Bool_1_argbuf_d;
  logic lizzieLet0_4MQNode_4QNode_Bool_4QNone_Bool_1_argbuf_r;
  Pointer_CTf_t lizzieLet0_4MQNode_4QNode_Bool_4QVal_Bool_1_argbuf_d;
  logic lizzieLet0_4MQNode_4QNode_Bool_4QVal_Bool_1_argbuf_r;
  Pointer_MaskQTree_t lizzieLet0_4MQNode_4QNode_Bool_5QNone_Bool_d;
  logic lizzieLet0_4MQNode_4QNode_Bool_5QNone_Bool_r;
  Pointer_MaskQTree_t _109_d;
  logic _109_r;
  assign _109_r = 1'd1;
  Pointer_MaskQTree_t lizzieLet0_4MQNode_4QNode_Bool_5QNode_Bool_d;
  logic lizzieLet0_4MQNode_4QNode_Bool_5QNode_Bool_r;
  Pointer_MaskQTree_t _108_d;
  logic _108_r;
  assign _108_r = 1'd1;
  Pointer_MaskQTree_t lizzieLet0_4MQNode_4QNode_Bool_5QNone_Bool_1_argbuf_d;
  logic lizzieLet0_4MQNode_4QNode_Bool_5QNone_Bool_1_argbuf_r;
  Pointer_MaskQTree_t lizzieLet0_4MQNode_4QNode_Bool_6QNone_Bool_d;
  logic lizzieLet0_4MQNode_4QNode_Bool_6QNone_Bool_r;
  Pointer_MaskQTree_t _107_d;
  logic _107_r;
  assign _107_r = 1'd1;
  Pointer_MaskQTree_t lizzieLet0_4MQNode_4QNode_Bool_6QNode_Bool_d;
  logic lizzieLet0_4MQNode_4QNode_Bool_6QNode_Bool_r;
  Pointer_MaskQTree_t _106_d;
  logic _106_r;
  assign _106_r = 1'd1;
  Pointer_MaskQTree_t lizzieLet0_4MQNode_4QNode_Bool_6QNone_Bool_1_argbuf_d;
  logic lizzieLet0_4MQNode_4QNode_Bool_6QNone_Bool_1_argbuf_r;
  Pointer_MaskQTree_t lizzieLet0_4MQNode_4QNode_Bool_7QNone_Bool_d;
  logic lizzieLet0_4MQNode_4QNode_Bool_7QNone_Bool_r;
  Pointer_MaskQTree_t _105_d;
  logic _105_r;
  assign _105_r = 1'd1;
  Pointer_MaskQTree_t lizzieLet0_4MQNode_4QNode_Bool_7QNode_Bool_d;
  logic lizzieLet0_4MQNode_4QNode_Bool_7QNode_Bool_r;
  Pointer_MaskQTree_t _104_d;
  logic _104_r;
  assign _104_r = 1'd1;
  Pointer_MaskQTree_t lizzieLet0_4MQNode_4QNode_Bool_7QNone_Bool_1_argbuf_d;
  logic lizzieLet0_4MQNode_4QNode_Bool_7QNone_Bool_1_argbuf_r;
  Pointer_MaskQTree_t lizzieLet0_4MQNode_4QNode_Bool_8QNone_Bool_d;
  logic lizzieLet0_4MQNode_4QNode_Bool_8QNone_Bool_r;
  Pointer_MaskQTree_t _103_d;
  logic _103_r;
  assign _103_r = 1'd1;
  Pointer_MaskQTree_t lizzieLet0_4MQNode_4QNode_Bool_8QNode_Bool_d;
  logic lizzieLet0_4MQNode_4QNode_Bool_8QNode_Bool_r;
  Pointer_MaskQTree_t _102_d;
  logic _102_r;
  assign _102_r = 1'd1;
  Pointer_MaskQTree_t lizzieLet0_4MQNode_4QNode_Bool_8QNode_Bool_1_argbuf_d;
  logic lizzieLet0_4MQNode_4QNode_Bool_8QNode_Bool_1_argbuf_r;
  Pointer_MaskQTree_t lizzieLet0_4MQNode_4QNode_Bool_8QNone_Bool_1_argbuf_d;
  logic lizzieLet0_4MQNode_4QNode_Bool_8QNone_Bool_1_argbuf_r;
  Pointer_QTree_Bool_t lizzieLet0_4MQNode_4QNode_Bool_9QNone_Bool_d;
  logic lizzieLet0_4MQNode_4QNode_Bool_9QNone_Bool_r;
  Pointer_QTree_Bool_t _101_d;
  logic _101_r;
  assign _101_r = 1'd1;
  Pointer_QTree_Bool_t lizzieLet0_4MQNode_4QNode_Bool_9QNode_Bool_d;
  logic lizzieLet0_4MQNode_4QNode_Bool_9QNode_Bool_r;
  Pointer_QTree_Bool_t _100_d;
  logic _100_r;
  assign _100_r = 1'd1;
  Pointer_QTree_Bool_t lizzieLet0_4MQNode_4QNode_Bool_9QNone_Bool_1_argbuf_d;
  logic lizzieLet0_4MQNode_4QNode_Bool_9QNone_Bool_1_argbuf_r;
  QTree_Bool_t lizzieLet0_4MQNode_4QNone_Bool_1_d;
  logic lizzieLet0_4MQNode_4QNone_Bool_1_r;
  QTree_Bool_t lizzieLet0_4MQNode_4QNone_Bool_2_d;
  logic lizzieLet0_4MQNode_4QNone_Bool_2_r;
  QTree_Bool_t lizzieLet0_4MQNode_4QNone_Bool_3_d;
  logic lizzieLet0_4MQNode_4QNone_Bool_3_r;
  QTree_Bool_t lizzieLet0_4MQNode_4QNone_Bool_4_d;
  logic lizzieLet0_4MQNode_4QNone_Bool_4_r;
  QTree_Bool_t lizzieLet0_4MQNode_4QNone_Bool_5_d;
  logic lizzieLet0_4MQNode_4QNone_Bool_5_r;
  QTree_Bool_t lizzieLet0_4MQNode_4QNone_Bool_6_d;
  logic lizzieLet0_4MQNode_4QNone_Bool_6_r;
  QTree_Bool_t lizzieLet0_4MQNode_4QNone_Bool_7_d;
  logic lizzieLet0_4MQNode_4QNone_Bool_7_r;
  QTree_Bool_t lizzieLet0_4MQNode_4QNone_Bool_8_d;
  logic lizzieLet0_4MQNode_4QNone_Bool_8_r;
  Pointer_QTree_Bool_t t1a8d_destruct_d;
  logic t1a8d_destruct_r;
  Pointer_QTree_Bool_t t2a8e_destruct_d;
  logic t2a8e_destruct_r;
  Pointer_QTree_Bool_t t3a8f_destruct_d;
  logic t3a8f_destruct_r;
  Pointer_QTree_Bool_t t4a8g_destruct_d;
  logic t4a8g_destruct_r;
  QTree_Bool_t _99_d;
  logic _99_r;
  assign _99_r = 1'd1;
  QTree_Bool_t _98_d;
  logic _98_r;
  assign _98_r = 1'd1;
  QTree_Bool_t lizzieLet0_4MQNode_4QNone_Bool_1QNode_Bool_d;
  logic lizzieLet0_4MQNode_4QNone_Bool_1QNode_Bool_r;
  QTree_Bool_t _97_d;
  logic _97_r;
  assign _97_r = 1'd1;
  Go_t lizzieLet0_4MQNode_4QNone_Bool_3QNone_Bool_d;
  logic lizzieLet0_4MQNode_4QNone_Bool_3QNone_Bool_r;
  Go_t lizzieLet0_4MQNode_4QNone_Bool_3QVal_Bool_d;
  logic lizzieLet0_4MQNode_4QNone_Bool_3QVal_Bool_r;
  Go_t lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_d;
  logic lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_r;
  Go_t lizzieLet0_4MQNode_4QNone_Bool_3QError_Bool_d;
  logic lizzieLet0_4MQNode_4QNone_Bool_3QError_Bool_r;
  Go_t lizzieLet0_4MQNode_4QNone_Bool_3QError_Bool_1_d;
  logic lizzieLet0_4MQNode_4QNone_Bool_3QError_Bool_1_r;
  Go_t lizzieLet0_4MQNode_4QNone_Bool_3QError_Bool_2_d;
  logic lizzieLet0_4MQNode_4QNone_Bool_3QError_Bool_2_r;
  QTree_Bool_t lizzieLet0_4MQNode_4QNone_Bool_3QError_Bool_1QError_Bool_d;
  logic lizzieLet0_4MQNode_4QNone_Bool_3QError_Bool_1QError_Bool_r;
  QTree_Bool_t lizzieLet7_1_argbuf_d;
  logic lizzieLet7_1_argbuf_r;
  Go_t lizzieLet0_4MQNode_4QNone_Bool_3QError_Bool_2_argbuf_d;
  logic lizzieLet0_4MQNode_4QNone_Bool_3QError_Bool_2_argbuf_r;
  Go_t lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_1_d;
  logic lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_1_r;
  Go_t lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_2_d;
  logic lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_2_r;
  Go_t lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_3_d;
  logic lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_3_r;
  Go_t lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_4_d;
  logic lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_4_r;
  Go_t lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_5_d;
  logic lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_5_r;
  Go_t lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_1_argbuf_d;
  logic lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_1_argbuf_r;
  TupGo___Pointer_MaskQTree___Pointer_QTree_Bool_t \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool_1_d ;
  logic \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool_1_r ;
  Go_t lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_2_argbuf_d;
  logic lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_2_argbuf_r;
  TupGo___Pointer_MaskQTree___Pointer_QTree_Bool_t \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool2_d ;
  logic \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool2_r ;
  Go_t lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_3_argbuf_d;
  logic lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_3_argbuf_r;
  TupGo___Pointer_MaskQTree___Pointer_QTree_Bool_t \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool3_d ;
  logic \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool3_r ;
  Go_t lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_4_argbuf_d;
  logic lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_4_argbuf_r;
  TupGo___Pointer_MaskQTree___Pointer_QTree_Bool_t \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool4_d ;
  logic \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool4_r ;
  Go_t lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_5_argbuf_d;
  logic lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_5_argbuf_r;
  Go_t lizzieLet0_4MQNode_4QNone_Bool_3QNone_Bool_1_d;
  logic lizzieLet0_4MQNode_4QNone_Bool_3QNone_Bool_1_r;
  Go_t lizzieLet0_4MQNode_4QNone_Bool_3QNone_Bool_2_d;
  logic lizzieLet0_4MQNode_4QNone_Bool_3QNone_Bool_2_r;
  QTree_Bool_t lizzieLet0_4MQNode_4QNone_Bool_3QNone_Bool_1QNone_Bool_d;
  logic lizzieLet0_4MQNode_4QNone_Bool_3QNone_Bool_1QNone_Bool_r;
  QTree_Bool_t lizzieLet4_1_argbuf_d;
  logic lizzieLet4_1_argbuf_r;
  Go_t lizzieLet0_4MQNode_4QNone_Bool_3QNone_Bool_2_argbuf_d;
  logic lizzieLet0_4MQNode_4QNone_Bool_3QNone_Bool_2_argbuf_r;
  Go_t lizzieLet0_4MQNode_4QNone_Bool_3QVal_Bool_1_d;
  logic lizzieLet0_4MQNode_4QNone_Bool_3QVal_Bool_1_r;
  Go_t lizzieLet0_4MQNode_4QNone_Bool_3QVal_Bool_2_d;
  logic lizzieLet0_4MQNode_4QNone_Bool_3QVal_Bool_2_r;
  QTree_Bool_t lizzieLet0_4MQNode_4QNone_Bool_3QVal_Bool_1QError_Bool_d;
  logic lizzieLet0_4MQNode_4QNone_Bool_3QVal_Bool_1QError_Bool_r;
  QTree_Bool_t lizzieLet5_1_argbuf_d;
  logic lizzieLet5_1_argbuf_r;
  Go_t lizzieLet0_4MQNode_4QNone_Bool_3QVal_Bool_2_argbuf_d;
  logic lizzieLet0_4MQNode_4QNone_Bool_3QVal_Bool_2_argbuf_r;
  Pointer_CTf_t lizzieLet0_4MQNode_4QNone_Bool_4QNone_Bool_d;
  logic lizzieLet0_4MQNode_4QNone_Bool_4QNone_Bool_r;
  Pointer_CTf_t lizzieLet0_4MQNode_4QNone_Bool_4QVal_Bool_d;
  logic lizzieLet0_4MQNode_4QNone_Bool_4QVal_Bool_r;
  Pointer_CTf_t lizzieLet0_4MQNode_4QNone_Bool_4QNode_Bool_d;
  logic lizzieLet0_4MQNode_4QNone_Bool_4QNode_Bool_r;
  Pointer_CTf_t lizzieLet0_4MQNode_4QNone_Bool_4QError_Bool_d;
  logic lizzieLet0_4MQNode_4QNone_Bool_4QError_Bool_r;
  Pointer_CTf_t lizzieLet0_4MQNode_4QNone_Bool_4QError_Bool_1_argbuf_d;
  logic lizzieLet0_4MQNode_4QNone_Bool_4QError_Bool_1_argbuf_r;
  Pointer_CTf_t lizzieLet0_4MQNode_4QNone_Bool_4QNode_Bool_1_argbuf_d;
  logic lizzieLet0_4MQNode_4QNone_Bool_4QNode_Bool_1_argbuf_r;
  Pointer_CTf_t lizzieLet0_4MQNode_4QNone_Bool_4QNone_Bool_1_argbuf_d;
  logic lizzieLet0_4MQNode_4QNone_Bool_4QNone_Bool_1_argbuf_r;
  Pointer_CTf_t lizzieLet0_4MQNode_4QNone_Bool_4QVal_Bool_1_argbuf_d;
  logic lizzieLet0_4MQNode_4QNone_Bool_4QVal_Bool_1_argbuf_r;
  Pointer_MaskQTree_t _96_d;
  logic _96_r;
  assign _96_r = 1'd1;
  Pointer_MaskQTree_t _95_d;
  logic _95_r;
  assign _95_r = 1'd1;
  Pointer_MaskQTree_t lizzieLet0_4MQNode_4QNone_Bool_5QNode_Bool_d;
  logic lizzieLet0_4MQNode_4QNone_Bool_5QNode_Bool_r;
  Pointer_MaskQTree_t _94_d;
  logic _94_r;
  assign _94_r = 1'd1;
  Pointer_MaskQTree_t lizzieLet0_4MQNode_4QNone_Bool_5QNode_Bool_1_argbuf_d;
  logic lizzieLet0_4MQNode_4QNone_Bool_5QNode_Bool_1_argbuf_r;
  Pointer_MaskQTree_t _93_d;
  logic _93_r;
  assign _93_r = 1'd1;
  Pointer_MaskQTree_t _92_d;
  logic _92_r;
  assign _92_r = 1'd1;
  Pointer_MaskQTree_t lizzieLet0_4MQNode_4QNone_Bool_6QNode_Bool_d;
  logic lizzieLet0_4MQNode_4QNone_Bool_6QNode_Bool_r;
  Pointer_MaskQTree_t _91_d;
  logic _91_r;
  assign _91_r = 1'd1;
  Pointer_MaskQTree_t lizzieLet0_4MQNode_4QNone_Bool_6QNode_Bool_1_argbuf_d;
  logic lizzieLet0_4MQNode_4QNone_Bool_6QNode_Bool_1_argbuf_r;
  Pointer_MaskQTree_t _90_d;
  logic _90_r;
  assign _90_r = 1'd1;
  Pointer_MaskQTree_t _89_d;
  logic _89_r;
  assign _89_r = 1'd1;
  Pointer_MaskQTree_t lizzieLet0_4MQNode_4QNone_Bool_7QNode_Bool_d;
  logic lizzieLet0_4MQNode_4QNone_Bool_7QNode_Bool_r;
  Pointer_MaskQTree_t _88_d;
  logic _88_r;
  assign _88_r = 1'd1;
  Pointer_MaskQTree_t lizzieLet0_4MQNode_4QNone_Bool_7QNode_Bool_1_argbuf_d;
  logic lizzieLet0_4MQNode_4QNone_Bool_7QNode_Bool_1_argbuf_r;
  Pointer_MaskQTree_t _87_d;
  logic _87_r;
  assign _87_r = 1'd1;
  Pointer_MaskQTree_t _86_d;
  logic _86_r;
  assign _86_r = 1'd1;
  Pointer_MaskQTree_t lizzieLet0_4MQNode_4QNone_Bool_8QNode_Bool_d;
  logic lizzieLet0_4MQNode_4QNone_Bool_8QNode_Bool_r;
  Pointer_MaskQTree_t _85_d;
  logic _85_r;
  assign _85_r = 1'd1;
  Pointer_MaskQTree_t lizzieLet0_4MQNode_4QNone_Bool_8QNode_Bool_1_argbuf_d;
  logic lizzieLet0_4MQNode_4QNone_Bool_8QNode_Bool_1_argbuf_r;
  QTree_Bool_t lizzieLet0_4MQNode_4QVal_Bool_1_d;
  logic lizzieLet0_4MQNode_4QVal_Bool_1_r;
  QTree_Bool_t lizzieLet0_4MQNode_4QVal_Bool_2_d;
  logic lizzieLet0_4MQNode_4QVal_Bool_2_r;
  QTree_Bool_t lizzieLet0_4MQNode_4QVal_Bool_3_d;
  logic lizzieLet0_4MQNode_4QVal_Bool_3_r;
  QTree_Bool_t lizzieLet0_4MQNode_4QVal_Bool_4_d;
  logic lizzieLet0_4MQNode_4QVal_Bool_4_r;
  QTree_Bool_t lizzieLet0_4MQNode_4QVal_Bool_5_d;
  logic lizzieLet0_4MQNode_4QVal_Bool_5_r;
  MyBool_t va8i_destruct_d;
  logic va8i_destruct_r;
  QTree_Bool_t _84_d;
  logic _84_r;
  assign _84_r = 1'd1;
  QTree_Bool_t lizzieLet0_4MQNode_4QVal_Bool_1QVal_Bool_d;
  logic lizzieLet0_4MQNode_4QVal_Bool_1QVal_Bool_r;
  QTree_Bool_t _83_d;
  logic _83_r;
  assign _83_r = 1'd1;
  QTree_Bool_t _82_d;
  logic _82_r;
  assign _82_r = 1'd1;
  Go_t lizzieLet0_4MQNode_4QVal_Bool_3QNone_Bool_d;
  logic lizzieLet0_4MQNode_4QVal_Bool_3QNone_Bool_r;
  Go_t lizzieLet0_4MQNode_4QVal_Bool_3QVal_Bool_d;
  logic lizzieLet0_4MQNode_4QVal_Bool_3QVal_Bool_r;
  Go_t lizzieLet0_4MQNode_4QVal_Bool_3QNode_Bool_d;
  logic lizzieLet0_4MQNode_4QVal_Bool_3QNode_Bool_r;
  Go_t lizzieLet0_4MQNode_4QVal_Bool_3QError_Bool_d;
  logic lizzieLet0_4MQNode_4QVal_Bool_3QError_Bool_r;
  Go_t lizzieLet0_4MQNode_4QVal_Bool_3QError_Bool_1_d;
  logic lizzieLet0_4MQNode_4QVal_Bool_3QError_Bool_1_r;
  Go_t lizzieLet0_4MQNode_4QVal_Bool_3QError_Bool_2_d;
  logic lizzieLet0_4MQNode_4QVal_Bool_3QError_Bool_2_r;
  QTree_Bool_t lizzieLet0_4MQNode_4QVal_Bool_3QError_Bool_1QError_Bool_d;
  logic lizzieLet0_4MQNode_4QVal_Bool_3QError_Bool_1QError_Bool_r;
  QTree_Bool_t lizzieLet9_1_1_argbuf_d;
  logic lizzieLet9_1_1_argbuf_r;
  Go_t lizzieLet0_4MQNode_4QVal_Bool_3QError_Bool_2_argbuf_d;
  logic lizzieLet0_4MQNode_4QVal_Bool_3QError_Bool_2_argbuf_r;
  Go_t lizzieLet0_4MQNode_4QVal_Bool_3QNode_Bool_1_d;
  logic lizzieLet0_4MQNode_4QVal_Bool_3QNode_Bool_1_r;
  Go_t lizzieLet0_4MQNode_4QVal_Bool_3QNode_Bool_2_d;
  logic lizzieLet0_4MQNode_4QVal_Bool_3QNode_Bool_2_r;
  QTree_Bool_t lizzieLet0_4MQNode_4QVal_Bool_3QNode_Bool_1QError_Bool_d;
  logic lizzieLet0_4MQNode_4QVal_Bool_3QNode_Bool_1QError_Bool_r;
  QTree_Bool_t lizzieLet13_1_1_argbuf_d;
  logic lizzieLet13_1_1_argbuf_r;
  Go_t lizzieLet0_4MQNode_4QVal_Bool_3QNode_Bool_2_argbuf_d;
  logic lizzieLet0_4MQNode_4QVal_Bool_3QNode_Bool_2_argbuf_r;
  Go_t lizzieLet0_4MQNode_4QVal_Bool_3QNone_Bool_1_d;
  logic lizzieLet0_4MQNode_4QVal_Bool_3QNone_Bool_1_r;
  Go_t lizzieLet0_4MQNode_4QVal_Bool_3QNone_Bool_2_d;
  logic lizzieLet0_4MQNode_4QVal_Bool_3QNone_Bool_2_r;
  QTree_Bool_t lizzieLet0_4MQNode_4QVal_Bool_3QNone_Bool_1QError_Bool_d;
  logic lizzieLet0_4MQNode_4QVal_Bool_3QNone_Bool_1QError_Bool_r;
  QTree_Bool_t lizzieLet9_1_argbuf_d;
  logic lizzieLet9_1_argbuf_r;
  Go_t lizzieLet0_4MQNode_4QVal_Bool_3QNone_Bool_2_argbuf_d;
  logic lizzieLet0_4MQNode_4QVal_Bool_3QNone_Bool_2_argbuf_r;
  Pointer_CTf_t lizzieLet0_4MQNode_4QVal_Bool_4QNone_Bool_d;
  logic lizzieLet0_4MQNode_4QVal_Bool_4QNone_Bool_r;
  Pointer_CTf_t lizzieLet0_4MQNode_4QVal_Bool_4QVal_Bool_d;
  logic lizzieLet0_4MQNode_4QVal_Bool_4QVal_Bool_r;
  Pointer_CTf_t lizzieLet0_4MQNode_4QVal_Bool_4QNode_Bool_d;
  logic lizzieLet0_4MQNode_4QVal_Bool_4QNode_Bool_r;
  Pointer_CTf_t lizzieLet0_4MQNode_4QVal_Bool_4QError_Bool_d;
  logic lizzieLet0_4MQNode_4QVal_Bool_4QError_Bool_r;
  Pointer_CTf_t lizzieLet0_4MQNode_4QVal_Bool_4QError_Bool_1_argbuf_d;
  logic lizzieLet0_4MQNode_4QVal_Bool_4QError_Bool_1_argbuf_r;
  Pointer_CTf_t lizzieLet0_4MQNode_4QVal_Bool_4QNode_Bool_1_argbuf_d;
  logic lizzieLet0_4MQNode_4QVal_Bool_4QNode_Bool_1_argbuf_r;
  Pointer_CTf_t lizzieLet0_4MQNode_4QVal_Bool_4QNone_Bool_1_argbuf_d;
  logic lizzieLet0_4MQNode_4QVal_Bool_4QNone_Bool_1_argbuf_r;
  MyBool_t _81_d;
  logic _81_r;
  assign _81_r = 1'd1;
  MyBool_t lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_d;
  logic lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_r;
  MyBool_t _80_d;
  logic _80_r;
  assign _80_r = 1'd1;
  MyBool_t _79_d;
  logic _79_r;
  assign _79_r = 1'd1;
  MyBool_t lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1_d;
  logic lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1_r;
  MyBool_t lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_2_d;
  logic lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_2_r;
  MyBool_t lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3_d;
  logic lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3_r;
  Go_t lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyFalse_d;
  logic lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyFalse_r;
  Go_t lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyTrue_d;
  logic lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyTrue_r;
  Go_t lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyTrue_1_d;
  logic lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyTrue_1_r;
  Go_t lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyTrue_2_d;
  logic lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyTrue_2_r;
  QTree_Bool_t lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyTrue_1QError_Bool_d;
  logic lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyTrue_1QError_Bool_r;
  QTree_Bool_t lizzieLet12_1_argbuf_d;
  logic lizzieLet12_1_argbuf_r;
  Go_t lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyTrue_2_argbuf_d;
  logic lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyTrue_2_argbuf_r;
  Pointer_CTf_t lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_2MyFalse_d;
  logic lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_2MyFalse_r;
  Pointer_CTf_t lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_2MyTrue_d;
  logic lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_2MyTrue_r;
  Pointer_CTf_t lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_2MyTrue_1_argbuf_d;
  logic lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_2MyTrue_1_argbuf_r;
  MyBool_t lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_d;
  logic lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_r;
  MyBool_t _78_d;
  logic _78_r;
  assign _78_r = 1'd1;
  MyBool_t lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1_d;
  logic lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1_r;
  MyBool_t lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_2_d;
  logic lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_2_r;
  Go_t lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyFalse_d;
  logic lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyFalse_r;
  Go_t lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyTrue_d;
  logic lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyTrue_r;
  Go_t lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyFalse_1_d;
  logic lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyFalse_1_r;
  Go_t lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyFalse_2_d;
  logic lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyFalse_2_r;
  QTree_Bool_t lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_d;
  logic lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_r;
  QTree_Bool_t lizzieLet10_1_argbuf_d;
  logic lizzieLet10_1_argbuf_r;
  Go_t lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyFalse_2_argbuf_d;
  logic lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyFalse_2_argbuf_r;
  Go_t lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyTrue_1_d;
  logic lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyTrue_1_r;
  Go_t lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyTrue_2_d;
  logic lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyTrue_2_r;
  QTree_Bool_t lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyTrue_1QError_Bool_d;
  logic lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyTrue_1QError_Bool_r;
  QTree_Bool_t lizzieLet11_1_argbuf_d;
  logic lizzieLet11_1_argbuf_r;
  Go_t lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyTrue_2_argbuf_d;
  logic lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyTrue_2_argbuf_r;
  Pointer_CTf_t lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_2MyFalse_d;
  logic lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_2MyFalse_r;
  Pointer_CTf_t lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_2MyTrue_d;
  logic lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_2MyTrue_r;
  Pointer_CTf_t lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_2MyFalse_1_argbuf_d;
  logic lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_2MyFalse_1_argbuf_r;
  Pointer_CTf_t lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_2MyTrue_1_argbuf_d;
  logic lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_2MyTrue_1_argbuf_r;
  Pointer_CTf_t lizzieLet0_4MQNode_5QNone_Bool_d;
  logic lizzieLet0_4MQNode_5QNone_Bool_r;
  Pointer_CTf_t lizzieLet0_4MQNode_5QVal_Bool_d;
  logic lizzieLet0_4MQNode_5QVal_Bool_r;
  Pointer_CTf_t lizzieLet0_4MQNode_5QNode_Bool_d;
  logic lizzieLet0_4MQNode_5QNode_Bool_r;
  Pointer_CTf_t lizzieLet0_4MQNode_5QError_Bool_d;
  logic lizzieLet0_4MQNode_5QError_Bool_r;
  Pointer_CTf_t lizzieLet0_4MQNode_5QError_Bool_1_argbuf_d;
  logic lizzieLet0_4MQNode_5QError_Bool_1_argbuf_r;
  Pointer_MaskQTree_t lizzieLet0_4MQNode_6QNone_Bool_d;
  logic lizzieLet0_4MQNode_6QNone_Bool_r;
  Pointer_MaskQTree_t _77_d;
  logic _77_r;
  assign _77_r = 1'd1;
  Pointer_MaskQTree_t lizzieLet0_4MQNode_6QNode_Bool_d;
  logic lizzieLet0_4MQNode_6QNode_Bool_r;
  Pointer_MaskQTree_t _76_d;
  logic _76_r;
  assign _76_r = 1'd1;
  Pointer_MaskQTree_t lizzieLet0_4MQNode_7QNone_Bool_d;
  logic lizzieLet0_4MQNode_7QNone_Bool_r;
  Pointer_MaskQTree_t _75_d;
  logic _75_r;
  assign _75_r = 1'd1;
  Pointer_MaskQTree_t lizzieLet0_4MQNode_7QNode_Bool_d;
  logic lizzieLet0_4MQNode_7QNode_Bool_r;
  Pointer_MaskQTree_t _74_d;
  logic _74_r;
  assign _74_r = 1'd1;
  Pointer_MaskQTree_t lizzieLet0_4MQNode_8QNone_Bool_d;
  logic lizzieLet0_4MQNode_8QNone_Bool_r;
  Pointer_MaskQTree_t _73_d;
  logic _73_r;
  assign _73_r = 1'd1;
  Pointer_MaskQTree_t lizzieLet0_4MQNode_8QNode_Bool_d;
  logic lizzieLet0_4MQNode_8QNode_Bool_r;
  Pointer_MaskQTree_t _72_d;
  logic _72_r;
  assign _72_r = 1'd1;
  Pointer_MaskQTree_t lizzieLet0_4MQNode_9QNone_Bool_d;
  logic lizzieLet0_4MQNode_9QNone_Bool_r;
  Pointer_MaskQTree_t _71_d;
  logic _71_r;
  assign _71_r = 1'd1;
  Pointer_MaskQTree_t lizzieLet0_4MQNode_9QNode_Bool_d;
  logic lizzieLet0_4MQNode_9QNode_Bool_r;
  Pointer_MaskQTree_t _70_d;
  logic _70_r;
  assign _70_r = 1'd1;
  QTree_Bool_t _69_d;
  logic _69_r;
  assign _69_r = 1'd1;
  QTree_Bool_t _68_d;
  logic _68_r;
  assign _68_r = 1'd1;
  QTree_Bool_t lizzieLet0_5MQNode_d;
  logic lizzieLet0_5MQNode_r;
  Pointer_QTree_Bool_t _67_d;
  logic _67_r;
  assign _67_r = 1'd1;
  Pointer_QTree_Bool_t lizzieLet0_6MQVal_d;
  logic lizzieLet0_6MQVal_r;
  Pointer_QTree_Bool_t _66_d;
  logic _66_r;
  assign _66_r = 1'd1;
  Pointer_QTree_Bool_t lizzieLet0_6MQVal_1_argbuf_d;
  logic lizzieLet0_6MQVal_1_argbuf_r;
  Pointer_QTree_Bool_t _65_d;
  logic _65_r;
  assign _65_r = 1'd1;
  Pointer_QTree_Bool_t lizzieLet0_7MQVal_d;
  logic lizzieLet0_7MQVal_r;
  Pointer_QTree_Bool_t _64_d;
  logic _64_r;
  assign _64_r = 1'd1;
  Pointer_QTree_Bool_t lizzieLet0_7MQVal_1_argbuf_d;
  logic lizzieLet0_7MQVal_1_argbuf_r;
  Pointer_CTf_t lizzieLet0_8MQNone_d;
  logic lizzieLet0_8MQNone_r;
  Pointer_CTf_t lizzieLet0_8MQVal_d;
  logic lizzieLet0_8MQVal_r;
  Pointer_CTf_t lizzieLet0_8MQNode_d;
  logic lizzieLet0_8MQNode_r;
  Pointer_CTf_t lizzieLet0_8MQNone_1_argbuf_d;
  logic lizzieLet0_8MQNone_1_argbuf_r;
  Pointer_CTf_t lizzieLet0_8MQVal_1_argbuf_d;
  logic lizzieLet0_8MQVal_1_argbuf_r;
  Pointer_QTree_Bool_t q1a8P_destruct_d;
  logic q1a8P_destruct_r;
  Pointer_QTree_Bool_t q2a8Q_destruct_d;
  logic q2a8Q_destruct_r;
  Pointer_QTree_Bool_t q3a8R_destruct_d;
  logic q3a8R_destruct_r;
  Pointer_QTree_Bool_t q4a8S_destruct_d;
  logic q4a8S_destruct_r;
  MyBool_t v1a8J_destruct_d;
  logic v1a8J_destruct_r;
  QTree_Bool_t _63_d;
  logic _63_r;
  assign _63_r = 1'd1;
  QTree_Bool_t lizzieLet20_1_1QVal_Bool_d;
  logic lizzieLet20_1_1QVal_Bool_r;
  QTree_Bool_t lizzieLet20_1_1QNode_Bool_d;
  logic lizzieLet20_1_1QNode_Bool_r;
  QTree_Bool_t _62_d;
  logic _62_r;
  assign _62_r = 1'd1;
  Go_t lizzieLet20_1_3QNone_Bool_d;
  logic lizzieLet20_1_3QNone_Bool_r;
  Go_t lizzieLet20_1_3QVal_Bool_d;
  logic lizzieLet20_1_3QVal_Bool_r;
  Go_t lizzieLet20_1_3QNode_Bool_d;
  logic lizzieLet20_1_3QNode_Bool_r;
  Go_t lizzieLet20_1_3QError_Bool_d;
  logic lizzieLet20_1_3QError_Bool_r;
  Go_t lizzieLet20_1_3QError_Bool_1_d;
  logic lizzieLet20_1_3QError_Bool_1_r;
  Go_t lizzieLet20_1_3QError_Bool_2_d;
  logic lizzieLet20_1_3QError_Bool_2_r;
  QTree_Bool_t lizzieLet20_1_3QError_Bool_1QError_Bool_d;
  logic lizzieLet20_1_3QError_Bool_1QError_Bool_r;
  QTree_Bool_t lizzieLet31_1_argbuf_d;
  logic lizzieLet31_1_argbuf_r;
  Go_t lizzieLet20_1_3QError_Bool_2_argbuf_d;
  logic lizzieLet20_1_3QError_Bool_2_argbuf_r;
  Go_t lizzieLet20_1_3QNone_Bool_1_argbuf_d;
  logic lizzieLet20_1_3QNone_Bool_1_argbuf_r;
  C12_t go_10_goMux_choice_d;
  logic go_10_goMux_choice_r;
  Go_t go_10_goMux_data_d;
  logic go_10_goMux_data_r;
  QTree_Bool_t _61_d;
  logic _61_r;
  assign _61_r = 1'd1;
  QTree_Bool_t lizzieLet20_1_4QVal_Bool_d;
  logic lizzieLet20_1_4QVal_Bool_r;
  QTree_Bool_t lizzieLet20_1_4QNode_Bool_d;
  logic lizzieLet20_1_4QNode_Bool_r;
  QTree_Bool_t _60_d;
  logic _60_r;
  assign _60_r = 1'd1;
  QTree_Bool_t lizzieLet20_1_4QNode_Bool_1_d;
  logic lizzieLet20_1_4QNode_Bool_1_r;
  QTree_Bool_t lizzieLet20_1_4QNode_Bool_2_d;
  logic lizzieLet20_1_4QNode_Bool_2_r;
  QTree_Bool_t lizzieLet20_1_4QNode_Bool_3_d;
  logic lizzieLet20_1_4QNode_Bool_3_r;
  QTree_Bool_t lizzieLet20_1_4QNode_Bool_4_d;
  logic lizzieLet20_1_4QNode_Bool_4_r;
  QTree_Bool_t lizzieLet20_1_4QNode_Bool_5_d;
  logic lizzieLet20_1_4QNode_Bool_5_r;
  QTree_Bool_t lizzieLet20_1_4QNode_Bool_6_d;
  logic lizzieLet20_1_4QNode_Bool_6_r;
  QTree_Bool_t lizzieLet20_1_4QNode_Bool_7_d;
  logic lizzieLet20_1_4QNode_Bool_7_r;
  QTree_Bool_t lizzieLet20_1_4QNode_Bool_8_d;
  logic lizzieLet20_1_4QNode_Bool_8_r;
  QTree_Bool_t lizzieLet20_1_4QNode_Bool_9_d;
  logic lizzieLet20_1_4QNode_Bool_9_r;
  Pointer_QTree_Bool_t t1a8U_destruct_d;
  logic t1a8U_destruct_r;
  Pointer_QTree_Bool_t t2a8V_destruct_d;
  logic t2a8V_destruct_r;
  Pointer_QTree_Bool_t t3a8W_destruct_d;
  logic t3a8W_destruct_r;
  Pointer_QTree_Bool_t t4a8X_destruct_d;
  logic t4a8X_destruct_r;
  QTree_Bool_t _59_d;
  logic _59_r;
  assign _59_r = 1'd1;
  QTree_Bool_t _58_d;
  logic _58_r;
  assign _58_r = 1'd1;
  QTree_Bool_t lizzieLet20_1_4QNode_Bool_1QNode_Bool_d;
  logic lizzieLet20_1_4QNode_Bool_1QNode_Bool_r;
  QTree_Bool_t _57_d;
  logic _57_r;
  assign _57_r = 1'd1;
  Go_t lizzieLet20_1_4QNode_Bool_3QNone_Bool_d;
  logic lizzieLet20_1_4QNode_Bool_3QNone_Bool_r;
  Go_t lizzieLet20_1_4QNode_Bool_3QVal_Bool_d;
  logic lizzieLet20_1_4QNode_Bool_3QVal_Bool_r;
  Go_t lizzieLet20_1_4QNode_Bool_3QNode_Bool_d;
  logic lizzieLet20_1_4QNode_Bool_3QNode_Bool_r;
  Go_t lizzieLet20_1_4QNode_Bool_3QError_Bool_d;
  logic lizzieLet20_1_4QNode_Bool_3QError_Bool_r;
  Go_t lizzieLet20_1_4QNode_Bool_3QError_Bool_1_d;
  logic lizzieLet20_1_4QNode_Bool_3QError_Bool_1_r;
  Go_t lizzieLet20_1_4QNode_Bool_3QError_Bool_2_d;
  logic lizzieLet20_1_4QNode_Bool_3QError_Bool_2_r;
  QTree_Bool_t lizzieLet20_1_4QNode_Bool_3QError_Bool_1QError_Bool_d;
  logic lizzieLet20_1_4QNode_Bool_3QError_Bool_1QError_Bool_r;
  QTree_Bool_t lizzieLet30_1_argbuf_d;
  logic lizzieLet30_1_argbuf_r;
  Go_t lizzieLet20_1_4QNode_Bool_3QError_Bool_2_argbuf_d;
  logic lizzieLet20_1_4QNode_Bool_3QError_Bool_2_argbuf_r;
  Go_t lizzieLet20_1_4QNode_Bool_3QNode_Bool_1_argbuf_d;
  logic lizzieLet20_1_4QNode_Bool_3QNode_Bool_1_argbuf_r;
  Go_t lizzieLet20_1_4QNode_Bool_3QNone_Bool_1_argbuf_d;
  logic lizzieLet20_1_4QNode_Bool_3QNone_Bool_1_argbuf_r;
  Go_t lizzieLet20_1_4QNode_Bool_3QVal_Bool_1_d;
  logic lizzieLet20_1_4QNode_Bool_3QVal_Bool_1_r;
  Go_t lizzieLet20_1_4QNode_Bool_3QVal_Bool_2_d;
  logic lizzieLet20_1_4QNode_Bool_3QVal_Bool_2_r;
  QTree_Bool_t lizzieLet20_1_4QNode_Bool_3QVal_Bool_1QError_Bool_d;
  logic lizzieLet20_1_4QNode_Bool_3QVal_Bool_1QError_Bool_r;
  QTree_Bool_t lizzieLet28_1_argbuf_d;
  logic lizzieLet28_1_argbuf_r;
  Go_t lizzieLet20_1_4QNode_Bool_3QVal_Bool_2_argbuf_d;
  logic lizzieLet20_1_4QNode_Bool_3QVal_Bool_2_argbuf_r;
  Pointer_QTree_Bool_t lizzieLet20_1_4QNode_Bool_4QNone_Bool_d;
  logic lizzieLet20_1_4QNode_Bool_4QNone_Bool_r;
  Pointer_QTree_Bool_t _56_d;
  logic _56_r;
  assign _56_r = 1'd1;
  Pointer_QTree_Bool_t _55_d;
  logic _55_r;
  assign _55_r = 1'd1;
  Pointer_QTree_Bool_t _54_d;
  logic _54_r;
  assign _54_r = 1'd1;
  Pointer_QTree_Bool_t lizzieLet20_1_4QNode_Bool_4QNone_Bool_1_argbuf_d;
  logic lizzieLet20_1_4QNode_Bool_4QNone_Bool_1_argbuf_r;
  \Pointer_CTf'_t  lizzieLet20_1_4QNode_Bool_5QNone_Bool_d;
  logic lizzieLet20_1_4QNode_Bool_5QNone_Bool_r;
  \Pointer_CTf'_t  lizzieLet20_1_4QNode_Bool_5QVal_Bool_d;
  logic lizzieLet20_1_4QNode_Bool_5QVal_Bool_r;
  \Pointer_CTf'_t  lizzieLet20_1_4QNode_Bool_5QNode_Bool_d;
  logic lizzieLet20_1_4QNode_Bool_5QNode_Bool_r;
  \Pointer_CTf'_t  lizzieLet20_1_4QNode_Bool_5QError_Bool_d;
  logic lizzieLet20_1_4QNode_Bool_5QError_Bool_r;
  \Pointer_CTf'_t  lizzieLet20_1_4QNode_Bool_5QError_Bool_1_argbuf_d;
  logic lizzieLet20_1_4QNode_Bool_5QError_Bool_1_argbuf_r;
  \CTf'_t  \lizzieLet20_1_4QNode_Bool_5QNode_Bool_1lizzieLet20_1_4QNode_Bool_6QNode_Bool_1t1a8U_1lizzieLet20_1_4QNode_Bool_7QNode_Bool_1t2a8V_1lizzieLet20_1_4QNode_Bool_8QNode_Bool_1t3a8W_1Lcall_f'3_d ;
  logic \lizzieLet20_1_4QNode_Bool_5QNode_Bool_1lizzieLet20_1_4QNode_Bool_6QNode_Bool_1t1a8U_1lizzieLet20_1_4QNode_Bool_7QNode_Bool_1t2a8V_1lizzieLet20_1_4QNode_Bool_8QNode_Bool_1t3a8W_1Lcall_f'3_r ;
  \CTf'_t  lizzieLet29_1_argbuf_d;
  logic lizzieLet29_1_argbuf_r;
  \Pointer_CTf'_t  lizzieLet20_1_4QNode_Bool_5QNone_Bool_1_argbuf_d;
  logic lizzieLet20_1_4QNode_Bool_5QNone_Bool_1_argbuf_r;
  \Pointer_CTf'_t  lizzieLet20_1_4QNode_Bool_5QVal_Bool_1_argbuf_d;
  logic lizzieLet20_1_4QNode_Bool_5QVal_Bool_1_argbuf_r;
  Pointer_QTree_Bool_t _53_d;
  logic _53_r;
  assign _53_r = 1'd1;
  Pointer_QTree_Bool_t _52_d;
  logic _52_r;
  assign _52_r = 1'd1;
  Pointer_QTree_Bool_t lizzieLet20_1_4QNode_Bool_6QNode_Bool_d;
  logic lizzieLet20_1_4QNode_Bool_6QNode_Bool_r;
  Pointer_QTree_Bool_t _51_d;
  logic _51_r;
  assign _51_r = 1'd1;
  Pointer_QTree_Bool_t _50_d;
  logic _50_r;
  assign _50_r = 1'd1;
  Pointer_QTree_Bool_t _49_d;
  logic _49_r;
  assign _49_r = 1'd1;
  Pointer_QTree_Bool_t lizzieLet20_1_4QNode_Bool_7QNode_Bool_d;
  logic lizzieLet20_1_4QNode_Bool_7QNode_Bool_r;
  Pointer_QTree_Bool_t _48_d;
  logic _48_r;
  assign _48_r = 1'd1;
  Pointer_QTree_Bool_t _47_d;
  logic _47_r;
  assign _47_r = 1'd1;
  Pointer_QTree_Bool_t _46_d;
  logic _46_r;
  assign _46_r = 1'd1;
  Pointer_QTree_Bool_t lizzieLet20_1_4QNode_Bool_8QNode_Bool_d;
  logic lizzieLet20_1_4QNode_Bool_8QNode_Bool_r;
  Pointer_QTree_Bool_t _45_d;
  logic _45_r;
  assign _45_r = 1'd1;
  Pointer_QTree_Bool_t _44_d;
  logic _44_r;
  assign _44_r = 1'd1;
  Pointer_QTree_Bool_t _43_d;
  logic _43_r;
  assign _43_r = 1'd1;
  Pointer_QTree_Bool_t lizzieLet20_1_4QNode_Bool_9QNode_Bool_d;
  logic lizzieLet20_1_4QNode_Bool_9QNode_Bool_r;
  Pointer_QTree_Bool_t _42_d;
  logic _42_r;
  assign _42_r = 1'd1;
  Pointer_QTree_Bool_t lizzieLet20_1_4QNode_Bool_9QNode_Bool_1_argbuf_d;
  logic lizzieLet20_1_4QNode_Bool_9QNode_Bool_1_argbuf_r;
  QTree_Bool_t lizzieLet20_1_4QVal_Bool_1_d;
  logic lizzieLet20_1_4QVal_Bool_1_r;
  QTree_Bool_t lizzieLet20_1_4QVal_Bool_2_d;
  logic lizzieLet20_1_4QVal_Bool_2_r;
  QTree_Bool_t lizzieLet20_1_4QVal_Bool_3_d;
  logic lizzieLet20_1_4QVal_Bool_3_r;
  QTree_Bool_t lizzieLet20_1_4QVal_Bool_4_d;
  logic lizzieLet20_1_4QVal_Bool_4_r;
  QTree_Bool_t lizzieLet20_1_4QVal_Bool_5_d;
  logic lizzieLet20_1_4QVal_Bool_5_r;
  QTree_Bool_t lizzieLet20_1_4QVal_Bool_6_d;
  logic lizzieLet20_1_4QVal_Bool_6_r;
  MyBool_t va8K_destruct_d;
  logic va8K_destruct_r;
  QTree_Bool_t _41_d;
  logic _41_r;
  assign _41_r = 1'd1;
  QTree_Bool_t lizzieLet20_1_4QVal_Bool_1QVal_Bool_d;
  logic lizzieLet20_1_4QVal_Bool_1QVal_Bool_r;
  QTree_Bool_t _40_d;
  logic _40_r;
  assign _40_r = 1'd1;
  QTree_Bool_t _39_d;
  logic _39_r;
  assign _39_r = 1'd1;
  Go_t lizzieLet20_1_4QVal_Bool_3QNone_Bool_d;
  logic lizzieLet20_1_4QVal_Bool_3QNone_Bool_r;
  Go_t lizzieLet20_1_4QVal_Bool_3QVal_Bool_d;
  logic lizzieLet20_1_4QVal_Bool_3QVal_Bool_r;
  Go_t lizzieLet20_1_4QVal_Bool_3QNode_Bool_d;
  logic lizzieLet20_1_4QVal_Bool_3QNode_Bool_r;
  Go_t lizzieLet20_1_4QVal_Bool_3QError_Bool_d;
  logic lizzieLet20_1_4QVal_Bool_3QError_Bool_r;
  Go_t lizzieLet20_1_4QVal_Bool_3QError_Bool_1_d;
  logic lizzieLet20_1_4QVal_Bool_3QError_Bool_1_r;
  Go_t lizzieLet20_1_4QVal_Bool_3QError_Bool_2_d;
  logic lizzieLet20_1_4QVal_Bool_3QError_Bool_2_r;
  QTree_Bool_t lizzieLet20_1_4QVal_Bool_3QError_Bool_1QError_Bool_d;
  logic lizzieLet20_1_4QVal_Bool_3QError_Bool_1QError_Bool_r;
  QTree_Bool_t lizzieLet26_1_1_argbuf_d;
  logic lizzieLet26_1_1_argbuf_r;
  Go_t lizzieLet20_1_4QVal_Bool_3QError_Bool_2_argbuf_d;
  logic lizzieLet20_1_4QVal_Bool_3QError_Bool_2_argbuf_r;
  Go_t lizzieLet20_1_4QVal_Bool_3QNode_Bool_1_d;
  logic lizzieLet20_1_4QVal_Bool_3QNode_Bool_1_r;
  Go_t lizzieLet20_1_4QVal_Bool_3QNode_Bool_2_d;
  logic lizzieLet20_1_4QVal_Bool_3QNode_Bool_2_r;
  QTree_Bool_t lizzieLet20_1_4QVal_Bool_3QNode_Bool_1QError_Bool_d;
  logic lizzieLet20_1_4QVal_Bool_3QNode_Bool_1QError_Bool_r;
  QTree_Bool_t lizzieLet25_1_1_argbuf_d;
  logic lizzieLet25_1_1_argbuf_r;
  Go_t lizzieLet20_1_4QVal_Bool_3QNode_Bool_2_argbuf_d;
  logic lizzieLet20_1_4QVal_Bool_3QNode_Bool_2_argbuf_r;
  Go_t lizzieLet20_1_4QVal_Bool_3QNone_Bool_1_argbuf_d;
  logic lizzieLet20_1_4QVal_Bool_3QNone_Bool_1_argbuf_r;
  Pointer_QTree_Bool_t lizzieLet20_1_4QVal_Bool_4QNone_Bool_d;
  logic lizzieLet20_1_4QVal_Bool_4QNone_Bool_r;
  Pointer_QTree_Bool_t _38_d;
  logic _38_r;
  assign _38_r = 1'd1;
  Pointer_QTree_Bool_t _37_d;
  logic _37_r;
  assign _37_r = 1'd1;
  Pointer_QTree_Bool_t _36_d;
  logic _36_r;
  assign _36_r = 1'd1;
  Pointer_QTree_Bool_t lizzieLet20_1_4QVal_Bool_4QNone_Bool_1_argbuf_d;
  logic lizzieLet20_1_4QVal_Bool_4QNone_Bool_1_argbuf_r;
  \Pointer_CTf'_t  lizzieLet20_1_4QVal_Bool_5QNone_Bool_d;
  logic lizzieLet20_1_4QVal_Bool_5QNone_Bool_r;
  \Pointer_CTf'_t  lizzieLet20_1_4QVal_Bool_5QVal_Bool_d;
  logic lizzieLet20_1_4QVal_Bool_5QVal_Bool_r;
  \Pointer_CTf'_t  lizzieLet20_1_4QVal_Bool_5QNode_Bool_d;
  logic lizzieLet20_1_4QVal_Bool_5QNode_Bool_r;
  \Pointer_CTf'_t  lizzieLet20_1_4QVal_Bool_5QError_Bool_d;
  logic lizzieLet20_1_4QVal_Bool_5QError_Bool_r;
  \Pointer_CTf'_t  lizzieLet20_1_4QVal_Bool_5QError_Bool_1_argbuf_d;
  logic lizzieLet20_1_4QVal_Bool_5QError_Bool_1_argbuf_r;
  \Pointer_CTf'_t  lizzieLet20_1_4QVal_Bool_5QNode_Bool_1_argbuf_d;
  logic lizzieLet20_1_4QVal_Bool_5QNode_Bool_1_argbuf_r;
  \Pointer_CTf'_t  lizzieLet20_1_4QVal_Bool_5QNone_Bool_1_argbuf_d;
  logic lizzieLet20_1_4QVal_Bool_5QNone_Bool_1_argbuf_r;
  MyBool_t _35_d;
  logic _35_r;
  assign _35_r = 1'd1;
  MyBool_t lizzieLet20_1_4QVal_Bool_6QVal_Bool_d;
  logic lizzieLet20_1_4QVal_Bool_6QVal_Bool_r;
  MyBool_t _34_d;
  logic _34_r;
  assign _34_r = 1'd1;
  MyBool_t _33_d;
  logic _33_r;
  assign _33_r = 1'd1;
  MyBool_t lizzieLet20_1_4QVal_Bool_6QVal_Bool_1_d;
  logic lizzieLet20_1_4QVal_Bool_6QVal_Bool_1_r;
  MyBool_t lizzieLet20_1_4QVal_Bool_6QVal_Bool_2_d;
  logic lizzieLet20_1_4QVal_Bool_6QVal_Bool_2_r;
  MyBool_t lizzieLet20_1_4QVal_Bool_6QVal_Bool_3_d;
  logic lizzieLet20_1_4QVal_Bool_6QVal_Bool_3_r;
  Go_t lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyFalse_d;
  logic lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyFalse_r;
  Go_t lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyTrue_d;
  logic lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyTrue_r;
  Go_t lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyTrue_1_d;
  logic lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyTrue_1_r;
  Go_t lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyTrue_2_d;
  logic lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyTrue_2_r;
  Go_t lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyTrue_1_argbuf_d;
  logic lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyTrue_1_argbuf_r;
  TupGo_t \lvlrcX-0TupGo2_d ;
  logic \lvlrcX-0TupGo2_r ;
  Go_t lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyTrue_2_argbuf_d;
  logic lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyTrue_2_argbuf_r;
  \Pointer_CTf'_t  lizzieLet20_1_4QVal_Bool_6QVal_Bool_2MyFalse_d;
  logic lizzieLet20_1_4QVal_Bool_6QVal_Bool_2MyFalse_r;
  \Pointer_CTf'_t  lizzieLet20_1_4QVal_Bool_6QVal_Bool_2MyTrue_d;
  logic lizzieLet20_1_4QVal_Bool_6QVal_Bool_2MyTrue_r;
  \Pointer_CTf'_t  lizzieLet20_1_4QVal_Bool_6QVal_Bool_2MyTrue_1_argbuf_d;
  logic lizzieLet20_1_4QVal_Bool_6QVal_Bool_2MyTrue_1_argbuf_r;
  MyBool_t lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_d;
  logic lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_r;
  MyBool_t _32_d;
  logic _32_r;
  assign _32_r = 1'd1;
  MyBool_t lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1_d;
  logic lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1_r;
  MyBool_t lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_2_d;
  logic lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_2_r;
  Go_t lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_d;
  logic lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_r;
  Go_t lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_d;
  logic lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_r;
  Go_t lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1_d;
  logic lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1_r;
  Go_t lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_d;
  logic lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_r;
  QTree_Bool_t lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_d;
  logic lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_r;
  QTree_Bool_t lizzieLet22_1_1_argbuf_d;
  logic lizzieLet22_1_1_argbuf_r;
  Go_t lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_argbuf_d;
  logic lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_argbuf_r;
  Go_t lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_d;
  logic lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_r;
  Go_t lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_d;
  logic lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_r;
  Go_t lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_argbuf_d;
  logic lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_argbuf_r;
  TupGo_t \lvlrcX-0TupGo_1_d ;
  logic \lvlrcX-0TupGo_1_r ;
  Go_t lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_argbuf_d;
  logic lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_argbuf_r;
  \Pointer_CTf'_t  lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_2MyFalse_d;
  logic lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_2MyFalse_r;
  \Pointer_CTf'_t  lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_2MyTrue_d;
  logic lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_2MyTrue_r;
  \Pointer_CTf'_t  lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_2MyFalse_1_argbuf_d;
  logic lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_2MyFalse_1_argbuf_r;
  \Pointer_CTf'_t  lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_2MyTrue_1_argbuf_d;
  logic lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_2MyTrue_1_argbuf_r;
  Pointer_QTree_Bool_t _31_d;
  logic _31_r;
  assign _31_r = 1'd1;
  Pointer_QTree_Bool_t lizzieLet20_1_5QVal_Bool_d;
  logic lizzieLet20_1_5QVal_Bool_r;
  Pointer_QTree_Bool_t lizzieLet20_1_5QNode_Bool_d;
  logic lizzieLet20_1_5QNode_Bool_r;
  Pointer_QTree_Bool_t _30_d;
  logic _30_r;
  assign _30_r = 1'd1;
  Pointer_QTree_Bool_t lizzieLet20_1_6QNone_Bool_d;
  logic lizzieLet20_1_6QNone_Bool_r;
  Pointer_QTree_Bool_t _29_d;
  logic _29_r;
  assign _29_r = 1'd1;
  Pointer_QTree_Bool_t _28_d;
  logic _28_r;
  assign _28_r = 1'd1;
  Pointer_QTree_Bool_t _27_d;
  logic _27_r;
  assign _27_r = 1'd1;
  Pointer_QTree_Bool_t lizzieLet20_1_6QNone_Bool_1_argbuf_d;
  logic lizzieLet20_1_6QNone_Bool_1_argbuf_r;
  \Pointer_CTf'_t  lizzieLet20_1_7QNone_Bool_d;
  logic lizzieLet20_1_7QNone_Bool_r;
  \Pointer_CTf'_t  lizzieLet20_1_7QVal_Bool_d;
  logic lizzieLet20_1_7QVal_Bool_r;
  \Pointer_CTf'_t  lizzieLet20_1_7QNode_Bool_d;
  logic lizzieLet20_1_7QNode_Bool_r;
  \Pointer_CTf'_t  lizzieLet20_1_7QError_Bool_d;
  logic lizzieLet20_1_7QError_Bool_r;
  \Pointer_CTf'_t  lizzieLet20_1_7QError_Bool_1_argbuf_d;
  logic lizzieLet20_1_7QError_Bool_1_argbuf_r;
  \Pointer_CTf'_t  lizzieLet20_1_7QNone_Bool_1_argbuf_d;
  logic lizzieLet20_1_7QNone_Bool_1_argbuf_r;
  Pointer_MaskQTree_t q1a8y_destruct_d;
  logic q1a8y_destruct_r;
  Pointer_MaskQTree_t q2a8z_destruct_d;
  logic q2a8z_destruct_r;
  Pointer_MaskQTree_t q3a8A_destruct_d;
  logic q3a8A_destruct_r;
  Pointer_MaskQTree_t q5a8B_destruct_d;
  logic q5a8B_destruct_r;
  MaskQTree_t _26_d;
  logic _26_r;
  assign _26_r = 1'd1;
  MaskQTree_t _25_d;
  logic _25_r;
  assign _25_r = 1'd1;
  MaskQTree_t lizzieLet32_1MQNode_d;
  logic lizzieLet32_1MQNode_r;
  Go_t lizzieLet32_3MQNone_d;
  logic lizzieLet32_3MQNone_r;
  Go_t lizzieLet32_3MQVal_d;
  logic lizzieLet32_3MQVal_r;
  Go_t lizzieLet32_3MQNode_d;
  logic lizzieLet32_3MQNode_r;
  Go_t lizzieLet32_3MQNone_1_d;
  logic lizzieLet32_3MQNone_1_r;
  Go_t lizzieLet32_3MQNone_2_d;
  logic lizzieLet32_3MQNone_2_r;
  QTree_Bool_t lizzieLet32_3MQNone_1QNone_Bool_d;
  logic lizzieLet32_3MQNone_1QNone_Bool_r;
  QTree_Bool_t lizzieLet33_1_argbuf_d;
  logic lizzieLet33_1_argbuf_r;
  Go_t lizzieLet32_3MQNone_2_argbuf_d;
  logic lizzieLet32_3MQNone_2_argbuf_r;
  C6_t go_11_goMux_choice_d;
  logic go_11_goMux_choice_r;
  Go_t go_11_goMux_data_d;
  logic go_11_goMux_data_r;
  Go_t lizzieLet32_3MQVal_1_argbuf_d;
  logic lizzieLet32_3MQVal_1_argbuf_r;
  QTree_Bool_t _24_d;
  logic _24_r;
  assign _24_r = 1'd1;
  QTree_Bool_t _23_d;
  logic _23_r;
  assign _23_r = 1'd1;
  QTree_Bool_t lizzieLet32_4MQNode_d;
  logic lizzieLet32_4MQNode_r;
  QTree_Bool_t lizzieLet32_4MQNode_1_d;
  logic lizzieLet32_4MQNode_1_r;
  QTree_Bool_t lizzieLet32_4MQNode_2_d;
  logic lizzieLet32_4MQNode_2_r;
  QTree_Bool_t lizzieLet32_4MQNode_3_d;
  logic lizzieLet32_4MQNode_3_r;
  QTree_Bool_t lizzieLet32_4MQNode_4_d;
  logic lizzieLet32_4MQNode_4_r;
  QTree_Bool_t lizzieLet32_4MQNode_5_d;
  logic lizzieLet32_4MQNode_5_r;
  QTree_Bool_t lizzieLet32_4MQNode_6_d;
  logic lizzieLet32_4MQNode_6_r;
  QTree_Bool_t lizzieLet32_4MQNode_7_d;
  logic lizzieLet32_4MQNode_7_r;
  QTree_Bool_t lizzieLet32_4MQNode_8_d;
  logic lizzieLet32_4MQNode_8_r;
  Pointer_QTree_Bool_t t1a8D_destruct_d;
  logic t1a8D_destruct_r;
  Pointer_QTree_Bool_t t2a8E_destruct_d;
  logic t2a8E_destruct_r;
  Pointer_QTree_Bool_t t3a8F_destruct_d;
  logic t3a8F_destruct_r;
  Pointer_QTree_Bool_t t4a8G_destruct_d;
  logic t4a8G_destruct_r;
  QTree_Bool_t _22_d;
  logic _22_r;
  assign _22_r = 1'd1;
  QTree_Bool_t _21_d;
  logic _21_r;
  assign _21_r = 1'd1;
  QTree_Bool_t lizzieLet32_4MQNode_1QNode_Bool_d;
  logic lizzieLet32_4MQNode_1QNode_Bool_r;
  QTree_Bool_t _20_d;
  logic _20_r;
  assign _20_r = 1'd1;
  Go_t lizzieLet32_4MQNode_3QNone_Bool_d;
  logic lizzieLet32_4MQNode_3QNone_Bool_r;
  Go_t lizzieLet32_4MQNode_3QVal_Bool_d;
  logic lizzieLet32_4MQNode_3QVal_Bool_r;
  Go_t lizzieLet32_4MQNode_3QNode_Bool_d;
  logic lizzieLet32_4MQNode_3QNode_Bool_r;
  Go_t lizzieLet32_4MQNode_3QError_Bool_d;
  logic lizzieLet32_4MQNode_3QError_Bool_r;
  Go_t lizzieLet32_4MQNode_3QError_Bool_1_d;
  logic lizzieLet32_4MQNode_3QError_Bool_1_r;
  Go_t lizzieLet32_4MQNode_3QError_Bool_2_d;
  logic lizzieLet32_4MQNode_3QError_Bool_2_r;
  QTree_Bool_t lizzieLet32_4MQNode_3QError_Bool_1QError_Bool_d;
  logic lizzieLet32_4MQNode_3QError_Bool_1QError_Bool_r;
  QTree_Bool_t lizzieLet38_1_argbuf_d;
  logic lizzieLet38_1_argbuf_r;
  Go_t lizzieLet32_4MQNode_3QError_Bool_2_argbuf_d;
  logic lizzieLet32_4MQNode_3QError_Bool_2_argbuf_r;
  Go_t lizzieLet32_4MQNode_3QNode_Bool_1_argbuf_d;
  logic lizzieLet32_4MQNode_3QNode_Bool_1_argbuf_r;
  Go_t lizzieLet32_4MQNode_3QNone_Bool_1_d;
  logic lizzieLet32_4MQNode_3QNone_Bool_1_r;
  Go_t lizzieLet32_4MQNode_3QNone_Bool_2_d;
  logic lizzieLet32_4MQNode_3QNone_Bool_2_r;
  QTree_Bool_t lizzieLet32_4MQNode_3QNone_Bool_1QNone_Bool_d;
  logic lizzieLet32_4MQNode_3QNone_Bool_1QNone_Bool_r;
  QTree_Bool_t lizzieLet35_1_argbuf_d;
  logic lizzieLet35_1_argbuf_r;
  Go_t lizzieLet32_4MQNode_3QNone_Bool_2_argbuf_d;
  logic lizzieLet32_4MQNode_3QNone_Bool_2_argbuf_r;
  Go_t lizzieLet32_4MQNode_3QVal_Bool_1_d;
  logic lizzieLet32_4MQNode_3QVal_Bool_1_r;
  Go_t lizzieLet32_4MQNode_3QVal_Bool_2_d;
  logic lizzieLet32_4MQNode_3QVal_Bool_2_r;
  QTree_Bool_t lizzieLet32_4MQNode_3QVal_Bool_1QError_Bool_d;
  logic lizzieLet32_4MQNode_3QVal_Bool_1QError_Bool_r;
  QTree_Bool_t lizzieLet36_1_argbuf_d;
  logic lizzieLet36_1_argbuf_r;
  Go_t lizzieLet32_4MQNode_3QVal_Bool_2_argbuf_d;
  logic lizzieLet32_4MQNode_3QVal_Bool_2_argbuf_r;
  \Pointer_CTf'''''''''_f'''''''''_Bool_t  lizzieLet32_4MQNode_4QNone_Bool_d;
  logic lizzieLet32_4MQNode_4QNone_Bool_r;
  \Pointer_CTf'''''''''_f'''''''''_Bool_t  lizzieLet32_4MQNode_4QVal_Bool_d;
  logic lizzieLet32_4MQNode_4QVal_Bool_r;
  \Pointer_CTf'''''''''_f'''''''''_Bool_t  lizzieLet32_4MQNode_4QNode_Bool_d;
  logic lizzieLet32_4MQNode_4QNode_Bool_r;
  \Pointer_CTf'''''''''_f'''''''''_Bool_t  lizzieLet32_4MQNode_4QError_Bool_d;
  logic lizzieLet32_4MQNode_4QError_Bool_r;
  \Pointer_CTf'''''''''_f'''''''''_Bool_t  lizzieLet32_4MQNode_4QError_Bool_1_argbuf_d;
  logic lizzieLet32_4MQNode_4QError_Bool_1_argbuf_r;
  \CTf'''''''''_f'''''''''_Bool_t  \lizzieLet32_4MQNode_4QNode_Bool_1lizzieLet32_4MQNode_5QNode_Bool_1t1a8D_1lizzieLet32_4MQNode_6QNode_Bool_1t2a8E_1lizzieLet32_4MQNode_7QNode_Bool_1t3a8F_1Lcall_f'''''''''_f'''''''''_Bool3_d ;
  logic \lizzieLet32_4MQNode_4QNode_Bool_1lizzieLet32_4MQNode_5QNode_Bool_1t1a8D_1lizzieLet32_4MQNode_6QNode_Bool_1t2a8E_1lizzieLet32_4MQNode_7QNode_Bool_1t3a8F_1Lcall_f'''''''''_f'''''''''_Bool3_r ;
  \CTf'''''''''_f'''''''''_Bool_t  lizzieLet37_1_argbuf_d;
  logic lizzieLet37_1_argbuf_r;
  \Pointer_CTf'''''''''_f'''''''''_Bool_t  lizzieLet32_4MQNode_4QNone_Bool_1_argbuf_d;
  logic lizzieLet32_4MQNode_4QNone_Bool_1_argbuf_r;
  \Pointer_CTf'''''''''_f'''''''''_Bool_t  lizzieLet32_4MQNode_4QVal_Bool_1_argbuf_d;
  logic lizzieLet32_4MQNode_4QVal_Bool_1_argbuf_r;
  Pointer_MaskQTree_t _19_d;
  logic _19_r;
  assign _19_r = 1'd1;
  Pointer_MaskQTree_t _18_d;
  logic _18_r;
  assign _18_r = 1'd1;
  Pointer_MaskQTree_t lizzieLet32_4MQNode_5QNode_Bool_d;
  logic lizzieLet32_4MQNode_5QNode_Bool_r;
  Pointer_MaskQTree_t _17_d;
  logic _17_r;
  assign _17_r = 1'd1;
  Pointer_MaskQTree_t _16_d;
  logic _16_r;
  assign _16_r = 1'd1;
  Pointer_MaskQTree_t _15_d;
  logic _15_r;
  assign _15_r = 1'd1;
  Pointer_MaskQTree_t lizzieLet32_4MQNode_6QNode_Bool_d;
  logic lizzieLet32_4MQNode_6QNode_Bool_r;
  Pointer_MaskQTree_t _14_d;
  logic _14_r;
  assign _14_r = 1'd1;
  Pointer_MaskQTree_t _13_d;
  logic _13_r;
  assign _13_r = 1'd1;
  Pointer_MaskQTree_t _12_d;
  logic _12_r;
  assign _12_r = 1'd1;
  Pointer_MaskQTree_t lizzieLet32_4MQNode_7QNode_Bool_d;
  logic lizzieLet32_4MQNode_7QNode_Bool_r;
  Pointer_MaskQTree_t _11_d;
  logic _11_r;
  assign _11_r = 1'd1;
  Pointer_MaskQTree_t _10_d;
  logic _10_r;
  assign _10_r = 1'd1;
  Pointer_MaskQTree_t _9_d;
  logic _9_r;
  assign _9_r = 1'd1;
  Pointer_MaskQTree_t lizzieLet32_4MQNode_8QNode_Bool_d;
  logic lizzieLet32_4MQNode_8QNode_Bool_r;
  Pointer_MaskQTree_t _8_d;
  logic _8_r;
  assign _8_r = 1'd1;
  Pointer_MaskQTree_t lizzieLet32_4MQNode_8QNode_Bool_1_argbuf_d;
  logic lizzieLet32_4MQNode_8QNode_Bool_1_argbuf_r;
  Pointer_QTree_Bool_t _7_d;
  logic _7_r;
  assign _7_r = 1'd1;
  Pointer_QTree_Bool_t lizzieLet32_5MQVal_d;
  logic lizzieLet32_5MQVal_r;
  Pointer_QTree_Bool_t _6_d;
  logic _6_r;
  assign _6_r = 1'd1;
  Pointer_QTree_Bool_t lizzieLet32_5MQVal_1_argbuf_d;
  logic lizzieLet32_5MQVal_1_argbuf_r;
  \Pointer_CTf'''''''''_f'''''''''_Bool_t  lizzieLet32_6MQNone_d;
  logic lizzieLet32_6MQNone_r;
  \Pointer_CTf'''''''''_f'''''''''_Bool_t  lizzieLet32_6MQVal_d;
  logic lizzieLet32_6MQVal_r;
  \Pointer_CTf'''''''''_f'''''''''_Bool_t  lizzieLet32_6MQNode_d;
  logic lizzieLet32_6MQNode_r;
  \Pointer_CTf'''''''''_f'''''''''_Bool_t  lizzieLet32_6MQNone_1_argbuf_d;
  logic lizzieLet32_6MQNone_1_argbuf_r;
  \Pointer_CTf'''''''''_f'''''''''_Bool_t  lizzieLet32_6MQVal_1_argbuf_d;
  logic lizzieLet32_6MQVal_1_argbuf_r;
  Pointer_QTree_Bool_t es_9_destruct_d;
  logic es_9_destruct_r;
  Pointer_QTree_Bool_t es_10_1_destruct_d;
  logic es_10_1_destruct_r;
  Pointer_QTree_Bool_t es_11_2_destruct_d;
  logic es_11_2_destruct_r;
  Pointer_CTf_t sc_0_6_destruct_d;
  logic sc_0_6_destruct_r;
  Pointer_QTree_Bool_t es_10_destruct_d;
  logic es_10_destruct_r;
  Pointer_QTree_Bool_t es_11_1_destruct_d;
  logic es_11_1_destruct_r;
  Pointer_CTf_t sc_0_5_destruct_d;
  logic sc_0_5_destruct_r;
  Pointer_MaskQTree_t q1a88_3_destruct_d;
  logic q1a88_3_destruct_r;
  Pointer_QTree_Bool_t \q1'a8n_3_destruct_d ;
  logic \q1'a8n_3_destruct_r ;
  Pointer_QTree_Bool_t t1a8s_3_destruct_d;
  logic t1a8s_3_destruct_r;
  Pointer_QTree_Bool_t es_11_destruct_d;
  logic es_11_destruct_r;
  Pointer_CTf_t sc_0_4_destruct_d;
  logic sc_0_4_destruct_r;
  Pointer_MaskQTree_t q1a88_2_destruct_d;
  logic q1a88_2_destruct_r;
  Pointer_QTree_Bool_t \q1'a8n_2_destruct_d ;
  logic \q1'a8n_2_destruct_r ;
  Pointer_QTree_Bool_t t1a8s_2_destruct_d;
  logic t1a8s_2_destruct_r;
  Pointer_MaskQTree_t q2a89_2_destruct_d;
  logic q2a89_2_destruct_r;
  Pointer_QTree_Bool_t \q2'a8o_2_destruct_d ;
  logic \q2'a8o_2_destruct_r ;
  Pointer_QTree_Bool_t t2a8t_2_destruct_d;
  logic t2a8t_2_destruct_r;
  Pointer_CTf_t sc_0_3_destruct_d;
  logic sc_0_3_destruct_r;
  Pointer_MaskQTree_t q1a88_1_destruct_d;
  logic q1a88_1_destruct_r;
  Pointer_QTree_Bool_t \q1'a8n_1_destruct_d ;
  logic \q1'a8n_1_destruct_r ;
  Pointer_QTree_Bool_t t1a8s_1_destruct_d;
  logic t1a8s_1_destruct_r;
  Pointer_MaskQTree_t q2a89_1_destruct_d;
  logic q2a89_1_destruct_r;
  Pointer_QTree_Bool_t \q2'a8o_1_destruct_d ;
  logic \q2'a8o_1_destruct_r ;
  Pointer_QTree_Bool_t t2a8t_1_destruct_d;
  logic t2a8t_1_destruct_r;
  Pointer_MaskQTree_t q3a8a_1_destruct_d;
  logic q3a8a_1_destruct_r;
  Pointer_QTree_Bool_t \q3'a8p_1_destruct_d ;
  logic \q3'a8p_1_destruct_r ;
  Pointer_QTree_Bool_t t3a8u_1_destruct_d;
  logic t3a8u_1_destruct_r;
  CTf_t _5_d;
  logic _5_r;
  assign _5_r = 1'd1;
  CTf_t lizzieLet43_1Lcall_f3_d;
  logic lizzieLet43_1Lcall_f3_r;
  CTf_t lizzieLet43_1Lcall_f2_d;
  logic lizzieLet43_1Lcall_f2_r;
  CTf_t lizzieLet43_1Lcall_f1_d;
  logic lizzieLet43_1Lcall_f1_r;
  CTf_t lizzieLet43_1Lcall_f0_d;
  logic lizzieLet43_1Lcall_f0_r;
  Go_t _4_d;
  logic _4_r;
  assign _4_r = 1'd1;
  Go_t lizzieLet43_3Lcall_f3_d;
  logic lizzieLet43_3Lcall_f3_r;
  Go_t lizzieLet43_3Lcall_f2_d;
  logic lizzieLet43_3Lcall_f2_r;
  Go_t lizzieLet43_3Lcall_f1_d;
  logic lizzieLet43_3Lcall_f1_r;
  Go_t lizzieLet43_3Lcall_f0_d;
  logic lizzieLet43_3Lcall_f0_r;
  Go_t lizzieLet43_3Lcall_f0_1_argbuf_d;
  logic lizzieLet43_3Lcall_f0_1_argbuf_r;
  Go_t lizzieLet43_3Lcall_f1_1_argbuf_d;
  logic lizzieLet43_3Lcall_f1_1_argbuf_r;
  Go_t lizzieLet43_3Lcall_f2_1_argbuf_d;
  logic lizzieLet43_3Lcall_f2_1_argbuf_r;
  Go_t lizzieLet43_3Lcall_f3_1_argbuf_d;
  logic lizzieLet43_3Lcall_f3_1_argbuf_r;
  Pointer_QTree_Bool_t lizzieLet43_4Lfsbos_d;
  logic lizzieLet43_4Lfsbos_r;
  Pointer_QTree_Bool_t lizzieLet43_4Lcall_f3_d;
  logic lizzieLet43_4Lcall_f3_r;
  Pointer_QTree_Bool_t lizzieLet43_4Lcall_f2_d;
  logic lizzieLet43_4Lcall_f2_r;
  Pointer_QTree_Bool_t lizzieLet43_4Lcall_f1_d;
  logic lizzieLet43_4Lcall_f1_r;
  Pointer_QTree_Bool_t lizzieLet43_4Lcall_f0_d;
  logic lizzieLet43_4Lcall_f0_r;
  QTree_Bool_t lizzieLet43_4Lcall_f0_1es_9_1es_10_1_1es_11_2_1QNode_Bool_d;
  logic lizzieLet43_4Lcall_f0_1es_9_1es_10_1_1es_11_2_1QNode_Bool_r;
  QTree_Bool_t lizzieLet47_1_argbuf_d;
  logic lizzieLet47_1_argbuf_r;
  CTf_t lizzieLet43_4Lcall_f1_1es_10_1es_11_1_1sc_0_5_1Lcall_f0_d;
  logic lizzieLet43_4Lcall_f1_1es_10_1es_11_1_1sc_0_5_1Lcall_f0_r;
  CTf_t lizzieLet46_1_argbuf_d;
  logic lizzieLet46_1_argbuf_r;
  CTf_t \lizzieLet43_4Lcall_f2_1es_11_1sc_0_4_1q1a88_2_1q1'a8n_2_1t1a8s_2_1Lcall_f1_d ;
  logic \lizzieLet43_4Lcall_f2_1es_11_1sc_0_4_1q1a88_2_1q1'a8n_2_1t1a8s_2_1Lcall_f1_r ;
  CTf_t lizzieLet45_1_argbuf_d;
  logic lizzieLet45_1_argbuf_r;
  CTf_t \lizzieLet43_4Lcall_f3_1sc_0_3_1q1a88_1_1q1'a8n_1_1t1a8s_1_1q2a89_1_1q2'a8o_1_1t2a8t_1_1Lcall_f2_d ;
  logic \lizzieLet43_4Lcall_f3_1sc_0_3_1q1a88_1_1q1'a8n_1_1t1a8s_1_1q2a89_1_1q2'a8o_1_1t2a8t_1_1Lcall_f2_r ;
  CTf_t lizzieLet44_1_argbuf_d;
  logic lizzieLet44_1_argbuf_r;
  Pointer_QTree_Bool_t lizzieLet43_4Lfsbos_1_merge_merge_fork_1_d;
  logic lizzieLet43_4Lfsbos_1_merge_merge_fork_1_r;
  Pointer_QTree_Bool_t lizzieLet43_4Lfsbos_1_merge_merge_fork_2_d;
  logic lizzieLet43_4Lfsbos_1_merge_merge_fork_2_r;
  Go_t call_f_goConst_d;
  logic call_f_goConst_r;
  Pointer_QTree_Bool_t f_resbuf_d;
  logic f_resbuf_r;
  Pointer_QTree_Bool_t es_1_1_destruct_d;
  logic es_1_1_destruct_r;
  Pointer_QTree_Bool_t es_2_2_destruct_d;
  logic es_2_2_destruct_r;
  Pointer_QTree_Bool_t es_3_3_destruct_d;
  logic es_3_3_destruct_r;
  \Pointer_CTf'_t  sc_0_10_destruct_d;
  logic sc_0_10_destruct_r;
  Pointer_QTree_Bool_t es_2_1_destruct_d;
  logic es_2_1_destruct_r;
  Pointer_QTree_Bool_t es_3_2_destruct_d;
  logic es_3_2_destruct_r;
  \Pointer_CTf'_t  sc_0_9_destruct_d;
  logic sc_0_9_destruct_r;
  Pointer_QTree_Bool_t q1a8P_3_destruct_d;
  logic q1a8P_3_destruct_r;
  Pointer_QTree_Bool_t t1a8U_3_destruct_d;
  logic t1a8U_3_destruct_r;
  Pointer_QTree_Bool_t es_3_1_destruct_d;
  logic es_3_1_destruct_r;
  \Pointer_CTf'_t  sc_0_8_destruct_d;
  logic sc_0_8_destruct_r;
  Pointer_QTree_Bool_t q1a8P_2_destruct_d;
  logic q1a8P_2_destruct_r;
  Pointer_QTree_Bool_t t1a8U_2_destruct_d;
  logic t1a8U_2_destruct_r;
  Pointer_QTree_Bool_t q2a8Q_2_destruct_d;
  logic q2a8Q_2_destruct_r;
  Pointer_QTree_Bool_t t2a8V_2_destruct_d;
  logic t2a8V_2_destruct_r;
  \Pointer_CTf'_t  sc_0_7_destruct_d;
  logic sc_0_7_destruct_r;
  Pointer_QTree_Bool_t q1a8P_1_destruct_d;
  logic q1a8P_1_destruct_r;
  Pointer_QTree_Bool_t t1a8U_1_destruct_d;
  logic t1a8U_1_destruct_r;
  Pointer_QTree_Bool_t q2a8Q_1_destruct_d;
  logic q2a8Q_1_destruct_r;
  Pointer_QTree_Bool_t t2a8V_1_destruct_d;
  logic t2a8V_1_destruct_r;
  Pointer_QTree_Bool_t q3a8R_1_destruct_d;
  logic q3a8R_1_destruct_r;
  Pointer_QTree_Bool_t t3a8W_1_destruct_d;
  logic t3a8W_1_destruct_r;
  \CTf'_t  _3_d;
  logic _3_r;
  assign _3_r = 1'd1;
  \CTf'_t  \lizzieLet48_1Lcall_f'3_d ;
  logic \lizzieLet48_1Lcall_f'3_r ;
  \CTf'_t  \lizzieLet48_1Lcall_f'2_d ;
  logic \lizzieLet48_1Lcall_f'2_r ;
  \CTf'_t  \lizzieLet48_1Lcall_f'1_d ;
  logic \lizzieLet48_1Lcall_f'1_r ;
  \CTf'_t  \lizzieLet48_1Lcall_f'0_d ;
  logic \lizzieLet48_1Lcall_f'0_r ;
  Go_t _2_d;
  logic _2_r;
  assign _2_r = 1'd1;
  Go_t \lizzieLet48_3Lcall_f'3_d ;
  logic \lizzieLet48_3Lcall_f'3_r ;
  Go_t \lizzieLet48_3Lcall_f'2_d ;
  logic \lizzieLet48_3Lcall_f'2_r ;
  Go_t \lizzieLet48_3Lcall_f'1_d ;
  logic \lizzieLet48_3Lcall_f'1_r ;
  Go_t \lizzieLet48_3Lcall_f'0_d ;
  logic \lizzieLet48_3Lcall_f'0_r ;
  Go_t \lizzieLet48_3Lcall_f'0_1_argbuf_d ;
  logic \lizzieLet48_3Lcall_f'0_1_argbuf_r ;
  Go_t \lizzieLet48_3Lcall_f'1_1_argbuf_d ;
  logic \lizzieLet48_3Lcall_f'1_1_argbuf_r ;
  Go_t \lizzieLet48_3Lcall_f'2_1_argbuf_d ;
  logic \lizzieLet48_3Lcall_f'2_1_argbuf_r ;
  Go_t \lizzieLet48_3Lcall_f'3_1_argbuf_d ;
  logic \lizzieLet48_3Lcall_f'3_1_argbuf_r ;
  Pointer_QTree_Bool_t \lizzieLet48_4Lf'sbos_d ;
  logic \lizzieLet48_4Lf'sbos_r ;
  Pointer_QTree_Bool_t \lizzieLet48_4Lcall_f'3_d ;
  logic \lizzieLet48_4Lcall_f'3_r ;
  Pointer_QTree_Bool_t \lizzieLet48_4Lcall_f'2_d ;
  logic \lizzieLet48_4Lcall_f'2_r ;
  Pointer_QTree_Bool_t \lizzieLet48_4Lcall_f'1_d ;
  logic \lizzieLet48_4Lcall_f'1_r ;
  Pointer_QTree_Bool_t \lizzieLet48_4Lcall_f'0_d ;
  logic \lizzieLet48_4Lcall_f'0_r ;
  QTree_Bool_t \lizzieLet48_4Lcall_f'0_1es_1_1_1es_2_2_1es_3_3_1QNode_Bool_d ;
  logic \lizzieLet48_4Lcall_f'0_1es_1_1_1es_2_2_1es_3_3_1QNode_Bool_r ;
  QTree_Bool_t lizzieLet52_1_argbuf_d;
  logic lizzieLet52_1_argbuf_r;
  \CTf'_t  \lizzieLet48_4Lcall_f'1_1es_2_1_1es_3_2_1sc_0_9_1Lcall_f'0_d ;
  logic \lizzieLet48_4Lcall_f'1_1es_2_1_1es_3_2_1sc_0_9_1Lcall_f'0_r ;
  \CTf'_t  lizzieLet51_1_argbuf_d;
  logic lizzieLet51_1_argbuf_r;
  \CTf'_t  \lizzieLet48_4Lcall_f'2_1es_3_1_1sc_0_8_1q1a8P_2_1t1a8U_2_1Lcall_f'1_d ;
  logic \lizzieLet48_4Lcall_f'2_1es_3_1_1sc_0_8_1q1a8P_2_1t1a8U_2_1Lcall_f'1_r ;
  \CTf'_t  lizzieLet50_1_argbuf_d;
  logic lizzieLet50_1_argbuf_r;
  \CTf'_t  \lizzieLet48_4Lcall_f'3_1sc_0_7_1q1a8P_1_1t1a8U_1_1q2a8Q_1_1t2a8V_1_1Lcall_f'2_d ;
  logic \lizzieLet48_4Lcall_f'3_1sc_0_7_1q1a8P_1_1t1a8U_1_1q2a8Q_1_1t2a8V_1_1Lcall_f'2_r ;
  \CTf'_t  lizzieLet49_1_argbuf_d;
  logic lizzieLet49_1_argbuf_r;
  Pointer_QTree_Bool_t \lizzieLet48_4Lf'sbos_1_merge_merge_fork_1_d ;
  logic \lizzieLet48_4Lf'sbos_1_merge_merge_fork_1_r ;
  Pointer_QTree_Bool_t \lizzieLet48_4Lf'sbos_1_merge_merge_fork_2_d ;
  logic \lizzieLet48_4Lf'sbos_1_merge_merge_fork_2_r ;
  Go_t \call_f'_goConst_d ;
  logic \call_f'_goConst_r ;
  Pointer_QTree_Bool_t \f'_resbuf_d ;
  logic \f'_resbuf_r ;
  Pointer_QTree_Bool_t es_1_2_destruct_d;
  logic es_1_2_destruct_r;
  Pointer_QTree_Bool_t es_2_4_destruct_d;
  logic es_2_4_destruct_r;
  Pointer_QTree_Bool_t es_3_6_destruct_d;
  logic es_3_6_destruct_r;
  \Pointer_CTf'''''''''_f'''''''''_Bool_t  sc_0_14_destruct_d;
  logic sc_0_14_destruct_r;
  Pointer_QTree_Bool_t es_2_3_destruct_d;
  logic es_2_3_destruct_r;
  Pointer_QTree_Bool_t es_3_5_destruct_d;
  logic es_3_5_destruct_r;
  \Pointer_CTf'''''''''_f'''''''''_Bool_t  sc_0_13_destruct_d;
  logic sc_0_13_destruct_r;
  Pointer_MaskQTree_t q1a8y_3_destruct_d;
  logic q1a8y_3_destruct_r;
  Pointer_QTree_Bool_t t1a8D_3_destruct_d;
  logic t1a8D_3_destruct_r;
  Pointer_QTree_Bool_t es_3_4_destruct_d;
  logic es_3_4_destruct_r;
  \Pointer_CTf'''''''''_f'''''''''_Bool_t  sc_0_12_destruct_d;
  logic sc_0_12_destruct_r;
  Pointer_MaskQTree_t q1a8y_2_destruct_d;
  logic q1a8y_2_destruct_r;
  Pointer_QTree_Bool_t t1a8D_2_destruct_d;
  logic t1a8D_2_destruct_r;
  Pointer_MaskQTree_t q2a8z_2_destruct_d;
  logic q2a8z_2_destruct_r;
  Pointer_QTree_Bool_t t2a8E_2_destruct_d;
  logic t2a8E_2_destruct_r;
  \Pointer_CTf'''''''''_f'''''''''_Bool_t  sc_0_11_destruct_d;
  logic sc_0_11_destruct_r;
  Pointer_MaskQTree_t q1a8y_1_destruct_d;
  logic q1a8y_1_destruct_r;
  Pointer_QTree_Bool_t t1a8D_1_destruct_d;
  logic t1a8D_1_destruct_r;
  Pointer_MaskQTree_t q2a8z_1_destruct_d;
  logic q2a8z_1_destruct_r;
  Pointer_QTree_Bool_t t2a8E_1_destruct_d;
  logic t2a8E_1_destruct_r;
  Pointer_MaskQTree_t q3a8A_1_destruct_d;
  logic q3a8A_1_destruct_r;
  Pointer_QTree_Bool_t t3a8F_1_destruct_d;
  logic t3a8F_1_destruct_r;
  \CTf'''''''''_f'''''''''_Bool_t  _1_d;
  logic _1_r;
  assign _1_r = 1'd1;
  \CTf'''''''''_f'''''''''_Bool_t  \lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool3_d ;
  logic \lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool3_r ;
  \CTf'''''''''_f'''''''''_Bool_t  \lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool2_d ;
  logic \lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool2_r ;
  \CTf'''''''''_f'''''''''_Bool_t  \lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool1_d ;
  logic \lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool1_r ;
  \CTf'''''''''_f'''''''''_Bool_t  \lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool0_d ;
  logic \lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool0_r ;
  Go_t _0_d;
  logic _0_r;
  assign _0_r = 1'd1;
  Go_t \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool3_d ;
  logic \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool3_r ;
  Go_t \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool2_d ;
  logic \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool2_r ;
  Go_t \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool1_d ;
  logic \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool1_r ;
  Go_t \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool0_d ;
  logic \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool0_r ;
  Go_t \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool0_1_argbuf_d ;
  logic \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool0_1_argbuf_r ;
  Go_t \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool1_1_argbuf_d ;
  logic \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool1_1_argbuf_r ;
  Go_t \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool2_1_argbuf_d ;
  logic \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool2_1_argbuf_r ;
  Go_t \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool3_1_argbuf_d ;
  logic \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool3_1_argbuf_r ;
  Pointer_QTree_Bool_t \lizzieLet53_4Lf'''''''''_f'''''''''_Boolsbos_d ;
  logic \lizzieLet53_4Lf'''''''''_f'''''''''_Boolsbos_r ;
  Pointer_QTree_Bool_t \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool3_d ;
  logic \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool3_r ;
  Pointer_QTree_Bool_t \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool2_d ;
  logic \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool2_r ;
  Pointer_QTree_Bool_t \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool1_d ;
  logic \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool1_r ;
  Pointer_QTree_Bool_t \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool0_d ;
  logic \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool0_r ;
  QTree_Bool_t \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool0_1es_1_2_1es_2_4_1es_3_6_1QNode_Bool_d ;
  logic \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool0_1es_1_2_1es_2_4_1es_3_6_1QNode_Bool_r ;
  QTree_Bool_t lizzieLet57_1_argbuf_d;
  logic lizzieLet57_1_argbuf_r;
  \CTf'''''''''_f'''''''''_Bool_t  \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool1_1es_2_3_1es_3_5_1sc_0_13_1Lcall_f'''''''''_f'''''''''_Bool0_d ;
  logic \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool1_1es_2_3_1es_3_5_1sc_0_13_1Lcall_f'''''''''_f'''''''''_Bool0_r ;
  \CTf'''''''''_f'''''''''_Bool_t  lizzieLet56_1_argbuf_d;
  logic lizzieLet56_1_argbuf_r;
  \CTf'''''''''_f'''''''''_Bool_t  \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool2_1es_3_4_1sc_0_12_1q1a8y_2_1t1a8D_2_1Lcall_f'''''''''_f'''''''''_Bool1_d ;
  logic \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool2_1es_3_4_1sc_0_12_1q1a8y_2_1t1a8D_2_1Lcall_f'''''''''_f'''''''''_Bool1_r ;
  \CTf'''''''''_f'''''''''_Bool_t  lizzieLet55_1_argbuf_d;
  logic lizzieLet55_1_argbuf_r;
  \CTf'''''''''_f'''''''''_Bool_t  \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool3_1sc_0_11_1q1a8y_1_1t1a8D_1_1q2a8z_1_1t2a8E_1_1Lcall_f'''''''''_f'''''''''_Bool2_d ;
  logic \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool3_1sc_0_11_1q1a8y_1_1t1a8D_1_1q2a8z_1_1t2a8E_1_1Lcall_f'''''''''_f'''''''''_Bool2_r ;
  \CTf'''''''''_f'''''''''_Bool_t  lizzieLet54_1_argbuf_d;
  logic lizzieLet54_1_argbuf_r;
  Pointer_QTree_Bool_t \lizzieLet53_4Lf'''''''''_f'''''''''_Boolsbos_1_merge_merge_fork_1_d ;
  logic \lizzieLet53_4Lf'''''''''_f'''''''''_Boolsbos_1_merge_merge_fork_1_r ;
  Pointer_QTree_Bool_t \lizzieLet53_4Lf'''''''''_f'''''''''_Boolsbos_1_merge_merge_fork_2_d ;
  logic \lizzieLet53_4Lf'''''''''_f'''''''''_Boolsbos_1_merge_merge_fork_2_r ;
  Go_t \call_f'''''''''_f'''''''''_Bool_goConst_d ;
  logic \call_f'''''''''_f'''''''''_Bool_goConst_r ;
  C2_t \lvlrcX-0_choice_d ;
  logic \lvlrcX-0_choice_r ;
  TupGo_t \lvlrcX-0_data_d ;
  logic \lvlrcX-0_data_r ;
  MyBool_t go_8_1MyTrue_d;
  logic go_8_1MyTrue_r;
  Pointer_QTree_Bool_t \lvlrcX-0_resbuf_d ;
  logic \lvlrcX-0_resbuf_r ;
  Pointer_QTree_Bool_t \lvlrcX-0_2_argbuf_d ;
  logic \lvlrcX-0_2_argbuf_r ;
  Pointer_QTree_Bool_t lizzieLet24_1_1_argbuf_d;
  logic lizzieLet24_1_1_argbuf_r;
  Pointer_QTree_Bool_t \lvlrcX-0_1_d ;
  logic \lvlrcX-0_1_r ;
  Pointer_QTree_Bool_t \lvlrcX-0_2_d ;
  logic \lvlrcX-0_2_r ;
  Go_t \lvlrcX-0TupGogo_8_d ;
  logic \lvlrcX-0TupGogo_8_r ;
  Pointer_QTree_Bool_t lizzieLet23_1_1_argbuf_d;
  logic lizzieLet23_1_1_argbuf_r;
  Pointer_MaskQTree_t m1a85_1_argbuf_d;
  logic m1a85_1_argbuf_r;
  Pointer_QTree_Bool_t m2a86_1_argbuf_d;
  logic m2a86_1_argbuf_r;
  Pointer_QTree_Bool_t m2a86_1_d;
  logic m2a86_1_r;
  Pointer_QTree_Bool_t m2a86_2_d;
  logic m2a86_2_r;
  Pointer_QTree_Bool_t m2a8H_1_argbuf_d;
  logic m2a8H_1_argbuf_r;
  Pointer_QTree_Bool_t m2a8H_1_d;
  logic m2a8H_1_r;
  Pointer_QTree_Bool_t m2a8H_2_d;
  logic m2a8H_2_r;
  Pointer_QTree_Bool_t m3a87_1_argbuf_d;
  logic m3a87_1_argbuf_r;
  Pointer_QTree_Bool_t m3a87_1_d;
  logic m3a87_1_r;
  Pointer_QTree_Bool_t m3a87_2_d;
  logic m3a87_2_r;
  Pointer_QTree_Bool_t m3a8I_1_argbuf_d;
  logic m3a8I_1_argbuf_r;
  Pointer_QTree_Bool_t m3a8I_1_d;
  logic m3a8I_1_r;
  Pointer_QTree_Bool_t m3a8I_2_d;
  logic m3a8I_2_r;
  Pointer_QTree_Bool_t \q1'a8n_3_1_argbuf_d ;
  logic \q1'a8n_3_1_argbuf_r ;
  Pointer_MaskQTree_t q1a88_3_1_argbuf_d;
  logic q1a88_3_1_argbuf_r;
  Pointer_QTree_Bool_t q1a8P_3_1_argbuf_d;
  logic q1a8P_3_1_argbuf_r;
  Pointer_MaskQTree_t q1a8y_3_1_argbuf_d;
  logic q1a8y_3_1_argbuf_r;
  Pointer_QTree_Bool_t \q2'a8o_2_1_argbuf_d ;
  logic \q2'a8o_2_1_argbuf_r ;
  Pointer_MaskQTree_t q2a89_2_1_argbuf_d;
  logic q2a89_2_1_argbuf_r;
  Pointer_QTree_Bool_t q2a8Q_2_1_argbuf_d;
  logic q2a8Q_2_1_argbuf_r;
  Pointer_MaskQTree_t q2a8z_2_1_argbuf_d;
  logic q2a8z_2_1_argbuf_r;
  Pointer_QTree_Bool_t \q3'a8p_1_1_argbuf_d ;
  logic \q3'a8p_1_1_argbuf_r ;
  Pointer_MaskQTree_t q3a8A_1_1_argbuf_d;
  logic q3a8A_1_1_argbuf_r;
  Pointer_QTree_Bool_t q3a8R_1_1_argbuf_d;
  logic q3a8R_1_1_argbuf_r;
  Pointer_MaskQTree_t q3a8a_1_1_argbuf_d;
  logic q3a8a_1_1_argbuf_r;
  Pointer_QTree_Bool_t \q4'a8x_1_argbuf_d ;
  logic \q4'a8x_1_argbuf_r ;
  Pointer_QTree_Bool_t \q4'a8x_1_d ;
  logic \q4'a8x_1_r ;
  Pointer_QTree_Bool_t \q4'a8x_2_d ;
  logic \q4'a8x_2_r ;
  Pointer_MaskQTree_t q4a8w_1_argbuf_d;
  logic q4a8w_1_argbuf_r;
  \CTf'''''''''_f'''''''''_Bool_t  \readPointer_CTf'''''''''_f'''''''''_Boolscfarg_0_2_1_argbuf_rwb_d ;
  logic \readPointer_CTf'''''''''_f'''''''''_Boolscfarg_0_2_1_argbuf_rwb_r ;
  \CTf'''''''''_f'''''''''_Bool_t  lizzieLet53_1_d;
  logic lizzieLet53_1_r;
  \CTf'''''''''_f'''''''''_Bool_t  lizzieLet53_2_d;
  logic lizzieLet53_2_r;
  \CTf'''''''''_f'''''''''_Bool_t  lizzieLet53_3_d;
  logic lizzieLet53_3_r;
  \CTf'''''''''_f'''''''''_Bool_t  lizzieLet53_4_d;
  logic lizzieLet53_4_r;
  \CTf'_t  \readPointer_CTf'scfarg_0_1_1_argbuf_rwb_d ;
  logic \readPointer_CTf'scfarg_0_1_1_argbuf_rwb_r ;
  \CTf'_t  lizzieLet48_1_d;
  logic lizzieLet48_1_r;
  \CTf'_t  lizzieLet48_2_d;
  logic lizzieLet48_2_r;
  \CTf'_t  lizzieLet48_3_d;
  logic lizzieLet48_3_r;
  \CTf'_t  lizzieLet48_4_d;
  logic lizzieLet48_4_r;
  CTf_t readPointer_CTfscfarg_0_1_argbuf_rwb_d;
  logic readPointer_CTfscfarg_0_1_argbuf_rwb_r;
  CTf_t lizzieLet43_1_d;
  logic lizzieLet43_1_r;
  CTf_t lizzieLet43_2_d;
  logic lizzieLet43_2_r;
  CTf_t lizzieLet43_3_d;
  logic lizzieLet43_3_r;
  CTf_t lizzieLet43_4_d;
  logic lizzieLet43_4_r;
  MaskQTree_t readPointer_MaskQTreem1a85_1_argbuf_rwb_d;
  logic readPointer_MaskQTreem1a85_1_argbuf_rwb_r;
  MaskQTree_t lizzieLet0_1_d;
  logic lizzieLet0_1_r;
  MaskQTree_t lizzieLet0_2_d;
  logic lizzieLet0_2_r;
  MaskQTree_t lizzieLet0_3_d;
  logic lizzieLet0_3_r;
  MaskQTree_t lizzieLet0_4_d;
  logic lizzieLet0_4_r;
  MaskQTree_t lizzieLet0_5_d;
  logic lizzieLet0_5_r;
  MaskQTree_t lizzieLet0_6_d;
  logic lizzieLet0_6_r;
  MaskQTree_t lizzieLet0_7_d;
  logic lizzieLet0_7_r;
  MaskQTree_t lizzieLet0_8_d;
  logic lizzieLet0_8_r;
  MaskQTree_t readPointer_MaskQTreeq4a8w_1_argbuf_rwb_d;
  logic readPointer_MaskQTreeq4a8w_1_argbuf_rwb_r;
  MaskQTree_t lizzieLet32_1_d;
  logic lizzieLet32_1_r;
  MaskQTree_t lizzieLet32_2_d;
  logic lizzieLet32_2_r;
  MaskQTree_t lizzieLet32_3_d;
  logic lizzieLet32_3_r;
  MaskQTree_t lizzieLet32_4_d;
  logic lizzieLet32_4_r;
  MaskQTree_t lizzieLet32_5_d;
  logic lizzieLet32_5_r;
  MaskQTree_t lizzieLet32_6_d;
  logic lizzieLet32_6_r;
  QTree_Bool_t readPointer_QTree_Boolm2a86_1_argbuf_rwb_d;
  logic readPointer_QTree_Boolm2a86_1_argbuf_rwb_r;
  QTree_Bool_t readPointer_QTree_Boolm2a8H_1_argbuf_rwb_d;
  logic readPointer_QTree_Boolm2a8H_1_argbuf_rwb_r;
  QTree_Bool_t lizzieLet20_1_1_d;
  logic lizzieLet20_1_1_r;
  QTree_Bool_t lizzieLet20_1_2_d;
  logic lizzieLet20_1_2_r;
  QTree_Bool_t lizzieLet20_1_3_d;
  logic lizzieLet20_1_3_r;
  QTree_Bool_t lizzieLet20_1_4_d;
  logic lizzieLet20_1_4_r;
  QTree_Bool_t lizzieLet20_1_5_d;
  logic lizzieLet20_1_5_r;
  QTree_Bool_t lizzieLet20_1_6_d;
  logic lizzieLet20_1_6_r;
  QTree_Bool_t lizzieLet20_1_7_d;
  logic lizzieLet20_1_7_r;
  QTree_Bool_t readPointer_QTree_Boolm3a87_1_argbuf_rwb_d;
  logic readPointer_QTree_Boolm3a87_1_argbuf_rwb_r;
  QTree_Bool_t readPointer_QTree_Boolm3a8I_1_argbuf_rwb_d;
  logic readPointer_QTree_Boolm3a8I_1_argbuf_rwb_r;
  QTree_Bool_t \readPointer_QTree_Boolq4'a8x_1_argbuf_rwb_d ;
  logic \readPointer_QTree_Boolq4'a8x_1_argbuf_rwb_r ;
  \Pointer_CTf'_t  sc_0_10_1_argbuf_d;
  logic sc_0_10_1_argbuf_r;
  \Pointer_CTf'''''''''_f'''''''''_Bool_t  sc_0_14_1_argbuf_d;
  logic sc_0_14_1_argbuf_r;
  Pointer_CTf_t sc_0_6_1_argbuf_d;
  logic sc_0_6_1_argbuf_r;
  \Pointer_CTf'_t  scfarg_0_1_1_argbuf_d;
  logic scfarg_0_1_1_argbuf_r;
  \Pointer_CTf'''''''''_f'''''''''_Bool_t  scfarg_0_2_1_argbuf_d;
  logic scfarg_0_2_1_argbuf_r;
  Pointer_CTf_t scfarg_0_1_argbuf_d;
  logic scfarg_0_1_argbuf_r;
  Pointer_QTree_Bool_t t1a8D_3_1_argbuf_d;
  logic t1a8D_3_1_argbuf_r;
  Pointer_QTree_Bool_t t1a8U_3_1_argbuf_d;
  logic t1a8U_3_1_argbuf_r;
  Pointer_QTree_Bool_t t1a8d_1_argbuf_d;
  logic t1a8d_1_argbuf_r;
  Pointer_QTree_Bool_t t1a8s_3_1_argbuf_d;
  logic t1a8s_3_1_argbuf_r;
  Pointer_QTree_Bool_t t2a8E_2_1_argbuf_d;
  logic t2a8E_2_1_argbuf_r;
  Pointer_QTree_Bool_t t2a8V_2_1_argbuf_d;
  logic t2a8V_2_1_argbuf_r;
  Pointer_QTree_Bool_t t2a8e_1_argbuf_d;
  logic t2a8e_1_argbuf_r;
  Pointer_QTree_Bool_t t2a8t_2_1_argbuf_d;
  logic t2a8t_2_1_argbuf_r;
  Pointer_QTree_Bool_t t3a8F_1_1_argbuf_d;
  logic t3a8F_1_1_argbuf_r;
  Pointer_QTree_Bool_t t3a8W_1_1_argbuf_d;
  logic t3a8W_1_1_argbuf_r;
  Pointer_QTree_Bool_t t3a8f_1_argbuf_d;
  logic t3a8f_1_argbuf_r;
  Pointer_QTree_Bool_t t3a8u_1_1_argbuf_d;
  logic t3a8u_1_1_argbuf_r;
  Pointer_QTree_Bool_t t4a8G_1_argbuf_d;
  logic t4a8G_1_argbuf_r;
  Pointer_QTree_Bool_t t4a8X_1_argbuf_d;
  logic t4a8X_1_argbuf_r;
  Pointer_QTree_Bool_t t4a8g_1_argbuf_d;
  logic t4a8g_1_argbuf_r;
  Pointer_QTree_Bool_t t4a8v_1_argbuf_d;
  logic t4a8v_1_argbuf_r;
  \Pointer_CTf'''''''''_f'''''''''_Bool_t  \writeCTf'''''''''_f'''''''''_BoollizzieLet37_1_argbuf_rwb_d ;
  logic \writeCTf'''''''''_f'''''''''_BoollizzieLet37_1_argbuf_rwb_r ;
  \Pointer_CTf'''''''''_f'''''''''_Bool_t  sca3_2_1_argbuf_d;
  logic sca3_2_1_argbuf_r;
  \Pointer_CTf'''''''''_f'''''''''_Bool_t  \writeCTf'''''''''_f'''''''''_BoollizzieLet41_1_argbuf_rwb_d ;
  logic \writeCTf'''''''''_f'''''''''_BoollizzieLet41_1_argbuf_rwb_r ;
  \Pointer_CTf'''''''''_f'''''''''_Bool_t  lizzieLet5_1_1_argbuf_d;
  logic lizzieLet5_1_1_argbuf_r;
  \Pointer_CTf'''''''''_f'''''''''_Bool_t  \writeCTf'''''''''_f'''''''''_BoollizzieLet54_1_argbuf_rwb_d ;
  logic \writeCTf'''''''''_f'''''''''_BoollizzieLet54_1_argbuf_rwb_r ;
  \Pointer_CTf'''''''''_f'''''''''_Bool_t  sca2_2_1_argbuf_d;
  logic sca2_2_1_argbuf_r;
  \Pointer_CTf'''''''''_f'''''''''_Bool_t  \writeCTf'''''''''_f'''''''''_BoollizzieLet55_1_argbuf_rwb_d ;
  logic \writeCTf'''''''''_f'''''''''_BoollizzieLet55_1_argbuf_rwb_r ;
  \Pointer_CTf'''''''''_f'''''''''_Bool_t  sca1_2_1_argbuf_d;
  logic sca1_2_1_argbuf_r;
  \Pointer_CTf'''''''''_f'''''''''_Bool_t  \writeCTf'''''''''_f'''''''''_BoollizzieLet56_1_argbuf_rwb_d ;
  logic \writeCTf'''''''''_f'''''''''_BoollizzieLet56_1_argbuf_rwb_r ;
  \Pointer_CTf'''''''''_f'''''''''_Bool_t  sca0_2_1_argbuf_d;
  logic sca0_2_1_argbuf_r;
  \Pointer_CTf'_t  \writeCTf'lizzieLet29_1_argbuf_rwb_d ;
  logic \writeCTf'lizzieLet29_1_argbuf_rwb_r ;
  \Pointer_CTf'_t  sca3_1_1_argbuf_d;
  logic sca3_1_1_argbuf_r;
  \Pointer_CTf'_t  \writeCTf'lizzieLet40_1_argbuf_rwb_d ;
  logic \writeCTf'lizzieLet40_1_argbuf_rwb_r ;
  \Pointer_CTf'_t  lizzieLet12_1_1_argbuf_d;
  logic lizzieLet12_1_1_argbuf_r;
  \Pointer_CTf'_t  \writeCTf'lizzieLet49_1_argbuf_rwb_d ;
  logic \writeCTf'lizzieLet49_1_argbuf_rwb_r ;
  \Pointer_CTf'_t  sca2_1_1_argbuf_d;
  logic sca2_1_1_argbuf_r;
  \Pointer_CTf'_t  \writeCTf'lizzieLet50_1_argbuf_rwb_d ;
  logic \writeCTf'lizzieLet50_1_argbuf_rwb_r ;
  \Pointer_CTf'_t  sca1_1_1_argbuf_d;
  logic sca1_1_1_argbuf_r;
  \Pointer_CTf'_t  \writeCTf'lizzieLet51_1_argbuf_rwb_d ;
  logic \writeCTf'lizzieLet51_1_argbuf_rwb_r ;
  \Pointer_CTf'_t  sca0_1_1_argbuf_d;
  logic sca0_1_1_argbuf_r;
  Pointer_CTf_t writeCTflizzieLet17_1_1_argbuf_rwb_d;
  logic writeCTflizzieLet17_1_1_argbuf_rwb_r;
  Pointer_CTf_t sca3_1_argbuf_d;
  logic sca3_1_argbuf_r;
  Pointer_CTf_t writeCTflizzieLet39_1_argbuf_rwb_d;
  logic writeCTflizzieLet39_1_argbuf_rwb_r;
  Pointer_CTf_t lizzieLet28_1_1_argbuf_d;
  logic lizzieLet28_1_1_argbuf_r;
  Pointer_CTf_t writeCTflizzieLet44_1_argbuf_rwb_d;
  logic writeCTflizzieLet44_1_argbuf_rwb_r;
  Pointer_CTf_t sca2_1_argbuf_d;
  logic sca2_1_argbuf_r;
  Pointer_CTf_t writeCTflizzieLet45_1_argbuf_rwb_d;
  logic writeCTflizzieLet45_1_argbuf_rwb_r;
  Pointer_CTf_t sca1_1_argbuf_d;
  logic sca1_1_argbuf_r;
  Pointer_CTf_t writeCTflizzieLet46_1_argbuf_rwb_d;
  logic writeCTflizzieLet46_1_argbuf_rwb_r;
  Pointer_CTf_t sca0_1_argbuf_d;
  logic sca0_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet10_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet10_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t lizzieLet20_1_argbuf_d;
  logic lizzieLet20_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet11_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet11_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t lizzieLet21_1_argbuf_d;
  logic lizzieLet21_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet12_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet12_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t lizzieLet22_1_argbuf_d;
  logic lizzieLet22_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet13_1_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet13_1_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t lizzieLet23_1_argbuf_d;
  logic lizzieLet23_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet15_1_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet15_1_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t lizzieLet24_1_argbuf_d;
  logic lizzieLet24_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet16_1_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet16_1_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t lizzieLet25_1_argbuf_d;
  logic lizzieLet25_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet18_1_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet18_1_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t lizzieLet26_1_argbuf_d;
  logic lizzieLet26_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet19_2_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet19_2_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t lizzieLet27_1_argbuf_d;
  logic lizzieLet27_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet1_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet1_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t lizzieLet13_1_argbuf_d;
  logic lizzieLet13_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet22_1_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet22_1_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t lizzieLet6_1_1_argbuf_d;
  logic lizzieLet6_1_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet25_1_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet25_1_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t lizzieLet7_1_1_argbuf_d;
  logic lizzieLet7_1_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet26_1_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet26_1_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t lizzieLet8_1_argbuf_d;
  logic lizzieLet8_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet28_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet28_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t lizzieLet9_2_1_argbuf_d;
  logic lizzieLet9_2_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet30_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet30_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t lizzieLet10_1_1_argbuf_d;
  logic lizzieLet10_1_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet31_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet31_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t lizzieLet11_1_1_argbuf_d;
  logic lizzieLet11_1_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet33_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet33_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t lizzieLet1_1_1_argbuf_d;
  logic lizzieLet1_1_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet35_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet35_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t lizzieLet2_1_1_argbuf_d;
  logic lizzieLet2_1_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet36_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet36_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t lizzieLet3_1_1_argbuf_d;
  logic lizzieLet3_1_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet38_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet38_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t lizzieLet4_1_1_argbuf_d;
  logic lizzieLet4_1_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet42_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet42_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet47_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet47_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t contRet_0_1_argbuf_d;
  logic contRet_0_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet4_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet4_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t lizzieLet15_1_argbuf_d;
  logic lizzieLet15_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet52_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet52_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t contRet_0_1_1_argbuf_d;
  logic contRet_0_1_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet57_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet57_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t contRet_0_2_1_argbuf_d;
  logic contRet_0_2_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet5_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet5_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t lizzieLet16_1_argbuf_d;
  logic lizzieLet16_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet6_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet6_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t lizzieLet17_1_argbuf_d;
  logic lizzieLet17_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet7_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet7_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t lizzieLet18_1_argbuf_d;
  logic lizzieLet18_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet9_1_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet9_1_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t lizzieLet19_1_1_argbuf_d;
  logic lizzieLet19_1_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet9_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet9_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t lizzieLet19_1_argbuf_d;
  logic lizzieLet19_1_argbuf_r;
  
  /* fork (Ty Go) : (sourceGo,Go) > [(goFork,Go),
                                (goFor_2,Go),
                                (goFor_3,Go),
                                (goFor_4,Go),
                                (goFor_5,Go),
                                (goFor_6,Go),
                                (goFor_7,Go)] */
  logic [6:0] sourceGo_emitted;
  logic [6:0] sourceGo_done;
  assign goFork_d = (sourceGo_d[0] && (! sourceGo_emitted[0]));
  assign goFor_2_d = (sourceGo_d[0] && (! sourceGo_emitted[1]));
  assign goFor_3_d = (sourceGo_d[0] && (! sourceGo_emitted[2]));
  assign goFor_4_d = (sourceGo_d[0] && (! sourceGo_emitted[3]));
  assign goFor_5_d = (sourceGo_d[0] && (! sourceGo_emitted[4]));
  assign goFor_6_d = (sourceGo_d[0] && (! sourceGo_emitted[5]));
  assign goFor_7_d = (sourceGo_d[0] && (! sourceGo_emitted[6]));
  assign sourceGo_done = (sourceGo_emitted | ({goFor_7_d[0],
                                               goFor_6_d[0],
                                               goFor_5_d[0],
                                               goFor_4_d[0],
                                               goFor_3_d[0],
                                               goFor_2_d[0],
                                               goFork_d[0]} & {goFor_7_r,
                                                               goFor_6_r,
                                                               goFor_5_r,
                                                               goFor_4_r,
                                                               goFor_3_r,
                                                               goFor_2_r,
                                                               goFork_r}));
  assign sourceGo_r = (& sourceGo_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) sourceGo_emitted <= 7'd0;
    else
      sourceGo_emitted <= (sourceGo_r ? 7'd0 :
                           sourceGo_done);
  
  /* const (Ty Word16#,
       Lit 0) : (go_1_dummy_write_QTree_Bool,Go) > (initHP_QTree_Bool,Word16#) */
  assign initHP_QTree_Bool_d = {16'd0,
                                go_1_dummy_write_QTree_Bool_d[0]};
  assign go_1_dummy_write_QTree_Bool_r = initHP_QTree_Bool_r;
  
  /* const (Ty Word16#,
       Lit 1) : (incrHP_QTree_Bool1,Go) > (incrHP_QTree_Bool,Word16#) */
  assign incrHP_QTree_Bool_d = {16'd1, incrHP_QTree_Bool1_d[0]};
  assign incrHP_QTree_Bool1_r = incrHP_QTree_Bool_r;
  
  /* merge (Ty Go) : [(go_2_dummy_write_QTree_Bool,Go),
                 (incrHP_QTree_Bool2,Go)] > (incrHP_mergeQTree_Bool,Go) */
  logic [1:0] incrHP_mergeQTree_Bool_selected;
  logic [1:0] incrHP_mergeQTree_Bool_select;
  always_comb
    begin
      incrHP_mergeQTree_Bool_selected = 2'd0;
      if ((| incrHP_mergeQTree_Bool_select))
        incrHP_mergeQTree_Bool_selected = incrHP_mergeQTree_Bool_select;
      else
        if (go_2_dummy_write_QTree_Bool_d[0])
          incrHP_mergeQTree_Bool_selected[0] = 1'd1;
        else if (incrHP_QTree_Bool2_d[0])
          incrHP_mergeQTree_Bool_selected[1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeQTree_Bool_select <= 2'd0;
    else
      incrHP_mergeQTree_Bool_select <= (incrHP_mergeQTree_Bool_r ? 2'd0 :
                                        incrHP_mergeQTree_Bool_selected);
  always_comb
    if (incrHP_mergeQTree_Bool_selected[0])
      incrHP_mergeQTree_Bool_d = go_2_dummy_write_QTree_Bool_d;
    else if (incrHP_mergeQTree_Bool_selected[1])
      incrHP_mergeQTree_Bool_d = incrHP_QTree_Bool2_d;
    else incrHP_mergeQTree_Bool_d = 1'd0;
  assign {incrHP_QTree_Bool2_r,
          go_2_dummy_write_QTree_Bool_r} = (incrHP_mergeQTree_Bool_r ? incrHP_mergeQTree_Bool_selected :
                                            2'd0);
  
  /* fork (Ty Go) : (incrHP_mergeQTree_Bool_buf,Go) > [(incrHP_QTree_Bool1,Go),
                                                  (incrHP_QTree_Bool2,Go)] */
  logic [1:0] incrHP_mergeQTree_Bool_buf_emitted;
  logic [1:0] incrHP_mergeQTree_Bool_buf_done;
  assign incrHP_QTree_Bool1_d = (incrHP_mergeQTree_Bool_buf_d[0] && (! incrHP_mergeQTree_Bool_buf_emitted[0]));
  assign incrHP_QTree_Bool2_d = (incrHP_mergeQTree_Bool_buf_d[0] && (! incrHP_mergeQTree_Bool_buf_emitted[1]));
  assign incrHP_mergeQTree_Bool_buf_done = (incrHP_mergeQTree_Bool_buf_emitted | ({incrHP_QTree_Bool2_d[0],
                                                                                   incrHP_QTree_Bool1_d[0]} & {incrHP_QTree_Bool2_r,
                                                                                                               incrHP_QTree_Bool1_r}));
  assign incrHP_mergeQTree_Bool_buf_r = (& incrHP_mergeQTree_Bool_buf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeQTree_Bool_buf_emitted <= 2'd0;
    else
      incrHP_mergeQTree_Bool_buf_emitted <= (incrHP_mergeQTree_Bool_buf_r ? 2'd0 :
                                             incrHP_mergeQTree_Bool_buf_done);
  
  /* op_add (Ty Word16#) : (incrHP_QTree_Bool,Word16#) (forkHP1_QTree_Bool,Word16#) > (addHP_QTree_Bool,Word16#) */
  assign addHP_QTree_Bool_d = {(incrHP_QTree_Bool_d[16:1] + forkHP1_QTree_Bool_d[16:1]),
                               (incrHP_QTree_Bool_d[0] && forkHP1_QTree_Bool_d[0])};
  assign {incrHP_QTree_Bool_r,
          forkHP1_QTree_Bool_r} = {2 {(addHP_QTree_Bool_r && addHP_QTree_Bool_d[0])}};
  
  /* merge (Ty Word16#) : [(initHP_QTree_Bool,Word16#),
                      (addHP_QTree_Bool,Word16#)] > (mergeHP_QTree_Bool,Word16#) */
  logic [1:0] mergeHP_QTree_Bool_selected;
  logic [1:0] mergeHP_QTree_Bool_select;
  always_comb
    begin
      mergeHP_QTree_Bool_selected = 2'd0;
      if ((| mergeHP_QTree_Bool_select))
        mergeHP_QTree_Bool_selected = mergeHP_QTree_Bool_select;
      else
        if (initHP_QTree_Bool_d[0]) mergeHP_QTree_Bool_selected[0] = 1'd1;
        else if (addHP_QTree_Bool_d[0])
          mergeHP_QTree_Bool_selected[1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_QTree_Bool_select <= 2'd0;
    else
      mergeHP_QTree_Bool_select <= (mergeHP_QTree_Bool_r ? 2'd0 :
                                    mergeHP_QTree_Bool_selected);
  always_comb
    if (mergeHP_QTree_Bool_selected[0])
      mergeHP_QTree_Bool_d = initHP_QTree_Bool_d;
    else if (mergeHP_QTree_Bool_selected[1])
      mergeHP_QTree_Bool_d = addHP_QTree_Bool_d;
    else mergeHP_QTree_Bool_d = {16'd0, 1'd0};
  assign {addHP_QTree_Bool_r,
          initHP_QTree_Bool_r} = (mergeHP_QTree_Bool_r ? mergeHP_QTree_Bool_selected :
                                  2'd0);
  
  /* buf (Ty Go) : (incrHP_mergeQTree_Bool,Go) > (incrHP_mergeQTree_Bool_buf,Go) */
  Go_t incrHP_mergeQTree_Bool_bufchan_d;
  logic incrHP_mergeQTree_Bool_bufchan_r;
  assign incrHP_mergeQTree_Bool_r = ((! incrHP_mergeQTree_Bool_bufchan_d[0]) || incrHP_mergeQTree_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeQTree_Bool_bufchan_d <= 1'd0;
    else
      if (incrHP_mergeQTree_Bool_r)
        incrHP_mergeQTree_Bool_bufchan_d <= incrHP_mergeQTree_Bool_d;
  Go_t incrHP_mergeQTree_Bool_bufchan_buf;
  assign incrHP_mergeQTree_Bool_bufchan_r = (! incrHP_mergeQTree_Bool_bufchan_buf[0]);
  assign incrHP_mergeQTree_Bool_buf_d = (incrHP_mergeQTree_Bool_bufchan_buf[0] ? incrHP_mergeQTree_Bool_bufchan_buf :
                                         incrHP_mergeQTree_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeQTree_Bool_bufchan_buf <= 1'd0;
    else
      if ((incrHP_mergeQTree_Bool_buf_r && incrHP_mergeQTree_Bool_bufchan_buf[0]))
        incrHP_mergeQTree_Bool_bufchan_buf <= 1'd0;
      else if (((! incrHP_mergeQTree_Bool_buf_r) && (! incrHP_mergeQTree_Bool_bufchan_buf[0])))
        incrHP_mergeQTree_Bool_bufchan_buf <= incrHP_mergeQTree_Bool_bufchan_d;
  
  /* buf (Ty Word16#) : (mergeHP_QTree_Bool,Word16#) > (mergeHP_QTree_Bool_buf,Word16#) */
  \Word16#_t  mergeHP_QTree_Bool_bufchan_d;
  logic mergeHP_QTree_Bool_bufchan_r;
  assign mergeHP_QTree_Bool_r = ((! mergeHP_QTree_Bool_bufchan_d[0]) || mergeHP_QTree_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_QTree_Bool_bufchan_d <= {16'd0, 1'd0};
    else
      if (mergeHP_QTree_Bool_r)
        mergeHP_QTree_Bool_bufchan_d <= mergeHP_QTree_Bool_d;
  \Word16#_t  mergeHP_QTree_Bool_bufchan_buf;
  assign mergeHP_QTree_Bool_bufchan_r = (! mergeHP_QTree_Bool_bufchan_buf[0]);
  assign mergeHP_QTree_Bool_buf_d = (mergeHP_QTree_Bool_bufchan_buf[0] ? mergeHP_QTree_Bool_bufchan_buf :
                                     mergeHP_QTree_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      mergeHP_QTree_Bool_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((mergeHP_QTree_Bool_buf_r && mergeHP_QTree_Bool_bufchan_buf[0]))
        mergeHP_QTree_Bool_bufchan_buf <= {16'd0, 1'd0};
      else if (((! mergeHP_QTree_Bool_buf_r) && (! mergeHP_QTree_Bool_bufchan_buf[0])))
        mergeHP_QTree_Bool_bufchan_buf <= mergeHP_QTree_Bool_bufchan_d;
  
  /* sink (Ty Word16#) : (forkHP1_QTree_Bool_snk,Word16#) > */
  assign {forkHP1_QTree_Bool_snk_r,
          forkHP1_QTree_Bool_snk_dout} = {forkHP1_QTree_Bool_snk_rout,
                                          forkHP1_QTree_Bool_snk_d};
  
  /* source (Ty Go) : > (\QTree_Bool_src,Go) */
  
  /* fork (Ty Go) : (\QTree_Bool_src,Go) > [(go_1_dummy_write_QTree_Bool,Go),
                                       (go_2_dummy_write_QTree_Bool,Go)] */
  logic [1:0] \\QTree_Bool_src_emitted ;
  logic [1:0] \\QTree_Bool_src_done ;
  assign go_1_dummy_write_QTree_Bool_d = (\\QTree_Bool_src_d [0] && (! \\QTree_Bool_src_emitted [0]));
  assign go_2_dummy_write_QTree_Bool_d = (\\QTree_Bool_src_d [0] && (! \\QTree_Bool_src_emitted [1]));
  assign \\QTree_Bool_src_done  = (\\QTree_Bool_src_emitted  | ({go_2_dummy_write_QTree_Bool_d[0],
                                                                 go_1_dummy_write_QTree_Bool_d[0]} & {go_2_dummy_write_QTree_Bool_r,
                                                                                                      go_1_dummy_write_QTree_Bool_r}));
  assign \\QTree_Bool_src_r  = (& \\QTree_Bool_src_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \\QTree_Bool_src_emitted  <= 2'd0;
    else
      \\QTree_Bool_src_emitted  <= (\\QTree_Bool_src_r  ? 2'd0 :
                                    \\QTree_Bool_src_done );
  
  /* source (Ty QTree_Bool) : > (dummy_write_QTree_Bool,QTree_Bool) */
  
  /* sink (Ty Pointer_QTree_Bool) : (dummy_write_QTree_Bool_sink,Pointer_QTree_Bool) > */
  assign {dummy_write_QTree_Bool_sink_r,
          dummy_write_QTree_Bool_sink_dout} = {dummy_write_QTree_Bool_sink_rout,
                                               dummy_write_QTree_Bool_sink_d};
  
  /* fork (Ty Word16#) : (mergeHP_QTree_Bool_buf,Word16#) > [(forkHP1_QTree_Bool,Word16#),
                                                        (forkHP1_QTree_Bool_snk,Word16#),
                                                        (forkHP1_QTree_Boo3,Word16#),
                                                        (forkHP1_QTree_Boo4,Word16#)] */
  logic [3:0] mergeHP_QTree_Bool_buf_emitted;
  logic [3:0] mergeHP_QTree_Bool_buf_done;
  assign forkHP1_QTree_Bool_d = {mergeHP_QTree_Bool_buf_d[16:1],
                                 (mergeHP_QTree_Bool_buf_d[0] && (! mergeHP_QTree_Bool_buf_emitted[0]))};
  assign forkHP1_QTree_Bool_snk_d = {mergeHP_QTree_Bool_buf_d[16:1],
                                     (mergeHP_QTree_Bool_buf_d[0] && (! mergeHP_QTree_Bool_buf_emitted[1]))};
  assign forkHP1_QTree_Boo3_d = {mergeHP_QTree_Bool_buf_d[16:1],
                                 (mergeHP_QTree_Bool_buf_d[0] && (! mergeHP_QTree_Bool_buf_emitted[2]))};
  assign forkHP1_QTree_Boo4_d = {mergeHP_QTree_Bool_buf_d[16:1],
                                 (mergeHP_QTree_Bool_buf_d[0] && (! mergeHP_QTree_Bool_buf_emitted[3]))};
  assign mergeHP_QTree_Bool_buf_done = (mergeHP_QTree_Bool_buf_emitted | ({forkHP1_QTree_Boo4_d[0],
                                                                           forkHP1_QTree_Boo3_d[0],
                                                                           forkHP1_QTree_Bool_snk_d[0],
                                                                           forkHP1_QTree_Bool_d[0]} & {forkHP1_QTree_Boo4_r,
                                                                                                       forkHP1_QTree_Boo3_r,
                                                                                                       forkHP1_QTree_Bool_snk_r,
                                                                                                       forkHP1_QTree_Bool_r}));
  assign mergeHP_QTree_Bool_buf_r = (& mergeHP_QTree_Bool_buf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_QTree_Bool_buf_emitted <= 4'd0;
    else
      mergeHP_QTree_Bool_buf_emitted <= (mergeHP_QTree_Bool_buf_r ? 4'd0 :
                                         mergeHP_QTree_Bool_buf_done);
  
  /* mergectrl (Ty C2,
           Ty MemIn_QTree_Bool) : [(dconReadIn_QTree_Bool,MemIn_QTree_Bool),
                                   (dconWriteIn_QTree_Bool,MemIn_QTree_Bool)] > (memMergeChoice_QTree_Bool,C2) (memMergeIn_QTree_Bool,MemIn_QTree_Bool) */
  logic [1:0] dconReadIn_QTree_Bool_select_d;
  assign dconReadIn_QTree_Bool_select_d = ((| dconReadIn_QTree_Bool_select_q) ? dconReadIn_QTree_Bool_select_q :
                                           (dconReadIn_QTree_Bool_d[0] ? 2'd1 :
                                            (dconWriteIn_QTree_Bool_d[0] ? 2'd2 :
                                             2'd0)));
  logic [1:0] dconReadIn_QTree_Bool_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) dconReadIn_QTree_Bool_select_q <= 2'd0;
    else
      dconReadIn_QTree_Bool_select_q <= (dconReadIn_QTree_Bool_done ? 2'd0 :
                                         dconReadIn_QTree_Bool_select_d);
  logic [1:0] dconReadIn_QTree_Bool_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) dconReadIn_QTree_Bool_emit_q <= 2'd0;
    else
      dconReadIn_QTree_Bool_emit_q <= (dconReadIn_QTree_Bool_done ? 2'd0 :
                                       dconReadIn_QTree_Bool_emit_d);
  logic [1:0] dconReadIn_QTree_Bool_emit_d;
  assign dconReadIn_QTree_Bool_emit_d = (dconReadIn_QTree_Bool_emit_q | ({memMergeChoice_QTree_Bool_d[0],
                                                                          memMergeIn_QTree_Bool_d[0]} & {memMergeChoice_QTree_Bool_r,
                                                                                                         memMergeIn_QTree_Bool_r}));
  logic dconReadIn_QTree_Bool_done;
  assign dconReadIn_QTree_Bool_done = (& dconReadIn_QTree_Bool_emit_d);
  assign {dconWriteIn_QTree_Bool_r,
          dconReadIn_QTree_Bool_r} = (dconReadIn_QTree_Bool_done ? dconReadIn_QTree_Bool_select_d :
                                      2'd0);
  assign memMergeIn_QTree_Bool_d = ((dconReadIn_QTree_Bool_select_d[0] && (! dconReadIn_QTree_Bool_emit_q[0])) ? dconReadIn_QTree_Bool_d :
                                    ((dconReadIn_QTree_Bool_select_d[1] && (! dconReadIn_QTree_Bool_emit_q[0])) ? dconWriteIn_QTree_Bool_d :
                                     {83'd0, 1'd0}));
  assign memMergeChoice_QTree_Bool_d = ((dconReadIn_QTree_Bool_select_d[0] && (! dconReadIn_QTree_Bool_emit_q[1])) ? C1_2_dc(1'd1) :
                                        ((dconReadIn_QTree_Bool_select_d[1] && (! dconReadIn_QTree_Bool_emit_q[1])) ? C2_2_dc(1'd1) :
                                         {1'd0, 1'd0}));
  
  /* bram (Ty MemIn_QTree_Bool,
      Ty MemOut_QTree_Bool) : (memMergeIn_QTree_Bool_dbuf,MemIn_QTree_Bool) > (memOut_QTree_Bool,MemOut_QTree_Bool) */
  logic [65:0] memMergeIn_QTree_Bool_dbuf_mem[65535:0];
  logic [15:0] memMergeIn_QTree_Bool_dbuf_address;
  logic [65:0] memMergeIn_QTree_Bool_dbuf_din;
  logic [65:0] memOut_QTree_Bool_q;
  logic memOut_QTree_Bool_valid;
  logic memMergeIn_QTree_Bool_dbuf_we;
  logic memOut_QTree_Bool_we;
  assign memMergeIn_QTree_Bool_dbuf_din = memMergeIn_QTree_Bool_dbuf_d[83:18];
  assign memMergeIn_QTree_Bool_dbuf_address = memMergeIn_QTree_Bool_dbuf_d[17:2];
  assign memMergeIn_QTree_Bool_dbuf_we = (memMergeIn_QTree_Bool_dbuf_d[1:1] && memMergeIn_QTree_Bool_dbuf_d[0]);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        memOut_QTree_Bool_we <= 1'd0;
        memOut_QTree_Bool_valid <= 1'd0;
      end
    else
      begin
        memOut_QTree_Bool_we <= memMergeIn_QTree_Bool_dbuf_we;
        memOut_QTree_Bool_valid <= memMergeIn_QTree_Bool_dbuf_d[0];
        if (memMergeIn_QTree_Bool_dbuf_we)
          begin
            memMergeIn_QTree_Bool_dbuf_mem[memMergeIn_QTree_Bool_dbuf_address] <= memMergeIn_QTree_Bool_dbuf_din;
            memOut_QTree_Bool_q <= memMergeIn_QTree_Bool_dbuf_din;
          end
        else
          memOut_QTree_Bool_q <= memMergeIn_QTree_Bool_dbuf_mem[memMergeIn_QTree_Bool_dbuf_address];
      end
  assign memOut_QTree_Bool_d = {memOut_QTree_Bool_q,
                                memOut_QTree_Bool_we,
                                memOut_QTree_Bool_valid};
  assign memMergeIn_QTree_Bool_dbuf_r = ((! memOut_QTree_Bool_valid) || memOut_QTree_Bool_r);
  logic [31:0] profiling_MemIn_QTree_Bool_read;
  logic [31:0] profiling_MemIn_QTree_Bool_write;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        profiling_MemIn_QTree_Bool_write <= 0;
        profiling_MemIn_QTree_Bool_read <= 0;
      end
    else
      if ((memMergeIn_QTree_Bool_dbuf_we == 1'd1))
        profiling_MemIn_QTree_Bool_write <= (profiling_MemIn_QTree_Bool_write + 1);
      else
        if ((memOut_QTree_Bool_valid == 1'd1))
          profiling_MemIn_QTree_Bool_read <= (profiling_MemIn_QTree_Bool_read + 1);
  
  /* demux (Ty C2,
       Ty MemOut_QTree_Bool) : (memMergeChoice_QTree_Bool,C2) (memOut_QTree_Bool_dbuf,MemOut_QTree_Bool) > [(memReadOut_QTree_Bool,MemOut_QTree_Bool),
                                                                                                            (memWriteOut_QTree_Bool,MemOut_QTree_Bool)] */
  logic [1:0] memOut_QTree_Bool_dbuf_onehotd;
  always_comb
    if ((memMergeChoice_QTree_Bool_d[0] && memOut_QTree_Bool_dbuf_d[0]))
      unique case (memMergeChoice_QTree_Bool_d[1:1])
        1'd0: memOut_QTree_Bool_dbuf_onehotd = 2'd1;
        1'd1: memOut_QTree_Bool_dbuf_onehotd = 2'd2;
        default: memOut_QTree_Bool_dbuf_onehotd = 2'd0;
      endcase
    else memOut_QTree_Bool_dbuf_onehotd = 2'd0;
  assign memReadOut_QTree_Bool_d = {memOut_QTree_Bool_dbuf_d[67:1],
                                    memOut_QTree_Bool_dbuf_onehotd[0]};
  assign memWriteOut_QTree_Bool_d = {memOut_QTree_Bool_dbuf_d[67:1],
                                     memOut_QTree_Bool_dbuf_onehotd[1]};
  assign memOut_QTree_Bool_dbuf_r = (| (memOut_QTree_Bool_dbuf_onehotd & {memWriteOut_QTree_Bool_r,
                                                                          memReadOut_QTree_Bool_r}));
  assign memMergeChoice_QTree_Bool_r = memOut_QTree_Bool_dbuf_r;
  
  /* dbuf (Ty MemIn_QTree_Bool) : (memMergeIn_QTree_Bool_rbuf,MemIn_QTree_Bool) > (memMergeIn_QTree_Bool_dbuf,MemIn_QTree_Bool) */
  assign memMergeIn_QTree_Bool_rbuf_r = ((! memMergeIn_QTree_Bool_dbuf_d[0]) || memMergeIn_QTree_Bool_dbuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memMergeIn_QTree_Bool_dbuf_d <= {83'd0, 1'd0};
    else
      if (memMergeIn_QTree_Bool_rbuf_r)
        memMergeIn_QTree_Bool_dbuf_d <= memMergeIn_QTree_Bool_rbuf_d;
  
  /* rbuf (Ty MemIn_QTree_Bool) : (memMergeIn_QTree_Bool,MemIn_QTree_Bool) > (memMergeIn_QTree_Bool_rbuf,MemIn_QTree_Bool) */
  MemIn_QTree_Bool_t memMergeIn_QTree_Bool_buf;
  assign memMergeIn_QTree_Bool_r = (! memMergeIn_QTree_Bool_buf[0]);
  assign memMergeIn_QTree_Bool_rbuf_d = (memMergeIn_QTree_Bool_buf[0] ? memMergeIn_QTree_Bool_buf :
                                         memMergeIn_QTree_Bool_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memMergeIn_QTree_Bool_buf <= {83'd0, 1'd0};
    else
      if ((memMergeIn_QTree_Bool_rbuf_r && memMergeIn_QTree_Bool_buf[0]))
        memMergeIn_QTree_Bool_buf <= {83'd0, 1'd0};
      else if (((! memMergeIn_QTree_Bool_rbuf_r) && (! memMergeIn_QTree_Bool_buf[0])))
        memMergeIn_QTree_Bool_buf <= memMergeIn_QTree_Bool_d;
  
  /* dbuf (Ty MemOut_QTree_Bool) : (memOut_QTree_Bool_rbuf,MemOut_QTree_Bool) > (memOut_QTree_Bool_dbuf,MemOut_QTree_Bool) */
  assign memOut_QTree_Bool_rbuf_r = ((! memOut_QTree_Bool_dbuf_d[0]) || memOut_QTree_Bool_dbuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memOut_QTree_Bool_dbuf_d <= {67'd0, 1'd0};
    else
      if (memOut_QTree_Bool_rbuf_r)
        memOut_QTree_Bool_dbuf_d <= memOut_QTree_Bool_rbuf_d;
  
  /* rbuf (Ty MemOut_QTree_Bool) : (memOut_QTree_Bool,MemOut_QTree_Bool) > (memOut_QTree_Bool_rbuf,MemOut_QTree_Bool) */
  MemOut_QTree_Bool_t memOut_QTree_Bool_buf;
  assign memOut_QTree_Bool_r = (! memOut_QTree_Bool_buf[0]);
  assign memOut_QTree_Bool_rbuf_d = (memOut_QTree_Bool_buf[0] ? memOut_QTree_Bool_buf :
                                     memOut_QTree_Bool_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memOut_QTree_Bool_buf <= {67'd0, 1'd0};
    else
      if ((memOut_QTree_Bool_rbuf_r && memOut_QTree_Bool_buf[0]))
        memOut_QTree_Bool_buf <= {67'd0, 1'd0};
      else if (((! memOut_QTree_Bool_rbuf_r) && (! memOut_QTree_Bool_buf[0])))
        memOut_QTree_Bool_buf <= memOut_QTree_Bool_d;
  
  /* mergectrl (Ty C5,
           Ty Pointer_QTree_Bool) : [(m2a86_1_argbuf,Pointer_QTree_Bool),
                                     (m2a8H_1_argbuf,Pointer_QTree_Bool),
                                     (m3a87_1_argbuf,Pointer_QTree_Bool),
                                     (m3a8I_1_argbuf,Pointer_QTree_Bool),
                                     (q4'a8x_1_argbuf,Pointer_QTree_Bool)] > (readMerge_choice_QTree_Bool,C5) (readMerge_data_QTree_Bool,Pointer_QTree_Bool) */
  logic [4:0] m2a86_1_argbuf_select_d;
  assign m2a86_1_argbuf_select_d = ((| m2a86_1_argbuf_select_q) ? m2a86_1_argbuf_select_q :
                                    (m2a86_1_argbuf_d[0] ? 5'd1 :
                                     (m2a8H_1_argbuf_d[0] ? 5'd2 :
                                      (m3a87_1_argbuf_d[0] ? 5'd4 :
                                       (m3a8I_1_argbuf_d[0] ? 5'd8 :
                                        (\q4'a8x_1_argbuf_d [0] ? 5'd16 :
                                         5'd0))))));
  logic [4:0] m2a86_1_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m2a86_1_argbuf_select_q <= 5'd0;
    else
      m2a86_1_argbuf_select_q <= (m2a86_1_argbuf_done ? 5'd0 :
                                  m2a86_1_argbuf_select_d);
  logic [1:0] m2a86_1_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m2a86_1_argbuf_emit_q <= 2'd0;
    else
      m2a86_1_argbuf_emit_q <= (m2a86_1_argbuf_done ? 2'd0 :
                                m2a86_1_argbuf_emit_d);
  logic [1:0] m2a86_1_argbuf_emit_d;
  assign m2a86_1_argbuf_emit_d = (m2a86_1_argbuf_emit_q | ({readMerge_choice_QTree_Bool_d[0],
                                                            readMerge_data_QTree_Bool_d[0]} & {readMerge_choice_QTree_Bool_r,
                                                                                               readMerge_data_QTree_Bool_r}));
  logic m2a86_1_argbuf_done;
  assign m2a86_1_argbuf_done = (& m2a86_1_argbuf_emit_d);
  assign {\q4'a8x_1_argbuf_r ,
          m3a8I_1_argbuf_r,
          m3a87_1_argbuf_r,
          m2a8H_1_argbuf_r,
          m2a86_1_argbuf_r} = (m2a86_1_argbuf_done ? m2a86_1_argbuf_select_d :
                               5'd0);
  assign readMerge_data_QTree_Bool_d = ((m2a86_1_argbuf_select_d[0] && (! m2a86_1_argbuf_emit_q[0])) ? m2a86_1_argbuf_d :
                                        ((m2a86_1_argbuf_select_d[1] && (! m2a86_1_argbuf_emit_q[0])) ? m2a8H_1_argbuf_d :
                                         ((m2a86_1_argbuf_select_d[2] && (! m2a86_1_argbuf_emit_q[0])) ? m3a87_1_argbuf_d :
                                          ((m2a86_1_argbuf_select_d[3] && (! m2a86_1_argbuf_emit_q[0])) ? m3a8I_1_argbuf_d :
                                           ((m2a86_1_argbuf_select_d[4] && (! m2a86_1_argbuf_emit_q[0])) ? \q4'a8x_1_argbuf_d  :
                                            {16'd0, 1'd0})))));
  assign readMerge_choice_QTree_Bool_d = ((m2a86_1_argbuf_select_d[0] && (! m2a86_1_argbuf_emit_q[1])) ? C1_5_dc(1'd1) :
                                          ((m2a86_1_argbuf_select_d[1] && (! m2a86_1_argbuf_emit_q[1])) ? C2_5_dc(1'd1) :
                                           ((m2a86_1_argbuf_select_d[2] && (! m2a86_1_argbuf_emit_q[1])) ? C3_5_dc(1'd1) :
                                            ((m2a86_1_argbuf_select_d[3] && (! m2a86_1_argbuf_emit_q[1])) ? C4_5_dc(1'd1) :
                                             ((m2a86_1_argbuf_select_d[4] && (! m2a86_1_argbuf_emit_q[1])) ? C5_5_dc(1'd1) :
                                              {3'd0, 1'd0})))));
  
  /* demux (Ty C5,
       Ty QTree_Bool) : (readMerge_choice_QTree_Bool,C5) (destructReadOut_QTree_Bool,QTree_Bool) > [(readPointer_QTree_Boolm2a86_1_argbuf,QTree_Bool),
                                                                                                    (readPointer_QTree_Boolm2a8H_1_argbuf,QTree_Bool),
                                                                                                    (readPointer_QTree_Boolm3a87_1_argbuf,QTree_Bool),
                                                                                                    (readPointer_QTree_Boolm3a8I_1_argbuf,QTree_Bool),
                                                                                                    (readPointer_QTree_Boolq4'a8x_1_argbuf,QTree_Bool)] */
  logic [4:0] destructReadOut_QTree_Bool_onehotd;
  always_comb
    if ((readMerge_choice_QTree_Bool_d[0] && destructReadOut_QTree_Bool_d[0]))
      unique case (readMerge_choice_QTree_Bool_d[3:1])
        3'd0: destructReadOut_QTree_Bool_onehotd = 5'd1;
        3'd1: destructReadOut_QTree_Bool_onehotd = 5'd2;
        3'd2: destructReadOut_QTree_Bool_onehotd = 5'd4;
        3'd3: destructReadOut_QTree_Bool_onehotd = 5'd8;
        3'd4: destructReadOut_QTree_Bool_onehotd = 5'd16;
        default: destructReadOut_QTree_Bool_onehotd = 5'd0;
      endcase
    else destructReadOut_QTree_Bool_onehotd = 5'd0;
  assign readPointer_QTree_Boolm2a86_1_argbuf_d = {destructReadOut_QTree_Bool_d[66:1],
                                                   destructReadOut_QTree_Bool_onehotd[0]};
  assign readPointer_QTree_Boolm2a8H_1_argbuf_d = {destructReadOut_QTree_Bool_d[66:1],
                                                   destructReadOut_QTree_Bool_onehotd[1]};
  assign readPointer_QTree_Boolm3a87_1_argbuf_d = {destructReadOut_QTree_Bool_d[66:1],
                                                   destructReadOut_QTree_Bool_onehotd[2]};
  assign readPointer_QTree_Boolm3a8I_1_argbuf_d = {destructReadOut_QTree_Bool_d[66:1],
                                                   destructReadOut_QTree_Bool_onehotd[3]};
  assign \readPointer_QTree_Boolq4'a8x_1_argbuf_d  = {destructReadOut_QTree_Bool_d[66:1],
                                                      destructReadOut_QTree_Bool_onehotd[4]};
  assign destructReadOut_QTree_Bool_r = (| (destructReadOut_QTree_Bool_onehotd & {\readPointer_QTree_Boolq4'a8x_1_argbuf_r ,
                                                                                  readPointer_QTree_Boolm3a8I_1_argbuf_r,
                                                                                  readPointer_QTree_Boolm3a87_1_argbuf_r,
                                                                                  readPointer_QTree_Boolm2a8H_1_argbuf_r,
                                                                                  readPointer_QTree_Boolm2a86_1_argbuf_r}));
  assign readMerge_choice_QTree_Bool_r = destructReadOut_QTree_Bool_r;
  
  /* destruct (Ty Pointer_QTree_Bool,
          Dcon Pointer_QTree_Bool) : (readMerge_data_QTree_Bool,Pointer_QTree_Bool) > [(destructReadIn_QTree_Bool,Word16#)] */
  assign destructReadIn_QTree_Bool_d = {readMerge_data_QTree_Bool_d[16:1],
                                        readMerge_data_QTree_Bool_d[0]};
  assign readMerge_data_QTree_Bool_r = destructReadIn_QTree_Bool_r;
  
  /* dcon (Ty MemIn_QTree_Bool,
      Dcon ReadIn_QTree_Bool) : [(destructReadIn_QTree_Bool,Word16#)] > (dconReadIn_QTree_Bool,MemIn_QTree_Bool) */
  assign dconReadIn_QTree_Bool_d = ReadIn_QTree_Bool_dc((& {destructReadIn_QTree_Bool_d[0]}), destructReadIn_QTree_Bool_d);
  assign {destructReadIn_QTree_Bool_r} = {1 {(dconReadIn_QTree_Bool_r && dconReadIn_QTree_Bool_d[0])}};
  
  /* destruct (Ty MemOut_QTree_Bool,
          Dcon ReadOut_QTree_Bool) : (memReadOut_QTree_Bool,MemOut_QTree_Bool) > [(destructReadOut_QTree_Bool,QTree_Bool)] */
  assign destructReadOut_QTree_Bool_d = {memReadOut_QTree_Bool_d[67:2],
                                         memReadOut_QTree_Bool_d[0]};
  assign memReadOut_QTree_Bool_r = destructReadOut_QTree_Bool_r;
  
  /* mergectrl (Ty C30,
           Ty QTree_Bool) : [(lizzieLet10_1_argbuf,QTree_Bool),
                             (lizzieLet11_1_argbuf,QTree_Bool),
                             (lizzieLet12_1_argbuf,QTree_Bool),
                             (lizzieLet13_1_1_argbuf,QTree_Bool),
                             (lizzieLet15_1_1_argbuf,QTree_Bool),
                             (lizzieLet16_1_1_argbuf,QTree_Bool),
                             (lizzieLet18_1_1_argbuf,QTree_Bool),
                             (lizzieLet19_2_1_argbuf,QTree_Bool),
                             (lizzieLet1_1_argbuf,QTree_Bool),
                             (lizzieLet22_1_1_argbuf,QTree_Bool),
                             (lizzieLet25_1_1_argbuf,QTree_Bool),
                             (lizzieLet26_1_1_argbuf,QTree_Bool),
                             (lizzieLet28_1_argbuf,QTree_Bool),
                             (lizzieLet30_1_argbuf,QTree_Bool),
                             (lizzieLet31_1_argbuf,QTree_Bool),
                             (lizzieLet33_1_argbuf,QTree_Bool),
                             (lizzieLet35_1_argbuf,QTree_Bool),
                             (lizzieLet36_1_argbuf,QTree_Bool),
                             (lizzieLet38_1_argbuf,QTree_Bool),
                             (lizzieLet42_1_argbuf,QTree_Bool),
                             (lizzieLet47_1_argbuf,QTree_Bool),
                             (lizzieLet4_1_argbuf,QTree_Bool),
                             (lizzieLet52_1_argbuf,QTree_Bool),
                             (lizzieLet57_1_argbuf,QTree_Bool),
                             (lizzieLet5_1_argbuf,QTree_Bool),
                             (lizzieLet6_1_argbuf,QTree_Bool),
                             (lizzieLet7_1_argbuf,QTree_Bool),
                             (lizzieLet9_1_1_argbuf,QTree_Bool),
                             (lizzieLet9_1_argbuf,QTree_Bool),
                             (dummy_write_QTree_Bool,QTree_Bool)] > (writeMerge_choice_QTree_Bool,C30) (writeMerge_data_QTree_Bool,QTree_Bool) */
  logic [29:0] lizzieLet10_1_argbuf_select_d;
  assign lizzieLet10_1_argbuf_select_d = ((| lizzieLet10_1_argbuf_select_q) ? lizzieLet10_1_argbuf_select_q :
                                          (lizzieLet10_1_argbuf_d[0] ? 30'd1 :
                                           (lizzieLet11_1_argbuf_d[0] ? 30'd2 :
                                            (lizzieLet12_1_argbuf_d[0] ? 30'd4 :
                                             (lizzieLet13_1_1_argbuf_d[0] ? 30'd8 :
                                              (lizzieLet15_1_1_argbuf_d[0] ? 30'd16 :
                                               (lizzieLet16_1_1_argbuf_d[0] ? 30'd32 :
                                                (lizzieLet18_1_1_argbuf_d[0] ? 30'd64 :
                                                 (lizzieLet19_2_1_argbuf_d[0] ? 30'd128 :
                                                  (lizzieLet1_1_argbuf_d[0] ? 30'd256 :
                                                   (lizzieLet22_1_1_argbuf_d[0] ? 30'd512 :
                                                    (lizzieLet25_1_1_argbuf_d[0] ? 30'd1024 :
                                                     (lizzieLet26_1_1_argbuf_d[0] ? 30'd2048 :
                                                      (lizzieLet28_1_argbuf_d[0] ? 30'd4096 :
                                                       (lizzieLet30_1_argbuf_d[0] ? 30'd8192 :
                                                        (lizzieLet31_1_argbuf_d[0] ? 30'd16384 :
                                                         (lizzieLet33_1_argbuf_d[0] ? 30'd32768 :
                                                          (lizzieLet35_1_argbuf_d[0] ? 30'd65536 :
                                                           (lizzieLet36_1_argbuf_d[0] ? 30'd131072 :
                                                            (lizzieLet38_1_argbuf_d[0] ? 30'd262144 :
                                                             (lizzieLet42_1_argbuf_d[0] ? 30'd524288 :
                                                              (lizzieLet47_1_argbuf_d[0] ? 30'd1048576 :
                                                               (lizzieLet4_1_argbuf_d[0] ? 30'd2097152 :
                                                                (lizzieLet52_1_argbuf_d[0] ? 30'd4194304 :
                                                                 (lizzieLet57_1_argbuf_d[0] ? 30'd8388608 :
                                                                  (lizzieLet5_1_argbuf_d[0] ? 30'd16777216 :
                                                                   (lizzieLet6_1_argbuf_d[0] ? 30'd33554432 :
                                                                    (lizzieLet7_1_argbuf_d[0] ? 30'd67108864 :
                                                                     (lizzieLet9_1_1_argbuf_d[0] ? 30'd134217728 :
                                                                      (lizzieLet9_1_argbuf_d[0] ? 30'd268435456 :
                                                                       (dummy_write_QTree_Bool_d[0] ? 30'd536870912 :
                                                                        30'd0)))))))))))))))))))))))))))))));
  logic [29:0] lizzieLet10_1_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet10_1_argbuf_select_q <= 30'd0;
    else
      lizzieLet10_1_argbuf_select_q <= (lizzieLet10_1_argbuf_done ? 30'd0 :
                                        lizzieLet10_1_argbuf_select_d);
  logic [1:0] lizzieLet10_1_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet10_1_argbuf_emit_q <= 2'd0;
    else
      lizzieLet10_1_argbuf_emit_q <= (lizzieLet10_1_argbuf_done ? 2'd0 :
                                      lizzieLet10_1_argbuf_emit_d);
  logic [1:0] lizzieLet10_1_argbuf_emit_d;
  assign lizzieLet10_1_argbuf_emit_d = (lizzieLet10_1_argbuf_emit_q | ({writeMerge_choice_QTree_Bool_d[0],
                                                                        writeMerge_data_QTree_Bool_d[0]} & {writeMerge_choice_QTree_Bool_r,
                                                                                                            writeMerge_data_QTree_Bool_r}));
  logic lizzieLet10_1_argbuf_done;
  assign lizzieLet10_1_argbuf_done = (& lizzieLet10_1_argbuf_emit_d);
  assign {dummy_write_QTree_Bool_r,
          lizzieLet9_1_argbuf_r,
          lizzieLet9_1_1_argbuf_r,
          lizzieLet7_1_argbuf_r,
          lizzieLet6_1_argbuf_r,
          lizzieLet5_1_argbuf_r,
          lizzieLet57_1_argbuf_r,
          lizzieLet52_1_argbuf_r,
          lizzieLet4_1_argbuf_r,
          lizzieLet47_1_argbuf_r,
          lizzieLet42_1_argbuf_r,
          lizzieLet38_1_argbuf_r,
          lizzieLet36_1_argbuf_r,
          lizzieLet35_1_argbuf_r,
          lizzieLet33_1_argbuf_r,
          lizzieLet31_1_argbuf_r,
          lizzieLet30_1_argbuf_r,
          lizzieLet28_1_argbuf_r,
          lizzieLet26_1_1_argbuf_r,
          lizzieLet25_1_1_argbuf_r,
          lizzieLet22_1_1_argbuf_r,
          lizzieLet1_1_argbuf_r,
          lizzieLet19_2_1_argbuf_r,
          lizzieLet18_1_1_argbuf_r,
          lizzieLet16_1_1_argbuf_r,
          lizzieLet15_1_1_argbuf_r,
          lizzieLet13_1_1_argbuf_r,
          lizzieLet12_1_argbuf_r,
          lizzieLet11_1_argbuf_r,
          lizzieLet10_1_argbuf_r} = (lizzieLet10_1_argbuf_done ? lizzieLet10_1_argbuf_select_d :
                                     30'd0);
  assign writeMerge_data_QTree_Bool_d = ((lizzieLet10_1_argbuf_select_d[0] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet10_1_argbuf_d :
                                         ((lizzieLet10_1_argbuf_select_d[1] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet11_1_argbuf_d :
                                          ((lizzieLet10_1_argbuf_select_d[2] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet12_1_argbuf_d :
                                           ((lizzieLet10_1_argbuf_select_d[3] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet13_1_1_argbuf_d :
                                            ((lizzieLet10_1_argbuf_select_d[4] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet15_1_1_argbuf_d :
                                             ((lizzieLet10_1_argbuf_select_d[5] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet16_1_1_argbuf_d :
                                              ((lizzieLet10_1_argbuf_select_d[6] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet18_1_1_argbuf_d :
                                               ((lizzieLet10_1_argbuf_select_d[7] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet19_2_1_argbuf_d :
                                                ((lizzieLet10_1_argbuf_select_d[8] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet1_1_argbuf_d :
                                                 ((lizzieLet10_1_argbuf_select_d[9] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet22_1_1_argbuf_d :
                                                  ((lizzieLet10_1_argbuf_select_d[10] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet25_1_1_argbuf_d :
                                                   ((lizzieLet10_1_argbuf_select_d[11] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet26_1_1_argbuf_d :
                                                    ((lizzieLet10_1_argbuf_select_d[12] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet28_1_argbuf_d :
                                                     ((lizzieLet10_1_argbuf_select_d[13] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet30_1_argbuf_d :
                                                      ((lizzieLet10_1_argbuf_select_d[14] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet31_1_argbuf_d :
                                                       ((lizzieLet10_1_argbuf_select_d[15] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet33_1_argbuf_d :
                                                        ((lizzieLet10_1_argbuf_select_d[16] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet35_1_argbuf_d :
                                                         ((lizzieLet10_1_argbuf_select_d[17] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet36_1_argbuf_d :
                                                          ((lizzieLet10_1_argbuf_select_d[18] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet38_1_argbuf_d :
                                                           ((lizzieLet10_1_argbuf_select_d[19] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet42_1_argbuf_d :
                                                            ((lizzieLet10_1_argbuf_select_d[20] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet47_1_argbuf_d :
                                                             ((lizzieLet10_1_argbuf_select_d[21] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet4_1_argbuf_d :
                                                              ((lizzieLet10_1_argbuf_select_d[22] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet52_1_argbuf_d :
                                                               ((lizzieLet10_1_argbuf_select_d[23] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet57_1_argbuf_d :
                                                                ((lizzieLet10_1_argbuf_select_d[24] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet5_1_argbuf_d :
                                                                 ((lizzieLet10_1_argbuf_select_d[25] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet6_1_argbuf_d :
                                                                  ((lizzieLet10_1_argbuf_select_d[26] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet7_1_argbuf_d :
                                                                   ((lizzieLet10_1_argbuf_select_d[27] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet9_1_1_argbuf_d :
                                                                    ((lizzieLet10_1_argbuf_select_d[28] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet9_1_argbuf_d :
                                                                     ((lizzieLet10_1_argbuf_select_d[29] && (! lizzieLet10_1_argbuf_emit_q[0])) ? dummy_write_QTree_Bool_d :
                                                                      {66'd0,
                                                                       1'd0}))))))))))))))))))))))))))))));
  assign writeMerge_choice_QTree_Bool_d = ((lizzieLet10_1_argbuf_select_d[0] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C1_30_dc(1'd1) :
                                           ((lizzieLet10_1_argbuf_select_d[1] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C2_30_dc(1'd1) :
                                            ((lizzieLet10_1_argbuf_select_d[2] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C3_30_dc(1'd1) :
                                             ((lizzieLet10_1_argbuf_select_d[3] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C4_30_dc(1'd1) :
                                              ((lizzieLet10_1_argbuf_select_d[4] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C5_30_dc(1'd1) :
                                               ((lizzieLet10_1_argbuf_select_d[5] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C6_30_dc(1'd1) :
                                                ((lizzieLet10_1_argbuf_select_d[6] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C7_30_dc(1'd1) :
                                                 ((lizzieLet10_1_argbuf_select_d[7] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C8_30_dc(1'd1) :
                                                  ((lizzieLet10_1_argbuf_select_d[8] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C9_30_dc(1'd1) :
                                                   ((lizzieLet10_1_argbuf_select_d[9] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C10_30_dc(1'd1) :
                                                    ((lizzieLet10_1_argbuf_select_d[10] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C11_30_dc(1'd1) :
                                                     ((lizzieLet10_1_argbuf_select_d[11] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C12_30_dc(1'd1) :
                                                      ((lizzieLet10_1_argbuf_select_d[12] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C13_30_dc(1'd1) :
                                                       ((lizzieLet10_1_argbuf_select_d[13] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C14_30_dc(1'd1) :
                                                        ((lizzieLet10_1_argbuf_select_d[14] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C15_30_dc(1'd1) :
                                                         ((lizzieLet10_1_argbuf_select_d[15] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C16_30_dc(1'd1) :
                                                          ((lizzieLet10_1_argbuf_select_d[16] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C17_30_dc(1'd1) :
                                                           ((lizzieLet10_1_argbuf_select_d[17] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C18_30_dc(1'd1) :
                                                            ((lizzieLet10_1_argbuf_select_d[18] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C19_30_dc(1'd1) :
                                                             ((lizzieLet10_1_argbuf_select_d[19] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C20_30_dc(1'd1) :
                                                              ((lizzieLet10_1_argbuf_select_d[20] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C21_30_dc(1'd1) :
                                                               ((lizzieLet10_1_argbuf_select_d[21] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C22_30_dc(1'd1) :
                                                                ((lizzieLet10_1_argbuf_select_d[22] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C23_30_dc(1'd1) :
                                                                 ((lizzieLet10_1_argbuf_select_d[23] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C24_30_dc(1'd1) :
                                                                  ((lizzieLet10_1_argbuf_select_d[24] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C25_30_dc(1'd1) :
                                                                   ((lizzieLet10_1_argbuf_select_d[25] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C26_30_dc(1'd1) :
                                                                    ((lizzieLet10_1_argbuf_select_d[26] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C27_30_dc(1'd1) :
                                                                     ((lizzieLet10_1_argbuf_select_d[27] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C28_30_dc(1'd1) :
                                                                      ((lizzieLet10_1_argbuf_select_d[28] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C29_30_dc(1'd1) :
                                                                       ((lizzieLet10_1_argbuf_select_d[29] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C30_30_dc(1'd1) :
                                                                        {5'd0,
                                                                         1'd0}))))))))))))))))))))))))))))));
  
  /* demux (Ty C30,
       Ty Pointer_QTree_Bool) : (writeMerge_choice_QTree_Bool,C30) (demuxWriteResult_QTree_Bool,Pointer_QTree_Bool) > [(writeQTree_BoollizzieLet10_1_argbuf,Pointer_QTree_Bool),
                                                                                                                       (writeQTree_BoollizzieLet11_1_argbuf,Pointer_QTree_Bool),
                                                                                                                       (writeQTree_BoollizzieLet12_1_argbuf,Pointer_QTree_Bool),
                                                                                                                       (writeQTree_BoollizzieLet13_1_1_argbuf,Pointer_QTree_Bool),
                                                                                                                       (writeQTree_BoollizzieLet15_1_1_argbuf,Pointer_QTree_Bool),
                                                                                                                       (writeQTree_BoollizzieLet16_1_1_argbuf,Pointer_QTree_Bool),
                                                                                                                       (writeQTree_BoollizzieLet18_1_1_argbuf,Pointer_QTree_Bool),
                                                                                                                       (writeQTree_BoollizzieLet19_2_1_argbuf,Pointer_QTree_Bool),
                                                                                                                       (writeQTree_BoollizzieLet1_1_argbuf,Pointer_QTree_Bool),
                                                                                                                       (writeQTree_BoollizzieLet22_1_1_argbuf,Pointer_QTree_Bool),
                                                                                                                       (writeQTree_BoollizzieLet25_1_1_argbuf,Pointer_QTree_Bool),
                                                                                                                       (writeQTree_BoollizzieLet26_1_1_argbuf,Pointer_QTree_Bool),
                                                                                                                       (writeQTree_BoollizzieLet28_1_argbuf,Pointer_QTree_Bool),
                                                                                                                       (writeQTree_BoollizzieLet30_1_argbuf,Pointer_QTree_Bool),
                                                                                                                       (writeQTree_BoollizzieLet31_1_argbuf,Pointer_QTree_Bool),
                                                                                                                       (writeQTree_BoollizzieLet33_1_argbuf,Pointer_QTree_Bool),
                                                                                                                       (writeQTree_BoollizzieLet35_1_argbuf,Pointer_QTree_Bool),
                                                                                                                       (writeQTree_BoollizzieLet36_1_argbuf,Pointer_QTree_Bool),
                                                                                                                       (writeQTree_BoollizzieLet38_1_argbuf,Pointer_QTree_Bool),
                                                                                                                       (writeQTree_BoollizzieLet42_1_argbuf,Pointer_QTree_Bool),
                                                                                                                       (writeQTree_BoollizzieLet47_1_argbuf,Pointer_QTree_Bool),
                                                                                                                       (writeQTree_BoollizzieLet4_1_argbuf,Pointer_QTree_Bool),
                                                                                                                       (writeQTree_BoollizzieLet52_1_argbuf,Pointer_QTree_Bool),
                                                                                                                       (writeQTree_BoollizzieLet57_1_argbuf,Pointer_QTree_Bool),
                                                                                                                       (writeQTree_BoollizzieLet5_1_argbuf,Pointer_QTree_Bool),
                                                                                                                       (writeQTree_BoollizzieLet6_1_argbuf,Pointer_QTree_Bool),
                                                                                                                       (writeQTree_BoollizzieLet7_1_argbuf,Pointer_QTree_Bool),
                                                                                                                       (writeQTree_BoollizzieLet9_1_1_argbuf,Pointer_QTree_Bool),
                                                                                                                       (writeQTree_BoollizzieLet9_1_argbuf,Pointer_QTree_Bool),
                                                                                                                       (dummy_write_QTree_Bool_sink,Pointer_QTree_Bool)] */
  logic [29:0] demuxWriteResult_QTree_Bool_onehotd;
  always_comb
    if ((writeMerge_choice_QTree_Bool_d[0] && demuxWriteResult_QTree_Bool_d[0]))
      unique case (writeMerge_choice_QTree_Bool_d[5:1])
        5'd0: demuxWriteResult_QTree_Bool_onehotd = 30'd1;
        5'd1: demuxWriteResult_QTree_Bool_onehotd = 30'd2;
        5'd2: demuxWriteResult_QTree_Bool_onehotd = 30'd4;
        5'd3: demuxWriteResult_QTree_Bool_onehotd = 30'd8;
        5'd4: demuxWriteResult_QTree_Bool_onehotd = 30'd16;
        5'd5: demuxWriteResult_QTree_Bool_onehotd = 30'd32;
        5'd6: demuxWriteResult_QTree_Bool_onehotd = 30'd64;
        5'd7: demuxWriteResult_QTree_Bool_onehotd = 30'd128;
        5'd8: demuxWriteResult_QTree_Bool_onehotd = 30'd256;
        5'd9: demuxWriteResult_QTree_Bool_onehotd = 30'd512;
        5'd10: demuxWriteResult_QTree_Bool_onehotd = 30'd1024;
        5'd11: demuxWriteResult_QTree_Bool_onehotd = 30'd2048;
        5'd12: demuxWriteResult_QTree_Bool_onehotd = 30'd4096;
        5'd13: demuxWriteResult_QTree_Bool_onehotd = 30'd8192;
        5'd14: demuxWriteResult_QTree_Bool_onehotd = 30'd16384;
        5'd15: demuxWriteResult_QTree_Bool_onehotd = 30'd32768;
        5'd16: demuxWriteResult_QTree_Bool_onehotd = 30'd65536;
        5'd17: demuxWriteResult_QTree_Bool_onehotd = 30'd131072;
        5'd18: demuxWriteResult_QTree_Bool_onehotd = 30'd262144;
        5'd19: demuxWriteResult_QTree_Bool_onehotd = 30'd524288;
        5'd20: demuxWriteResult_QTree_Bool_onehotd = 30'd1048576;
        5'd21: demuxWriteResult_QTree_Bool_onehotd = 30'd2097152;
        5'd22: demuxWriteResult_QTree_Bool_onehotd = 30'd4194304;
        5'd23: demuxWriteResult_QTree_Bool_onehotd = 30'd8388608;
        5'd24: demuxWriteResult_QTree_Bool_onehotd = 30'd16777216;
        5'd25: demuxWriteResult_QTree_Bool_onehotd = 30'd33554432;
        5'd26: demuxWriteResult_QTree_Bool_onehotd = 30'd67108864;
        5'd27: demuxWriteResult_QTree_Bool_onehotd = 30'd134217728;
        5'd28: demuxWriteResult_QTree_Bool_onehotd = 30'd268435456;
        5'd29: demuxWriteResult_QTree_Bool_onehotd = 30'd536870912;
        default: demuxWriteResult_QTree_Bool_onehotd = 30'd0;
      endcase
    else demuxWriteResult_QTree_Bool_onehotd = 30'd0;
  assign writeQTree_BoollizzieLet10_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                  demuxWriteResult_QTree_Bool_onehotd[0]};
  assign writeQTree_BoollizzieLet11_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                  demuxWriteResult_QTree_Bool_onehotd[1]};
  assign writeQTree_BoollizzieLet12_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                  demuxWriteResult_QTree_Bool_onehotd[2]};
  assign writeQTree_BoollizzieLet13_1_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                    demuxWriteResult_QTree_Bool_onehotd[3]};
  assign writeQTree_BoollizzieLet15_1_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                    demuxWriteResult_QTree_Bool_onehotd[4]};
  assign writeQTree_BoollizzieLet16_1_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                    demuxWriteResult_QTree_Bool_onehotd[5]};
  assign writeQTree_BoollizzieLet18_1_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                    demuxWriteResult_QTree_Bool_onehotd[6]};
  assign writeQTree_BoollizzieLet19_2_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                    demuxWriteResult_QTree_Bool_onehotd[7]};
  assign writeQTree_BoollizzieLet1_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                 demuxWriteResult_QTree_Bool_onehotd[8]};
  assign writeQTree_BoollizzieLet22_1_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                    demuxWriteResult_QTree_Bool_onehotd[9]};
  assign writeQTree_BoollizzieLet25_1_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                    demuxWriteResult_QTree_Bool_onehotd[10]};
  assign writeQTree_BoollizzieLet26_1_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                    demuxWriteResult_QTree_Bool_onehotd[11]};
  assign writeQTree_BoollizzieLet28_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                  demuxWriteResult_QTree_Bool_onehotd[12]};
  assign writeQTree_BoollizzieLet30_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                  demuxWriteResult_QTree_Bool_onehotd[13]};
  assign writeQTree_BoollizzieLet31_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                  demuxWriteResult_QTree_Bool_onehotd[14]};
  assign writeQTree_BoollizzieLet33_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                  demuxWriteResult_QTree_Bool_onehotd[15]};
  assign writeQTree_BoollizzieLet35_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                  demuxWriteResult_QTree_Bool_onehotd[16]};
  assign writeQTree_BoollizzieLet36_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                  demuxWriteResult_QTree_Bool_onehotd[17]};
  assign writeQTree_BoollizzieLet38_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                  demuxWriteResult_QTree_Bool_onehotd[18]};
  assign writeQTree_BoollizzieLet42_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                  demuxWriteResult_QTree_Bool_onehotd[19]};
  assign writeQTree_BoollizzieLet47_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                  demuxWriteResult_QTree_Bool_onehotd[20]};
  assign writeQTree_BoollizzieLet4_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                 demuxWriteResult_QTree_Bool_onehotd[21]};
  assign writeQTree_BoollizzieLet52_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                  demuxWriteResult_QTree_Bool_onehotd[22]};
  assign writeQTree_BoollizzieLet57_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                  demuxWriteResult_QTree_Bool_onehotd[23]};
  assign writeQTree_BoollizzieLet5_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                 demuxWriteResult_QTree_Bool_onehotd[24]};
  assign writeQTree_BoollizzieLet6_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                 demuxWriteResult_QTree_Bool_onehotd[25]};
  assign writeQTree_BoollizzieLet7_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                 demuxWriteResult_QTree_Bool_onehotd[26]};
  assign writeQTree_BoollizzieLet9_1_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                   demuxWriteResult_QTree_Bool_onehotd[27]};
  assign writeQTree_BoollizzieLet9_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                 demuxWriteResult_QTree_Bool_onehotd[28]};
  assign dummy_write_QTree_Bool_sink_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                          demuxWriteResult_QTree_Bool_onehotd[29]};
  assign demuxWriteResult_QTree_Bool_r = (| (demuxWriteResult_QTree_Bool_onehotd & {dummy_write_QTree_Bool_sink_r,
                                                                                    writeQTree_BoollizzieLet9_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet9_1_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet7_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet6_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet5_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet57_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet52_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet4_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet47_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet42_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet38_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet36_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet35_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet33_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet31_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet30_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet28_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet26_1_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet25_1_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet22_1_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet1_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet19_2_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet18_1_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet16_1_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet15_1_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet13_1_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet12_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet11_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet10_1_argbuf_r}));
  assign writeMerge_choice_QTree_Bool_r = demuxWriteResult_QTree_Bool_r;
  
  /* dcon (Ty MemIn_QTree_Bool,
      Dcon WriteIn_QTree_Bool) : [(forkHP1_QTree_Boo3,Word16#),
                                  (writeMerge_data_QTree_Bool,QTree_Bool)] > (dconWriteIn_QTree_Bool,MemIn_QTree_Bool) */
  assign dconWriteIn_QTree_Bool_d = WriteIn_QTree_Bool_dc((& {forkHP1_QTree_Boo3_d[0],
                                                              writeMerge_data_QTree_Bool_d[0]}), forkHP1_QTree_Boo3_d, writeMerge_data_QTree_Bool_d);
  assign {forkHP1_QTree_Boo3_r,
          writeMerge_data_QTree_Bool_r} = {2 {(dconWriteIn_QTree_Bool_r && dconWriteIn_QTree_Bool_d[0])}};
  
  /* dcon (Ty Pointer_QTree_Bool,
      Dcon Pointer_QTree_Bool) : [(forkHP1_QTree_Boo4,Word16#)] > (dconPtr_QTree_Bool,Pointer_QTree_Bool) */
  assign dconPtr_QTree_Bool_d = Pointer_QTree_Bool_dc((& {forkHP1_QTree_Boo4_d[0]}), forkHP1_QTree_Boo4_d);
  assign {forkHP1_QTree_Boo4_r} = {1 {(dconPtr_QTree_Bool_r && dconPtr_QTree_Bool_d[0])}};
  
  /* demux (Ty MemOut_QTree_Bool,
       Ty Pointer_QTree_Bool) : (memWriteOut_QTree_Bool,MemOut_QTree_Bool) (dconPtr_QTree_Bool,Pointer_QTree_Bool) > [(_130,Pointer_QTree_Bool),
                                                                                                                      (demuxWriteResult_QTree_Bool,Pointer_QTree_Bool)] */
  logic [1:0] dconPtr_QTree_Bool_onehotd;
  always_comb
    if ((memWriteOut_QTree_Bool_d[0] && dconPtr_QTree_Bool_d[0]))
      unique case (memWriteOut_QTree_Bool_d[1:1])
        1'd0: dconPtr_QTree_Bool_onehotd = 2'd1;
        1'd1: dconPtr_QTree_Bool_onehotd = 2'd2;
        default: dconPtr_QTree_Bool_onehotd = 2'd0;
      endcase
    else dconPtr_QTree_Bool_onehotd = 2'd0;
  assign _130_d = {dconPtr_QTree_Bool_d[16:1],
                   dconPtr_QTree_Bool_onehotd[0]};
  assign demuxWriteResult_QTree_Bool_d = {dconPtr_QTree_Bool_d[16:1],
                                          dconPtr_QTree_Bool_onehotd[1]};
  assign dconPtr_QTree_Bool_r = (| (dconPtr_QTree_Bool_onehotd & {demuxWriteResult_QTree_Bool_r,
                                                                  _130_r}));
  assign memWriteOut_QTree_Bool_r = dconPtr_QTree_Bool_r;
  
  /* const (Ty Word16#,Lit 0) : (goFor_2,Go) > (initHP_CTf,Word16#) */
  assign initHP_CTf_d = {16'd0, goFor_2_d[0]};
  assign goFor_2_r = initHP_CTf_r;
  
  /* const (Ty Word16#,Lit 1) : (incrHP_CTf1,Go) > (incrHP_CTf,Word16#) */
  assign incrHP_CTf_d = {16'd1, incrHP_CTf1_d[0]};
  assign incrHP_CTf1_r = incrHP_CTf_r;
  
  /* merge (Ty Go) : [(goFor_3,Go),
                 (incrHP_CTf2,Go)] > (incrHP_mergeCTf,Go) */
  logic [1:0] incrHP_mergeCTf_selected;
  logic [1:0] incrHP_mergeCTf_select;
  always_comb
    begin
      incrHP_mergeCTf_selected = 2'd0;
      if ((| incrHP_mergeCTf_select))
        incrHP_mergeCTf_selected = incrHP_mergeCTf_select;
      else
        if (goFor_3_d[0]) incrHP_mergeCTf_selected[0] = 1'd1;
        else if (incrHP_CTf2_d[0]) incrHP_mergeCTf_selected[1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeCTf_select <= 2'd0;
    else
      incrHP_mergeCTf_select <= (incrHP_mergeCTf_r ? 2'd0 :
                                 incrHP_mergeCTf_selected);
  always_comb
    if (incrHP_mergeCTf_selected[0]) incrHP_mergeCTf_d = goFor_3_d;
    else if (incrHP_mergeCTf_selected[1])
      incrHP_mergeCTf_d = incrHP_CTf2_d;
    else incrHP_mergeCTf_d = 1'd0;
  assign {incrHP_CTf2_r,
          goFor_3_r} = (incrHP_mergeCTf_r ? incrHP_mergeCTf_selected :
                        2'd0);
  
  /* fork (Ty Go) : (incrHP_mergeCTf_buf,Go) > [(incrHP_CTf1,Go),
                                           (incrHP_CTf2,Go)] */
  logic [1:0] incrHP_mergeCTf_buf_emitted;
  logic [1:0] incrHP_mergeCTf_buf_done;
  assign incrHP_CTf1_d = (incrHP_mergeCTf_buf_d[0] && (! incrHP_mergeCTf_buf_emitted[0]));
  assign incrHP_CTf2_d = (incrHP_mergeCTf_buf_d[0] && (! incrHP_mergeCTf_buf_emitted[1]));
  assign incrHP_mergeCTf_buf_done = (incrHP_mergeCTf_buf_emitted | ({incrHP_CTf2_d[0],
                                                                     incrHP_CTf1_d[0]} & {incrHP_CTf2_r,
                                                                                          incrHP_CTf1_r}));
  assign incrHP_mergeCTf_buf_r = (& incrHP_mergeCTf_buf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeCTf_buf_emitted <= 2'd0;
    else
      incrHP_mergeCTf_buf_emitted <= (incrHP_mergeCTf_buf_r ? 2'd0 :
                                      incrHP_mergeCTf_buf_done);
  
  /* op_add (Ty Word16#) : (incrHP_CTf,Word16#) (forkHP1_CTf,Word16#) > (addHP_CTf,Word16#) */
  assign addHP_CTf_d = {(incrHP_CTf_d[16:1] + forkHP1_CTf_d[16:1]),
                        (incrHP_CTf_d[0] && forkHP1_CTf_d[0])};
  assign {incrHP_CTf_r,
          forkHP1_CTf_r} = {2 {(addHP_CTf_r && addHP_CTf_d[0])}};
  
  /* merge (Ty Word16#) : [(initHP_CTf,Word16#),
                      (addHP_CTf,Word16#)] > (mergeHP_CTf,Word16#) */
  logic [1:0] mergeHP_CTf_selected;
  logic [1:0] mergeHP_CTf_select;
  always_comb
    begin
      mergeHP_CTf_selected = 2'd0;
      if ((| mergeHP_CTf_select))
        mergeHP_CTf_selected = mergeHP_CTf_select;
      else
        if (initHP_CTf_d[0]) mergeHP_CTf_selected[0] = 1'd1;
        else if (addHP_CTf_d[0]) mergeHP_CTf_selected[1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_CTf_select <= 2'd0;
    else
      mergeHP_CTf_select <= (mergeHP_CTf_r ? 2'd0 :
                             mergeHP_CTf_selected);
  always_comb
    if (mergeHP_CTf_selected[0]) mergeHP_CTf_d = initHP_CTf_d;
    else if (mergeHP_CTf_selected[1]) mergeHP_CTf_d = addHP_CTf_d;
    else mergeHP_CTf_d = {16'd0, 1'd0};
  assign {addHP_CTf_r,
          initHP_CTf_r} = (mergeHP_CTf_r ? mergeHP_CTf_selected :
                           2'd0);
  
  /* buf (Ty Go) : (incrHP_mergeCTf,Go) > (incrHP_mergeCTf_buf,Go) */
  Go_t incrHP_mergeCTf_bufchan_d;
  logic incrHP_mergeCTf_bufchan_r;
  assign incrHP_mergeCTf_r = ((! incrHP_mergeCTf_bufchan_d[0]) || incrHP_mergeCTf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeCTf_bufchan_d <= 1'd0;
    else
      if (incrHP_mergeCTf_r)
        incrHP_mergeCTf_bufchan_d <= incrHP_mergeCTf_d;
  Go_t incrHP_mergeCTf_bufchan_buf;
  assign incrHP_mergeCTf_bufchan_r = (! incrHP_mergeCTf_bufchan_buf[0]);
  assign incrHP_mergeCTf_buf_d = (incrHP_mergeCTf_bufchan_buf[0] ? incrHP_mergeCTf_bufchan_buf :
                                  incrHP_mergeCTf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeCTf_bufchan_buf <= 1'd0;
    else
      if ((incrHP_mergeCTf_buf_r && incrHP_mergeCTf_bufchan_buf[0]))
        incrHP_mergeCTf_bufchan_buf <= 1'd0;
      else if (((! incrHP_mergeCTf_buf_r) && (! incrHP_mergeCTf_bufchan_buf[0])))
        incrHP_mergeCTf_bufchan_buf <= incrHP_mergeCTf_bufchan_d;
  
  /* buf (Ty Word16#) : (mergeHP_CTf,Word16#) > (mergeHP_CTf_buf,Word16#) */
  \Word16#_t  mergeHP_CTf_bufchan_d;
  logic mergeHP_CTf_bufchan_r;
  assign mergeHP_CTf_r = ((! mergeHP_CTf_bufchan_d[0]) || mergeHP_CTf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_CTf_bufchan_d <= {16'd0, 1'd0};
    else if (mergeHP_CTf_r) mergeHP_CTf_bufchan_d <= mergeHP_CTf_d;
  \Word16#_t  mergeHP_CTf_bufchan_buf;
  assign mergeHP_CTf_bufchan_r = (! mergeHP_CTf_bufchan_buf[0]);
  assign mergeHP_CTf_buf_d = (mergeHP_CTf_bufchan_buf[0] ? mergeHP_CTf_bufchan_buf :
                              mergeHP_CTf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_CTf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((mergeHP_CTf_buf_r && mergeHP_CTf_bufchan_buf[0]))
        mergeHP_CTf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! mergeHP_CTf_buf_r) && (! mergeHP_CTf_bufchan_buf[0])))
        mergeHP_CTf_bufchan_buf <= mergeHP_CTf_bufchan_d;
  
  /* fork (Ty Word16#) : (mergeHP_CTf_buf,Word16#) > [(forkHP1_CTf,Word16#),
                                                 (forkHP1_CT2,Word16#),
                                                 (forkHP1_CT3,Word16#)] */
  logic [2:0] mergeHP_CTf_buf_emitted;
  logic [2:0] mergeHP_CTf_buf_done;
  assign forkHP1_CTf_d = {mergeHP_CTf_buf_d[16:1],
                          (mergeHP_CTf_buf_d[0] && (! mergeHP_CTf_buf_emitted[0]))};
  assign forkHP1_CT2_d = {mergeHP_CTf_buf_d[16:1],
                          (mergeHP_CTf_buf_d[0] && (! mergeHP_CTf_buf_emitted[1]))};
  assign forkHP1_CT3_d = {mergeHP_CTf_buf_d[16:1],
                          (mergeHP_CTf_buf_d[0] && (! mergeHP_CTf_buf_emitted[2]))};
  assign mergeHP_CTf_buf_done = (mergeHP_CTf_buf_emitted | ({forkHP1_CT3_d[0],
                                                             forkHP1_CT2_d[0],
                                                             forkHP1_CTf_d[0]} & {forkHP1_CT3_r,
                                                                                  forkHP1_CT2_r,
                                                                                  forkHP1_CTf_r}));
  assign mergeHP_CTf_buf_r = (& mergeHP_CTf_buf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_CTf_buf_emitted <= 3'd0;
    else
      mergeHP_CTf_buf_emitted <= (mergeHP_CTf_buf_r ? 3'd0 :
                                  mergeHP_CTf_buf_done);
  
  /* mergectrl (Ty C2,Ty MemIn_CTf) : [(dconReadIn_CTf,MemIn_CTf),
                                  (dconWriteIn_CTf,MemIn_CTf)] > (memMergeChoice_CTf,C2) (memMergeIn_CTf,MemIn_CTf) */
  logic [1:0] dconReadIn_CTf_select_d;
  assign dconReadIn_CTf_select_d = ((| dconReadIn_CTf_select_q) ? dconReadIn_CTf_select_q :
                                    (dconReadIn_CTf_d[0] ? 2'd1 :
                                     (dconWriteIn_CTf_d[0] ? 2'd2 :
                                      2'd0)));
  logic [1:0] dconReadIn_CTf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) dconReadIn_CTf_select_q <= 2'd0;
    else
      dconReadIn_CTf_select_q <= (dconReadIn_CTf_done ? 2'd0 :
                                  dconReadIn_CTf_select_d);
  logic [1:0] dconReadIn_CTf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) dconReadIn_CTf_emit_q <= 2'd0;
    else
      dconReadIn_CTf_emit_q <= (dconReadIn_CTf_done ? 2'd0 :
                                dconReadIn_CTf_emit_d);
  logic [1:0] dconReadIn_CTf_emit_d;
  assign dconReadIn_CTf_emit_d = (dconReadIn_CTf_emit_q | ({memMergeChoice_CTf_d[0],
                                                            memMergeIn_CTf_d[0]} & {memMergeChoice_CTf_r,
                                                                                    memMergeIn_CTf_r}));
  logic dconReadIn_CTf_done;
  assign dconReadIn_CTf_done = (& dconReadIn_CTf_emit_d);
  assign {dconWriteIn_CTf_r,
          dconReadIn_CTf_r} = (dconReadIn_CTf_done ? dconReadIn_CTf_select_d :
                               2'd0);
  assign memMergeIn_CTf_d = ((dconReadIn_CTf_select_d[0] && (! dconReadIn_CTf_emit_q[0])) ? dconReadIn_CTf_d :
                             ((dconReadIn_CTf_select_d[1] && (! dconReadIn_CTf_emit_q[0])) ? dconWriteIn_CTf_d :
                              {180'd0, 1'd0}));
  assign memMergeChoice_CTf_d = ((dconReadIn_CTf_select_d[0] && (! dconReadIn_CTf_emit_q[1])) ? C1_2_dc(1'd1) :
                                 ((dconReadIn_CTf_select_d[1] && (! dconReadIn_CTf_emit_q[1])) ? C2_2_dc(1'd1) :
                                  {1'd0, 1'd0}));
  
  /* bram (Ty MemIn_CTf,
      Ty MemOut_CTf) : (memMergeIn_CTf_dbuf,MemIn_CTf) > (memOut_CTf,MemOut_CTf) */
  logic [162:0] memMergeIn_CTf_dbuf_mem[65535:0];
  logic [15:0] memMergeIn_CTf_dbuf_address;
  logic [162:0] memMergeIn_CTf_dbuf_din;
  logic [162:0] memOut_CTf_q;
  logic memOut_CTf_valid;
  logic memMergeIn_CTf_dbuf_we;
  logic memOut_CTf_we;
  assign memMergeIn_CTf_dbuf_din = memMergeIn_CTf_dbuf_d[180:18];
  assign memMergeIn_CTf_dbuf_address = memMergeIn_CTf_dbuf_d[17:2];
  assign memMergeIn_CTf_dbuf_we = (memMergeIn_CTf_dbuf_d[1:1] && memMergeIn_CTf_dbuf_d[0]);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        memOut_CTf_we <= 1'd0;
        memOut_CTf_valid <= 1'd0;
      end
    else
      begin
        memOut_CTf_we <= memMergeIn_CTf_dbuf_we;
        memOut_CTf_valid <= memMergeIn_CTf_dbuf_d[0];
        if (memMergeIn_CTf_dbuf_we)
          begin
            memMergeIn_CTf_dbuf_mem[memMergeIn_CTf_dbuf_address] <= memMergeIn_CTf_dbuf_din;
            memOut_CTf_q <= memMergeIn_CTf_dbuf_din;
          end
        else
          memOut_CTf_q <= memMergeIn_CTf_dbuf_mem[memMergeIn_CTf_dbuf_address];
      end
  assign memOut_CTf_d = {memOut_CTf_q,
                         memOut_CTf_we,
                         memOut_CTf_valid};
  assign memMergeIn_CTf_dbuf_r = ((! memOut_CTf_valid) || memOut_CTf_r);
  logic [31:0] profiling_MemIn_CTf_read;
  logic [31:0] profiling_MemIn_CTf_write;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        profiling_MemIn_CTf_write <= 0;
        profiling_MemIn_CTf_read <= 0;
      end
    else
      if ((memMergeIn_CTf_dbuf_we == 1'd1))
        profiling_MemIn_CTf_write <= (profiling_MemIn_CTf_write + 1);
      else
        if ((memOut_CTf_valid == 1'd1))
          profiling_MemIn_CTf_read <= (profiling_MemIn_CTf_read + 1);
  
  /* demux (Ty C2,
       Ty MemOut_CTf) : (memMergeChoice_CTf,C2) (memOut_CTf_dbuf,MemOut_CTf) > [(memReadOut_CTf,MemOut_CTf),
                                                                                (memWriteOut_CTf,MemOut_CTf)] */
  logic [1:0] memOut_CTf_dbuf_onehotd;
  always_comb
    if ((memMergeChoice_CTf_d[0] && memOut_CTf_dbuf_d[0]))
      unique case (memMergeChoice_CTf_d[1:1])
        1'd0: memOut_CTf_dbuf_onehotd = 2'd1;
        1'd1: memOut_CTf_dbuf_onehotd = 2'd2;
        default: memOut_CTf_dbuf_onehotd = 2'd0;
      endcase
    else memOut_CTf_dbuf_onehotd = 2'd0;
  assign memReadOut_CTf_d = {memOut_CTf_dbuf_d[164:1],
                             memOut_CTf_dbuf_onehotd[0]};
  assign memWriteOut_CTf_d = {memOut_CTf_dbuf_d[164:1],
                              memOut_CTf_dbuf_onehotd[1]};
  assign memOut_CTf_dbuf_r = (| (memOut_CTf_dbuf_onehotd & {memWriteOut_CTf_r,
                                                            memReadOut_CTf_r}));
  assign memMergeChoice_CTf_r = memOut_CTf_dbuf_r;
  
  /* dbuf (Ty MemIn_CTf) : (memMergeIn_CTf_rbuf,MemIn_CTf) > (memMergeIn_CTf_dbuf,MemIn_CTf) */
  assign memMergeIn_CTf_rbuf_r = ((! memMergeIn_CTf_dbuf_d[0]) || memMergeIn_CTf_dbuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memMergeIn_CTf_dbuf_d <= {180'd0, 1'd0};
    else
      if (memMergeIn_CTf_rbuf_r)
        memMergeIn_CTf_dbuf_d <= memMergeIn_CTf_rbuf_d;
  
  /* rbuf (Ty MemIn_CTf) : (memMergeIn_CTf,MemIn_CTf) > (memMergeIn_CTf_rbuf,MemIn_CTf) */
  MemIn_CTf_t memMergeIn_CTf_buf;
  assign memMergeIn_CTf_r = (! memMergeIn_CTf_buf[0]);
  assign memMergeIn_CTf_rbuf_d = (memMergeIn_CTf_buf[0] ? memMergeIn_CTf_buf :
                                  memMergeIn_CTf_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memMergeIn_CTf_buf <= {180'd0, 1'd0};
    else
      if ((memMergeIn_CTf_rbuf_r && memMergeIn_CTf_buf[0]))
        memMergeIn_CTf_buf <= {180'd0, 1'd0};
      else if (((! memMergeIn_CTf_rbuf_r) && (! memMergeIn_CTf_buf[0])))
        memMergeIn_CTf_buf <= memMergeIn_CTf_d;
  
  /* dbuf (Ty MemOut_CTf) : (memOut_CTf_rbuf,MemOut_CTf) > (memOut_CTf_dbuf,MemOut_CTf) */
  assign memOut_CTf_rbuf_r = ((! memOut_CTf_dbuf_d[0]) || memOut_CTf_dbuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memOut_CTf_dbuf_d <= {164'd0, 1'd0};
    else if (memOut_CTf_rbuf_r) memOut_CTf_dbuf_d <= memOut_CTf_rbuf_d;
  
  /* rbuf (Ty MemOut_CTf) : (memOut_CTf,MemOut_CTf) > (memOut_CTf_rbuf,MemOut_CTf) */
  MemOut_CTf_t memOut_CTf_buf;
  assign memOut_CTf_r = (! memOut_CTf_buf[0]);
  assign memOut_CTf_rbuf_d = (memOut_CTf_buf[0] ? memOut_CTf_buf :
                              memOut_CTf_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memOut_CTf_buf <= {164'd0, 1'd0};
    else
      if ((memOut_CTf_rbuf_r && memOut_CTf_buf[0]))
        memOut_CTf_buf <= {164'd0, 1'd0};
      else if (((! memOut_CTf_rbuf_r) && (! memOut_CTf_buf[0])))
        memOut_CTf_buf <= memOut_CTf_d;
  
  /* destruct (Ty Pointer_CTf,
          Dcon Pointer_CTf) : (scfarg_0_1_argbuf,Pointer_CTf) > [(destructReadIn_CTf,Word16#)] */
  assign destructReadIn_CTf_d = {scfarg_0_1_argbuf_d[16:1],
                                 scfarg_0_1_argbuf_d[0]};
  assign scfarg_0_1_argbuf_r = destructReadIn_CTf_r;
  
  /* dcon (Ty MemIn_CTf,
      Dcon ReadIn_CTf) : [(destructReadIn_CTf,Word16#)] > (dconReadIn_CTf,MemIn_CTf) */
  assign dconReadIn_CTf_d = ReadIn_CTf_dc((& {destructReadIn_CTf_d[0]}), destructReadIn_CTf_d);
  assign {destructReadIn_CTf_r} = {1 {(dconReadIn_CTf_r && dconReadIn_CTf_d[0])}};
  
  /* destruct (Ty MemOut_CTf,
          Dcon ReadOut_CTf) : (memReadOut_CTf,MemOut_CTf) > [(readPointer_CTfscfarg_0_1_argbuf,CTf)] */
  assign readPointer_CTfscfarg_0_1_argbuf_d = {memReadOut_CTf_d[164:2],
                                               memReadOut_CTf_d[0]};
  assign memReadOut_CTf_r = readPointer_CTfscfarg_0_1_argbuf_r;
  
  /* mergectrl (Ty C5,Ty CTf) : [(lizzieLet17_1_1_argbuf,CTf),
                            (lizzieLet39_1_argbuf,CTf),
                            (lizzieLet44_1_argbuf,CTf),
                            (lizzieLet45_1_argbuf,CTf),
                            (lizzieLet46_1_argbuf,CTf)] > (writeMerge_choice_CTf,C5) (writeMerge_data_CTf,CTf) */
  logic [4:0] lizzieLet17_1_1_argbuf_select_d;
  assign lizzieLet17_1_1_argbuf_select_d = ((| lizzieLet17_1_1_argbuf_select_q) ? lizzieLet17_1_1_argbuf_select_q :
                                            (lizzieLet17_1_1_argbuf_d[0] ? 5'd1 :
                                             (lizzieLet39_1_argbuf_d[0] ? 5'd2 :
                                              (lizzieLet44_1_argbuf_d[0] ? 5'd4 :
                                               (lizzieLet45_1_argbuf_d[0] ? 5'd8 :
                                                (lizzieLet46_1_argbuf_d[0] ? 5'd16 :
                                                 5'd0))))));
  logic [4:0] lizzieLet17_1_1_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet17_1_1_argbuf_select_q <= 5'd0;
    else
      lizzieLet17_1_1_argbuf_select_q <= (lizzieLet17_1_1_argbuf_done ? 5'd0 :
                                          lizzieLet17_1_1_argbuf_select_d);
  logic [1:0] lizzieLet17_1_1_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet17_1_1_argbuf_emit_q <= 2'd0;
    else
      lizzieLet17_1_1_argbuf_emit_q <= (lizzieLet17_1_1_argbuf_done ? 2'd0 :
                                        lizzieLet17_1_1_argbuf_emit_d);
  logic [1:0] lizzieLet17_1_1_argbuf_emit_d;
  assign lizzieLet17_1_1_argbuf_emit_d = (lizzieLet17_1_1_argbuf_emit_q | ({writeMerge_choice_CTf_d[0],
                                                                            writeMerge_data_CTf_d[0]} & {writeMerge_choice_CTf_r,
                                                                                                         writeMerge_data_CTf_r}));
  logic lizzieLet17_1_1_argbuf_done;
  assign lizzieLet17_1_1_argbuf_done = (& lizzieLet17_1_1_argbuf_emit_d);
  assign {lizzieLet46_1_argbuf_r,
          lizzieLet45_1_argbuf_r,
          lizzieLet44_1_argbuf_r,
          lizzieLet39_1_argbuf_r,
          lizzieLet17_1_1_argbuf_r} = (lizzieLet17_1_1_argbuf_done ? lizzieLet17_1_1_argbuf_select_d :
                                       5'd0);
  assign writeMerge_data_CTf_d = ((lizzieLet17_1_1_argbuf_select_d[0] && (! lizzieLet17_1_1_argbuf_emit_q[0])) ? lizzieLet17_1_1_argbuf_d :
                                  ((lizzieLet17_1_1_argbuf_select_d[1] && (! lizzieLet17_1_1_argbuf_emit_q[0])) ? lizzieLet39_1_argbuf_d :
                                   ((lizzieLet17_1_1_argbuf_select_d[2] && (! lizzieLet17_1_1_argbuf_emit_q[0])) ? lizzieLet44_1_argbuf_d :
                                    ((lizzieLet17_1_1_argbuf_select_d[3] && (! lizzieLet17_1_1_argbuf_emit_q[0])) ? lizzieLet45_1_argbuf_d :
                                     ((lizzieLet17_1_1_argbuf_select_d[4] && (! lizzieLet17_1_1_argbuf_emit_q[0])) ? lizzieLet46_1_argbuf_d :
                                      {163'd0, 1'd0})))));
  assign writeMerge_choice_CTf_d = ((lizzieLet17_1_1_argbuf_select_d[0] && (! lizzieLet17_1_1_argbuf_emit_q[1])) ? C1_5_dc(1'd1) :
                                    ((lizzieLet17_1_1_argbuf_select_d[1] && (! lizzieLet17_1_1_argbuf_emit_q[1])) ? C2_5_dc(1'd1) :
                                     ((lizzieLet17_1_1_argbuf_select_d[2] && (! lizzieLet17_1_1_argbuf_emit_q[1])) ? C3_5_dc(1'd1) :
                                      ((lizzieLet17_1_1_argbuf_select_d[3] && (! lizzieLet17_1_1_argbuf_emit_q[1])) ? C4_5_dc(1'd1) :
                                       ((lizzieLet17_1_1_argbuf_select_d[4] && (! lizzieLet17_1_1_argbuf_emit_q[1])) ? C5_5_dc(1'd1) :
                                        {3'd0, 1'd0})))));
  
  /* demux (Ty C5,
       Ty Pointer_CTf) : (writeMerge_choice_CTf,C5) (demuxWriteResult_CTf,Pointer_CTf) > [(writeCTflizzieLet17_1_1_argbuf,Pointer_CTf),
                                                                                          (writeCTflizzieLet39_1_argbuf,Pointer_CTf),
                                                                                          (writeCTflizzieLet44_1_argbuf,Pointer_CTf),
                                                                                          (writeCTflizzieLet45_1_argbuf,Pointer_CTf),
                                                                                          (writeCTflizzieLet46_1_argbuf,Pointer_CTf)] */
  logic [4:0] demuxWriteResult_CTf_onehotd;
  always_comb
    if ((writeMerge_choice_CTf_d[0] && demuxWriteResult_CTf_d[0]))
      unique case (writeMerge_choice_CTf_d[3:1])
        3'd0: demuxWriteResult_CTf_onehotd = 5'd1;
        3'd1: demuxWriteResult_CTf_onehotd = 5'd2;
        3'd2: demuxWriteResult_CTf_onehotd = 5'd4;
        3'd3: demuxWriteResult_CTf_onehotd = 5'd8;
        3'd4: demuxWriteResult_CTf_onehotd = 5'd16;
        default: demuxWriteResult_CTf_onehotd = 5'd0;
      endcase
    else demuxWriteResult_CTf_onehotd = 5'd0;
  assign writeCTflizzieLet17_1_1_argbuf_d = {demuxWriteResult_CTf_d[16:1],
                                             demuxWriteResult_CTf_onehotd[0]};
  assign writeCTflizzieLet39_1_argbuf_d = {demuxWriteResult_CTf_d[16:1],
                                           demuxWriteResult_CTf_onehotd[1]};
  assign writeCTflizzieLet44_1_argbuf_d = {demuxWriteResult_CTf_d[16:1],
                                           demuxWriteResult_CTf_onehotd[2]};
  assign writeCTflizzieLet45_1_argbuf_d = {demuxWriteResult_CTf_d[16:1],
                                           demuxWriteResult_CTf_onehotd[3]};
  assign writeCTflizzieLet46_1_argbuf_d = {demuxWriteResult_CTf_d[16:1],
                                           demuxWriteResult_CTf_onehotd[4]};
  assign demuxWriteResult_CTf_r = (| (demuxWriteResult_CTf_onehotd & {writeCTflizzieLet46_1_argbuf_r,
                                                                      writeCTflizzieLet45_1_argbuf_r,
                                                                      writeCTflizzieLet44_1_argbuf_r,
                                                                      writeCTflizzieLet39_1_argbuf_r,
                                                                      writeCTflizzieLet17_1_1_argbuf_r}));
  assign writeMerge_choice_CTf_r = demuxWriteResult_CTf_r;
  
  /* dcon (Ty MemIn_CTf,Dcon WriteIn_CTf) : [(forkHP1_CT2,Word16#),
                                        (writeMerge_data_CTf,CTf)] > (dconWriteIn_CTf,MemIn_CTf) */
  assign dconWriteIn_CTf_d = WriteIn_CTf_dc((& {forkHP1_CT2_d[0],
                                                writeMerge_data_CTf_d[0]}), forkHP1_CT2_d, writeMerge_data_CTf_d);
  assign {forkHP1_CT2_r,
          writeMerge_data_CTf_r} = {2 {(dconWriteIn_CTf_r && dconWriteIn_CTf_d[0])}};
  
  /* dcon (Ty Pointer_CTf,
      Dcon Pointer_CTf) : [(forkHP1_CT3,Word16#)] > (dconPtr_CTf,Pointer_CTf) */
  assign dconPtr_CTf_d = Pointer_CTf_dc((& {forkHP1_CT3_d[0]}), forkHP1_CT3_d);
  assign {forkHP1_CT3_r} = {1 {(dconPtr_CTf_r && dconPtr_CTf_d[0])}};
  
  /* demux (Ty MemOut_CTf,
       Ty Pointer_CTf) : (memWriteOut_CTf,MemOut_CTf) (dconPtr_CTf,Pointer_CTf) > [(_129,Pointer_CTf),
                                                                                   (demuxWriteResult_CTf,Pointer_CTf)] */
  logic [1:0] dconPtr_CTf_onehotd;
  always_comb
    if ((memWriteOut_CTf_d[0] && dconPtr_CTf_d[0]))
      unique case (memWriteOut_CTf_d[1:1])
        1'd0: dconPtr_CTf_onehotd = 2'd1;
        1'd1: dconPtr_CTf_onehotd = 2'd2;
        default: dconPtr_CTf_onehotd = 2'd0;
      endcase
    else dconPtr_CTf_onehotd = 2'd0;
  assign _129_d = {dconPtr_CTf_d[16:1], dconPtr_CTf_onehotd[0]};
  assign demuxWriteResult_CTf_d = {dconPtr_CTf_d[16:1],
                                   dconPtr_CTf_onehotd[1]};
  assign dconPtr_CTf_r = (| (dconPtr_CTf_onehotd & {demuxWriteResult_CTf_r,
                                                    _129_r}));
  assign memWriteOut_CTf_r = dconPtr_CTf_r;
  
  /* const (Ty Word16#,Lit 0) : (goFor_4,Go) > (initHP_CTf',Word16#) */
  assign \initHP_CTf'_d  = {16'd0, goFor_4_d[0]};
  assign goFor_4_r = \initHP_CTf'_r ;
  
  /* const (Ty Word16#,
       Lit 1) : (incrHP_CTf'1,Go) > (incrHP_CTf',Word16#) */
  assign \incrHP_CTf'_d  = {16'd1, \incrHP_CTf'1_d [0]};
  assign \incrHP_CTf'1_r  = \incrHP_CTf'_r ;
  
  /* merge (Ty Go) : [(goFor_5,Go),
                 (incrHP_CTf'2,Go)] > (incrHP_mergeCTf',Go) */
  logic [1:0] \incrHP_mergeCTf'_selected ;
  logic [1:0] \incrHP_mergeCTf'_select ;
  always_comb
    begin
      \incrHP_mergeCTf'_selected  = 2'd0;
      if ((| \incrHP_mergeCTf'_select ))
        \incrHP_mergeCTf'_selected  = \incrHP_mergeCTf'_select ;
      else
        if (goFor_5_d[0]) \incrHP_mergeCTf'_selected [0] = 1'd1;
        else if (\incrHP_CTf'2_d [0])
          \incrHP_mergeCTf'_selected [1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \incrHP_mergeCTf'_select  <= 2'd0;
    else
      \incrHP_mergeCTf'_select  <= (\incrHP_mergeCTf'_r  ? 2'd0 :
                                    \incrHP_mergeCTf'_selected );
  always_comb
    if (\incrHP_mergeCTf'_selected [0])
      \incrHP_mergeCTf'_d  = goFor_5_d;
    else if (\incrHP_mergeCTf'_selected [1])
      \incrHP_mergeCTf'_d  = \incrHP_CTf'2_d ;
    else \incrHP_mergeCTf'_d  = 1'd0;
  assign {\incrHP_CTf'2_r ,
          goFor_5_r} = (\incrHP_mergeCTf'_r  ? \incrHP_mergeCTf'_selected  :
                        2'd0);
  
  /* fork (Ty Go) : (incrHP_mergeCTf'_buf,Go) > [(incrHP_CTf'1,Go),
                                            (incrHP_CTf'2,Go)] */
  logic [1:0] \incrHP_mergeCTf'_buf_emitted ;
  logic [1:0] \incrHP_mergeCTf'_buf_done ;
  assign \incrHP_CTf'1_d  = (\incrHP_mergeCTf'_buf_d [0] && (! \incrHP_mergeCTf'_buf_emitted [0]));
  assign \incrHP_CTf'2_d  = (\incrHP_mergeCTf'_buf_d [0] && (! \incrHP_mergeCTf'_buf_emitted [1]));
  assign \incrHP_mergeCTf'_buf_done  = (\incrHP_mergeCTf'_buf_emitted  | ({\incrHP_CTf'2_d [0],
                                                                           \incrHP_CTf'1_d [0]} & {\incrHP_CTf'2_r ,
                                                                                                   \incrHP_CTf'1_r }));
  assign \incrHP_mergeCTf'_buf_r  = (& \incrHP_mergeCTf'_buf_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \incrHP_mergeCTf'_buf_emitted  <= 2'd0;
    else
      \incrHP_mergeCTf'_buf_emitted  <= (\incrHP_mergeCTf'_buf_r  ? 2'd0 :
                                         \incrHP_mergeCTf'_buf_done );
  
  /* op_add (Ty Word16#) : (incrHP_CTf',Word16#) (forkHP1_CTf',Word16#) > (addHP_CTf',Word16#) */
  assign \addHP_CTf'_d  = {(\incrHP_CTf'_d [16:1] + \forkHP1_CTf'_d [16:1]),
                           (\incrHP_CTf'_d [0] && \forkHP1_CTf'_d [0])};
  assign {\incrHP_CTf'_r ,
          \forkHP1_CTf'_r } = {2 {(\addHP_CTf'_r  && \addHP_CTf'_d [0])}};
  
  /* merge (Ty Word16#) : [(initHP_CTf',Word16#),
                      (addHP_CTf',Word16#)] > (mergeHP_CTf',Word16#) */
  logic [1:0] \mergeHP_CTf'_selected ;
  logic [1:0] \mergeHP_CTf'_select ;
  always_comb
    begin
      \mergeHP_CTf'_selected  = 2'd0;
      if ((| \mergeHP_CTf'_select ))
        \mergeHP_CTf'_selected  = \mergeHP_CTf'_select ;
      else
        if (\initHP_CTf'_d [0]) \mergeHP_CTf'_selected [0] = 1'd1;
        else if (\addHP_CTf'_d [0]) \mergeHP_CTf'_selected [1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \mergeHP_CTf'_select  <= 2'd0;
    else
      \mergeHP_CTf'_select  <= (\mergeHP_CTf'_r  ? 2'd0 :
                                \mergeHP_CTf'_selected );
  always_comb
    if (\mergeHP_CTf'_selected [0]) \mergeHP_CTf'_d  = \initHP_CTf'_d ;
    else if (\mergeHP_CTf'_selected [1])
      \mergeHP_CTf'_d  = \addHP_CTf'_d ;
    else \mergeHP_CTf'_d  = {16'd0, 1'd0};
  assign {\addHP_CTf'_r ,
          \initHP_CTf'_r } = (\mergeHP_CTf'_r  ? \mergeHP_CTf'_selected  :
                              2'd0);
  
  /* buf (Ty Go) : (incrHP_mergeCTf',Go) > (incrHP_mergeCTf'_buf,Go) */
  Go_t \incrHP_mergeCTf'_bufchan_d ;
  logic \incrHP_mergeCTf'_bufchan_r ;
  assign \incrHP_mergeCTf'_r  = ((! \incrHP_mergeCTf'_bufchan_d [0]) || \incrHP_mergeCTf'_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \incrHP_mergeCTf'_bufchan_d  <= 1'd0;
    else
      if (\incrHP_mergeCTf'_r )
        \incrHP_mergeCTf'_bufchan_d  <= \incrHP_mergeCTf'_d ;
  Go_t \incrHP_mergeCTf'_bufchan_buf ;
  assign \incrHP_mergeCTf'_bufchan_r  = (! \incrHP_mergeCTf'_bufchan_buf [0]);
  assign \incrHP_mergeCTf'_buf_d  = (\incrHP_mergeCTf'_bufchan_buf [0] ? \incrHP_mergeCTf'_bufchan_buf  :
                                     \incrHP_mergeCTf'_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \incrHP_mergeCTf'_bufchan_buf  <= 1'd0;
    else
      if ((\incrHP_mergeCTf'_buf_r  && \incrHP_mergeCTf'_bufchan_buf [0]))
        \incrHP_mergeCTf'_bufchan_buf  <= 1'd0;
      else if (((! \incrHP_mergeCTf'_buf_r ) && (! \incrHP_mergeCTf'_bufchan_buf [0])))
        \incrHP_mergeCTf'_bufchan_buf  <= \incrHP_mergeCTf'_bufchan_d ;
  
  /* buf (Ty Word16#) : (mergeHP_CTf',Word16#) > (mergeHP_CTf'_buf,Word16#) */
  \Word16#_t  \mergeHP_CTf'_bufchan_d ;
  logic \mergeHP_CTf'_bufchan_r ;
  assign \mergeHP_CTf'_r  = ((! \mergeHP_CTf'_bufchan_d [0]) || \mergeHP_CTf'_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \mergeHP_CTf'_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\mergeHP_CTf'_r ) \mergeHP_CTf'_bufchan_d  <= \mergeHP_CTf'_d ;
  \Word16#_t  \mergeHP_CTf'_bufchan_buf ;
  assign \mergeHP_CTf'_bufchan_r  = (! \mergeHP_CTf'_bufchan_buf [0]);
  assign \mergeHP_CTf'_buf_d  = (\mergeHP_CTf'_bufchan_buf [0] ? \mergeHP_CTf'_bufchan_buf  :
                                 \mergeHP_CTf'_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \mergeHP_CTf'_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((\mergeHP_CTf'_buf_r  && \mergeHP_CTf'_bufchan_buf [0]))
        \mergeHP_CTf'_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! \mergeHP_CTf'_buf_r ) && (! \mergeHP_CTf'_bufchan_buf [0])))
        \mergeHP_CTf'_bufchan_buf  <= \mergeHP_CTf'_bufchan_d ;
  
  /* fork (Ty Word16#) : (mergeHP_CTf'_buf,Word16#) > [(forkHP1_CTf',Word16#),
                                                  (forkHP1_CTf2,Word16#),
                                                  (forkHP1_CTf3,Word16#)] */
  logic [2:0] \mergeHP_CTf'_buf_emitted ;
  logic [2:0] \mergeHP_CTf'_buf_done ;
  assign \forkHP1_CTf'_d  = {\mergeHP_CTf'_buf_d [16:1],
                             (\mergeHP_CTf'_buf_d [0] && (! \mergeHP_CTf'_buf_emitted [0]))};
  assign forkHP1_CTf2_d = {\mergeHP_CTf'_buf_d [16:1],
                           (\mergeHP_CTf'_buf_d [0] && (! \mergeHP_CTf'_buf_emitted [1]))};
  assign forkHP1_CTf3_d = {\mergeHP_CTf'_buf_d [16:1],
                           (\mergeHP_CTf'_buf_d [0] && (! \mergeHP_CTf'_buf_emitted [2]))};
  assign \mergeHP_CTf'_buf_done  = (\mergeHP_CTf'_buf_emitted  | ({forkHP1_CTf3_d[0],
                                                                   forkHP1_CTf2_d[0],
                                                                   \forkHP1_CTf'_d [0]} & {forkHP1_CTf3_r,
                                                                                           forkHP1_CTf2_r,
                                                                                           \forkHP1_CTf'_r }));
  assign \mergeHP_CTf'_buf_r  = (& \mergeHP_CTf'_buf_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \mergeHP_CTf'_buf_emitted  <= 3'd0;
    else
      \mergeHP_CTf'_buf_emitted  <= (\mergeHP_CTf'_buf_r  ? 3'd0 :
                                     \mergeHP_CTf'_buf_done );
  
  /* mergectrl (Ty C2,Ty MemIn_CTf') : [(dconReadIn_CTf',MemIn_CTf'),
                                   (dconWriteIn_CTf',MemIn_CTf')] > (memMergeChoice_CTf',C2) (memMergeIn_CTf',MemIn_CTf') */
  logic [1:0] \dconReadIn_CTf'_select_d ;
  assign \dconReadIn_CTf'_select_d  = ((| \dconReadIn_CTf'_select_q ) ? \dconReadIn_CTf'_select_q  :
                                       (\dconReadIn_CTf'_d [0] ? 2'd1 :
                                        (\dconWriteIn_CTf'_d [0] ? 2'd2 :
                                         2'd0)));
  logic [1:0] \dconReadIn_CTf'_select_q ;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \dconReadIn_CTf'_select_q  <= 2'd0;
    else
      \dconReadIn_CTf'_select_q  <= (\dconReadIn_CTf'_done  ? 2'd0 :
                                     \dconReadIn_CTf'_select_d );
  logic [1:0] \dconReadIn_CTf'_emit_q ;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \dconReadIn_CTf'_emit_q  <= 2'd0;
    else
      \dconReadIn_CTf'_emit_q  <= (\dconReadIn_CTf'_done  ? 2'd0 :
                                   \dconReadIn_CTf'_emit_d );
  logic [1:0] \dconReadIn_CTf'_emit_d ;
  assign \dconReadIn_CTf'_emit_d  = (\dconReadIn_CTf'_emit_q  | ({\memMergeChoice_CTf'_d [0],
                                                                  \memMergeIn_CTf'_d [0]} & {\memMergeChoice_CTf'_r ,
                                                                                             \memMergeIn_CTf'_r }));
  logic \dconReadIn_CTf'_done ;
  assign \dconReadIn_CTf'_done  = (& \dconReadIn_CTf'_emit_d );
  assign {\dconWriteIn_CTf'_r ,
          \dconReadIn_CTf'_r } = (\dconReadIn_CTf'_done  ? \dconReadIn_CTf'_select_d  :
                                  2'd0);
  assign \memMergeIn_CTf'_d  = ((\dconReadIn_CTf'_select_d [0] && (! \dconReadIn_CTf'_emit_q [0])) ? \dconReadIn_CTf'_d  :
                                ((\dconReadIn_CTf'_select_d [1] && (! \dconReadIn_CTf'_emit_q [0])) ? \dconWriteIn_CTf'_d  :
                                 {132'd0, 1'd0}));
  assign \memMergeChoice_CTf'_d  = ((\dconReadIn_CTf'_select_d [0] && (! \dconReadIn_CTf'_emit_q [1])) ? C1_2_dc(1'd1) :
                                    ((\dconReadIn_CTf'_select_d [1] && (! \dconReadIn_CTf'_emit_q [1])) ? C2_2_dc(1'd1) :
                                     {1'd0, 1'd0}));
  
  /* bram (Ty MemIn_CTf',
      Ty MemOut_CTf') : (memMergeIn_CTf'_dbuf,MemIn_CTf') > (memOut_CTf',MemOut_CTf') */
  logic [114:0] \memMergeIn_CTf'_dbuf_mem [65535:0];
  logic [15:0] \memMergeIn_CTf'_dbuf_address ;
  logic [114:0] \memMergeIn_CTf'_dbuf_din ;
  logic [114:0] \memOut_CTf'_q ;
  logic \memOut_CTf'_valid ;
  logic \memMergeIn_CTf'_dbuf_we ;
  logic \memOut_CTf'_we ;
  assign \memMergeIn_CTf'_dbuf_din  = \memMergeIn_CTf'_dbuf_d [132:18];
  assign \memMergeIn_CTf'_dbuf_address  = \memMergeIn_CTf'_dbuf_d [17:2];
  assign \memMergeIn_CTf'_dbuf_we  = (\memMergeIn_CTf'_dbuf_d [1:1] && \memMergeIn_CTf'_dbuf_d [0]);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        \memOut_CTf'_we  <= 1'd0;
        \memOut_CTf'_valid  <= 1'd0;
      end
    else
      begin
        \memOut_CTf'_we  <= \memMergeIn_CTf'_dbuf_we ;
        \memOut_CTf'_valid  <= \memMergeIn_CTf'_dbuf_d [0];
        if (\memMergeIn_CTf'_dbuf_we )
          begin
            \memMergeIn_CTf'_dbuf_mem [\memMergeIn_CTf'_dbuf_address ] <= \memMergeIn_CTf'_dbuf_din ;
            \memOut_CTf'_q  <= \memMergeIn_CTf'_dbuf_din ;
          end
        else
          \memOut_CTf'_q  <= \memMergeIn_CTf'_dbuf_mem [\memMergeIn_CTf'_dbuf_address ];
      end
  assign \memOut_CTf'_d  = {\memOut_CTf'_q ,
                            \memOut_CTf'_we ,
                            \memOut_CTf'_valid };
  assign \memMergeIn_CTf'_dbuf_r  = ((! \memOut_CTf'_valid ) || \memOut_CTf'_r );
  logic [31:0] \profiling_MemIn_CTf'_read ;
  logic [31:0] \profiling_MemIn_CTf'_write ;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        \profiling_MemIn_CTf'_write  <= 0;
        \profiling_MemIn_CTf'_read  <= 0;
      end
    else
      if ((\memMergeIn_CTf'_dbuf_we  == 1'd1))
        \profiling_MemIn_CTf'_write  <= (\profiling_MemIn_CTf'_write  + 1);
      else
        if ((\memOut_CTf'_valid  == 1'd1))
          \profiling_MemIn_CTf'_read  <= (\profiling_MemIn_CTf'_read  + 1);
  
  /* demux (Ty C2,
       Ty MemOut_CTf') : (memMergeChoice_CTf',C2) (memOut_CTf'_dbuf,MemOut_CTf') > [(memReadOut_CTf',MemOut_CTf'),
                                                                                    (memWriteOut_CTf',MemOut_CTf')] */
  logic [1:0] \memOut_CTf'_dbuf_onehotd ;
  always_comb
    if ((\memMergeChoice_CTf'_d [0] && \memOut_CTf'_dbuf_d [0]))
      unique case (\memMergeChoice_CTf'_d [1:1])
        1'd0: \memOut_CTf'_dbuf_onehotd  = 2'd1;
        1'd1: \memOut_CTf'_dbuf_onehotd  = 2'd2;
        default: \memOut_CTf'_dbuf_onehotd  = 2'd0;
      endcase
    else \memOut_CTf'_dbuf_onehotd  = 2'd0;
  assign \memReadOut_CTf'_d  = {\memOut_CTf'_dbuf_d [116:1],
                                \memOut_CTf'_dbuf_onehotd [0]};
  assign \memWriteOut_CTf'_d  = {\memOut_CTf'_dbuf_d [116:1],
                                 \memOut_CTf'_dbuf_onehotd [1]};
  assign \memOut_CTf'_dbuf_r  = (| (\memOut_CTf'_dbuf_onehotd  & {\memWriteOut_CTf'_r ,
                                                                  \memReadOut_CTf'_r }));
  assign \memMergeChoice_CTf'_r  = \memOut_CTf'_dbuf_r ;
  
  /* dbuf (Ty MemIn_CTf') : (memMergeIn_CTf'_rbuf,MemIn_CTf') > (memMergeIn_CTf'_dbuf,MemIn_CTf') */
  assign \memMergeIn_CTf'_rbuf_r  = ((! \memMergeIn_CTf'_dbuf_d [0]) || \memMergeIn_CTf'_dbuf_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \memMergeIn_CTf'_dbuf_d  <= {132'd0, 1'd0};
    else
      if (\memMergeIn_CTf'_rbuf_r )
        \memMergeIn_CTf'_dbuf_d  <= \memMergeIn_CTf'_rbuf_d ;
  
  /* rbuf (Ty MemIn_CTf') : (memMergeIn_CTf',MemIn_CTf') > (memMergeIn_CTf'_rbuf,MemIn_CTf') */
  \MemIn_CTf'_t  \memMergeIn_CTf'_buf ;
  assign \memMergeIn_CTf'_r  = (! \memMergeIn_CTf'_buf [0]);
  assign \memMergeIn_CTf'_rbuf_d  = (\memMergeIn_CTf'_buf [0] ? \memMergeIn_CTf'_buf  :
                                     \memMergeIn_CTf'_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \memMergeIn_CTf'_buf  <= {132'd0, 1'd0};
    else
      if ((\memMergeIn_CTf'_rbuf_r  && \memMergeIn_CTf'_buf [0]))
        \memMergeIn_CTf'_buf  <= {132'd0, 1'd0};
      else if (((! \memMergeIn_CTf'_rbuf_r ) && (! \memMergeIn_CTf'_buf [0])))
        \memMergeIn_CTf'_buf  <= \memMergeIn_CTf'_d ;
  
  /* dbuf (Ty MemOut_CTf') : (memOut_CTf'_rbuf,MemOut_CTf') > (memOut_CTf'_dbuf,MemOut_CTf') */
  assign \memOut_CTf'_rbuf_r  = ((! \memOut_CTf'_dbuf_d [0]) || \memOut_CTf'_dbuf_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \memOut_CTf'_dbuf_d  <= {116'd0, 1'd0};
    else
      if (\memOut_CTf'_rbuf_r )
        \memOut_CTf'_dbuf_d  <= \memOut_CTf'_rbuf_d ;
  
  /* rbuf (Ty MemOut_CTf') : (memOut_CTf',MemOut_CTf') > (memOut_CTf'_rbuf,MemOut_CTf') */
  \MemOut_CTf'_t  \memOut_CTf'_buf ;
  assign \memOut_CTf'_r  = (! \memOut_CTf'_buf [0]);
  assign \memOut_CTf'_rbuf_d  = (\memOut_CTf'_buf [0] ? \memOut_CTf'_buf  :
                                 \memOut_CTf'_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \memOut_CTf'_buf  <= {116'd0, 1'd0};
    else
      if ((\memOut_CTf'_rbuf_r  && \memOut_CTf'_buf [0]))
        \memOut_CTf'_buf  <= {116'd0, 1'd0};
      else if (((! \memOut_CTf'_rbuf_r ) && (! \memOut_CTf'_buf [0])))
        \memOut_CTf'_buf  <= \memOut_CTf'_d ;
  
  /* destruct (Ty Pointer_CTf',
          Dcon Pointer_CTf') : (scfarg_0_1_1_argbuf,Pointer_CTf') > [(destructReadIn_CTf',Word16#)] */
  assign \destructReadIn_CTf'_d  = {scfarg_0_1_1_argbuf_d[16:1],
                                    scfarg_0_1_1_argbuf_d[0]};
  assign scfarg_0_1_1_argbuf_r = \destructReadIn_CTf'_r ;
  
  /* dcon (Ty MemIn_CTf',
      Dcon ReadIn_CTf') : [(destructReadIn_CTf',Word16#)] > (dconReadIn_CTf',MemIn_CTf') */
  assign \dconReadIn_CTf'_d  = \ReadIn_CTf'_dc ((& {\destructReadIn_CTf'_d [0]}), \destructReadIn_CTf'_d );
  assign {\destructReadIn_CTf'_r } = {1 {(\dconReadIn_CTf'_r  && \dconReadIn_CTf'_d [0])}};
  
  /* destruct (Ty MemOut_CTf',
          Dcon ReadOut_CTf') : (memReadOut_CTf',MemOut_CTf') > [(readPointer_CTf'scfarg_0_1_1_argbuf,CTf')] */
  assign \readPointer_CTf'scfarg_0_1_1_argbuf_d  = {\memReadOut_CTf'_d [116:2],
                                                    \memReadOut_CTf'_d [0]};
  assign \memReadOut_CTf'_r  = \readPointer_CTf'scfarg_0_1_1_argbuf_r ;
  
  /* mergectrl (Ty C5,Ty CTf') : [(lizzieLet29_1_argbuf,CTf'),
                             (lizzieLet40_1_argbuf,CTf'),
                             (lizzieLet49_1_argbuf,CTf'),
                             (lizzieLet50_1_argbuf,CTf'),
                             (lizzieLet51_1_argbuf,CTf')] > (writeMerge_choice_CTf',C5) (writeMerge_data_CTf',CTf') */
  logic [4:0] lizzieLet29_1_argbuf_select_d;
  assign lizzieLet29_1_argbuf_select_d = ((| lizzieLet29_1_argbuf_select_q) ? lizzieLet29_1_argbuf_select_q :
                                          (lizzieLet29_1_argbuf_d[0] ? 5'd1 :
                                           (lizzieLet40_1_argbuf_d[0] ? 5'd2 :
                                            (lizzieLet49_1_argbuf_d[0] ? 5'd4 :
                                             (lizzieLet50_1_argbuf_d[0] ? 5'd8 :
                                              (lizzieLet51_1_argbuf_d[0] ? 5'd16 :
                                               5'd0))))));
  logic [4:0] lizzieLet29_1_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet29_1_argbuf_select_q <= 5'd0;
    else
      lizzieLet29_1_argbuf_select_q <= (lizzieLet29_1_argbuf_done ? 5'd0 :
                                        lizzieLet29_1_argbuf_select_d);
  logic [1:0] lizzieLet29_1_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet29_1_argbuf_emit_q <= 2'd0;
    else
      lizzieLet29_1_argbuf_emit_q <= (lizzieLet29_1_argbuf_done ? 2'd0 :
                                      lizzieLet29_1_argbuf_emit_d);
  logic [1:0] lizzieLet29_1_argbuf_emit_d;
  assign lizzieLet29_1_argbuf_emit_d = (lizzieLet29_1_argbuf_emit_q | ({\writeMerge_choice_CTf'_d [0],
                                                                        \writeMerge_data_CTf'_d [0]} & {\writeMerge_choice_CTf'_r ,
                                                                                                        \writeMerge_data_CTf'_r }));
  logic lizzieLet29_1_argbuf_done;
  assign lizzieLet29_1_argbuf_done = (& lizzieLet29_1_argbuf_emit_d);
  assign {lizzieLet51_1_argbuf_r,
          lizzieLet50_1_argbuf_r,
          lizzieLet49_1_argbuf_r,
          lizzieLet40_1_argbuf_r,
          lizzieLet29_1_argbuf_r} = (lizzieLet29_1_argbuf_done ? lizzieLet29_1_argbuf_select_d :
                                     5'd0);
  assign \writeMerge_data_CTf'_d  = ((lizzieLet29_1_argbuf_select_d[0] && (! lizzieLet29_1_argbuf_emit_q[0])) ? lizzieLet29_1_argbuf_d :
                                     ((lizzieLet29_1_argbuf_select_d[1] && (! lizzieLet29_1_argbuf_emit_q[0])) ? lizzieLet40_1_argbuf_d :
                                      ((lizzieLet29_1_argbuf_select_d[2] && (! lizzieLet29_1_argbuf_emit_q[0])) ? lizzieLet49_1_argbuf_d :
                                       ((lizzieLet29_1_argbuf_select_d[3] && (! lizzieLet29_1_argbuf_emit_q[0])) ? lizzieLet50_1_argbuf_d :
                                        ((lizzieLet29_1_argbuf_select_d[4] && (! lizzieLet29_1_argbuf_emit_q[0])) ? lizzieLet51_1_argbuf_d :
                                         {115'd0, 1'd0})))));
  assign \writeMerge_choice_CTf'_d  = ((lizzieLet29_1_argbuf_select_d[0] && (! lizzieLet29_1_argbuf_emit_q[1])) ? C1_5_dc(1'd1) :
                                       ((lizzieLet29_1_argbuf_select_d[1] && (! lizzieLet29_1_argbuf_emit_q[1])) ? C2_5_dc(1'd1) :
                                        ((lizzieLet29_1_argbuf_select_d[2] && (! lizzieLet29_1_argbuf_emit_q[1])) ? C3_5_dc(1'd1) :
                                         ((lizzieLet29_1_argbuf_select_d[3] && (! lizzieLet29_1_argbuf_emit_q[1])) ? C4_5_dc(1'd1) :
                                          ((lizzieLet29_1_argbuf_select_d[4] && (! lizzieLet29_1_argbuf_emit_q[1])) ? C5_5_dc(1'd1) :
                                           {3'd0, 1'd0})))));
  
  /* demux (Ty C5,
       Ty Pointer_CTf') : (writeMerge_choice_CTf',C5) (demuxWriteResult_CTf',Pointer_CTf') > [(writeCTf'lizzieLet29_1_argbuf,Pointer_CTf'),
                                                                                              (writeCTf'lizzieLet40_1_argbuf,Pointer_CTf'),
                                                                                              (writeCTf'lizzieLet49_1_argbuf,Pointer_CTf'),
                                                                                              (writeCTf'lizzieLet50_1_argbuf,Pointer_CTf'),
                                                                                              (writeCTf'lizzieLet51_1_argbuf,Pointer_CTf')] */
  logic [4:0] \demuxWriteResult_CTf'_onehotd ;
  always_comb
    if ((\writeMerge_choice_CTf'_d [0] && \demuxWriteResult_CTf'_d [0]))
      unique case (\writeMerge_choice_CTf'_d [3:1])
        3'd0: \demuxWriteResult_CTf'_onehotd  = 5'd1;
        3'd1: \demuxWriteResult_CTf'_onehotd  = 5'd2;
        3'd2: \demuxWriteResult_CTf'_onehotd  = 5'd4;
        3'd3: \demuxWriteResult_CTf'_onehotd  = 5'd8;
        3'd4: \demuxWriteResult_CTf'_onehotd  = 5'd16;
        default: \demuxWriteResult_CTf'_onehotd  = 5'd0;
      endcase
    else \demuxWriteResult_CTf'_onehotd  = 5'd0;
  assign \writeCTf'lizzieLet29_1_argbuf_d  = {\demuxWriteResult_CTf'_d [16:1],
                                              \demuxWriteResult_CTf'_onehotd [0]};
  assign \writeCTf'lizzieLet40_1_argbuf_d  = {\demuxWriteResult_CTf'_d [16:1],
                                              \demuxWriteResult_CTf'_onehotd [1]};
  assign \writeCTf'lizzieLet49_1_argbuf_d  = {\demuxWriteResult_CTf'_d [16:1],
                                              \demuxWriteResult_CTf'_onehotd [2]};
  assign \writeCTf'lizzieLet50_1_argbuf_d  = {\demuxWriteResult_CTf'_d [16:1],
                                              \demuxWriteResult_CTf'_onehotd [3]};
  assign \writeCTf'lizzieLet51_1_argbuf_d  = {\demuxWriteResult_CTf'_d [16:1],
                                              \demuxWriteResult_CTf'_onehotd [4]};
  assign \demuxWriteResult_CTf'_r  = (| (\demuxWriteResult_CTf'_onehotd  & {\writeCTf'lizzieLet51_1_argbuf_r ,
                                                                            \writeCTf'lizzieLet50_1_argbuf_r ,
                                                                            \writeCTf'lizzieLet49_1_argbuf_r ,
                                                                            \writeCTf'lizzieLet40_1_argbuf_r ,
                                                                            \writeCTf'lizzieLet29_1_argbuf_r }));
  assign \writeMerge_choice_CTf'_r  = \demuxWriteResult_CTf'_r ;
  
  /* dcon (Ty MemIn_CTf',Dcon WriteIn_CTf') : [(forkHP1_CTf2,Word16#),
                                          (writeMerge_data_CTf',CTf')] > (dconWriteIn_CTf',MemIn_CTf') */
  assign \dconWriteIn_CTf'_d  = \WriteIn_CTf'_dc ((& {forkHP1_CTf2_d[0],
                                                      \writeMerge_data_CTf'_d [0]}), forkHP1_CTf2_d, \writeMerge_data_CTf'_d );
  assign {forkHP1_CTf2_r,
          \writeMerge_data_CTf'_r } = {2 {(\dconWriteIn_CTf'_r  && \dconWriteIn_CTf'_d [0])}};
  
  /* dcon (Ty Pointer_CTf',
      Dcon Pointer_CTf') : [(forkHP1_CTf3,Word16#)] > (dconPtr_CTf',Pointer_CTf') */
  assign \dconPtr_CTf'_d  = \Pointer_CTf'_dc ((& {forkHP1_CTf3_d[0]}), forkHP1_CTf3_d);
  assign {forkHP1_CTf3_r} = {1 {(\dconPtr_CTf'_r  && \dconPtr_CTf'_d [0])}};
  
  /* demux (Ty MemOut_CTf',
       Ty Pointer_CTf') : (memWriteOut_CTf',MemOut_CTf') (dconPtr_CTf',Pointer_CTf') > [(_128,Pointer_CTf'),
                                                                                        (demuxWriteResult_CTf',Pointer_CTf')] */
  logic [1:0] \dconPtr_CTf'_onehotd ;
  always_comb
    if ((\memWriteOut_CTf'_d [0] && \dconPtr_CTf'_d [0]))
      unique case (\memWriteOut_CTf'_d [1:1])
        1'd0: \dconPtr_CTf'_onehotd  = 2'd1;
        1'd1: \dconPtr_CTf'_onehotd  = 2'd2;
        default: \dconPtr_CTf'_onehotd  = 2'd0;
      endcase
    else \dconPtr_CTf'_onehotd  = 2'd0;
  assign _128_d = {\dconPtr_CTf'_d [16:1],
                   \dconPtr_CTf'_onehotd [0]};
  assign \demuxWriteResult_CTf'_d  = {\dconPtr_CTf'_d [16:1],
                                      \dconPtr_CTf'_onehotd [1]};
  assign \dconPtr_CTf'_r  = (| (\dconPtr_CTf'_onehotd  & {\demuxWriteResult_CTf'_r ,
                                                          _128_r}));
  assign \memWriteOut_CTf'_r  = \dconPtr_CTf'_r ;
  
  /* const (Ty Word16#,
       Lit 0) : (goFor_6,Go) > (initHP_CTf'''''''''_f'''''''''_Bool,Word16#) */
  assign \initHP_CTf'''''''''_f'''''''''_Bool_d  = {16'd0,
                                                    goFor_6_d[0]};
  assign goFor_6_r = \initHP_CTf'''''''''_f'''''''''_Bool_r ;
  
  /* const (Ty Word16#,
       Lit 1) : (incrHP_CTf'''''''''_f'''''''''_Bool1,Go) > (incrHP_CTf'''''''''_f'''''''''_Bool,Word16#) */
  assign \incrHP_CTf'''''''''_f'''''''''_Bool_d  = {16'd1,
                                                    \incrHP_CTf'''''''''_f'''''''''_Bool1_d [0]};
  assign \incrHP_CTf'''''''''_f'''''''''_Bool1_r  = \incrHP_CTf'''''''''_f'''''''''_Bool_r ;
  
  /* merge (Ty Go) : [(goFor_7,Go),
                 (incrHP_CTf'''''''''_f'''''''''_Bool2,Go)] > (incrHP_mergeCTf'''''''''_f'''''''''_Bool,Go) */
  logic [1:0] \incrHP_mergeCTf'''''''''_f'''''''''_Bool_selected ;
  logic [1:0] \incrHP_mergeCTf'''''''''_f'''''''''_Bool_select ;
  always_comb
    begin
      \incrHP_mergeCTf'''''''''_f'''''''''_Bool_selected  = 2'd0;
      if ((| \incrHP_mergeCTf'''''''''_f'''''''''_Bool_select ))
        \incrHP_mergeCTf'''''''''_f'''''''''_Bool_selected  = \incrHP_mergeCTf'''''''''_f'''''''''_Bool_select ;
      else
        if (goFor_7_d[0])
          \incrHP_mergeCTf'''''''''_f'''''''''_Bool_selected [0] = 1'd1;
        else if (\incrHP_CTf'''''''''_f'''''''''_Bool2_d [0])
          \incrHP_mergeCTf'''''''''_f'''''''''_Bool_selected [1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \incrHP_mergeCTf'''''''''_f'''''''''_Bool_select  <= 2'd0;
    else
      \incrHP_mergeCTf'''''''''_f'''''''''_Bool_select  <= (\incrHP_mergeCTf'''''''''_f'''''''''_Bool_r  ? 2'd0 :
                                                            \incrHP_mergeCTf'''''''''_f'''''''''_Bool_selected );
  always_comb
    if (\incrHP_mergeCTf'''''''''_f'''''''''_Bool_selected [0])
      \incrHP_mergeCTf'''''''''_f'''''''''_Bool_d  = goFor_7_d;
    else if (\incrHP_mergeCTf'''''''''_f'''''''''_Bool_selected [1])
      \incrHP_mergeCTf'''''''''_f'''''''''_Bool_d  = \incrHP_CTf'''''''''_f'''''''''_Bool2_d ;
    else \incrHP_mergeCTf'''''''''_f'''''''''_Bool_d  = 1'd0;
  assign {\incrHP_CTf'''''''''_f'''''''''_Bool2_r ,
          goFor_7_r} = (\incrHP_mergeCTf'''''''''_f'''''''''_Bool_r  ? \incrHP_mergeCTf'''''''''_f'''''''''_Bool_selected  :
                        2'd0);
  
  /* fork (Ty Go) : (incrHP_mergeCTf'''''''''_f'''''''''_Bool_buf,Go) > [(incrHP_CTf'''''''''_f'''''''''_Bool1,Go),
                                                                    (incrHP_CTf'''''''''_f'''''''''_Bool2,Go)] */
  logic [1:0] \incrHP_mergeCTf'''''''''_f'''''''''_Bool_buf_emitted ;
  logic [1:0] \incrHP_mergeCTf'''''''''_f'''''''''_Bool_buf_done ;
  assign \incrHP_CTf'''''''''_f'''''''''_Bool1_d  = (\incrHP_mergeCTf'''''''''_f'''''''''_Bool_buf_d [0] && (! \incrHP_mergeCTf'''''''''_f'''''''''_Bool_buf_emitted [0]));
  assign \incrHP_CTf'''''''''_f'''''''''_Bool2_d  = (\incrHP_mergeCTf'''''''''_f'''''''''_Bool_buf_d [0] && (! \incrHP_mergeCTf'''''''''_f'''''''''_Bool_buf_emitted [1]));
  assign \incrHP_mergeCTf'''''''''_f'''''''''_Bool_buf_done  = (\incrHP_mergeCTf'''''''''_f'''''''''_Bool_buf_emitted  | ({\incrHP_CTf'''''''''_f'''''''''_Bool2_d [0],
                                                                                                                           \incrHP_CTf'''''''''_f'''''''''_Bool1_d [0]} & {\incrHP_CTf'''''''''_f'''''''''_Bool2_r ,
                                                                                                                                                                           \incrHP_CTf'''''''''_f'''''''''_Bool1_r }));
  assign \incrHP_mergeCTf'''''''''_f'''''''''_Bool_buf_r  = (& \incrHP_mergeCTf'''''''''_f'''''''''_Bool_buf_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \incrHP_mergeCTf'''''''''_f'''''''''_Bool_buf_emitted  <= 2'd0;
    else
      \incrHP_mergeCTf'''''''''_f'''''''''_Bool_buf_emitted  <= (\incrHP_mergeCTf'''''''''_f'''''''''_Bool_buf_r  ? 2'd0 :
                                                                 \incrHP_mergeCTf'''''''''_f'''''''''_Bool_buf_done );
  
  /* op_add (Ty Word16#) : (incrHP_CTf'''''''''_f'''''''''_Bool,Word16#) (forkHP1_CTf'''''''''_f'''''''''_Bool,Word16#) > (addHP_CTf'''''''''_f'''''''''_Bool,Word16#) */
  assign \addHP_CTf'''''''''_f'''''''''_Bool_d  = {(\incrHP_CTf'''''''''_f'''''''''_Bool_d [16:1] + \forkHP1_CTf'''''''''_f'''''''''_Bool_d [16:1]),
                                                   (\incrHP_CTf'''''''''_f'''''''''_Bool_d [0] && \forkHP1_CTf'''''''''_f'''''''''_Bool_d [0])};
  assign {\incrHP_CTf'''''''''_f'''''''''_Bool_r ,
          \forkHP1_CTf'''''''''_f'''''''''_Bool_r } = {2 {(\addHP_CTf'''''''''_f'''''''''_Bool_r  && \addHP_CTf'''''''''_f'''''''''_Bool_d [0])}};
  
  /* merge (Ty Word16#) : [(initHP_CTf'''''''''_f'''''''''_Bool,Word16#),
                      (addHP_CTf'''''''''_f'''''''''_Bool,Word16#)] > (mergeHP_CTf'''''''''_f'''''''''_Bool,Word16#) */
  logic [1:0] \mergeHP_CTf'''''''''_f'''''''''_Bool_selected ;
  logic [1:0] \mergeHP_CTf'''''''''_f'''''''''_Bool_select ;
  always_comb
    begin
      \mergeHP_CTf'''''''''_f'''''''''_Bool_selected  = 2'd0;
      if ((| \mergeHP_CTf'''''''''_f'''''''''_Bool_select ))
        \mergeHP_CTf'''''''''_f'''''''''_Bool_selected  = \mergeHP_CTf'''''''''_f'''''''''_Bool_select ;
      else
        if (\initHP_CTf'''''''''_f'''''''''_Bool_d [0])
          \mergeHP_CTf'''''''''_f'''''''''_Bool_selected [0] = 1'd1;
        else if (\addHP_CTf'''''''''_f'''''''''_Bool_d [0])
          \mergeHP_CTf'''''''''_f'''''''''_Bool_selected [1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \mergeHP_CTf'''''''''_f'''''''''_Bool_select  <= 2'd0;
    else
      \mergeHP_CTf'''''''''_f'''''''''_Bool_select  <= (\mergeHP_CTf'''''''''_f'''''''''_Bool_r  ? 2'd0 :
                                                        \mergeHP_CTf'''''''''_f'''''''''_Bool_selected );
  always_comb
    if (\mergeHP_CTf'''''''''_f'''''''''_Bool_selected [0])
      \mergeHP_CTf'''''''''_f'''''''''_Bool_d  = \initHP_CTf'''''''''_f'''''''''_Bool_d ;
    else if (\mergeHP_CTf'''''''''_f'''''''''_Bool_selected [1])
      \mergeHP_CTf'''''''''_f'''''''''_Bool_d  = \addHP_CTf'''''''''_f'''''''''_Bool_d ;
    else \mergeHP_CTf'''''''''_f'''''''''_Bool_d  = {16'd0, 1'd0};
  assign {\addHP_CTf'''''''''_f'''''''''_Bool_r ,
          \initHP_CTf'''''''''_f'''''''''_Bool_r } = (\mergeHP_CTf'''''''''_f'''''''''_Bool_r  ? \mergeHP_CTf'''''''''_f'''''''''_Bool_selected  :
                                                      2'd0);
  
  /* buf (Ty Go) : (incrHP_mergeCTf'''''''''_f'''''''''_Bool,Go) > (incrHP_mergeCTf'''''''''_f'''''''''_Bool_buf,Go) */
  Go_t \incrHP_mergeCTf'''''''''_f'''''''''_Bool_bufchan_d ;
  logic \incrHP_mergeCTf'''''''''_f'''''''''_Bool_bufchan_r ;
  assign \incrHP_mergeCTf'''''''''_f'''''''''_Bool_r  = ((! \incrHP_mergeCTf'''''''''_f'''''''''_Bool_bufchan_d [0]) || \incrHP_mergeCTf'''''''''_f'''''''''_Bool_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \incrHP_mergeCTf'''''''''_f'''''''''_Bool_bufchan_d  <= 1'd0;
    else
      if (\incrHP_mergeCTf'''''''''_f'''''''''_Bool_r )
        \incrHP_mergeCTf'''''''''_f'''''''''_Bool_bufchan_d  <= \incrHP_mergeCTf'''''''''_f'''''''''_Bool_d ;
  Go_t \incrHP_mergeCTf'''''''''_f'''''''''_Bool_bufchan_buf ;
  assign \incrHP_mergeCTf'''''''''_f'''''''''_Bool_bufchan_r  = (! \incrHP_mergeCTf'''''''''_f'''''''''_Bool_bufchan_buf [0]);
  assign \incrHP_mergeCTf'''''''''_f'''''''''_Bool_buf_d  = (\incrHP_mergeCTf'''''''''_f'''''''''_Bool_bufchan_buf [0] ? \incrHP_mergeCTf'''''''''_f'''''''''_Bool_bufchan_buf  :
                                                             \incrHP_mergeCTf'''''''''_f'''''''''_Bool_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \incrHP_mergeCTf'''''''''_f'''''''''_Bool_bufchan_buf  <= 1'd0;
    else
      if ((\incrHP_mergeCTf'''''''''_f'''''''''_Bool_buf_r  && \incrHP_mergeCTf'''''''''_f'''''''''_Bool_bufchan_buf [0]))
        \incrHP_mergeCTf'''''''''_f'''''''''_Bool_bufchan_buf  <= 1'd0;
      else if (((! \incrHP_mergeCTf'''''''''_f'''''''''_Bool_buf_r ) && (! \incrHP_mergeCTf'''''''''_f'''''''''_Bool_bufchan_buf [0])))
        \incrHP_mergeCTf'''''''''_f'''''''''_Bool_bufchan_buf  <= \incrHP_mergeCTf'''''''''_f'''''''''_Bool_bufchan_d ;
  
  /* buf (Ty Word16#) : (mergeHP_CTf'''''''''_f'''''''''_Bool,Word16#) > (mergeHP_CTf'''''''''_f'''''''''_Bool_buf,Word16#) */
  \Word16#_t  \mergeHP_CTf'''''''''_f'''''''''_Bool_bufchan_d ;
  logic \mergeHP_CTf'''''''''_f'''''''''_Bool_bufchan_r ;
  assign \mergeHP_CTf'''''''''_f'''''''''_Bool_r  = ((! \mergeHP_CTf'''''''''_f'''''''''_Bool_bufchan_d [0]) || \mergeHP_CTf'''''''''_f'''''''''_Bool_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \mergeHP_CTf'''''''''_f'''''''''_Bool_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\mergeHP_CTf'''''''''_f'''''''''_Bool_r )
        \mergeHP_CTf'''''''''_f'''''''''_Bool_bufchan_d  <= \mergeHP_CTf'''''''''_f'''''''''_Bool_d ;
  \Word16#_t  \mergeHP_CTf'''''''''_f'''''''''_Bool_bufchan_buf ;
  assign \mergeHP_CTf'''''''''_f'''''''''_Bool_bufchan_r  = (! \mergeHP_CTf'''''''''_f'''''''''_Bool_bufchan_buf [0]);
  assign \mergeHP_CTf'''''''''_f'''''''''_Bool_buf_d  = (\mergeHP_CTf'''''''''_f'''''''''_Bool_bufchan_buf [0] ? \mergeHP_CTf'''''''''_f'''''''''_Bool_bufchan_buf  :
                                                         \mergeHP_CTf'''''''''_f'''''''''_Bool_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \mergeHP_CTf'''''''''_f'''''''''_Bool_bufchan_buf  <= {16'd0,
                                                             1'd0};
    else
      if ((\mergeHP_CTf'''''''''_f'''''''''_Bool_buf_r  && \mergeHP_CTf'''''''''_f'''''''''_Bool_bufchan_buf [0]))
        \mergeHP_CTf'''''''''_f'''''''''_Bool_bufchan_buf  <= {16'd0,
                                                               1'd0};
      else if (((! \mergeHP_CTf'''''''''_f'''''''''_Bool_buf_r ) && (! \mergeHP_CTf'''''''''_f'''''''''_Bool_bufchan_buf [0])))
        \mergeHP_CTf'''''''''_f'''''''''_Bool_bufchan_buf  <= \mergeHP_CTf'''''''''_f'''''''''_Bool_bufchan_d ;
  
  /* fork (Ty Word16#) : (mergeHP_CTf'''''''''_f'''''''''_Bool_buf,Word16#) > [(forkHP1_CTf'''''''''_f'''''''''_Bool,Word16#),
                                                                          (forkHP1_CTf'''''''''_f'''''''''_Boo2,Word16#),
                                                                          (forkHP1_CTf'''''''''_f'''''''''_Boo3,Word16#)] */
  logic [2:0] \mergeHP_CTf'''''''''_f'''''''''_Bool_buf_emitted ;
  logic [2:0] \mergeHP_CTf'''''''''_f'''''''''_Bool_buf_done ;
  assign \forkHP1_CTf'''''''''_f'''''''''_Bool_d  = {\mergeHP_CTf'''''''''_f'''''''''_Bool_buf_d [16:1],
                                                     (\mergeHP_CTf'''''''''_f'''''''''_Bool_buf_d [0] && (! \mergeHP_CTf'''''''''_f'''''''''_Bool_buf_emitted [0]))};
  assign \forkHP1_CTf'''''''''_f'''''''''_Boo2_d  = {\mergeHP_CTf'''''''''_f'''''''''_Bool_buf_d [16:1],
                                                     (\mergeHP_CTf'''''''''_f'''''''''_Bool_buf_d [0] && (! \mergeHP_CTf'''''''''_f'''''''''_Bool_buf_emitted [1]))};
  assign \forkHP1_CTf'''''''''_f'''''''''_Boo3_d  = {\mergeHP_CTf'''''''''_f'''''''''_Bool_buf_d [16:1],
                                                     (\mergeHP_CTf'''''''''_f'''''''''_Bool_buf_d [0] && (! \mergeHP_CTf'''''''''_f'''''''''_Bool_buf_emitted [2]))};
  assign \mergeHP_CTf'''''''''_f'''''''''_Bool_buf_done  = (\mergeHP_CTf'''''''''_f'''''''''_Bool_buf_emitted  | ({\forkHP1_CTf'''''''''_f'''''''''_Boo3_d [0],
                                                                                                                   \forkHP1_CTf'''''''''_f'''''''''_Boo2_d [0],
                                                                                                                   \forkHP1_CTf'''''''''_f'''''''''_Bool_d [0]} & {\forkHP1_CTf'''''''''_f'''''''''_Boo3_r ,
                                                                                                                                                                   \forkHP1_CTf'''''''''_f'''''''''_Boo2_r ,
                                                                                                                                                                   \forkHP1_CTf'''''''''_f'''''''''_Bool_r }));
  assign \mergeHP_CTf'''''''''_f'''''''''_Bool_buf_r  = (& \mergeHP_CTf'''''''''_f'''''''''_Bool_buf_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \mergeHP_CTf'''''''''_f'''''''''_Bool_buf_emitted  <= 3'd0;
    else
      \mergeHP_CTf'''''''''_f'''''''''_Bool_buf_emitted  <= (\mergeHP_CTf'''''''''_f'''''''''_Bool_buf_r  ? 3'd0 :
                                                             \mergeHP_CTf'''''''''_f'''''''''_Bool_buf_done );
  
  /* mergectrl (Ty C2,
           Ty MemIn_CTf'''''''''_f'''''''''_Bool) : [(dconReadIn_CTf'''''''''_f'''''''''_Bool,MemIn_CTf'''''''''_f'''''''''_Bool),
                                                     (dconWriteIn_CTf'''''''''_f'''''''''_Bool,MemIn_CTf'''''''''_f'''''''''_Bool)] > (memMergeChoice_CTf'''''''''_f'''''''''_Bool,C2) (memMergeIn_CTf'''''''''_f'''''''''_Bool,MemIn_CTf'''''''''_f'''''''''_Bool) */
  logic [1:0] \dconReadIn_CTf'''''''''_f'''''''''_Bool_select_d ;
  assign \dconReadIn_CTf'''''''''_f'''''''''_Bool_select_d  = ((| \dconReadIn_CTf'''''''''_f'''''''''_Bool_select_q ) ? \dconReadIn_CTf'''''''''_f'''''''''_Bool_select_q  :
                                                               (\dconReadIn_CTf'''''''''_f'''''''''_Bool_d [0] ? 2'd1 :
                                                                (\dconWriteIn_CTf'''''''''_f'''''''''_Bool_d [0] ? 2'd2 :
                                                                 2'd0)));
  logic [1:0] \dconReadIn_CTf'''''''''_f'''''''''_Bool_select_q ;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \dconReadIn_CTf'''''''''_f'''''''''_Bool_select_q  <= 2'd0;
    else
      \dconReadIn_CTf'''''''''_f'''''''''_Bool_select_q  <= (\dconReadIn_CTf'''''''''_f'''''''''_Bool_done  ? 2'd0 :
                                                             \dconReadIn_CTf'''''''''_f'''''''''_Bool_select_d );
  logic [1:0] \dconReadIn_CTf'''''''''_f'''''''''_Bool_emit_q ;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \dconReadIn_CTf'''''''''_f'''''''''_Bool_emit_q  <= 2'd0;
    else
      \dconReadIn_CTf'''''''''_f'''''''''_Bool_emit_q  <= (\dconReadIn_CTf'''''''''_f'''''''''_Bool_done  ? 2'd0 :
                                                           \dconReadIn_CTf'''''''''_f'''''''''_Bool_emit_d );
  logic [1:0] \dconReadIn_CTf'''''''''_f'''''''''_Bool_emit_d ;
  assign \dconReadIn_CTf'''''''''_f'''''''''_Bool_emit_d  = (\dconReadIn_CTf'''''''''_f'''''''''_Bool_emit_q  | ({\memMergeChoice_CTf'''''''''_f'''''''''_Bool_d [0],
                                                                                                                  \memMergeIn_CTf'''''''''_f'''''''''_Bool_d [0]} & {\memMergeChoice_CTf'''''''''_f'''''''''_Bool_r ,
                                                                                                                                                                     \memMergeIn_CTf'''''''''_f'''''''''_Bool_r }));
  logic \dconReadIn_CTf'''''''''_f'''''''''_Bool_done ;
  assign \dconReadIn_CTf'''''''''_f'''''''''_Bool_done  = (& \dconReadIn_CTf'''''''''_f'''''''''_Bool_emit_d );
  assign {\dconWriteIn_CTf'''''''''_f'''''''''_Bool_r ,
          \dconReadIn_CTf'''''''''_f'''''''''_Bool_r } = (\dconReadIn_CTf'''''''''_f'''''''''_Bool_done  ? \dconReadIn_CTf'''''''''_f'''''''''_Bool_select_d  :
                                                          2'd0);
  assign \memMergeIn_CTf'''''''''_f'''''''''_Bool_d  = ((\dconReadIn_CTf'''''''''_f'''''''''_Bool_select_d [0] && (! \dconReadIn_CTf'''''''''_f'''''''''_Bool_emit_q [0])) ? \dconReadIn_CTf'''''''''_f'''''''''_Bool_d  :
                                                        ((\dconReadIn_CTf'''''''''_f'''''''''_Bool_select_d [1] && (! \dconReadIn_CTf'''''''''_f'''''''''_Bool_emit_q [0])) ? \dconWriteIn_CTf'''''''''_f'''''''''_Bool_d  :
                                                         {132'd0, 1'd0}));
  assign \memMergeChoice_CTf'''''''''_f'''''''''_Bool_d  = ((\dconReadIn_CTf'''''''''_f'''''''''_Bool_select_d [0] && (! \dconReadIn_CTf'''''''''_f'''''''''_Bool_emit_q [1])) ? C1_2_dc(1'd1) :
                                                            ((\dconReadIn_CTf'''''''''_f'''''''''_Bool_select_d [1] && (! \dconReadIn_CTf'''''''''_f'''''''''_Bool_emit_q [1])) ? C2_2_dc(1'd1) :
                                                             {1'd0, 1'd0}));
  
  /* bram (Ty MemIn_CTf'''''''''_f'''''''''_Bool,
      Ty MemOut_CTf'''''''''_f'''''''''_Bool) : (memMergeIn_CTf'''''''''_f'''''''''_Bool_dbuf,MemIn_CTf'''''''''_f'''''''''_Bool) > (memOut_CTf'''''''''_f'''''''''_Bool,MemOut_CTf'''''''''_f'''''''''_Bool) */
  logic [114:0] \memMergeIn_CTf'''''''''_f'''''''''_Bool_dbuf_mem [65535:0];
  logic [15:0] \memMergeIn_CTf'''''''''_f'''''''''_Bool_dbuf_address ;
  logic [114:0] \memMergeIn_CTf'''''''''_f'''''''''_Bool_dbuf_din ;
  logic [114:0] \memOut_CTf'''''''''_f'''''''''_Bool_q ;
  logic \memOut_CTf'''''''''_f'''''''''_Bool_valid ;
  logic \memMergeIn_CTf'''''''''_f'''''''''_Bool_dbuf_we ;
  logic \memOut_CTf'''''''''_f'''''''''_Bool_we ;
  assign \memMergeIn_CTf'''''''''_f'''''''''_Bool_dbuf_din  = \memMergeIn_CTf'''''''''_f'''''''''_Bool_dbuf_d [132:18];
  assign \memMergeIn_CTf'''''''''_f'''''''''_Bool_dbuf_address  = \memMergeIn_CTf'''''''''_f'''''''''_Bool_dbuf_d [17:2];
  assign \memMergeIn_CTf'''''''''_f'''''''''_Bool_dbuf_we  = (\memMergeIn_CTf'''''''''_f'''''''''_Bool_dbuf_d [1:1] && \memMergeIn_CTf'''''''''_f'''''''''_Bool_dbuf_d [0]);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        \memOut_CTf'''''''''_f'''''''''_Bool_we  <= 1'd0;
        \memOut_CTf'''''''''_f'''''''''_Bool_valid  <= 1'd0;
      end
    else
      begin
        \memOut_CTf'''''''''_f'''''''''_Bool_we  <= \memMergeIn_CTf'''''''''_f'''''''''_Bool_dbuf_we ;
        \memOut_CTf'''''''''_f'''''''''_Bool_valid  <= \memMergeIn_CTf'''''''''_f'''''''''_Bool_dbuf_d [0];
        if (\memMergeIn_CTf'''''''''_f'''''''''_Bool_dbuf_we )
          begin
            \memMergeIn_CTf'''''''''_f'''''''''_Bool_dbuf_mem [\memMergeIn_CTf'''''''''_f'''''''''_Bool_dbuf_address ] <= \memMergeIn_CTf'''''''''_f'''''''''_Bool_dbuf_din ;
            \memOut_CTf'''''''''_f'''''''''_Bool_q  <= \memMergeIn_CTf'''''''''_f'''''''''_Bool_dbuf_din ;
          end
        else
          \memOut_CTf'''''''''_f'''''''''_Bool_q  <= \memMergeIn_CTf'''''''''_f'''''''''_Bool_dbuf_mem [\memMergeIn_CTf'''''''''_f'''''''''_Bool_dbuf_address ];
      end
  assign \memOut_CTf'''''''''_f'''''''''_Bool_d  = {\memOut_CTf'''''''''_f'''''''''_Bool_q ,
                                                    \memOut_CTf'''''''''_f'''''''''_Bool_we ,
                                                    \memOut_CTf'''''''''_f'''''''''_Bool_valid };
  assign \memMergeIn_CTf'''''''''_f'''''''''_Bool_dbuf_r  = ((! \memOut_CTf'''''''''_f'''''''''_Bool_valid ) || \memOut_CTf'''''''''_f'''''''''_Bool_r );
  logic [31:0] \profiling_MemIn_CTf'''''''''_f'''''''''_Bool_read ;
  logic [31:0] \profiling_MemIn_CTf'''''''''_f'''''''''_Bool_write ;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        \profiling_MemIn_CTf'''''''''_f'''''''''_Bool_write  <= 0;
        \profiling_MemIn_CTf'''''''''_f'''''''''_Bool_read  <= 0;
      end
    else
      if ((\memMergeIn_CTf'''''''''_f'''''''''_Bool_dbuf_we  == 1'd1))
        \profiling_MemIn_CTf'''''''''_f'''''''''_Bool_write  <= (\profiling_MemIn_CTf'''''''''_f'''''''''_Bool_write  + 1);
      else
        if ((\memOut_CTf'''''''''_f'''''''''_Bool_valid  == 1'd1))
          \profiling_MemIn_CTf'''''''''_f'''''''''_Bool_read  <= (\profiling_MemIn_CTf'''''''''_f'''''''''_Bool_read  + 1);
  
  /* demux (Ty C2,
       Ty MemOut_CTf'''''''''_f'''''''''_Bool) : (memMergeChoice_CTf'''''''''_f'''''''''_Bool,C2) (memOut_CTf'''''''''_f'''''''''_Bool_dbuf,MemOut_CTf'''''''''_f'''''''''_Bool) > [(memReadOut_CTf'''''''''_f'''''''''_Bool,MemOut_CTf'''''''''_f'''''''''_Bool),
                                                                                                                                                                                    (memWriteOut_CTf'''''''''_f'''''''''_Bool,MemOut_CTf'''''''''_f'''''''''_Bool)] */
  logic [1:0] \memOut_CTf'''''''''_f'''''''''_Bool_dbuf_onehotd ;
  always_comb
    if ((\memMergeChoice_CTf'''''''''_f'''''''''_Bool_d [0] && \memOut_CTf'''''''''_f'''''''''_Bool_dbuf_d [0]))
      unique case (\memMergeChoice_CTf'''''''''_f'''''''''_Bool_d [1:1])
        1'd0: \memOut_CTf'''''''''_f'''''''''_Bool_dbuf_onehotd  = 2'd1;
        1'd1: \memOut_CTf'''''''''_f'''''''''_Bool_dbuf_onehotd  = 2'd2;
        default: \memOut_CTf'''''''''_f'''''''''_Bool_dbuf_onehotd  = 2'd0;
      endcase
    else \memOut_CTf'''''''''_f'''''''''_Bool_dbuf_onehotd  = 2'd0;
  assign \memReadOut_CTf'''''''''_f'''''''''_Bool_d  = {\memOut_CTf'''''''''_f'''''''''_Bool_dbuf_d [116:1],
                                                        \memOut_CTf'''''''''_f'''''''''_Bool_dbuf_onehotd [0]};
  assign \memWriteOut_CTf'''''''''_f'''''''''_Bool_d  = {\memOut_CTf'''''''''_f'''''''''_Bool_dbuf_d [116:1],
                                                         \memOut_CTf'''''''''_f'''''''''_Bool_dbuf_onehotd [1]};
  assign \memOut_CTf'''''''''_f'''''''''_Bool_dbuf_r  = (| (\memOut_CTf'''''''''_f'''''''''_Bool_dbuf_onehotd  & {\memWriteOut_CTf'''''''''_f'''''''''_Bool_r ,
                                                                                                                  \memReadOut_CTf'''''''''_f'''''''''_Bool_r }));
  assign \memMergeChoice_CTf'''''''''_f'''''''''_Bool_r  = \memOut_CTf'''''''''_f'''''''''_Bool_dbuf_r ;
  
  /* dbuf (Ty MemIn_CTf'''''''''_f'''''''''_Bool) : (memMergeIn_CTf'''''''''_f'''''''''_Bool_rbuf,MemIn_CTf'''''''''_f'''''''''_Bool) > (memMergeIn_CTf'''''''''_f'''''''''_Bool_dbuf,MemIn_CTf'''''''''_f'''''''''_Bool) */
  assign \memMergeIn_CTf'''''''''_f'''''''''_Bool_rbuf_r  = ((! \memMergeIn_CTf'''''''''_f'''''''''_Bool_dbuf_d [0]) || \memMergeIn_CTf'''''''''_f'''''''''_Bool_dbuf_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \memMergeIn_CTf'''''''''_f'''''''''_Bool_dbuf_d  <= {132'd0, 1'd0};
    else
      if (\memMergeIn_CTf'''''''''_f'''''''''_Bool_rbuf_r )
        \memMergeIn_CTf'''''''''_f'''''''''_Bool_dbuf_d  <= \memMergeIn_CTf'''''''''_f'''''''''_Bool_rbuf_d ;
  
  /* rbuf (Ty MemIn_CTf'''''''''_f'''''''''_Bool) : (memMergeIn_CTf'''''''''_f'''''''''_Bool,MemIn_CTf'''''''''_f'''''''''_Bool) > (memMergeIn_CTf'''''''''_f'''''''''_Bool_rbuf,MemIn_CTf'''''''''_f'''''''''_Bool) */
  \MemIn_CTf'''''''''_f'''''''''_Bool_t  \memMergeIn_CTf'''''''''_f'''''''''_Bool_buf ;
  assign \memMergeIn_CTf'''''''''_f'''''''''_Bool_r  = (! \memMergeIn_CTf'''''''''_f'''''''''_Bool_buf [0]);
  assign \memMergeIn_CTf'''''''''_f'''''''''_Bool_rbuf_d  = (\memMergeIn_CTf'''''''''_f'''''''''_Bool_buf [0] ? \memMergeIn_CTf'''''''''_f'''''''''_Bool_buf  :
                                                             \memMergeIn_CTf'''''''''_f'''''''''_Bool_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \memMergeIn_CTf'''''''''_f'''''''''_Bool_buf  <= {132'd0, 1'd0};
    else
      if ((\memMergeIn_CTf'''''''''_f'''''''''_Bool_rbuf_r  && \memMergeIn_CTf'''''''''_f'''''''''_Bool_buf [0]))
        \memMergeIn_CTf'''''''''_f'''''''''_Bool_buf  <= {132'd0, 1'd0};
      else if (((! \memMergeIn_CTf'''''''''_f'''''''''_Bool_rbuf_r ) && (! \memMergeIn_CTf'''''''''_f'''''''''_Bool_buf [0])))
        \memMergeIn_CTf'''''''''_f'''''''''_Bool_buf  <= \memMergeIn_CTf'''''''''_f'''''''''_Bool_d ;
  
  /* dbuf (Ty MemOut_CTf'''''''''_f'''''''''_Bool) : (memOut_CTf'''''''''_f'''''''''_Bool_rbuf,MemOut_CTf'''''''''_f'''''''''_Bool) > (memOut_CTf'''''''''_f'''''''''_Bool_dbuf,MemOut_CTf'''''''''_f'''''''''_Bool) */
  assign \memOut_CTf'''''''''_f'''''''''_Bool_rbuf_r  = ((! \memOut_CTf'''''''''_f'''''''''_Bool_dbuf_d [0]) || \memOut_CTf'''''''''_f'''''''''_Bool_dbuf_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \memOut_CTf'''''''''_f'''''''''_Bool_dbuf_d  <= {116'd0, 1'd0};
    else
      if (\memOut_CTf'''''''''_f'''''''''_Bool_rbuf_r )
        \memOut_CTf'''''''''_f'''''''''_Bool_dbuf_d  <= \memOut_CTf'''''''''_f'''''''''_Bool_rbuf_d ;
  
  /* rbuf (Ty MemOut_CTf'''''''''_f'''''''''_Bool) : (memOut_CTf'''''''''_f'''''''''_Bool,MemOut_CTf'''''''''_f'''''''''_Bool) > (memOut_CTf'''''''''_f'''''''''_Bool_rbuf,MemOut_CTf'''''''''_f'''''''''_Bool) */
  \MemOut_CTf'''''''''_f'''''''''_Bool_t  \memOut_CTf'''''''''_f'''''''''_Bool_buf ;
  assign \memOut_CTf'''''''''_f'''''''''_Bool_r  = (! \memOut_CTf'''''''''_f'''''''''_Bool_buf [0]);
  assign \memOut_CTf'''''''''_f'''''''''_Bool_rbuf_d  = (\memOut_CTf'''''''''_f'''''''''_Bool_buf [0] ? \memOut_CTf'''''''''_f'''''''''_Bool_buf  :
                                                         \memOut_CTf'''''''''_f'''''''''_Bool_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \memOut_CTf'''''''''_f'''''''''_Bool_buf  <= {116'd0, 1'd0};
    else
      if ((\memOut_CTf'''''''''_f'''''''''_Bool_rbuf_r  && \memOut_CTf'''''''''_f'''''''''_Bool_buf [0]))
        \memOut_CTf'''''''''_f'''''''''_Bool_buf  <= {116'd0, 1'd0};
      else if (((! \memOut_CTf'''''''''_f'''''''''_Bool_rbuf_r ) && (! \memOut_CTf'''''''''_f'''''''''_Bool_buf [0])))
        \memOut_CTf'''''''''_f'''''''''_Bool_buf  <= \memOut_CTf'''''''''_f'''''''''_Bool_d ;
  
  /* destruct (Ty Pointer_CTf'''''''''_f'''''''''_Bool,
          Dcon Pointer_CTf'''''''''_f'''''''''_Bool) : (scfarg_0_2_1_argbuf,Pointer_CTf'''''''''_f'''''''''_Bool) > [(destructReadIn_CTf'''''''''_f'''''''''_Bool,Word16#)] */
  assign \destructReadIn_CTf'''''''''_f'''''''''_Bool_d  = {scfarg_0_2_1_argbuf_d[16:1],
                                                            scfarg_0_2_1_argbuf_d[0]};
  assign scfarg_0_2_1_argbuf_r = \destructReadIn_CTf'''''''''_f'''''''''_Bool_r ;
  
  /* dcon (Ty MemIn_CTf'''''''''_f'''''''''_Bool,
      Dcon ReadIn_CTf'''''''''_f'''''''''_Bool) : [(destructReadIn_CTf'''''''''_f'''''''''_Bool,Word16#)] > (dconReadIn_CTf'''''''''_f'''''''''_Bool,MemIn_CTf'''''''''_f'''''''''_Bool) */
  assign \dconReadIn_CTf'''''''''_f'''''''''_Bool_d  = \ReadIn_CTf'''''''''_f'''''''''_Bool_dc ((& {\destructReadIn_CTf'''''''''_f'''''''''_Bool_d [0]}), \destructReadIn_CTf'''''''''_f'''''''''_Bool_d );
  assign {\destructReadIn_CTf'''''''''_f'''''''''_Bool_r } = {1 {(\dconReadIn_CTf'''''''''_f'''''''''_Bool_r  && \dconReadIn_CTf'''''''''_f'''''''''_Bool_d [0])}};
  
  /* destruct (Ty MemOut_CTf'''''''''_f'''''''''_Bool,
          Dcon ReadOut_CTf'''''''''_f'''''''''_Bool) : (memReadOut_CTf'''''''''_f'''''''''_Bool,MemOut_CTf'''''''''_f'''''''''_Bool) > [(readPointer_CTf'''''''''_f'''''''''_Boolscfarg_0_2_1_argbuf,CTf'''''''''_f'''''''''_Bool)] */
  assign \readPointer_CTf'''''''''_f'''''''''_Boolscfarg_0_2_1_argbuf_d  = {\memReadOut_CTf'''''''''_f'''''''''_Bool_d [116:2],
                                                                            \memReadOut_CTf'''''''''_f'''''''''_Bool_d [0]};
  assign \memReadOut_CTf'''''''''_f'''''''''_Bool_r  = \readPointer_CTf'''''''''_f'''''''''_Boolscfarg_0_2_1_argbuf_r ;
  
  /* mergectrl (Ty C5,
           Ty CTf'''''''''_f'''''''''_Bool) : [(lizzieLet37_1_argbuf,CTf'''''''''_f'''''''''_Bool),
                                               (lizzieLet41_1_argbuf,CTf'''''''''_f'''''''''_Bool),
                                               (lizzieLet54_1_argbuf,CTf'''''''''_f'''''''''_Bool),
                                               (lizzieLet55_1_argbuf,CTf'''''''''_f'''''''''_Bool),
                                               (lizzieLet56_1_argbuf,CTf'''''''''_f'''''''''_Bool)] > (writeMerge_choice_CTf'''''''''_f'''''''''_Bool,C5) (writeMerge_data_CTf'''''''''_f'''''''''_Bool,CTf'''''''''_f'''''''''_Bool) */
  logic [4:0] lizzieLet37_1_argbuf_select_d;
  assign lizzieLet37_1_argbuf_select_d = ((| lizzieLet37_1_argbuf_select_q) ? lizzieLet37_1_argbuf_select_q :
                                          (lizzieLet37_1_argbuf_d[0] ? 5'd1 :
                                           (lizzieLet41_1_argbuf_d[0] ? 5'd2 :
                                            (lizzieLet54_1_argbuf_d[0] ? 5'd4 :
                                             (lizzieLet55_1_argbuf_d[0] ? 5'd8 :
                                              (lizzieLet56_1_argbuf_d[0] ? 5'd16 :
                                               5'd0))))));
  logic [4:0] lizzieLet37_1_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet37_1_argbuf_select_q <= 5'd0;
    else
      lizzieLet37_1_argbuf_select_q <= (lizzieLet37_1_argbuf_done ? 5'd0 :
                                        lizzieLet37_1_argbuf_select_d);
  logic [1:0] lizzieLet37_1_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet37_1_argbuf_emit_q <= 2'd0;
    else
      lizzieLet37_1_argbuf_emit_q <= (lizzieLet37_1_argbuf_done ? 2'd0 :
                                      lizzieLet37_1_argbuf_emit_d);
  logic [1:0] lizzieLet37_1_argbuf_emit_d;
  assign lizzieLet37_1_argbuf_emit_d = (lizzieLet37_1_argbuf_emit_q | ({\writeMerge_choice_CTf'''''''''_f'''''''''_Bool_d [0],
                                                                        \writeMerge_data_CTf'''''''''_f'''''''''_Bool_d [0]} & {\writeMerge_choice_CTf'''''''''_f'''''''''_Bool_r ,
                                                                                                                                \writeMerge_data_CTf'''''''''_f'''''''''_Bool_r }));
  logic lizzieLet37_1_argbuf_done;
  assign lizzieLet37_1_argbuf_done = (& lizzieLet37_1_argbuf_emit_d);
  assign {lizzieLet56_1_argbuf_r,
          lizzieLet55_1_argbuf_r,
          lizzieLet54_1_argbuf_r,
          lizzieLet41_1_argbuf_r,
          lizzieLet37_1_argbuf_r} = (lizzieLet37_1_argbuf_done ? lizzieLet37_1_argbuf_select_d :
                                     5'd0);
  assign \writeMerge_data_CTf'''''''''_f'''''''''_Bool_d  = ((lizzieLet37_1_argbuf_select_d[0] && (! lizzieLet37_1_argbuf_emit_q[0])) ? lizzieLet37_1_argbuf_d :
                                                             ((lizzieLet37_1_argbuf_select_d[1] && (! lizzieLet37_1_argbuf_emit_q[0])) ? lizzieLet41_1_argbuf_d :
                                                              ((lizzieLet37_1_argbuf_select_d[2] && (! lizzieLet37_1_argbuf_emit_q[0])) ? lizzieLet54_1_argbuf_d :
                                                               ((lizzieLet37_1_argbuf_select_d[3] && (! lizzieLet37_1_argbuf_emit_q[0])) ? lizzieLet55_1_argbuf_d :
                                                                ((lizzieLet37_1_argbuf_select_d[4] && (! lizzieLet37_1_argbuf_emit_q[0])) ? lizzieLet56_1_argbuf_d :
                                                                 {115'd0, 1'd0})))));
  assign \writeMerge_choice_CTf'''''''''_f'''''''''_Bool_d  = ((lizzieLet37_1_argbuf_select_d[0] && (! lizzieLet37_1_argbuf_emit_q[1])) ? C1_5_dc(1'd1) :
                                                               ((lizzieLet37_1_argbuf_select_d[1] && (! lizzieLet37_1_argbuf_emit_q[1])) ? C2_5_dc(1'd1) :
                                                                ((lizzieLet37_1_argbuf_select_d[2] && (! lizzieLet37_1_argbuf_emit_q[1])) ? C3_5_dc(1'd1) :
                                                                 ((lizzieLet37_1_argbuf_select_d[3] && (! lizzieLet37_1_argbuf_emit_q[1])) ? C4_5_dc(1'd1) :
                                                                  ((lizzieLet37_1_argbuf_select_d[4] && (! lizzieLet37_1_argbuf_emit_q[1])) ? C5_5_dc(1'd1) :
                                                                   {3'd0, 1'd0})))));
  
  /* demux (Ty C5,
       Ty Pointer_CTf'''''''''_f'''''''''_Bool) : (writeMerge_choice_CTf'''''''''_f'''''''''_Bool,C5) (demuxWriteResult_CTf'''''''''_f'''''''''_Bool,Pointer_CTf'''''''''_f'''''''''_Bool) > [(writeCTf'''''''''_f'''''''''_BoollizzieLet37_1_argbuf,Pointer_CTf'''''''''_f'''''''''_Bool),
                                                                                                                                                                                              (writeCTf'''''''''_f'''''''''_BoollizzieLet41_1_argbuf,Pointer_CTf'''''''''_f'''''''''_Bool),
                                                                                                                                                                                              (writeCTf'''''''''_f'''''''''_BoollizzieLet54_1_argbuf,Pointer_CTf'''''''''_f'''''''''_Bool),
                                                                                                                                                                                              (writeCTf'''''''''_f'''''''''_BoollizzieLet55_1_argbuf,Pointer_CTf'''''''''_f'''''''''_Bool),
                                                                                                                                                                                              (writeCTf'''''''''_f'''''''''_BoollizzieLet56_1_argbuf,Pointer_CTf'''''''''_f'''''''''_Bool)] */
  logic [4:0] \demuxWriteResult_CTf'''''''''_f'''''''''_Bool_onehotd ;
  always_comb
    if ((\writeMerge_choice_CTf'''''''''_f'''''''''_Bool_d [0] && \demuxWriteResult_CTf'''''''''_f'''''''''_Bool_d [0]))
      unique case (\writeMerge_choice_CTf'''''''''_f'''''''''_Bool_d [3:1])
        3'd0:
          \demuxWriteResult_CTf'''''''''_f'''''''''_Bool_onehotd  = 5'd1;
        3'd1:
          \demuxWriteResult_CTf'''''''''_f'''''''''_Bool_onehotd  = 5'd2;
        3'd2:
          \demuxWriteResult_CTf'''''''''_f'''''''''_Bool_onehotd  = 5'd4;
        3'd3:
          \demuxWriteResult_CTf'''''''''_f'''''''''_Bool_onehotd  = 5'd8;
        3'd4:
          \demuxWriteResult_CTf'''''''''_f'''''''''_Bool_onehotd  = 5'd16;
        default:
          \demuxWriteResult_CTf'''''''''_f'''''''''_Bool_onehotd  = 5'd0;
      endcase
    else
      \demuxWriteResult_CTf'''''''''_f'''''''''_Bool_onehotd  = 5'd0;
  assign \writeCTf'''''''''_f'''''''''_BoollizzieLet37_1_argbuf_d  = {\demuxWriteResult_CTf'''''''''_f'''''''''_Bool_d [16:1],
                                                                      \demuxWriteResult_CTf'''''''''_f'''''''''_Bool_onehotd [0]};
  assign \writeCTf'''''''''_f'''''''''_BoollizzieLet41_1_argbuf_d  = {\demuxWriteResult_CTf'''''''''_f'''''''''_Bool_d [16:1],
                                                                      \demuxWriteResult_CTf'''''''''_f'''''''''_Bool_onehotd [1]};
  assign \writeCTf'''''''''_f'''''''''_BoollizzieLet54_1_argbuf_d  = {\demuxWriteResult_CTf'''''''''_f'''''''''_Bool_d [16:1],
                                                                      \demuxWriteResult_CTf'''''''''_f'''''''''_Bool_onehotd [2]};
  assign \writeCTf'''''''''_f'''''''''_BoollizzieLet55_1_argbuf_d  = {\demuxWriteResult_CTf'''''''''_f'''''''''_Bool_d [16:1],
                                                                      \demuxWriteResult_CTf'''''''''_f'''''''''_Bool_onehotd [3]};
  assign \writeCTf'''''''''_f'''''''''_BoollizzieLet56_1_argbuf_d  = {\demuxWriteResult_CTf'''''''''_f'''''''''_Bool_d [16:1],
                                                                      \demuxWriteResult_CTf'''''''''_f'''''''''_Bool_onehotd [4]};
  assign \demuxWriteResult_CTf'''''''''_f'''''''''_Bool_r  = (| (\demuxWriteResult_CTf'''''''''_f'''''''''_Bool_onehotd  & {\writeCTf'''''''''_f'''''''''_BoollizzieLet56_1_argbuf_r ,
                                                                                                                            \writeCTf'''''''''_f'''''''''_BoollizzieLet55_1_argbuf_r ,
                                                                                                                            \writeCTf'''''''''_f'''''''''_BoollizzieLet54_1_argbuf_r ,
                                                                                                                            \writeCTf'''''''''_f'''''''''_BoollizzieLet41_1_argbuf_r ,
                                                                                                                            \writeCTf'''''''''_f'''''''''_BoollizzieLet37_1_argbuf_r }));
  assign \writeMerge_choice_CTf'''''''''_f'''''''''_Bool_r  = \demuxWriteResult_CTf'''''''''_f'''''''''_Bool_r ;
  
  /* dcon (Ty MemIn_CTf'''''''''_f'''''''''_Bool,
      Dcon WriteIn_CTf'''''''''_f'''''''''_Bool) : [(forkHP1_CTf'''''''''_f'''''''''_Boo2,Word16#),
                                                    (writeMerge_data_CTf'''''''''_f'''''''''_Bool,CTf'''''''''_f'''''''''_Bool)] > (dconWriteIn_CTf'''''''''_f'''''''''_Bool,MemIn_CTf'''''''''_f'''''''''_Bool) */
  assign \dconWriteIn_CTf'''''''''_f'''''''''_Bool_d  = \WriteIn_CTf'''''''''_f'''''''''_Bool_dc ((& {\forkHP1_CTf'''''''''_f'''''''''_Boo2_d [0],
                                                                                                      \writeMerge_data_CTf'''''''''_f'''''''''_Bool_d [0]}), \forkHP1_CTf'''''''''_f'''''''''_Boo2_d , \writeMerge_data_CTf'''''''''_f'''''''''_Bool_d );
  assign {\forkHP1_CTf'''''''''_f'''''''''_Boo2_r ,
          \writeMerge_data_CTf'''''''''_f'''''''''_Bool_r } = {2 {(\dconWriteIn_CTf'''''''''_f'''''''''_Bool_r  && \dconWriteIn_CTf'''''''''_f'''''''''_Bool_d [0])}};
  
  /* dcon (Ty Pointer_CTf'''''''''_f'''''''''_Bool,
      Dcon Pointer_CTf'''''''''_f'''''''''_Bool) : [(forkHP1_CTf'''''''''_f'''''''''_Boo3,Word16#)] > (dconPtr_CTf'''''''''_f'''''''''_Bool,Pointer_CTf'''''''''_f'''''''''_Bool) */
  assign \dconPtr_CTf'''''''''_f'''''''''_Bool_d  = \Pointer_CTf'''''''''_f'''''''''_Bool_dc ((& {\forkHP1_CTf'''''''''_f'''''''''_Boo3_d [0]}), \forkHP1_CTf'''''''''_f'''''''''_Boo3_d );
  assign {\forkHP1_CTf'''''''''_f'''''''''_Boo3_r } = {1 {(\dconPtr_CTf'''''''''_f'''''''''_Bool_r  && \dconPtr_CTf'''''''''_f'''''''''_Bool_d [0])}};
  
  /* demux (Ty MemOut_CTf'''''''''_f'''''''''_Bool,
       Ty Pointer_CTf'''''''''_f'''''''''_Bool) : (memWriteOut_CTf'''''''''_f'''''''''_Bool,MemOut_CTf'''''''''_f'''''''''_Bool) (dconPtr_CTf'''''''''_f'''''''''_Bool,Pointer_CTf'''''''''_f'''''''''_Bool) > [(_127,Pointer_CTf'''''''''_f'''''''''_Bool),
                                                                                                                                                                                                                (demuxWriteResult_CTf'''''''''_f'''''''''_Bool,Pointer_CTf'''''''''_f'''''''''_Bool)] */
  logic [1:0] \dconPtr_CTf'''''''''_f'''''''''_Bool_onehotd ;
  always_comb
    if ((\memWriteOut_CTf'''''''''_f'''''''''_Bool_d [0] && \dconPtr_CTf'''''''''_f'''''''''_Bool_d [0]))
      unique case (\memWriteOut_CTf'''''''''_f'''''''''_Bool_d [1:1])
        1'd0: \dconPtr_CTf'''''''''_f'''''''''_Bool_onehotd  = 2'd1;
        1'd1: \dconPtr_CTf'''''''''_f'''''''''_Bool_onehotd  = 2'd2;
        default: \dconPtr_CTf'''''''''_f'''''''''_Bool_onehotd  = 2'd0;
      endcase
    else \dconPtr_CTf'''''''''_f'''''''''_Bool_onehotd  = 2'd0;
  assign _127_d = {\dconPtr_CTf'''''''''_f'''''''''_Bool_d [16:1],
                   \dconPtr_CTf'''''''''_f'''''''''_Bool_onehotd [0]};
  assign \demuxWriteResult_CTf'''''''''_f'''''''''_Bool_d  = {\dconPtr_CTf'''''''''_f'''''''''_Bool_d [16:1],
                                                              \dconPtr_CTf'''''''''_f'''''''''_Bool_onehotd [1]};
  assign \dconPtr_CTf'''''''''_f'''''''''_Bool_r  = (| (\dconPtr_CTf'''''''''_f'''''''''_Bool_onehotd  & {\demuxWriteResult_CTf'''''''''_f'''''''''_Bool_r ,
                                                                                                          _127_r}));
  assign \memWriteOut_CTf'''''''''_f'''''''''_Bool_r  = \dconPtr_CTf'''''''''_f'''''''''_Bool_r ;
  
  /* const (Ty Word16#,
       Lit 0) : (go_1_dummy_write_MaskQTree,Go) > (initHP_MaskQTree,Word16#) */
  assign initHP_MaskQTree_d = {16'd0,
                               go_1_dummy_write_MaskQTree_d[0]};
  assign go_1_dummy_write_MaskQTree_r = initHP_MaskQTree_r;
  
  /* const (Ty Word16#,
       Lit 1) : (incrHP_MaskQTree1,Go) > (incrHP_MaskQTree,Word16#) */
  assign incrHP_MaskQTree_d = {16'd1, incrHP_MaskQTree1_d[0]};
  assign incrHP_MaskQTree1_r = incrHP_MaskQTree_r;
  
  /* merge (Ty Go) : [(go_2_dummy_write_MaskQTree,Go),
                 (incrHP_MaskQTree2,Go)] > (incrHP_mergeMaskQTree,Go) */
  logic [1:0] incrHP_mergeMaskQTree_selected;
  logic [1:0] incrHP_mergeMaskQTree_select;
  always_comb
    begin
      incrHP_mergeMaskQTree_selected = 2'd0;
      if ((| incrHP_mergeMaskQTree_select))
        incrHP_mergeMaskQTree_selected = incrHP_mergeMaskQTree_select;
      else
        if (go_2_dummy_write_MaskQTree_d[0])
          incrHP_mergeMaskQTree_selected[0] = 1'd1;
        else if (incrHP_MaskQTree2_d[0])
          incrHP_mergeMaskQTree_selected[1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeMaskQTree_select <= 2'd0;
    else
      incrHP_mergeMaskQTree_select <= (incrHP_mergeMaskQTree_r ? 2'd0 :
                                       incrHP_mergeMaskQTree_selected);
  always_comb
    if (incrHP_mergeMaskQTree_selected[0])
      incrHP_mergeMaskQTree_d = go_2_dummy_write_MaskQTree_d;
    else if (incrHP_mergeMaskQTree_selected[1])
      incrHP_mergeMaskQTree_d = incrHP_MaskQTree2_d;
    else incrHP_mergeMaskQTree_d = 1'd0;
  assign {incrHP_MaskQTree2_r,
          go_2_dummy_write_MaskQTree_r} = (incrHP_mergeMaskQTree_r ? incrHP_mergeMaskQTree_selected :
                                           2'd0);
  
  /* fork (Ty Go) : (incrHP_mergeMaskQTree_buf,Go) > [(incrHP_MaskQTree1,Go),
                                                 (incrHP_MaskQTree2,Go)] */
  logic [1:0] incrHP_mergeMaskQTree_buf_emitted;
  logic [1:0] incrHP_mergeMaskQTree_buf_done;
  assign incrHP_MaskQTree1_d = (incrHP_mergeMaskQTree_buf_d[0] && (! incrHP_mergeMaskQTree_buf_emitted[0]));
  assign incrHP_MaskQTree2_d = (incrHP_mergeMaskQTree_buf_d[0] && (! incrHP_mergeMaskQTree_buf_emitted[1]));
  assign incrHP_mergeMaskQTree_buf_done = (incrHP_mergeMaskQTree_buf_emitted | ({incrHP_MaskQTree2_d[0],
                                                                                 incrHP_MaskQTree1_d[0]} & {incrHP_MaskQTree2_r,
                                                                                                            incrHP_MaskQTree1_r}));
  assign incrHP_mergeMaskQTree_buf_r = (& incrHP_mergeMaskQTree_buf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeMaskQTree_buf_emitted <= 2'd0;
    else
      incrHP_mergeMaskQTree_buf_emitted <= (incrHP_mergeMaskQTree_buf_r ? 2'd0 :
                                            incrHP_mergeMaskQTree_buf_done);
  
  /* op_add (Ty Word16#) : (incrHP_MaskQTree,Word16#) (forkHP1_MaskQTree,Word16#) > (addHP_MaskQTree,Word16#) */
  assign addHP_MaskQTree_d = {(incrHP_MaskQTree_d[16:1] + forkHP1_MaskQTree_d[16:1]),
                              (incrHP_MaskQTree_d[0] && forkHP1_MaskQTree_d[0])};
  assign {incrHP_MaskQTree_r,
          forkHP1_MaskQTree_r} = {2 {(addHP_MaskQTree_r && addHP_MaskQTree_d[0])}};
  
  /* merge (Ty Word16#) : [(initHP_MaskQTree,Word16#),
                      (addHP_MaskQTree,Word16#)] > (mergeHP_MaskQTree,Word16#) */
  logic [1:0] mergeHP_MaskQTree_selected;
  logic [1:0] mergeHP_MaskQTree_select;
  always_comb
    begin
      mergeHP_MaskQTree_selected = 2'd0;
      if ((| mergeHP_MaskQTree_select))
        mergeHP_MaskQTree_selected = mergeHP_MaskQTree_select;
      else
        if (initHP_MaskQTree_d[0]) mergeHP_MaskQTree_selected[0] = 1'd1;
        else if (addHP_MaskQTree_d[0])
          mergeHP_MaskQTree_selected[1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_MaskQTree_select <= 2'd0;
    else
      mergeHP_MaskQTree_select <= (mergeHP_MaskQTree_r ? 2'd0 :
                                   mergeHP_MaskQTree_selected);
  always_comb
    if (mergeHP_MaskQTree_selected[0])
      mergeHP_MaskQTree_d = initHP_MaskQTree_d;
    else if (mergeHP_MaskQTree_selected[1])
      mergeHP_MaskQTree_d = addHP_MaskQTree_d;
    else mergeHP_MaskQTree_d = {16'd0, 1'd0};
  assign {addHP_MaskQTree_r,
          initHP_MaskQTree_r} = (mergeHP_MaskQTree_r ? mergeHP_MaskQTree_selected :
                                 2'd0);
  
  /* buf (Ty Go) : (incrHP_mergeMaskQTree,Go) > (incrHP_mergeMaskQTree_buf,Go) */
  Go_t incrHP_mergeMaskQTree_bufchan_d;
  logic incrHP_mergeMaskQTree_bufchan_r;
  assign incrHP_mergeMaskQTree_r = ((! incrHP_mergeMaskQTree_bufchan_d[0]) || incrHP_mergeMaskQTree_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeMaskQTree_bufchan_d <= 1'd0;
    else
      if (incrHP_mergeMaskQTree_r)
        incrHP_mergeMaskQTree_bufchan_d <= incrHP_mergeMaskQTree_d;
  Go_t incrHP_mergeMaskQTree_bufchan_buf;
  assign incrHP_mergeMaskQTree_bufchan_r = (! incrHP_mergeMaskQTree_bufchan_buf[0]);
  assign incrHP_mergeMaskQTree_buf_d = (incrHP_mergeMaskQTree_bufchan_buf[0] ? incrHP_mergeMaskQTree_bufchan_buf :
                                        incrHP_mergeMaskQTree_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeMaskQTree_bufchan_buf <= 1'd0;
    else
      if ((incrHP_mergeMaskQTree_buf_r && incrHP_mergeMaskQTree_bufchan_buf[0]))
        incrHP_mergeMaskQTree_bufchan_buf <= 1'd0;
      else if (((! incrHP_mergeMaskQTree_buf_r) && (! incrHP_mergeMaskQTree_bufchan_buf[0])))
        incrHP_mergeMaskQTree_bufchan_buf <= incrHP_mergeMaskQTree_bufchan_d;
  
  /* buf (Ty Word16#) : (mergeHP_MaskQTree,Word16#) > (mergeHP_MaskQTree_buf,Word16#) */
  \Word16#_t  mergeHP_MaskQTree_bufchan_d;
  logic mergeHP_MaskQTree_bufchan_r;
  assign mergeHP_MaskQTree_r = ((! mergeHP_MaskQTree_bufchan_d[0]) || mergeHP_MaskQTree_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_MaskQTree_bufchan_d <= {16'd0, 1'd0};
    else
      if (mergeHP_MaskQTree_r)
        mergeHP_MaskQTree_bufchan_d <= mergeHP_MaskQTree_d;
  \Word16#_t  mergeHP_MaskQTree_bufchan_buf;
  assign mergeHP_MaskQTree_bufchan_r = (! mergeHP_MaskQTree_bufchan_buf[0]);
  assign mergeHP_MaskQTree_buf_d = (mergeHP_MaskQTree_bufchan_buf[0] ? mergeHP_MaskQTree_bufchan_buf :
                                    mergeHP_MaskQTree_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      mergeHP_MaskQTree_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((mergeHP_MaskQTree_buf_r && mergeHP_MaskQTree_bufchan_buf[0]))
        mergeHP_MaskQTree_bufchan_buf <= {16'd0, 1'd0};
      else if (((! mergeHP_MaskQTree_buf_r) && (! mergeHP_MaskQTree_bufchan_buf[0])))
        mergeHP_MaskQTree_bufchan_buf <= mergeHP_MaskQTree_bufchan_d;
  
  /* sink (Ty Word16#) : (forkHP1_MaskQTree_snk,Word16#) > */
  assign {forkHP1_MaskQTree_snk_r,
          forkHP1_MaskQTree_snk_dout} = {forkHP1_MaskQTree_snk_rout,
                                         forkHP1_MaskQTree_snk_d};
  
  /* source (Ty Go) : > (\MaskQTree_src,Go) */
  
  /* fork (Ty Go) : (\MaskQTree_src,Go) > [(go_1_dummy_write_MaskQTree,Go),
                                      (go_2_dummy_write_MaskQTree,Go)] */
  logic [1:0] \\MaskQTree_src_emitted ;
  logic [1:0] \\MaskQTree_src_done ;
  assign go_1_dummy_write_MaskQTree_d = (\\MaskQTree_src_d [0] && (! \\MaskQTree_src_emitted [0]));
  assign go_2_dummy_write_MaskQTree_d = (\\MaskQTree_src_d [0] && (! \\MaskQTree_src_emitted [1]));
  assign \\MaskQTree_src_done  = (\\MaskQTree_src_emitted  | ({go_2_dummy_write_MaskQTree_d[0],
                                                               go_1_dummy_write_MaskQTree_d[0]} & {go_2_dummy_write_MaskQTree_r,
                                                                                                   go_1_dummy_write_MaskQTree_r}));
  assign \\MaskQTree_src_r  = (& \\MaskQTree_src_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \\MaskQTree_src_emitted  <= 2'd0;
    else
      \\MaskQTree_src_emitted  <= (\\MaskQTree_src_r  ? 2'd0 :
                                   \\MaskQTree_src_done );
  
  /* source (Ty MaskQTree) : > (dummy_write_MaskQTree,MaskQTree) */
  
  /* sink (Ty Pointer_MaskQTree) : (dummy_write_MaskQTree_sink,Pointer_MaskQTree) > */
  assign {dummy_write_MaskQTree_sink_r,
          dummy_write_MaskQTree_sink_dout} = {dummy_write_MaskQTree_sink_rout,
                                              dummy_write_MaskQTree_sink_d};
  
  /* fork (Ty Word16#) : (mergeHP_MaskQTree_buf,Word16#) > [(forkHP1_MaskQTree,Word16#),
                                                       (forkHP1_MaskQTree_snk,Word16#),
                                                       (forkHP1_MaskQTre3,Word16#),
                                                       (forkHP1_MaskQTre4,Word16#)] */
  logic [3:0] mergeHP_MaskQTree_buf_emitted;
  logic [3:0] mergeHP_MaskQTree_buf_done;
  assign forkHP1_MaskQTree_d = {mergeHP_MaskQTree_buf_d[16:1],
                                (mergeHP_MaskQTree_buf_d[0] && (! mergeHP_MaskQTree_buf_emitted[0]))};
  assign forkHP1_MaskQTree_snk_d = {mergeHP_MaskQTree_buf_d[16:1],
                                    (mergeHP_MaskQTree_buf_d[0] && (! mergeHP_MaskQTree_buf_emitted[1]))};
  assign forkHP1_MaskQTre3_d = {mergeHP_MaskQTree_buf_d[16:1],
                                (mergeHP_MaskQTree_buf_d[0] && (! mergeHP_MaskQTree_buf_emitted[2]))};
  assign forkHP1_MaskQTre4_d = {mergeHP_MaskQTree_buf_d[16:1],
                                (mergeHP_MaskQTree_buf_d[0] && (! mergeHP_MaskQTree_buf_emitted[3]))};
  assign mergeHP_MaskQTree_buf_done = (mergeHP_MaskQTree_buf_emitted | ({forkHP1_MaskQTre4_d[0],
                                                                         forkHP1_MaskQTre3_d[0],
                                                                         forkHP1_MaskQTree_snk_d[0],
                                                                         forkHP1_MaskQTree_d[0]} & {forkHP1_MaskQTre4_r,
                                                                                                    forkHP1_MaskQTre3_r,
                                                                                                    forkHP1_MaskQTree_snk_r,
                                                                                                    forkHP1_MaskQTree_r}));
  assign mergeHP_MaskQTree_buf_r = (& mergeHP_MaskQTree_buf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_MaskQTree_buf_emitted <= 4'd0;
    else
      mergeHP_MaskQTree_buf_emitted <= (mergeHP_MaskQTree_buf_r ? 4'd0 :
                                        mergeHP_MaskQTree_buf_done);
  
  /* mergectrl (Ty C2,
           Ty MemIn_MaskQTree) : [(dconReadIn_MaskQTree,MemIn_MaskQTree),
                                  (dconWriteIn_MaskQTree,MemIn_MaskQTree)] > (memMergeChoice_MaskQTree,C2) (memMergeIn_MaskQTree,MemIn_MaskQTree) */
  logic [1:0] dconReadIn_MaskQTree_select_d;
  assign dconReadIn_MaskQTree_select_d = ((| dconReadIn_MaskQTree_select_q) ? dconReadIn_MaskQTree_select_q :
                                          (dconReadIn_MaskQTree_d[0] ? 2'd1 :
                                           (dconWriteIn_MaskQTree_d[0] ? 2'd2 :
                                            2'd0)));
  logic [1:0] dconReadIn_MaskQTree_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) dconReadIn_MaskQTree_select_q <= 2'd0;
    else
      dconReadIn_MaskQTree_select_q <= (dconReadIn_MaskQTree_done ? 2'd0 :
                                        dconReadIn_MaskQTree_select_d);
  logic [1:0] dconReadIn_MaskQTree_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) dconReadIn_MaskQTree_emit_q <= 2'd0;
    else
      dconReadIn_MaskQTree_emit_q <= (dconReadIn_MaskQTree_done ? 2'd0 :
                                      dconReadIn_MaskQTree_emit_d);
  logic [1:0] dconReadIn_MaskQTree_emit_d;
  assign dconReadIn_MaskQTree_emit_d = (dconReadIn_MaskQTree_emit_q | ({memMergeChoice_MaskQTree_d[0],
                                                                        memMergeIn_MaskQTree_d[0]} & {memMergeChoice_MaskQTree_r,
                                                                                                      memMergeIn_MaskQTree_r}));
  logic dconReadIn_MaskQTree_done;
  assign dconReadIn_MaskQTree_done = (& dconReadIn_MaskQTree_emit_d);
  assign {dconWriteIn_MaskQTree_r,
          dconReadIn_MaskQTree_r} = (dconReadIn_MaskQTree_done ? dconReadIn_MaskQTree_select_d :
                                     2'd0);
  assign memMergeIn_MaskQTree_d = ((dconReadIn_MaskQTree_select_d[0] && (! dconReadIn_MaskQTree_emit_q[0])) ? dconReadIn_MaskQTree_d :
                                   ((dconReadIn_MaskQTree_select_d[1] && (! dconReadIn_MaskQTree_emit_q[0])) ? dconWriteIn_MaskQTree_d :
                                    {83'd0, 1'd0}));
  assign memMergeChoice_MaskQTree_d = ((dconReadIn_MaskQTree_select_d[0] && (! dconReadIn_MaskQTree_emit_q[1])) ? C1_2_dc(1'd1) :
                                       ((dconReadIn_MaskQTree_select_d[1] && (! dconReadIn_MaskQTree_emit_q[1])) ? C2_2_dc(1'd1) :
                                        {1'd0, 1'd0}));
  
  /* bram (Ty MemIn_MaskQTree,
      Ty MemOut_MaskQTree) : (memMergeIn_MaskQTree_dbuf,MemIn_MaskQTree) > (memOut_MaskQTree,MemOut_MaskQTree) */
  logic [65:0] memMergeIn_MaskQTree_dbuf_mem[65535:0];
  logic [15:0] memMergeIn_MaskQTree_dbuf_address;
  logic [65:0] memMergeIn_MaskQTree_dbuf_din;
  logic [65:0] memOut_MaskQTree_q;
  logic memOut_MaskQTree_valid;
  logic memMergeIn_MaskQTree_dbuf_we;
  logic memOut_MaskQTree_we;
  assign memMergeIn_MaskQTree_dbuf_din = memMergeIn_MaskQTree_dbuf_d[83:18];
  assign memMergeIn_MaskQTree_dbuf_address = memMergeIn_MaskQTree_dbuf_d[17:2];
  assign memMergeIn_MaskQTree_dbuf_we = (memMergeIn_MaskQTree_dbuf_d[1:1] && memMergeIn_MaskQTree_dbuf_d[0]);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        memOut_MaskQTree_we <= 1'd0;
        memOut_MaskQTree_valid <= 1'd0;
      end
    else
      begin
        memOut_MaskQTree_we <= memMergeIn_MaskQTree_dbuf_we;
        memOut_MaskQTree_valid <= memMergeIn_MaskQTree_dbuf_d[0];
        if (memMergeIn_MaskQTree_dbuf_we)
          begin
            memMergeIn_MaskQTree_dbuf_mem[memMergeIn_MaskQTree_dbuf_address] <= memMergeIn_MaskQTree_dbuf_din;
            memOut_MaskQTree_q <= memMergeIn_MaskQTree_dbuf_din;
          end
        else
          memOut_MaskQTree_q <= memMergeIn_MaskQTree_dbuf_mem[memMergeIn_MaskQTree_dbuf_address];
      end
  assign memOut_MaskQTree_d = {memOut_MaskQTree_q,
                               memOut_MaskQTree_we,
                               memOut_MaskQTree_valid};
  assign memMergeIn_MaskQTree_dbuf_r = ((! memOut_MaskQTree_valid) || memOut_MaskQTree_r);
  logic [31:0] profiling_MemIn_MaskQTree_read;
  logic [31:0] profiling_MemIn_MaskQTree_write;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        profiling_MemIn_MaskQTree_write <= 0;
        profiling_MemIn_MaskQTree_read <= 0;
      end
    else
      if ((memMergeIn_MaskQTree_dbuf_we == 1'd1))
        profiling_MemIn_MaskQTree_write <= (profiling_MemIn_MaskQTree_write + 1);
      else
        if ((memOut_MaskQTree_valid == 1'd1))
          profiling_MemIn_MaskQTree_read <= (profiling_MemIn_MaskQTree_read + 1);
  
  /* demux (Ty C2,
       Ty MemOut_MaskQTree) : (memMergeChoice_MaskQTree,C2) (memOut_MaskQTree_dbuf,MemOut_MaskQTree) > [(memReadOut_MaskQTree,MemOut_MaskQTree),
                                                                                                        (memWriteOut_MaskQTree,MemOut_MaskQTree)] */
  logic [1:0] memOut_MaskQTree_dbuf_onehotd;
  always_comb
    if ((memMergeChoice_MaskQTree_d[0] && memOut_MaskQTree_dbuf_d[0]))
      unique case (memMergeChoice_MaskQTree_d[1:1])
        1'd0: memOut_MaskQTree_dbuf_onehotd = 2'd1;
        1'd1: memOut_MaskQTree_dbuf_onehotd = 2'd2;
        default: memOut_MaskQTree_dbuf_onehotd = 2'd0;
      endcase
    else memOut_MaskQTree_dbuf_onehotd = 2'd0;
  assign memReadOut_MaskQTree_d = {memOut_MaskQTree_dbuf_d[67:1],
                                   memOut_MaskQTree_dbuf_onehotd[0]};
  assign memWriteOut_MaskQTree_d = {memOut_MaskQTree_dbuf_d[67:1],
                                    memOut_MaskQTree_dbuf_onehotd[1]};
  assign memOut_MaskQTree_dbuf_r = (| (memOut_MaskQTree_dbuf_onehotd & {memWriteOut_MaskQTree_r,
                                                                        memReadOut_MaskQTree_r}));
  assign memMergeChoice_MaskQTree_r = memOut_MaskQTree_dbuf_r;
  
  /* dbuf (Ty MemIn_MaskQTree) : (memMergeIn_MaskQTree_rbuf,MemIn_MaskQTree) > (memMergeIn_MaskQTree_dbuf,MemIn_MaskQTree) */
  assign memMergeIn_MaskQTree_rbuf_r = ((! memMergeIn_MaskQTree_dbuf_d[0]) || memMergeIn_MaskQTree_dbuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memMergeIn_MaskQTree_dbuf_d <= {83'd0, 1'd0};
    else
      if (memMergeIn_MaskQTree_rbuf_r)
        memMergeIn_MaskQTree_dbuf_d <= memMergeIn_MaskQTree_rbuf_d;
  
  /* rbuf (Ty MemIn_MaskQTree) : (memMergeIn_MaskQTree,MemIn_MaskQTree) > (memMergeIn_MaskQTree_rbuf,MemIn_MaskQTree) */
  MemIn_MaskQTree_t memMergeIn_MaskQTree_buf;
  assign memMergeIn_MaskQTree_r = (! memMergeIn_MaskQTree_buf[0]);
  assign memMergeIn_MaskQTree_rbuf_d = (memMergeIn_MaskQTree_buf[0] ? memMergeIn_MaskQTree_buf :
                                        memMergeIn_MaskQTree_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memMergeIn_MaskQTree_buf <= {83'd0, 1'd0};
    else
      if ((memMergeIn_MaskQTree_rbuf_r && memMergeIn_MaskQTree_buf[0]))
        memMergeIn_MaskQTree_buf <= {83'd0, 1'd0};
      else if (((! memMergeIn_MaskQTree_rbuf_r) && (! memMergeIn_MaskQTree_buf[0])))
        memMergeIn_MaskQTree_buf <= memMergeIn_MaskQTree_d;
  
  /* dbuf (Ty MemOut_MaskQTree) : (memOut_MaskQTree_rbuf,MemOut_MaskQTree) > (memOut_MaskQTree_dbuf,MemOut_MaskQTree) */
  assign memOut_MaskQTree_rbuf_r = ((! memOut_MaskQTree_dbuf_d[0]) || memOut_MaskQTree_dbuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memOut_MaskQTree_dbuf_d <= {67'd0, 1'd0};
    else
      if (memOut_MaskQTree_rbuf_r)
        memOut_MaskQTree_dbuf_d <= memOut_MaskQTree_rbuf_d;
  
  /* rbuf (Ty MemOut_MaskQTree) : (memOut_MaskQTree,MemOut_MaskQTree) > (memOut_MaskQTree_rbuf,MemOut_MaskQTree) */
  MemOut_MaskQTree_t memOut_MaskQTree_buf;
  assign memOut_MaskQTree_r = (! memOut_MaskQTree_buf[0]);
  assign memOut_MaskQTree_rbuf_d = (memOut_MaskQTree_buf[0] ? memOut_MaskQTree_buf :
                                    memOut_MaskQTree_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memOut_MaskQTree_buf <= {67'd0, 1'd0};
    else
      if ((memOut_MaskQTree_rbuf_r && memOut_MaskQTree_buf[0]))
        memOut_MaskQTree_buf <= {67'd0, 1'd0};
      else if (((! memOut_MaskQTree_rbuf_r) && (! memOut_MaskQTree_buf[0])))
        memOut_MaskQTree_buf <= memOut_MaskQTree_d;
  
  /* mergectrl (Ty C2,
           Ty Pointer_MaskQTree) : [(m1a85_1_argbuf,Pointer_MaskQTree),
                                    (q4a8w_1_argbuf,Pointer_MaskQTree)] > (readMerge_choice_MaskQTree,C2) (readMerge_data_MaskQTree,Pointer_MaskQTree) */
  logic [1:0] m1a85_1_argbuf_select_d;
  assign m1a85_1_argbuf_select_d = ((| m1a85_1_argbuf_select_q) ? m1a85_1_argbuf_select_q :
                                    (m1a85_1_argbuf_d[0] ? 2'd1 :
                                     (q4a8w_1_argbuf_d[0] ? 2'd2 :
                                      2'd0)));
  logic [1:0] m1a85_1_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m1a85_1_argbuf_select_q <= 2'd0;
    else
      m1a85_1_argbuf_select_q <= (m1a85_1_argbuf_done ? 2'd0 :
                                  m1a85_1_argbuf_select_d);
  logic [1:0] m1a85_1_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m1a85_1_argbuf_emit_q <= 2'd0;
    else
      m1a85_1_argbuf_emit_q <= (m1a85_1_argbuf_done ? 2'd0 :
                                m1a85_1_argbuf_emit_d);
  logic [1:0] m1a85_1_argbuf_emit_d;
  assign m1a85_1_argbuf_emit_d = (m1a85_1_argbuf_emit_q | ({readMerge_choice_MaskQTree_d[0],
                                                            readMerge_data_MaskQTree_d[0]} & {readMerge_choice_MaskQTree_r,
                                                                                              readMerge_data_MaskQTree_r}));
  logic m1a85_1_argbuf_done;
  assign m1a85_1_argbuf_done = (& m1a85_1_argbuf_emit_d);
  assign {q4a8w_1_argbuf_r,
          m1a85_1_argbuf_r} = (m1a85_1_argbuf_done ? m1a85_1_argbuf_select_d :
                               2'd0);
  assign readMerge_data_MaskQTree_d = ((m1a85_1_argbuf_select_d[0] && (! m1a85_1_argbuf_emit_q[0])) ? m1a85_1_argbuf_d :
                                       ((m1a85_1_argbuf_select_d[1] && (! m1a85_1_argbuf_emit_q[0])) ? q4a8w_1_argbuf_d :
                                        {16'd0, 1'd0}));
  assign readMerge_choice_MaskQTree_d = ((m1a85_1_argbuf_select_d[0] && (! m1a85_1_argbuf_emit_q[1])) ? C1_2_dc(1'd1) :
                                         ((m1a85_1_argbuf_select_d[1] && (! m1a85_1_argbuf_emit_q[1])) ? C2_2_dc(1'd1) :
                                          {1'd0, 1'd0}));
  
  /* demux (Ty C2,
       Ty MaskQTree) : (readMerge_choice_MaskQTree,C2) (destructReadOut_MaskQTree,MaskQTree) > [(readPointer_MaskQTreem1a85_1_argbuf,MaskQTree),
                                                                                                (readPointer_MaskQTreeq4a8w_1_argbuf,MaskQTree)] */
  logic [1:0] destructReadOut_MaskQTree_onehotd;
  always_comb
    if ((readMerge_choice_MaskQTree_d[0] && destructReadOut_MaskQTree_d[0]))
      unique case (readMerge_choice_MaskQTree_d[1:1])
        1'd0: destructReadOut_MaskQTree_onehotd = 2'd1;
        1'd1: destructReadOut_MaskQTree_onehotd = 2'd2;
        default: destructReadOut_MaskQTree_onehotd = 2'd0;
      endcase
    else destructReadOut_MaskQTree_onehotd = 2'd0;
  assign readPointer_MaskQTreem1a85_1_argbuf_d = {destructReadOut_MaskQTree_d[66:1],
                                                  destructReadOut_MaskQTree_onehotd[0]};
  assign readPointer_MaskQTreeq4a8w_1_argbuf_d = {destructReadOut_MaskQTree_d[66:1],
                                                  destructReadOut_MaskQTree_onehotd[1]};
  assign destructReadOut_MaskQTree_r = (| (destructReadOut_MaskQTree_onehotd & {readPointer_MaskQTreeq4a8w_1_argbuf_r,
                                                                                readPointer_MaskQTreem1a85_1_argbuf_r}));
  assign readMerge_choice_MaskQTree_r = destructReadOut_MaskQTree_r;
  
  /* destruct (Ty Pointer_MaskQTree,
          Dcon Pointer_MaskQTree) : (readMerge_data_MaskQTree,Pointer_MaskQTree) > [(destructReadIn_MaskQTree,Word16#)] */
  assign destructReadIn_MaskQTree_d = {readMerge_data_MaskQTree_d[16:1],
                                       readMerge_data_MaskQTree_d[0]};
  assign readMerge_data_MaskQTree_r = destructReadIn_MaskQTree_r;
  
  /* dcon (Ty MemIn_MaskQTree,
      Dcon ReadIn_MaskQTree) : [(destructReadIn_MaskQTree,Word16#)] > (dconReadIn_MaskQTree,MemIn_MaskQTree) */
  assign dconReadIn_MaskQTree_d = ReadIn_MaskQTree_dc((& {destructReadIn_MaskQTree_d[0]}), destructReadIn_MaskQTree_d);
  assign {destructReadIn_MaskQTree_r} = {1 {(dconReadIn_MaskQTree_r && dconReadIn_MaskQTree_d[0])}};
  
  /* destruct (Ty MemOut_MaskQTree,
          Dcon ReadOut_MaskQTree) : (memReadOut_MaskQTree,MemOut_MaskQTree) > [(destructReadOut_MaskQTree,MaskQTree)] */
  assign destructReadOut_MaskQTree_d = {memReadOut_MaskQTree_d[67:2],
                                        memReadOut_MaskQTree_d[0]};
  assign memReadOut_MaskQTree_r = destructReadOut_MaskQTree_r;
  
  /* dcon (Ty MemIn_MaskQTree,
      Dcon WriteIn_MaskQTree) : [(forkHP1_MaskQTre3,Word16#),
                                 (dummy_write_MaskQTree,MaskQTree)] > (dconWriteIn_MaskQTree,MemIn_MaskQTree) */
  assign dconWriteIn_MaskQTree_d = WriteIn_MaskQTree_dc((& {forkHP1_MaskQTre3_d[0],
                                                            dummy_write_MaskQTree_d[0]}), forkHP1_MaskQTre3_d, dummy_write_MaskQTree_d);
  assign {forkHP1_MaskQTre3_r,
          dummy_write_MaskQTree_r} = {2 {(dconWriteIn_MaskQTree_r && dconWriteIn_MaskQTree_d[0])}};
  
  /* dcon (Ty Pointer_MaskQTree,
      Dcon Pointer_MaskQTree) : [(forkHP1_MaskQTre4,Word16#)] > (dconPtr_MaskQTree,Pointer_MaskQTree) */
  assign dconPtr_MaskQTree_d = Pointer_MaskQTree_dc((& {forkHP1_MaskQTre4_d[0]}), forkHP1_MaskQTre4_d);
  assign {forkHP1_MaskQTre4_r} = {1 {(dconPtr_MaskQTree_r && dconPtr_MaskQTree_d[0])}};
  
  /* demux (Ty MemOut_MaskQTree,
       Ty Pointer_MaskQTree) : (memWriteOut_MaskQTree,MemOut_MaskQTree) (dconPtr_MaskQTree,Pointer_MaskQTree) > [(_126,Pointer_MaskQTree),
                                                                                                                 (dummy_write_MaskQTree_sink,Pointer_MaskQTree)] */
  logic [1:0] dconPtr_MaskQTree_onehotd;
  always_comb
    if ((memWriteOut_MaskQTree_d[0] && dconPtr_MaskQTree_d[0]))
      unique case (memWriteOut_MaskQTree_d[1:1])
        1'd0: dconPtr_MaskQTree_onehotd = 2'd1;
        1'd1: dconPtr_MaskQTree_onehotd = 2'd2;
        default: dconPtr_MaskQTree_onehotd = 2'd0;
      endcase
    else dconPtr_MaskQTree_onehotd = 2'd0;
  assign _126_d = {dconPtr_MaskQTree_d[16:1],
                   dconPtr_MaskQTree_onehotd[0]};
  assign dummy_write_MaskQTree_sink_d = {dconPtr_MaskQTree_d[16:1],
                                         dconPtr_MaskQTree_onehotd[1]};
  assign dconPtr_MaskQTree_r = (| (dconPtr_MaskQTree_onehotd & {dummy_write_MaskQTree_sink_r,
                                                                _126_r}));
  assign memWriteOut_MaskQTree_r = dconPtr_MaskQTree_r;
  
  /* buf (Ty Go) : (goFork,Go) > (go_1_argbuf,Go) */
  Go_t goFork_bufchan_d;
  logic goFork_bufchan_r;
  assign goFork_r = ((! goFork_bufchan_d[0]) || goFork_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) goFork_bufchan_d <= 1'd0;
    else if (goFork_r) goFork_bufchan_d <= goFork_d;
  Go_t goFork_bufchan_buf;
  assign goFork_bufchan_r = (! goFork_bufchan_buf[0]);
  assign go_1_argbuf_d = (goFork_bufchan_buf[0] ? goFork_bufchan_buf :
                          goFork_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) goFork_bufchan_buf <= 1'd0;
    else
      if ((go_1_argbuf_r && goFork_bufchan_buf[0]))
        goFork_bufchan_buf <= 1'd0;
      else if (((! go_1_argbuf_r) && (! goFork_bufchan_buf[0])))
        goFork_bufchan_buf <= goFork_bufchan_d;
  
  /* source (Ty Go) : > (sourceGo,Go) */
  
  /* source (Ty Pointer_MaskQTree) : > (m1a82_0,Pointer_MaskQTree) */
  
  /* source (Ty Pointer_QTree_Bool) : > (m2a83_1,Pointer_QTree_Bool) */
  
  /* source (Ty Pointer_QTree_Bool) : > (m3a84_2,Pointer_QTree_Bool) */
  
  /* destruct (Ty TupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_CTf'''''''''_f'''''''''_Bool,
          Dcon TupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_CTf'''''''''_f'''''''''_Bool) : (call_f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_CTf'''''''''_f'''''''''_Bool_1,TupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_CTf'''''''''_f'''''''''_Bool) > [(call_f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_CTf'''''''''_f'''''''''_Boolgo_4,Go),
                                                                                                                                                                                                                                                                                                                          (call_f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_CTf'''''''''_f'''''''''_Boolq4a8w,Pointer_MaskQTree),
                                                                                                                                                                                                                                                                                                                          (call_f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_CTf'''''''''_f'''''''''_Boolq4'a8x,Pointer_QTree_Bool),
                                                                                                                                                                                                                                                                                                                          (call_f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_CTf'''''''''_f'''''''''_Boolsc_0_2,Pointer_CTf'''''''''_f'''''''''_Bool)] */
  logic [3:0] \call_f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_CTf'''''''''_f'''''''''_Bool_1_emitted ;
  logic [3:0] \call_f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_CTf'''''''''_f'''''''''_Bool_1_done ;
  assign \call_f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_CTf'''''''''_f'''''''''_Boolgo_4_d  = (\call_f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_CTf'''''''''_f'''''''''_Bool_1_d [0] && (! \call_f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_CTf'''''''''_f'''''''''_Bool_1_emitted [0]));
  assign \call_f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_CTf'''''''''_f'''''''''_Boolq4a8w_d  = {\call_f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_CTf'''''''''_f'''''''''_Bool_1_d [16:1],
                                                                                                                                          (\call_f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_CTf'''''''''_f'''''''''_Bool_1_d [0] && (! \call_f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_CTf'''''''''_f'''''''''_Bool_1_emitted [1]))};
  assign \call_f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_CTf'''''''''_f'''''''''_Boolq4'a8x_d  = {\call_f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_CTf'''''''''_f'''''''''_Bool_1_d [32:17],
                                                                                                                                           (\call_f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_CTf'''''''''_f'''''''''_Bool_1_d [0] && (! \call_f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_CTf'''''''''_f'''''''''_Bool_1_emitted [2]))};
  assign \call_f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_CTf'''''''''_f'''''''''_Boolsc_0_2_d  = {\call_f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_CTf'''''''''_f'''''''''_Bool_1_d [48:33],
                                                                                                                                           (\call_f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_CTf'''''''''_f'''''''''_Bool_1_d [0] && (! \call_f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_CTf'''''''''_f'''''''''_Bool_1_emitted [3]))};
  assign \call_f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_CTf'''''''''_f'''''''''_Bool_1_done  = (\call_f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_CTf'''''''''_f'''''''''_Bool_1_emitted  | ({\call_f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_CTf'''''''''_f'''''''''_Boolsc_0_2_d [0],
                                                                                                                                                                                                                                                                               \call_f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_CTf'''''''''_f'''''''''_Boolq4'a8x_d [0],
                                                                                                                                                                                                                                                                               \call_f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_CTf'''''''''_f'''''''''_Boolq4a8w_d [0],
                                                                                                                                                                                                                                                                               \call_f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_CTf'''''''''_f'''''''''_Boolgo_4_d [0]} & {\call_f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_CTf'''''''''_f'''''''''_Boolsc_0_2_r ,
                                                                                                                                                                                                                                                                                                                                                                                                                   \call_f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_CTf'''''''''_f'''''''''_Boolq4'a8x_r ,
                                                                                                                                                                                                                                                                                                                                                                                                                   \call_f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_CTf'''''''''_f'''''''''_Boolq4a8w_r ,
                                                                                                                                                                                                                                                                                                                                                                                                                   \call_f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_CTf'''''''''_f'''''''''_Boolgo_4_r }));
  assign \call_f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_CTf'''''''''_f'''''''''_Bool_1_r  = (& \call_f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_CTf'''''''''_f'''''''''_Bool_1_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \call_f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_CTf'''''''''_f'''''''''_Bool_1_emitted  <= 4'd0;
    else
      \call_f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_CTf'''''''''_f'''''''''_Bool_1_emitted  <= (\call_f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_CTf'''''''''_f'''''''''_Bool_1_r  ? 4'd0 :
                                                                                                                                           \call_f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_CTf'''''''''_f'''''''''_Bool_1_done );
  
  /* rbuf (Ty Go) : (call_f'''''''''_f'''''''''_Bool_goConst,Go) > (call_f'''''''''_f'''''''''_Bool_initBufi,Go) */
  Go_t \call_f'''''''''_f'''''''''_Bool_goConst_buf ;
  assign \call_f'''''''''_f'''''''''_Bool_goConst_r  = (! \call_f'''''''''_f'''''''''_Bool_goConst_buf [0]);
  assign \call_f'''''''''_f'''''''''_Bool_initBufi_d  = (\call_f'''''''''_f'''''''''_Bool_goConst_buf [0] ? \call_f'''''''''_f'''''''''_Bool_goConst_buf  :
                                                         \call_f'''''''''_f'''''''''_Bool_goConst_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \call_f'''''''''_f'''''''''_Bool_goConst_buf  <= 1'd0;
    else
      if ((\call_f'''''''''_f'''''''''_Bool_initBufi_r  && \call_f'''''''''_f'''''''''_Bool_goConst_buf [0]))
        \call_f'''''''''_f'''''''''_Bool_goConst_buf  <= 1'd0;
      else if (((! \call_f'''''''''_f'''''''''_Bool_initBufi_r ) && (! \call_f'''''''''_f'''''''''_Bool_goConst_buf [0])))
        \call_f'''''''''_f'''''''''_Bool_goConst_buf  <= \call_f'''''''''_f'''''''''_Bool_goConst_d ;
  
  /* mergectrl (Ty C5,
           Ty Go) : [(call_f'''''''''_f'''''''''_Bool_goMux1,Go),
                     (lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool3_1_argbuf,Go),
                     (lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool2_1_argbuf,Go),
                     (lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool1_1_argbuf,Go),
                     (lizzieLet32_4MQNode_3QNode_Bool_1_argbuf,Go)] > (go_4_goMux_choice,C5) (go_4_goMux_data,Go) */
  logic [4:0] \call_f'''''''''_f'''''''''_Bool_goMux1_select_d ;
  assign \call_f'''''''''_f'''''''''_Bool_goMux1_select_d  = ((| \call_f'''''''''_f'''''''''_Bool_goMux1_select_q ) ? \call_f'''''''''_f'''''''''_Bool_goMux1_select_q  :
                                                              (\call_f'''''''''_f'''''''''_Bool_goMux1_d [0] ? 5'd1 :
                                                               (\lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool3_1_argbuf_d [0] ? 5'd2 :
                                                                (\lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool2_1_argbuf_d [0] ? 5'd4 :
                                                                 (\lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool1_1_argbuf_d [0] ? 5'd8 :
                                                                  (lizzieLet32_4MQNode_3QNode_Bool_1_argbuf_d[0] ? 5'd16 :
                                                                   5'd0))))));
  logic [4:0] \call_f'''''''''_f'''''''''_Bool_goMux1_select_q ;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \call_f'''''''''_f'''''''''_Bool_goMux1_select_q  <= 5'd0;
    else
      \call_f'''''''''_f'''''''''_Bool_goMux1_select_q  <= (\call_f'''''''''_f'''''''''_Bool_goMux1_done  ? 5'd0 :
                                                            \call_f'''''''''_f'''''''''_Bool_goMux1_select_d );
  logic [1:0] \call_f'''''''''_f'''''''''_Bool_goMux1_emit_q ;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \call_f'''''''''_f'''''''''_Bool_goMux1_emit_q  <= 2'd0;
    else
      \call_f'''''''''_f'''''''''_Bool_goMux1_emit_q  <= (\call_f'''''''''_f'''''''''_Bool_goMux1_done  ? 2'd0 :
                                                          \call_f'''''''''_f'''''''''_Bool_goMux1_emit_d );
  logic [1:0] \call_f'''''''''_f'''''''''_Bool_goMux1_emit_d ;
  assign \call_f'''''''''_f'''''''''_Bool_goMux1_emit_d  = (\call_f'''''''''_f'''''''''_Bool_goMux1_emit_q  | ({go_4_goMux_choice_d[0],
                                                                                                                go_4_goMux_data_d[0]} & {go_4_goMux_choice_r,
                                                                                                                                         go_4_goMux_data_r}));
  logic \call_f'''''''''_f'''''''''_Bool_goMux1_done ;
  assign \call_f'''''''''_f'''''''''_Bool_goMux1_done  = (& \call_f'''''''''_f'''''''''_Bool_goMux1_emit_d );
  assign {lizzieLet32_4MQNode_3QNode_Bool_1_argbuf_r,
          \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool1_1_argbuf_r ,
          \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool2_1_argbuf_r ,
          \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool3_1_argbuf_r ,
          \call_f'''''''''_f'''''''''_Bool_goMux1_r } = (\call_f'''''''''_f'''''''''_Bool_goMux1_done  ? \call_f'''''''''_f'''''''''_Bool_goMux1_select_d  :
                                                         5'd0);
  assign go_4_goMux_data_d = ((\call_f'''''''''_f'''''''''_Bool_goMux1_select_d [0] && (! \call_f'''''''''_f'''''''''_Bool_goMux1_emit_q [0])) ? \call_f'''''''''_f'''''''''_Bool_goMux1_d  :
                              ((\call_f'''''''''_f'''''''''_Bool_goMux1_select_d [1] && (! \call_f'''''''''_f'''''''''_Bool_goMux1_emit_q [0])) ? \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool3_1_argbuf_d  :
                               ((\call_f'''''''''_f'''''''''_Bool_goMux1_select_d [2] && (! \call_f'''''''''_f'''''''''_Bool_goMux1_emit_q [0])) ? \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool2_1_argbuf_d  :
                                ((\call_f'''''''''_f'''''''''_Bool_goMux1_select_d [3] && (! \call_f'''''''''_f'''''''''_Bool_goMux1_emit_q [0])) ? \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool1_1_argbuf_d  :
                                 ((\call_f'''''''''_f'''''''''_Bool_goMux1_select_d [4] && (! \call_f'''''''''_f'''''''''_Bool_goMux1_emit_q [0])) ? lizzieLet32_4MQNode_3QNode_Bool_1_argbuf_d :
                                  1'd0)))));
  assign go_4_goMux_choice_d = ((\call_f'''''''''_f'''''''''_Bool_goMux1_select_d [0] && (! \call_f'''''''''_f'''''''''_Bool_goMux1_emit_q [1])) ? C1_5_dc(1'd1) :
                                ((\call_f'''''''''_f'''''''''_Bool_goMux1_select_d [1] && (! \call_f'''''''''_f'''''''''_Bool_goMux1_emit_q [1])) ? C2_5_dc(1'd1) :
                                 ((\call_f'''''''''_f'''''''''_Bool_goMux1_select_d [2] && (! \call_f'''''''''_f'''''''''_Bool_goMux1_emit_q [1])) ? C3_5_dc(1'd1) :
                                  ((\call_f'''''''''_f'''''''''_Bool_goMux1_select_d [3] && (! \call_f'''''''''_f'''''''''_Bool_goMux1_emit_q [1])) ? C4_5_dc(1'd1) :
                                   ((\call_f'''''''''_f'''''''''_Bool_goMux1_select_d [4] && (! \call_f'''''''''_f'''''''''_Bool_goMux1_emit_q [1])) ? C5_5_dc(1'd1) :
                                    {3'd0, 1'd0})))));
  
  /* fork (Ty Go) : (call_f'''''''''_f'''''''''_Bool_initBuf,Go) > [(call_f'''''''''_f'''''''''_Bool_unlockFork1,Go),
                                                               (call_f'''''''''_f'''''''''_Bool_unlockFork2,Go),
                                                               (call_f'''''''''_f'''''''''_Bool_unlockFork3,Go),
                                                               (call_f'''''''''_f'''''''''_Bool_unlockFork4,Go)] */
  logic [3:0] \call_f'''''''''_f'''''''''_Bool_initBuf_emitted ;
  logic [3:0] \call_f'''''''''_f'''''''''_Bool_initBuf_done ;
  assign \call_f'''''''''_f'''''''''_Bool_unlockFork1_d  = (\call_f'''''''''_f'''''''''_Bool_initBuf_d [0] && (! \call_f'''''''''_f'''''''''_Bool_initBuf_emitted [0]));
  assign \call_f'''''''''_f'''''''''_Bool_unlockFork2_d  = (\call_f'''''''''_f'''''''''_Bool_initBuf_d [0] && (! \call_f'''''''''_f'''''''''_Bool_initBuf_emitted [1]));
  assign \call_f'''''''''_f'''''''''_Bool_unlockFork3_d  = (\call_f'''''''''_f'''''''''_Bool_initBuf_d [0] && (! \call_f'''''''''_f'''''''''_Bool_initBuf_emitted [2]));
  assign \call_f'''''''''_f'''''''''_Bool_unlockFork4_d  = (\call_f'''''''''_f'''''''''_Bool_initBuf_d [0] && (! \call_f'''''''''_f'''''''''_Bool_initBuf_emitted [3]));
  assign \call_f'''''''''_f'''''''''_Bool_initBuf_done  = (\call_f'''''''''_f'''''''''_Bool_initBuf_emitted  | ({\call_f'''''''''_f'''''''''_Bool_unlockFork4_d [0],
                                                                                                                 \call_f'''''''''_f'''''''''_Bool_unlockFork3_d [0],
                                                                                                                 \call_f'''''''''_f'''''''''_Bool_unlockFork2_d [0],
                                                                                                                 \call_f'''''''''_f'''''''''_Bool_unlockFork1_d [0]} & {\call_f'''''''''_f'''''''''_Bool_unlockFork4_r ,
                                                                                                                                                                        \call_f'''''''''_f'''''''''_Bool_unlockFork3_r ,
                                                                                                                                                                        \call_f'''''''''_f'''''''''_Bool_unlockFork2_r ,
                                                                                                                                                                        \call_f'''''''''_f'''''''''_Bool_unlockFork1_r }));
  assign \call_f'''''''''_f'''''''''_Bool_initBuf_r  = (& \call_f'''''''''_f'''''''''_Bool_initBuf_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \call_f'''''''''_f'''''''''_Bool_initBuf_emitted  <= 4'd0;
    else
      \call_f'''''''''_f'''''''''_Bool_initBuf_emitted  <= (\call_f'''''''''_f'''''''''_Bool_initBuf_r  ? 4'd0 :
                                                            \call_f'''''''''_f'''''''''_Bool_initBuf_done );
  
  /* initbuf (Ty Go,
         Dcon Go) : (call_f'''''''''_f'''''''''_Bool_initBufi,Go) > (call_f'''''''''_f'''''''''_Bool_initBuf,Go) */
  assign \call_f'''''''''_f'''''''''_Bool_initBufi_r  = ((! \call_f'''''''''_f'''''''''_Bool_initBuf_d [0]) || \call_f'''''''''_f'''''''''_Bool_initBuf_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \call_f'''''''''_f'''''''''_Bool_initBuf_d  <= Go_dc(1'd1);
    else
      if (\call_f'''''''''_f'''''''''_Bool_initBufi_r )
        \call_f'''''''''_f'''''''''_Bool_initBuf_d  <= \call_f'''''''''_f'''''''''_Bool_initBufi_d ;
  
  /* mux (Ty Go,
     Ty Go) : (call_f'''''''''_f'''''''''_Bool_unlockFork1,Go) [(call_f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_CTf'''''''''_f'''''''''_Boolgo_4,Go)] > (call_f'''''''''_f'''''''''_Bool_goMux1,Go) */
  assign \call_f'''''''''_f'''''''''_Bool_goMux1_d  = (\call_f'''''''''_f'''''''''_Bool_unlockFork1_d [0] && \call_f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_CTf'''''''''_f'''''''''_Boolgo_4_d [0]);
  assign \call_f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_CTf'''''''''_f'''''''''_Boolgo_4_r  = (\call_f'''''''''_f'''''''''_Bool_goMux1_r  && (\call_f'''''''''_f'''''''''_Bool_unlockFork1_d [0] && \call_f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_CTf'''''''''_f'''''''''_Boolgo_4_d [0]));
  assign \call_f'''''''''_f'''''''''_Bool_unlockFork1_r  = (\call_f'''''''''_f'''''''''_Bool_goMux1_r  && (\call_f'''''''''_f'''''''''_Bool_unlockFork1_d [0] && \call_f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_CTf'''''''''_f'''''''''_Boolgo_4_d [0]));
  
  /* mux (Ty Go,
     Ty Pointer_MaskQTree) : (call_f'''''''''_f'''''''''_Bool_unlockFork2,Go) [(call_f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_CTf'''''''''_f'''''''''_Boolq4a8w,Pointer_MaskQTree)] > (call_f'''''''''_f'''''''''_Bool_goMux2,Pointer_MaskQTree) */
  assign \call_f'''''''''_f'''''''''_Bool_goMux2_d  = {\call_f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_CTf'''''''''_f'''''''''_Boolq4a8w_d [16:1],
                                                       (\call_f'''''''''_f'''''''''_Bool_unlockFork2_d [0] && \call_f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_CTf'''''''''_f'''''''''_Boolq4a8w_d [0])};
  assign \call_f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_CTf'''''''''_f'''''''''_Boolq4a8w_r  = (\call_f'''''''''_f'''''''''_Bool_goMux2_r  && (\call_f'''''''''_f'''''''''_Bool_unlockFork2_d [0] && \call_f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_CTf'''''''''_f'''''''''_Boolq4a8w_d [0]));
  assign \call_f'''''''''_f'''''''''_Bool_unlockFork2_r  = (\call_f'''''''''_f'''''''''_Bool_goMux2_r  && (\call_f'''''''''_f'''''''''_Bool_unlockFork2_d [0] && \call_f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_CTf'''''''''_f'''''''''_Boolq4a8w_d [0]));
  
  /* mux (Ty Go,
     Ty Pointer_QTree_Bool) : (call_f'''''''''_f'''''''''_Bool_unlockFork3,Go) [(call_f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_CTf'''''''''_f'''''''''_Boolq4'a8x,Pointer_QTree_Bool)] > (call_f'''''''''_f'''''''''_Bool_goMux3,Pointer_QTree_Bool) */
  assign \call_f'''''''''_f'''''''''_Bool_goMux3_d  = {\call_f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_CTf'''''''''_f'''''''''_Boolq4'a8x_d [16:1],
                                                       (\call_f'''''''''_f'''''''''_Bool_unlockFork3_d [0] && \call_f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_CTf'''''''''_f'''''''''_Boolq4'a8x_d [0])};
  assign \call_f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_CTf'''''''''_f'''''''''_Boolq4'a8x_r  = (\call_f'''''''''_f'''''''''_Bool_goMux3_r  && (\call_f'''''''''_f'''''''''_Bool_unlockFork3_d [0] && \call_f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_CTf'''''''''_f'''''''''_Boolq4'a8x_d [0]));
  assign \call_f'''''''''_f'''''''''_Bool_unlockFork3_r  = (\call_f'''''''''_f'''''''''_Bool_goMux3_r  && (\call_f'''''''''_f'''''''''_Bool_unlockFork3_d [0] && \call_f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_CTf'''''''''_f'''''''''_Boolq4'a8x_d [0]));
  
  /* mux (Ty Go,
     Ty Pointer_CTf'''''''''_f'''''''''_Bool) : (call_f'''''''''_f'''''''''_Bool_unlockFork4,Go) [(call_f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_CTf'''''''''_f'''''''''_Boolsc_0_2,Pointer_CTf'''''''''_f'''''''''_Bool)] > (call_f'''''''''_f'''''''''_Bool_goMux4,Pointer_CTf'''''''''_f'''''''''_Bool) */
  assign \call_f'''''''''_f'''''''''_Bool_goMux4_d  = {\call_f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_CTf'''''''''_f'''''''''_Boolsc_0_2_d [16:1],
                                                       (\call_f'''''''''_f'''''''''_Bool_unlockFork4_d [0] && \call_f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_CTf'''''''''_f'''''''''_Boolsc_0_2_d [0])};
  assign \call_f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_CTf'''''''''_f'''''''''_Boolsc_0_2_r  = (\call_f'''''''''_f'''''''''_Bool_goMux4_r  && (\call_f'''''''''_f'''''''''_Bool_unlockFork4_d [0] && \call_f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_CTf'''''''''_f'''''''''_Boolsc_0_2_d [0]));
  assign \call_f'''''''''_f'''''''''_Bool_unlockFork4_r  = (\call_f'''''''''_f'''''''''_Bool_goMux4_r  && (\call_f'''''''''_f'''''''''_Bool_unlockFork4_d [0] && \call_f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_CTf'''''''''_f'''''''''_Boolsc_0_2_d [0]));
  
  /* destruct (Ty TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf',
          Dcon TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf') : (call_f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf'_1,TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf') > [(call_f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf'go_3,Go),
                                                                                                                                                                                                                             (call_f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf'm2a8H,Pointer_QTree_Bool),
                                                                                                                                                                                                                             (call_f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf'm3a8I,Pointer_QTree_Bool),
                                                                                                                                                                                                                             (call_f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf'sc_0_1,Pointer_CTf')] */
  logic [3:0] \call_f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf'_1_emitted ;
  logic [3:0] \call_f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf'_1_done ;
  assign \call_f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf'go_3_d  = (\call_f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf'_1_d [0] && (! \call_f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf'_1_emitted [0]));
  assign \call_f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf'm2a8H_d  = {\call_f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf'_1_d [16:1],
                                                                                           (\call_f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf'_1_d [0] && (! \call_f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf'_1_emitted [1]))};
  assign \call_f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf'm3a8I_d  = {\call_f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf'_1_d [32:17],
                                                                                           (\call_f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf'_1_d [0] && (! \call_f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf'_1_emitted [2]))};
  assign \call_f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf'sc_0_1_d  = {\call_f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf'_1_d [48:33],
                                                                                            (\call_f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf'_1_d [0] && (! \call_f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf'_1_emitted [3]))};
  assign \call_f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf'_1_done  = (\call_f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf'_1_emitted  | ({\call_f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf'sc_0_1_d [0],
                                                                                                                                                                                 \call_f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf'm3a8I_d [0],
                                                                                                                                                                                 \call_f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf'm2a8H_d [0],
                                                                                                                                                                                 \call_f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf'go_3_d [0]} & {\call_f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf'sc_0_1_r ,
                                                                                                                                                                                                                                                                      \call_f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf'm3a8I_r ,
                                                                                                                                                                                                                                                                      \call_f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf'm2a8H_r ,
                                                                                                                                                                                                                                                                      \call_f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf'go_3_r }));
  assign \call_f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf'_1_r  = (& \call_f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf'_1_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \call_f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf'_1_emitted  <= 4'd0;
    else
      \call_f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf'_1_emitted  <= (\call_f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf'_1_r  ? 4'd0 :
                                                                                            \call_f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf'_1_done );
  
  /* rbuf (Ty Go) : (call_f'_goConst,Go) > (call_f'_initBufi,Go) */
  Go_t \call_f'_goConst_buf ;
  assign \call_f'_goConst_r  = (! \call_f'_goConst_buf [0]);
  assign \call_f'_initBufi_d  = (\call_f'_goConst_buf [0] ? \call_f'_goConst_buf  :
                                 \call_f'_goConst_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \call_f'_goConst_buf  <= 1'd0;
    else
      if ((\call_f'_initBufi_r  && \call_f'_goConst_buf [0]))
        \call_f'_goConst_buf  <= 1'd0;
      else if (((! \call_f'_initBufi_r ) && (! \call_f'_goConst_buf [0])))
        \call_f'_goConst_buf  <= \call_f'_goConst_d ;
  
  /* mergectrl (Ty C5,Ty Go) : [(call_f'_goMux1,Go),
                           (lizzieLet48_3Lcall_f'3_1_argbuf,Go),
                           (lizzieLet48_3Lcall_f'2_1_argbuf,Go),
                           (lizzieLet48_3Lcall_f'1_1_argbuf,Go),
                           (lizzieLet20_1_4QNode_Bool_3QNode_Bool_1_argbuf,Go)] > (go_3_goMux_choice,C5) (go_3_goMux_data,Go) */
  logic [4:0] \call_f'_goMux1_select_d ;
  assign \call_f'_goMux1_select_d  = ((| \call_f'_goMux1_select_q ) ? \call_f'_goMux1_select_q  :
                                      (\call_f'_goMux1_d [0] ? 5'd1 :
                                       (\lizzieLet48_3Lcall_f'3_1_argbuf_d [0] ? 5'd2 :
                                        (\lizzieLet48_3Lcall_f'2_1_argbuf_d [0] ? 5'd4 :
                                         (\lizzieLet48_3Lcall_f'1_1_argbuf_d [0] ? 5'd8 :
                                          (lizzieLet20_1_4QNode_Bool_3QNode_Bool_1_argbuf_d[0] ? 5'd16 :
                                           5'd0))))));
  logic [4:0] \call_f'_goMux1_select_q ;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \call_f'_goMux1_select_q  <= 5'd0;
    else
      \call_f'_goMux1_select_q  <= (\call_f'_goMux1_done  ? 5'd0 :
                                    \call_f'_goMux1_select_d );
  logic [1:0] \call_f'_goMux1_emit_q ;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \call_f'_goMux1_emit_q  <= 2'd0;
    else
      \call_f'_goMux1_emit_q  <= (\call_f'_goMux1_done  ? 2'd0 :
                                  \call_f'_goMux1_emit_d );
  logic [1:0] \call_f'_goMux1_emit_d ;
  assign \call_f'_goMux1_emit_d  = (\call_f'_goMux1_emit_q  | ({go_3_goMux_choice_d[0],
                                                                go_3_goMux_data_d[0]} & {go_3_goMux_choice_r,
                                                                                         go_3_goMux_data_r}));
  logic \call_f'_goMux1_done ;
  assign \call_f'_goMux1_done  = (& \call_f'_goMux1_emit_d );
  assign {lizzieLet20_1_4QNode_Bool_3QNode_Bool_1_argbuf_r,
          \lizzieLet48_3Lcall_f'1_1_argbuf_r ,
          \lizzieLet48_3Lcall_f'2_1_argbuf_r ,
          \lizzieLet48_3Lcall_f'3_1_argbuf_r ,
          \call_f'_goMux1_r } = (\call_f'_goMux1_done  ? \call_f'_goMux1_select_d  :
                                 5'd0);
  assign go_3_goMux_data_d = ((\call_f'_goMux1_select_d [0] && (! \call_f'_goMux1_emit_q [0])) ? \call_f'_goMux1_d  :
                              ((\call_f'_goMux1_select_d [1] && (! \call_f'_goMux1_emit_q [0])) ? \lizzieLet48_3Lcall_f'3_1_argbuf_d  :
                               ((\call_f'_goMux1_select_d [2] && (! \call_f'_goMux1_emit_q [0])) ? \lizzieLet48_3Lcall_f'2_1_argbuf_d  :
                                ((\call_f'_goMux1_select_d [3] && (! \call_f'_goMux1_emit_q [0])) ? \lizzieLet48_3Lcall_f'1_1_argbuf_d  :
                                 ((\call_f'_goMux1_select_d [4] && (! \call_f'_goMux1_emit_q [0])) ? lizzieLet20_1_4QNode_Bool_3QNode_Bool_1_argbuf_d :
                                  1'd0)))));
  assign go_3_goMux_choice_d = ((\call_f'_goMux1_select_d [0] && (! \call_f'_goMux1_emit_q [1])) ? C1_5_dc(1'd1) :
                                ((\call_f'_goMux1_select_d [1] && (! \call_f'_goMux1_emit_q [1])) ? C2_5_dc(1'd1) :
                                 ((\call_f'_goMux1_select_d [2] && (! \call_f'_goMux1_emit_q [1])) ? C3_5_dc(1'd1) :
                                  ((\call_f'_goMux1_select_d [3] && (! \call_f'_goMux1_emit_q [1])) ? C4_5_dc(1'd1) :
                                   ((\call_f'_goMux1_select_d [4] && (! \call_f'_goMux1_emit_q [1])) ? C5_5_dc(1'd1) :
                                    {3'd0, 1'd0})))));
  
  /* fork (Ty Go) : (call_f'_initBuf,Go) > [(call_f'_unlockFork1,Go),
                                       (call_f'_unlockFork2,Go),
                                       (call_f'_unlockFork3,Go),
                                       (call_f'_unlockFork4,Go)] */
  logic [3:0] \call_f'_initBuf_emitted ;
  logic [3:0] \call_f'_initBuf_done ;
  assign \call_f'_unlockFork1_d  = (\call_f'_initBuf_d [0] && (! \call_f'_initBuf_emitted [0]));
  assign \call_f'_unlockFork2_d  = (\call_f'_initBuf_d [0] && (! \call_f'_initBuf_emitted [1]));
  assign \call_f'_unlockFork3_d  = (\call_f'_initBuf_d [0] && (! \call_f'_initBuf_emitted [2]));
  assign \call_f'_unlockFork4_d  = (\call_f'_initBuf_d [0] && (! \call_f'_initBuf_emitted [3]));
  assign \call_f'_initBuf_done  = (\call_f'_initBuf_emitted  | ({\call_f'_unlockFork4_d [0],
                                                                 \call_f'_unlockFork3_d [0],
                                                                 \call_f'_unlockFork2_d [0],
                                                                 \call_f'_unlockFork1_d [0]} & {\call_f'_unlockFork4_r ,
                                                                                                \call_f'_unlockFork3_r ,
                                                                                                \call_f'_unlockFork2_r ,
                                                                                                \call_f'_unlockFork1_r }));
  assign \call_f'_initBuf_r  = (& \call_f'_initBuf_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \call_f'_initBuf_emitted  <= 4'd0;
    else
      \call_f'_initBuf_emitted  <= (\call_f'_initBuf_r  ? 4'd0 :
                                    \call_f'_initBuf_done );
  
  /* initbuf (Ty Go,
         Dcon Go) : (call_f'_initBufi,Go) > (call_f'_initBuf,Go) */
  assign \call_f'_initBufi_r  = ((! \call_f'_initBuf_d [0]) || \call_f'_initBuf_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \call_f'_initBuf_d  <= Go_dc(1'd1);
    else
      if (\call_f'_initBufi_r )
        \call_f'_initBuf_d  <= \call_f'_initBufi_d ;
  
  /* mux (Ty Go,
     Ty Go) : (call_f'_unlockFork1,Go) [(call_f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf'go_3,Go)] > (call_f'_goMux1,Go) */
  assign \call_f'_goMux1_d  = (\call_f'_unlockFork1_d [0] && \call_f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf'go_3_d [0]);
  assign \call_f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf'go_3_r  = (\call_f'_goMux1_r  && (\call_f'_unlockFork1_d [0] && \call_f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf'go_3_d [0]));
  assign \call_f'_unlockFork1_r  = (\call_f'_goMux1_r  && (\call_f'_unlockFork1_d [0] && \call_f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf'go_3_d [0]));
  
  /* mux (Ty Go,
     Ty Pointer_QTree_Bool) : (call_f'_unlockFork2,Go) [(call_f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf'm2a8H,Pointer_QTree_Bool)] > (call_f'_goMux2,Pointer_QTree_Bool) */
  assign \call_f'_goMux2_d  = {\call_f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf'm2a8H_d [16:1],
                               (\call_f'_unlockFork2_d [0] && \call_f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf'm2a8H_d [0])};
  assign \call_f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf'm2a8H_r  = (\call_f'_goMux2_r  && (\call_f'_unlockFork2_d [0] && \call_f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf'm2a8H_d [0]));
  assign \call_f'_unlockFork2_r  = (\call_f'_goMux2_r  && (\call_f'_unlockFork2_d [0] && \call_f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf'm2a8H_d [0]));
  
  /* mux (Ty Go,
     Ty Pointer_QTree_Bool) : (call_f'_unlockFork3,Go) [(call_f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf'm3a8I,Pointer_QTree_Bool)] > (call_f'_goMux3,Pointer_QTree_Bool) */
  assign \call_f'_goMux3_d  = {\call_f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf'm3a8I_d [16:1],
                               (\call_f'_unlockFork3_d [0] && \call_f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf'm3a8I_d [0])};
  assign \call_f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf'm3a8I_r  = (\call_f'_goMux3_r  && (\call_f'_unlockFork3_d [0] && \call_f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf'm3a8I_d [0]));
  assign \call_f'_unlockFork3_r  = (\call_f'_goMux3_r  && (\call_f'_unlockFork3_d [0] && \call_f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf'm3a8I_d [0]));
  
  /* mux (Ty Go,
     Ty Pointer_CTf') : (call_f'_unlockFork4,Go) [(call_f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf'sc_0_1,Pointer_CTf')] > (call_f'_goMux4,Pointer_CTf') */
  assign \call_f'_goMux4_d  = {\call_f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf'sc_0_1_d [16:1],
                               (\call_f'_unlockFork4_d [0] && \call_f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf'sc_0_1_d [0])};
  assign \call_f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf'sc_0_1_r  = (\call_f'_goMux4_r  && (\call_f'_unlockFork4_d [0] && \call_f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf'sc_0_1_d [0]));
  assign \call_f'_unlockFork4_r  = (\call_f'_goMux4_r  && (\call_f'_unlockFork4_d [0] && \call_f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf'sc_0_1_d [0]));
  
  /* destruct (Ty TupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf,
          Dcon TupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf) : (call_fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf_1,TupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf) > [(call_fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfgo_2,Go),
                                                                                                                                                                                                                                                                                     (call_fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfm1a85,Pointer_MaskQTree),
                                                                                                                                                                                                                                                                                     (call_fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfm2a86,Pointer_QTree_Bool),
                                                                                                                                                                                                                                                                                     (call_fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfm3a87,Pointer_QTree_Bool),
                                                                                                                                                                                                                                                                                     (call_fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfsc_0,Pointer_CTf)] */
  logic [4:0] call_fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf_1_emitted;
  logic [4:0] call_fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf_1_done;
  assign call_fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfgo_2_d = (call_fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf_1_d[0] && (! call_fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf_1_emitted[0]));
  assign call_fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfm1a85_d = {call_fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf_1_d[16:1],
                                                                                                           (call_fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf_1_d[0] && (! call_fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf_1_emitted[1]))};
  assign call_fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfm2a86_d = {call_fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf_1_d[32:17],
                                                                                                           (call_fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf_1_d[0] && (! call_fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf_1_emitted[2]))};
  assign call_fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfm3a87_d = {call_fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf_1_d[48:33],
                                                                                                           (call_fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf_1_d[0] && (! call_fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf_1_emitted[3]))};
  assign call_fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfsc_0_d = {call_fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf_1_d[64:49],
                                                                                                          (call_fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf_1_d[0] && (! call_fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf_1_emitted[4]))};
  assign call_fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf_1_done = (call_fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf_1_emitted | ({call_fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfsc_0_d[0],
                                                                                                                                                                                                                 call_fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfm3a87_d[0],
                                                                                                                                                                                                                 call_fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfm2a86_d[0],
                                                                                                                                                                                                                 call_fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfm1a85_d[0],
                                                                                                                                                                                                                 call_fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfgo_2_d[0]} & {call_fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfsc_0_r,
                                                                                                                                                                                                                                                                                                                      call_fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfm3a87_r,
                                                                                                                                                                                                                                                                                                                      call_fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfm2a86_r,
                                                                                                                                                                                                                                                                                                                      call_fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfm1a85_r,
                                                                                                                                                                                                                                                                                                                      call_fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfgo_2_r}));
  assign call_fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf_1_r = (& call_fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf_1_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      call_fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf_1_emitted <= 5'd0;
    else
      call_fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf_1_emitted <= (call_fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf_1_r ? 5'd0 :
                                                                                                            call_fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf_1_done);
  
  /* rbuf (Ty Go) : (call_f_goConst,Go) > (call_f_initBufi,Go) */
  Go_t call_f_goConst_buf;
  assign call_f_goConst_r = (! call_f_goConst_buf[0]);
  assign call_f_initBufi_d = (call_f_goConst_buf[0] ? call_f_goConst_buf :
                              call_f_goConst_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_f_goConst_buf <= 1'd0;
    else
      if ((call_f_initBufi_r && call_f_goConst_buf[0]))
        call_f_goConst_buf <= 1'd0;
      else if (((! call_f_initBufi_r) && (! call_f_goConst_buf[0])))
        call_f_goConst_buf <= call_f_goConst_d;
  
  /* mergectrl (Ty C5,Ty Go) : [(call_f_goMux1,Go),
                           (lizzieLet43_3Lcall_f3_1_argbuf,Go),
                           (lizzieLet43_3Lcall_f2_1_argbuf,Go),
                           (lizzieLet43_3Lcall_f1_1_argbuf,Go),
                           (lizzieLet0_4MQNode_4QNode_Bool_3QNode_Bool_1_argbuf,Go)] > (go_2_goMux_choice,C5) (go_2_goMux_data,Go) */
  logic [4:0] call_f_goMux1_select_d;
  assign call_f_goMux1_select_d = ((| call_f_goMux1_select_q) ? call_f_goMux1_select_q :
                                   (call_f_goMux1_d[0] ? 5'd1 :
                                    (lizzieLet43_3Lcall_f3_1_argbuf_d[0] ? 5'd2 :
                                     (lizzieLet43_3Lcall_f2_1_argbuf_d[0] ? 5'd4 :
                                      (lizzieLet43_3Lcall_f1_1_argbuf_d[0] ? 5'd8 :
                                       (lizzieLet0_4MQNode_4QNode_Bool_3QNode_Bool_1_argbuf_d[0] ? 5'd16 :
                                        5'd0))))));
  logic [4:0] call_f_goMux1_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_f_goMux1_select_q <= 5'd0;
    else
      call_f_goMux1_select_q <= (call_f_goMux1_done ? 5'd0 :
                                 call_f_goMux1_select_d);
  logic [1:0] call_f_goMux1_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_f_goMux1_emit_q <= 2'd0;
    else
      call_f_goMux1_emit_q <= (call_f_goMux1_done ? 2'd0 :
                               call_f_goMux1_emit_d);
  logic [1:0] call_f_goMux1_emit_d;
  assign call_f_goMux1_emit_d = (call_f_goMux1_emit_q | ({go_2_goMux_choice_d[0],
                                                          go_2_goMux_data_d[0]} & {go_2_goMux_choice_r,
                                                                                   go_2_goMux_data_r}));
  logic call_f_goMux1_done;
  assign call_f_goMux1_done = (& call_f_goMux1_emit_d);
  assign {lizzieLet0_4MQNode_4QNode_Bool_3QNode_Bool_1_argbuf_r,
          lizzieLet43_3Lcall_f1_1_argbuf_r,
          lizzieLet43_3Lcall_f2_1_argbuf_r,
          lizzieLet43_3Lcall_f3_1_argbuf_r,
          call_f_goMux1_r} = (call_f_goMux1_done ? call_f_goMux1_select_d :
                              5'd0);
  assign go_2_goMux_data_d = ((call_f_goMux1_select_d[0] && (! call_f_goMux1_emit_q[0])) ? call_f_goMux1_d :
                              ((call_f_goMux1_select_d[1] && (! call_f_goMux1_emit_q[0])) ? lizzieLet43_3Lcall_f3_1_argbuf_d :
                               ((call_f_goMux1_select_d[2] && (! call_f_goMux1_emit_q[0])) ? lizzieLet43_3Lcall_f2_1_argbuf_d :
                                ((call_f_goMux1_select_d[3] && (! call_f_goMux1_emit_q[0])) ? lizzieLet43_3Lcall_f1_1_argbuf_d :
                                 ((call_f_goMux1_select_d[4] && (! call_f_goMux1_emit_q[0])) ? lizzieLet0_4MQNode_4QNode_Bool_3QNode_Bool_1_argbuf_d :
                                  1'd0)))));
  assign go_2_goMux_choice_d = ((call_f_goMux1_select_d[0] && (! call_f_goMux1_emit_q[1])) ? C1_5_dc(1'd1) :
                                ((call_f_goMux1_select_d[1] && (! call_f_goMux1_emit_q[1])) ? C2_5_dc(1'd1) :
                                 ((call_f_goMux1_select_d[2] && (! call_f_goMux1_emit_q[1])) ? C3_5_dc(1'd1) :
                                  ((call_f_goMux1_select_d[3] && (! call_f_goMux1_emit_q[1])) ? C4_5_dc(1'd1) :
                                   ((call_f_goMux1_select_d[4] && (! call_f_goMux1_emit_q[1])) ? C5_5_dc(1'd1) :
                                    {3'd0, 1'd0})))));
  
  /* fork (Ty Go) : (call_f_initBuf,Go) > [(call_f_unlockFork1,Go),
                                      (call_f_unlockFork2,Go),
                                      (call_f_unlockFork3,Go),
                                      (call_f_unlockFork4,Go),
                                      (call_f_unlockFork5,Go)] */
  logic [4:0] call_f_initBuf_emitted;
  logic [4:0] call_f_initBuf_done;
  assign call_f_unlockFork1_d = (call_f_initBuf_d[0] && (! call_f_initBuf_emitted[0]));
  assign call_f_unlockFork2_d = (call_f_initBuf_d[0] && (! call_f_initBuf_emitted[1]));
  assign call_f_unlockFork3_d = (call_f_initBuf_d[0] && (! call_f_initBuf_emitted[2]));
  assign call_f_unlockFork4_d = (call_f_initBuf_d[0] && (! call_f_initBuf_emitted[3]));
  assign call_f_unlockFork5_d = (call_f_initBuf_d[0] && (! call_f_initBuf_emitted[4]));
  assign call_f_initBuf_done = (call_f_initBuf_emitted | ({call_f_unlockFork5_d[0],
                                                           call_f_unlockFork4_d[0],
                                                           call_f_unlockFork3_d[0],
                                                           call_f_unlockFork2_d[0],
                                                           call_f_unlockFork1_d[0]} & {call_f_unlockFork5_r,
                                                                                       call_f_unlockFork4_r,
                                                                                       call_f_unlockFork3_r,
                                                                                       call_f_unlockFork2_r,
                                                                                       call_f_unlockFork1_r}));
  assign call_f_initBuf_r = (& call_f_initBuf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_f_initBuf_emitted <= 5'd0;
    else
      call_f_initBuf_emitted <= (call_f_initBuf_r ? 5'd0 :
                                 call_f_initBuf_done);
  
  /* initbuf (Ty Go,
         Dcon Go) : (call_f_initBufi,Go) > (call_f_initBuf,Go) */
  assign call_f_initBufi_r = ((! call_f_initBuf_d[0]) || call_f_initBuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_f_initBuf_d <= Go_dc(1'd1);
    else if (call_f_initBufi_r) call_f_initBuf_d <= call_f_initBufi_d;
  
  /* mux (Ty Go,
     Ty Go) : (call_f_unlockFork1,Go) [(call_fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfgo_2,Go)] > (call_f_goMux1,Go) */
  assign call_f_goMux1_d = (call_f_unlockFork1_d[0] && call_fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfgo_2_d[0]);
  assign call_fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfgo_2_r = (call_f_goMux1_r && (call_f_unlockFork1_d[0] && call_fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfgo_2_d[0]));
  assign call_f_unlockFork1_r = (call_f_goMux1_r && (call_f_unlockFork1_d[0] && call_fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfgo_2_d[0]));
  
  /* mux (Ty Go,
     Ty Pointer_MaskQTree) : (call_f_unlockFork2,Go) [(call_fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfm1a85,Pointer_MaskQTree)] > (call_f_goMux2,Pointer_MaskQTree) */
  assign call_f_goMux2_d = {call_fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfm1a85_d[16:1],
                            (call_f_unlockFork2_d[0] && call_fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfm1a85_d[0])};
  assign call_fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfm1a85_r = (call_f_goMux2_r && (call_f_unlockFork2_d[0] && call_fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfm1a85_d[0]));
  assign call_f_unlockFork2_r = (call_f_goMux2_r && (call_f_unlockFork2_d[0] && call_fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfm1a85_d[0]));
  
  /* mux (Ty Go,
     Ty Pointer_QTree_Bool) : (call_f_unlockFork3,Go) [(call_fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfm2a86,Pointer_QTree_Bool)] > (call_f_goMux3,Pointer_QTree_Bool) */
  assign call_f_goMux3_d = {call_fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfm2a86_d[16:1],
                            (call_f_unlockFork3_d[0] && call_fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfm2a86_d[0])};
  assign call_fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfm2a86_r = (call_f_goMux3_r && (call_f_unlockFork3_d[0] && call_fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfm2a86_d[0]));
  assign call_f_unlockFork3_r = (call_f_goMux3_r && (call_f_unlockFork3_d[0] && call_fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfm2a86_d[0]));
  
  /* mux (Ty Go,
     Ty Pointer_QTree_Bool) : (call_f_unlockFork4,Go) [(call_fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfm3a87,Pointer_QTree_Bool)] > (call_f_goMux4,Pointer_QTree_Bool) */
  assign call_f_goMux4_d = {call_fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfm3a87_d[16:1],
                            (call_f_unlockFork4_d[0] && call_fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfm3a87_d[0])};
  assign call_fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfm3a87_r = (call_f_goMux4_r && (call_f_unlockFork4_d[0] && call_fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfm3a87_d[0]));
  assign call_f_unlockFork4_r = (call_f_goMux4_r && (call_f_unlockFork4_d[0] && call_fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfm3a87_d[0]));
  
  /* mux (Ty Go,
     Ty Pointer_CTf) : (call_f_unlockFork5,Go) [(call_fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfsc_0,Pointer_CTf)] > (call_f_goMux5,Pointer_CTf) */
  assign call_f_goMux5_d = {call_fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfsc_0_d[16:1],
                            (call_f_unlockFork5_d[0] && call_fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfsc_0_d[0])};
  assign call_fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfsc_0_r = (call_f_goMux5_r && (call_f_unlockFork5_d[0] && call_fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfsc_0_d[0]));
  assign call_f_unlockFork5_r = (call_f_goMux5_r && (call_f_unlockFork5_d[0] && call_fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTfsc_0_d[0]));
  
  /* buf (Ty QTree_Bool) : (es_0_1es_1_1es_2_1es_3_1QNode_Bool,QTree_Bool) > (lizzieLet6_1_argbuf,QTree_Bool) */
  QTree_Bool_t es_0_1es_1_1es_2_1es_3_1QNode_Bool_bufchan_d;
  logic es_0_1es_1_1es_2_1es_3_1QNode_Bool_bufchan_r;
  assign es_0_1es_1_1es_2_1es_3_1QNode_Bool_r = ((! es_0_1es_1_1es_2_1es_3_1QNode_Bool_bufchan_d[0]) || es_0_1es_1_1es_2_1es_3_1QNode_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_0_1es_1_1es_2_1es_3_1QNode_Bool_bufchan_d <= {66'd0, 1'd0};
    else
      if (es_0_1es_1_1es_2_1es_3_1QNode_Bool_r)
        es_0_1es_1_1es_2_1es_3_1QNode_Bool_bufchan_d <= es_0_1es_1_1es_2_1es_3_1QNode_Bool_d;
  QTree_Bool_t es_0_1es_1_1es_2_1es_3_1QNode_Bool_bufchan_buf;
  assign es_0_1es_1_1es_2_1es_3_1QNode_Bool_bufchan_r = (! es_0_1es_1_1es_2_1es_3_1QNode_Bool_bufchan_buf[0]);
  assign lizzieLet6_1_argbuf_d = (es_0_1es_1_1es_2_1es_3_1QNode_Bool_bufchan_buf[0] ? es_0_1es_1_1es_2_1es_3_1QNode_Bool_bufchan_buf :
                                  es_0_1es_1_1es_2_1es_3_1QNode_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_0_1es_1_1es_2_1es_3_1QNode_Bool_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((lizzieLet6_1_argbuf_r && es_0_1es_1_1es_2_1es_3_1QNode_Bool_bufchan_buf[0]))
        es_0_1es_1_1es_2_1es_3_1QNode_Bool_bufchan_buf <= {66'd0, 1'd0};
      else if (((! lizzieLet6_1_argbuf_r) && (! es_0_1es_1_1es_2_1es_3_1QNode_Bool_bufchan_buf[0])))
        es_0_1es_1_1es_2_1es_3_1QNode_Bool_bufchan_buf <= es_0_1es_1_1es_2_1es_3_1QNode_Bool_bufchan_d;
  
  /* buf (Ty QTree_Bool) : (es_4_1es_5_1es_6_1es_7_1QNode_Bool,QTree_Bool) > (lizzieLet15_1_1_argbuf,QTree_Bool) */
  QTree_Bool_t es_4_1es_5_1es_6_1es_7_1QNode_Bool_bufchan_d;
  logic es_4_1es_5_1es_6_1es_7_1QNode_Bool_bufchan_r;
  assign es_4_1es_5_1es_6_1es_7_1QNode_Bool_r = ((! es_4_1es_5_1es_6_1es_7_1QNode_Bool_bufchan_d[0]) || es_4_1es_5_1es_6_1es_7_1QNode_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_4_1es_5_1es_6_1es_7_1QNode_Bool_bufchan_d <= {66'd0, 1'd0};
    else
      if (es_4_1es_5_1es_6_1es_7_1QNode_Bool_r)
        es_4_1es_5_1es_6_1es_7_1QNode_Bool_bufchan_d <= es_4_1es_5_1es_6_1es_7_1QNode_Bool_d;
  QTree_Bool_t es_4_1es_5_1es_6_1es_7_1QNode_Bool_bufchan_buf;
  assign es_4_1es_5_1es_6_1es_7_1QNode_Bool_bufchan_r = (! es_4_1es_5_1es_6_1es_7_1QNode_Bool_bufchan_buf[0]);
  assign lizzieLet15_1_1_argbuf_d = (es_4_1es_5_1es_6_1es_7_1QNode_Bool_bufchan_buf[0] ? es_4_1es_5_1es_6_1es_7_1QNode_Bool_bufchan_buf :
                                     es_4_1es_5_1es_6_1es_7_1QNode_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_4_1es_5_1es_6_1es_7_1QNode_Bool_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((lizzieLet15_1_1_argbuf_r && es_4_1es_5_1es_6_1es_7_1QNode_Bool_bufchan_buf[0]))
        es_4_1es_5_1es_6_1es_7_1QNode_Bool_bufchan_buf <= {66'd0, 1'd0};
      else if (((! lizzieLet15_1_1_argbuf_r) && (! es_4_1es_5_1es_6_1es_7_1QNode_Bool_bufchan_buf[0])))
        es_4_1es_5_1es_6_1es_7_1QNode_Bool_bufchan_buf <= es_4_1es_5_1es_6_1es_7_1QNode_Bool_bufchan_d;
  
  /* mergectrl (Ty C8,
           Ty TupGo___Pointer_MaskQTree___Pointer_QTree_Bool) : [(f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool_1,TupGo___Pointer_MaskQTree___Pointer_QTree_Bool),
                                                                 (f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool2,TupGo___Pointer_MaskQTree___Pointer_QTree_Bool),
                                                                 (f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool3,TupGo___Pointer_MaskQTree___Pointer_QTree_Bool),
                                                                 (f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool4,TupGo___Pointer_MaskQTree___Pointer_QTree_Bool),
                                                                 (f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool5,TupGo___Pointer_MaskQTree___Pointer_QTree_Bool),
                                                                 (f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool6,TupGo___Pointer_MaskQTree___Pointer_QTree_Bool),
                                                                 (f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool7,TupGo___Pointer_MaskQTree___Pointer_QTree_Bool),
                                                                 (f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool8,TupGo___Pointer_MaskQTree___Pointer_QTree_Bool)] > (f'''''''''_f'''''''''_Bool_choice,C8) (f'''''''''_f'''''''''_Bool_data,TupGo___Pointer_MaskQTree___Pointer_QTree_Bool) */
  logic [7:0] \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool_1_select_d ;
  assign \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool_1_select_d  = ((| \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool_1_select_q ) ? \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool_1_select_q  :
                                                                                                  (\f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool_1_d [0] ? 8'd1 :
                                                                                                   (\f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool2_d [0] ? 8'd2 :
                                                                                                    (\f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool3_d [0] ? 8'd4 :
                                                                                                     (\f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool4_d [0] ? 8'd8 :
                                                                                                      (\f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool5_d [0] ? 8'd16 :
                                                                                                       (\f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool6_d [0] ? 8'd32 :
                                                                                                        (\f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool7_d [0] ? 8'd64 :
                                                                                                         (\f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool8_d [0] ? 8'd128 :
                                                                                                          8'd0)))))))));
  logic [7:0] \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool_1_select_q ;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool_1_select_q  <= 8'd0;
    else
      \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool_1_select_q  <= (\f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool_1_done  ? 8'd0 :
                                                                                                \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool_1_select_d );
  logic [1:0] \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool_1_emit_q ;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool_1_emit_q  <= 2'd0;
    else
      \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool_1_emit_q  <= (\f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool_1_done  ? 2'd0 :
                                                                                              \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool_1_emit_d );
  logic [1:0] \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool_1_emit_d ;
  assign \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool_1_emit_d  = (\f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool_1_emit_q  | ({\f'''''''''_f'''''''''_Bool_choice_d [0],
                                                                                                                                                                                        \f'''''''''_f'''''''''_Bool_data_d [0]} & {\f'''''''''_f'''''''''_Bool_choice_r ,
                                                                                                                                                                                                                                   \f'''''''''_f'''''''''_Bool_data_r }));
  logic \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool_1_done ;
  assign \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool_1_done  = (& \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool_1_emit_d );
  assign {\f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool8_r ,
          \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool7_r ,
          \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool6_r ,
          \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool5_r ,
          \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool4_r ,
          \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool3_r ,
          \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool2_r ,
          \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool_1_r } = (\f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool_1_done  ? \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool_1_select_d  :
                                                                                             8'd0);
  assign \f'''''''''_f'''''''''_Bool_data_d  = ((\f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool_1_select_d [0] && (! \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool_1_emit_q [0])) ? \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool_1_d  :
                                                ((\f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool_1_select_d [1] && (! \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool_1_emit_q [0])) ? \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool2_d  :
                                                 ((\f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool_1_select_d [2] && (! \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool_1_emit_q [0])) ? \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool3_d  :
                                                  ((\f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool_1_select_d [3] && (! \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool_1_emit_q [0])) ? \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool4_d  :
                                                   ((\f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool_1_select_d [4] && (! \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool_1_emit_q [0])) ? \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool5_d  :
                                                    ((\f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool_1_select_d [5] && (! \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool_1_emit_q [0])) ? \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool6_d  :
                                                     ((\f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool_1_select_d [6] && (! \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool_1_emit_q [0])) ? \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool7_d  :
                                                      ((\f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool_1_select_d [7] && (! \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool_1_emit_q [0])) ? \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool8_d  :
                                                       {32'd0, 1'd0}))))))));
  assign \f'''''''''_f'''''''''_Bool_choice_d  = ((\f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool_1_select_d [0] && (! \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool_1_emit_q [1])) ? C1_8_dc(1'd1) :
                                                  ((\f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool_1_select_d [1] && (! \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool_1_emit_q [1])) ? C2_8_dc(1'd1) :
                                                   ((\f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool_1_select_d [2] && (! \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool_1_emit_q [1])) ? C3_8_dc(1'd1) :
                                                    ((\f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool_1_select_d [3] && (! \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool_1_emit_q [1])) ? C4_8_dc(1'd1) :
                                                     ((\f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool_1_select_d [4] && (! \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool_1_emit_q [1])) ? C5_8_dc(1'd1) :
                                                      ((\f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool_1_select_d [5] && (! \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool_1_emit_q [1])) ? C6_8_dc(1'd1) :
                                                       ((\f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool_1_select_d [6] && (! \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool_1_emit_q [1])) ? C7_8_dc(1'd1) :
                                                        ((\f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool_1_select_d [7] && (! \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool_1_emit_q [1])) ? C8_8_dc(1'd1) :
                                                         {3'd0, 1'd0}))))))));
  
  /* fork (Ty Go) : (f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Boolgo_7,Go) > [(go_7_1,Go),
                                                                                                    (go_7_2,Go)] */
  logic [1:0] \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Boolgo_7_emitted ;
  logic [1:0] \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Boolgo_7_done ;
  assign go_7_1_d = (\f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Boolgo_7_d [0] && (! \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Boolgo_7_emitted [0]));
  assign go_7_2_d = (\f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Boolgo_7_d [0] && (! \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Boolgo_7_emitted [1]));
  assign \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Boolgo_7_done  = (\f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Boolgo_7_emitted  | ({go_7_2_d[0],
                                                                                                                                                                                           go_7_1_d[0]} & {go_7_2_r,
                                                                                                                                                                                                           go_7_1_r}));
  assign \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Boolgo_7_r  = (& \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Boolgo_7_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Boolgo_7_emitted  <= 2'd0;
    else
      \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Boolgo_7_emitted  <= (\f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Boolgo_7_r  ? 2'd0 :
                                                                                                 \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Boolgo_7_done );
  
  /* buf (Ty Pointer_QTree_Bool) : (f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Boolq4'a8x_1,Pointer_QTree_Bool) > (q4'a8x_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Boolq4'a8x_1_bufchan_d ;
  logic \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Boolq4'a8x_1_bufchan_r ;
  assign \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Boolq4'a8x_1_r  = ((! \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Boolq4'a8x_1_bufchan_d [0]) || \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Boolq4'a8x_1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Boolq4'a8x_1_bufchan_d  <= {16'd0,
                                                                                                       1'd0};
    else
      if (\f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Boolq4'a8x_1_r )
        \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Boolq4'a8x_1_bufchan_d  <= \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Boolq4'a8x_1_d ;
  Pointer_QTree_Bool_t \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Boolq4'a8x_1_bufchan_buf ;
  assign \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Boolq4'a8x_1_bufchan_r  = (! \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Boolq4'a8x_1_bufchan_buf [0]);
  assign \q4'a8x_1_1_argbuf_d  = (\f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Boolq4'a8x_1_bufchan_buf [0] ? \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Boolq4'a8x_1_bufchan_buf  :
                                  \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Boolq4'a8x_1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Boolq4'a8x_1_bufchan_buf  <= {16'd0,
                                                                                                         1'd0};
    else
      if ((\q4'a8x_1_1_argbuf_r  && \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Boolq4'a8x_1_bufchan_buf [0]))
        \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Boolq4'a8x_1_bufchan_buf  <= {16'd0,
                                                                                                           1'd0};
      else if (((! \q4'a8x_1_1_argbuf_r ) && (! \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Boolq4'a8x_1_bufchan_buf [0])))
        \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Boolq4'a8x_1_bufchan_buf  <= \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Boolq4'a8x_1_bufchan_d ;
  
  /* buf (Ty Pointer_MaskQTree) : (f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Boolq4a8w_1,Pointer_MaskQTree) > (q4a8w_1_1_argbuf,Pointer_MaskQTree) */
  Pointer_MaskQTree_t \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Boolq4a8w_1_bufchan_d ;
  logic \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Boolq4a8w_1_bufchan_r ;
  assign \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Boolq4a8w_1_r  = ((! \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Boolq4a8w_1_bufchan_d [0]) || \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Boolq4a8w_1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Boolq4a8w_1_bufchan_d  <= {16'd0,
                                                                                                      1'd0};
    else
      if (\f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Boolq4a8w_1_r )
        \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Boolq4a8w_1_bufchan_d  <= \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Boolq4a8w_1_d ;
  Pointer_MaskQTree_t \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Boolq4a8w_1_bufchan_buf ;
  assign \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Boolq4a8w_1_bufchan_r  = (! \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Boolq4a8w_1_bufchan_buf [0]);
  assign q4a8w_1_1_argbuf_d = (\f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Boolq4a8w_1_bufchan_buf [0] ? \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Boolq4a8w_1_bufchan_buf  :
                               \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Boolq4a8w_1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Boolq4a8w_1_bufchan_buf  <= {16'd0,
                                                                                                        1'd0};
    else
      if ((q4a8w_1_1_argbuf_r && \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Boolq4a8w_1_bufchan_buf [0]))
        \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Boolq4a8w_1_bufchan_buf  <= {16'd0,
                                                                                                          1'd0};
      else if (((! q4a8w_1_1_argbuf_r) && (! \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Boolq4a8w_1_bufchan_buf [0])))
        \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Boolq4a8w_1_bufchan_buf  <= \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Boolq4a8w_1_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Bool) : (f'''''''''_f'''''''''_Bool_1,Pointer_QTree_Bool) > (f'''''''''_f'''''''''_Bool_resbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t \f'''''''''_f'''''''''_Bool_1_bufchan_d ;
  logic \f'''''''''_f'''''''''_Bool_1_bufchan_r ;
  assign \f'''''''''_f'''''''''_Bool_1_r  = ((! \f'''''''''_f'''''''''_Bool_1_bufchan_d [0]) || \f'''''''''_f'''''''''_Bool_1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f'''''''''_f'''''''''_Bool_1_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\f'''''''''_f'''''''''_Bool_1_r )
        \f'''''''''_f'''''''''_Bool_1_bufchan_d  <= \f'''''''''_f'''''''''_Bool_1_d ;
  Pointer_QTree_Bool_t \f'''''''''_f'''''''''_Bool_1_bufchan_buf ;
  assign \f'''''''''_f'''''''''_Bool_1_bufchan_r  = (! \f'''''''''_f'''''''''_Bool_1_bufchan_buf [0]);
  assign \f'''''''''_f'''''''''_Bool_resbuf_d  = (\f'''''''''_f'''''''''_Bool_1_bufchan_buf [0] ? \f'''''''''_f'''''''''_Bool_1_bufchan_buf  :
                                                  \f'''''''''_f'''''''''_Bool_1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f'''''''''_f'''''''''_Bool_1_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((\f'''''''''_f'''''''''_Bool_resbuf_r  && \f'''''''''_f'''''''''_Bool_1_bufchan_buf [0]))
        \f'''''''''_f'''''''''_Bool_1_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! \f'''''''''_f'''''''''_Bool_resbuf_r ) && (! \f'''''''''_f'''''''''_Bool_1_bufchan_buf [0])))
        \f'''''''''_f'''''''''_Bool_1_bufchan_buf  <= \f'''''''''_f'''''''''_Bool_1_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Bool) : (f'''''''''_f'''''''''_Bool_2,Pointer_QTree_Bool) > (f'''''''''_f'''''''''_Bool_2_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t \f'''''''''_f'''''''''_Bool_2_bufchan_d ;
  logic \f'''''''''_f'''''''''_Bool_2_bufchan_r ;
  assign \f'''''''''_f'''''''''_Bool_2_r  = ((! \f'''''''''_f'''''''''_Bool_2_bufchan_d [0]) || \f'''''''''_f'''''''''_Bool_2_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f'''''''''_f'''''''''_Bool_2_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\f'''''''''_f'''''''''_Bool_2_r )
        \f'''''''''_f'''''''''_Bool_2_bufchan_d  <= \f'''''''''_f'''''''''_Bool_2_d ;
  Pointer_QTree_Bool_t \f'''''''''_f'''''''''_Bool_2_bufchan_buf ;
  assign \f'''''''''_f'''''''''_Bool_2_bufchan_r  = (! \f'''''''''_f'''''''''_Bool_2_bufchan_buf [0]);
  assign \f'''''''''_f'''''''''_Bool_2_argbuf_d  = (\f'''''''''_f'''''''''_Bool_2_bufchan_buf [0] ? \f'''''''''_f'''''''''_Bool_2_bufchan_buf  :
                                                    \f'''''''''_f'''''''''_Bool_2_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f'''''''''_f'''''''''_Bool_2_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((\f'''''''''_f'''''''''_Bool_2_argbuf_r  && \f'''''''''_f'''''''''_Bool_2_bufchan_buf [0]))
        \f'''''''''_f'''''''''_Bool_2_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! \f'''''''''_f'''''''''_Bool_2_argbuf_r ) && (! \f'''''''''_f'''''''''_Bool_2_bufchan_buf [0])))
        \f'''''''''_f'''''''''_Bool_2_bufchan_buf  <= \f'''''''''_f'''''''''_Bool_2_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Bool) : (f'''''''''_f'''''''''_Bool_3,Pointer_QTree_Bool) > (f'''''''''_f'''''''''_Bool_3_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t \f'''''''''_f'''''''''_Bool_3_bufchan_d ;
  logic \f'''''''''_f'''''''''_Bool_3_bufchan_r ;
  assign \f'''''''''_f'''''''''_Bool_3_r  = ((! \f'''''''''_f'''''''''_Bool_3_bufchan_d [0]) || \f'''''''''_f'''''''''_Bool_3_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f'''''''''_f'''''''''_Bool_3_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\f'''''''''_f'''''''''_Bool_3_r )
        \f'''''''''_f'''''''''_Bool_3_bufchan_d  <= \f'''''''''_f'''''''''_Bool_3_d ;
  Pointer_QTree_Bool_t \f'''''''''_f'''''''''_Bool_3_bufchan_buf ;
  assign \f'''''''''_f'''''''''_Bool_3_bufchan_r  = (! \f'''''''''_f'''''''''_Bool_3_bufchan_buf [0]);
  assign \f'''''''''_f'''''''''_Bool_3_argbuf_d  = (\f'''''''''_f'''''''''_Bool_3_bufchan_buf [0] ? \f'''''''''_f'''''''''_Bool_3_bufchan_buf  :
                                                    \f'''''''''_f'''''''''_Bool_3_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f'''''''''_f'''''''''_Bool_3_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((\f'''''''''_f'''''''''_Bool_3_argbuf_r  && \f'''''''''_f'''''''''_Bool_3_bufchan_buf [0]))
        \f'''''''''_f'''''''''_Bool_3_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! \f'''''''''_f'''''''''_Bool_3_argbuf_r ) && (! \f'''''''''_f'''''''''_Bool_3_bufchan_buf [0])))
        \f'''''''''_f'''''''''_Bool_3_bufchan_buf  <= \f'''''''''_f'''''''''_Bool_3_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Bool) : (f'''''''''_f'''''''''_Bool_4,Pointer_QTree_Bool) > (f'''''''''_f'''''''''_Bool_4_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t \f'''''''''_f'''''''''_Bool_4_bufchan_d ;
  logic \f'''''''''_f'''''''''_Bool_4_bufchan_r ;
  assign \f'''''''''_f'''''''''_Bool_4_r  = ((! \f'''''''''_f'''''''''_Bool_4_bufchan_d [0]) || \f'''''''''_f'''''''''_Bool_4_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f'''''''''_f'''''''''_Bool_4_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\f'''''''''_f'''''''''_Bool_4_r )
        \f'''''''''_f'''''''''_Bool_4_bufchan_d  <= \f'''''''''_f'''''''''_Bool_4_d ;
  Pointer_QTree_Bool_t \f'''''''''_f'''''''''_Bool_4_bufchan_buf ;
  assign \f'''''''''_f'''''''''_Bool_4_bufchan_r  = (! \f'''''''''_f'''''''''_Bool_4_bufchan_buf [0]);
  assign \f'''''''''_f'''''''''_Bool_4_argbuf_d  = (\f'''''''''_f'''''''''_Bool_4_bufchan_buf [0] ? \f'''''''''_f'''''''''_Bool_4_bufchan_buf  :
                                                    \f'''''''''_f'''''''''_Bool_4_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f'''''''''_f'''''''''_Bool_4_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((\f'''''''''_f'''''''''_Bool_4_argbuf_r  && \f'''''''''_f'''''''''_Bool_4_bufchan_buf [0]))
        \f'''''''''_f'''''''''_Bool_4_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! \f'''''''''_f'''''''''_Bool_4_argbuf_r ) && (! \f'''''''''_f'''''''''_Bool_4_bufchan_buf [0])))
        \f'''''''''_f'''''''''_Bool_4_bufchan_buf  <= \f'''''''''_f'''''''''_Bool_4_bufchan_d ;
  
  /* dcon (Ty QTree_Bool,
      Dcon QNode_Bool) : [(f'''''''''_f'''''''''_Bool_4_argbuf,Pointer_QTree_Bool),
                          (f'''''''''_f'''''''''_Bool_3_argbuf,Pointer_QTree_Bool),
                          (f'''''''''_f'''''''''_Bool_2_argbuf,Pointer_QTree_Bool),
                          (f'''''''''_f'''''''''_Bool_resbuf,Pointer_QTree_Bool)] > (es_0_1es_1_1es_2_1es_3_1QNode_Bool,QTree_Bool) */
  assign es_0_1es_1_1es_2_1es_3_1QNode_Bool_d = QNode_Bool_dc((& {\f'''''''''_f'''''''''_Bool_4_argbuf_d [0],
                                                                  \f'''''''''_f'''''''''_Bool_3_argbuf_d [0],
                                                                  \f'''''''''_f'''''''''_Bool_2_argbuf_d [0],
                                                                  \f'''''''''_f'''''''''_Bool_resbuf_d [0]}), \f'''''''''_f'''''''''_Bool_4_argbuf_d , \f'''''''''_f'''''''''_Bool_3_argbuf_d , \f'''''''''_f'''''''''_Bool_2_argbuf_d , \f'''''''''_f'''''''''_Bool_resbuf_d );
  assign {\f'''''''''_f'''''''''_Bool_4_argbuf_r ,
          \f'''''''''_f'''''''''_Bool_3_argbuf_r ,
          \f'''''''''_f'''''''''_Bool_2_argbuf_r ,
          \f'''''''''_f'''''''''_Bool_resbuf_r } = {4 {(es_0_1es_1_1es_2_1es_3_1QNode_Bool_r && es_0_1es_1_1es_2_1es_3_1QNode_Bool_d[0])}};
  
  /* buf (Ty Pointer_QTree_Bool) : (f'''''''''_f'''''''''_Bool_5,Pointer_QTree_Bool) > (f'''''''''_f'''''''''_Bool_5_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t \f'''''''''_f'''''''''_Bool_5_bufchan_d ;
  logic \f'''''''''_f'''''''''_Bool_5_bufchan_r ;
  assign \f'''''''''_f'''''''''_Bool_5_r  = ((! \f'''''''''_f'''''''''_Bool_5_bufchan_d [0]) || \f'''''''''_f'''''''''_Bool_5_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f'''''''''_f'''''''''_Bool_5_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\f'''''''''_f'''''''''_Bool_5_r )
        \f'''''''''_f'''''''''_Bool_5_bufchan_d  <= \f'''''''''_f'''''''''_Bool_5_d ;
  Pointer_QTree_Bool_t \f'''''''''_f'''''''''_Bool_5_bufchan_buf ;
  assign \f'''''''''_f'''''''''_Bool_5_bufchan_r  = (! \f'''''''''_f'''''''''_Bool_5_bufchan_buf [0]);
  assign \f'''''''''_f'''''''''_Bool_5_argbuf_d  = (\f'''''''''_f'''''''''_Bool_5_bufchan_buf [0] ? \f'''''''''_f'''''''''_Bool_5_bufchan_buf  :
                                                    \f'''''''''_f'''''''''_Bool_5_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f'''''''''_f'''''''''_Bool_5_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((\f'''''''''_f'''''''''_Bool_5_argbuf_r  && \f'''''''''_f'''''''''_Bool_5_bufchan_buf [0]))
        \f'''''''''_f'''''''''_Bool_5_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! \f'''''''''_f'''''''''_Bool_5_argbuf_r ) && (! \f'''''''''_f'''''''''_Bool_5_bufchan_buf [0])))
        \f'''''''''_f'''''''''_Bool_5_bufchan_buf  <= \f'''''''''_f'''''''''_Bool_5_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Bool) : (f'''''''''_f'''''''''_Bool_6,Pointer_QTree_Bool) > (f'''''''''_f'''''''''_Bool_6_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t \f'''''''''_f'''''''''_Bool_6_bufchan_d ;
  logic \f'''''''''_f'''''''''_Bool_6_bufchan_r ;
  assign \f'''''''''_f'''''''''_Bool_6_r  = ((! \f'''''''''_f'''''''''_Bool_6_bufchan_d [0]) || \f'''''''''_f'''''''''_Bool_6_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f'''''''''_f'''''''''_Bool_6_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\f'''''''''_f'''''''''_Bool_6_r )
        \f'''''''''_f'''''''''_Bool_6_bufchan_d  <= \f'''''''''_f'''''''''_Bool_6_d ;
  Pointer_QTree_Bool_t \f'''''''''_f'''''''''_Bool_6_bufchan_buf ;
  assign \f'''''''''_f'''''''''_Bool_6_bufchan_r  = (! \f'''''''''_f'''''''''_Bool_6_bufchan_buf [0]);
  assign \f'''''''''_f'''''''''_Bool_6_argbuf_d  = (\f'''''''''_f'''''''''_Bool_6_bufchan_buf [0] ? \f'''''''''_f'''''''''_Bool_6_bufchan_buf  :
                                                    \f'''''''''_f'''''''''_Bool_6_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f'''''''''_f'''''''''_Bool_6_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((\f'''''''''_f'''''''''_Bool_6_argbuf_r  && \f'''''''''_f'''''''''_Bool_6_bufchan_buf [0]))
        \f'''''''''_f'''''''''_Bool_6_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! \f'''''''''_f'''''''''_Bool_6_argbuf_r ) && (! \f'''''''''_f'''''''''_Bool_6_bufchan_buf [0])))
        \f'''''''''_f'''''''''_Bool_6_bufchan_buf  <= \f'''''''''_f'''''''''_Bool_6_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Bool) : (f'''''''''_f'''''''''_Bool_7,Pointer_QTree_Bool) > (f'''''''''_f'''''''''_Bool_7_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t \f'''''''''_f'''''''''_Bool_7_bufchan_d ;
  logic \f'''''''''_f'''''''''_Bool_7_bufchan_r ;
  assign \f'''''''''_f'''''''''_Bool_7_r  = ((! \f'''''''''_f'''''''''_Bool_7_bufchan_d [0]) || \f'''''''''_f'''''''''_Bool_7_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f'''''''''_f'''''''''_Bool_7_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\f'''''''''_f'''''''''_Bool_7_r )
        \f'''''''''_f'''''''''_Bool_7_bufchan_d  <= \f'''''''''_f'''''''''_Bool_7_d ;
  Pointer_QTree_Bool_t \f'''''''''_f'''''''''_Bool_7_bufchan_buf ;
  assign \f'''''''''_f'''''''''_Bool_7_bufchan_r  = (! \f'''''''''_f'''''''''_Bool_7_bufchan_buf [0]);
  assign \f'''''''''_f'''''''''_Bool_7_argbuf_d  = (\f'''''''''_f'''''''''_Bool_7_bufchan_buf [0] ? \f'''''''''_f'''''''''_Bool_7_bufchan_buf  :
                                                    \f'''''''''_f'''''''''_Bool_7_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f'''''''''_f'''''''''_Bool_7_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((\f'''''''''_f'''''''''_Bool_7_argbuf_r  && \f'''''''''_f'''''''''_Bool_7_bufchan_buf [0]))
        \f'''''''''_f'''''''''_Bool_7_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! \f'''''''''_f'''''''''_Bool_7_argbuf_r ) && (! \f'''''''''_f'''''''''_Bool_7_bufchan_buf [0])))
        \f'''''''''_f'''''''''_Bool_7_bufchan_buf  <= \f'''''''''_f'''''''''_Bool_7_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Bool) : (f'''''''''_f'''''''''_Bool_8,Pointer_QTree_Bool) > (f'''''''''_f'''''''''_Bool_8_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t \f'''''''''_f'''''''''_Bool_8_bufchan_d ;
  logic \f'''''''''_f'''''''''_Bool_8_bufchan_r ;
  assign \f'''''''''_f'''''''''_Bool_8_r  = ((! \f'''''''''_f'''''''''_Bool_8_bufchan_d [0]) || \f'''''''''_f'''''''''_Bool_8_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f'''''''''_f'''''''''_Bool_8_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\f'''''''''_f'''''''''_Bool_8_r )
        \f'''''''''_f'''''''''_Bool_8_bufchan_d  <= \f'''''''''_f'''''''''_Bool_8_d ;
  Pointer_QTree_Bool_t \f'''''''''_f'''''''''_Bool_8_bufchan_buf ;
  assign \f'''''''''_f'''''''''_Bool_8_bufchan_r  = (! \f'''''''''_f'''''''''_Bool_8_bufchan_buf [0]);
  assign \f'''''''''_f'''''''''_Bool_8_argbuf_d  = (\f'''''''''_f'''''''''_Bool_8_bufchan_buf [0] ? \f'''''''''_f'''''''''_Bool_8_bufchan_buf  :
                                                    \f'''''''''_f'''''''''_Bool_8_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f'''''''''_f'''''''''_Bool_8_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((\f'''''''''_f'''''''''_Bool_8_argbuf_r  && \f'''''''''_f'''''''''_Bool_8_bufchan_buf [0]))
        \f'''''''''_f'''''''''_Bool_8_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! \f'''''''''_f'''''''''_Bool_8_argbuf_r ) && (! \f'''''''''_f'''''''''_Bool_8_bufchan_buf [0])))
        \f'''''''''_f'''''''''_Bool_8_bufchan_buf  <= \f'''''''''_f'''''''''_Bool_8_bufchan_d ;
  
  /* dcon (Ty QTree_Bool,
      Dcon QNode_Bool) : [(f'''''''''_f'''''''''_Bool_8_argbuf,Pointer_QTree_Bool),
                          (f'''''''''_f'''''''''_Bool_7_argbuf,Pointer_QTree_Bool),
                          (f'''''''''_f'''''''''_Bool_6_argbuf,Pointer_QTree_Bool),
                          (f'''''''''_f'''''''''_Bool_5_argbuf,Pointer_QTree_Bool)] > (es_4_1es_5_1es_6_1es_7_1QNode_Bool,QTree_Bool) */
  assign es_4_1es_5_1es_6_1es_7_1QNode_Bool_d = QNode_Bool_dc((& {\f'''''''''_f'''''''''_Bool_8_argbuf_d [0],
                                                                  \f'''''''''_f'''''''''_Bool_7_argbuf_d [0],
                                                                  \f'''''''''_f'''''''''_Bool_6_argbuf_d [0],
                                                                  \f'''''''''_f'''''''''_Bool_5_argbuf_d [0]}), \f'''''''''_f'''''''''_Bool_8_argbuf_d , \f'''''''''_f'''''''''_Bool_7_argbuf_d , \f'''''''''_f'''''''''_Bool_6_argbuf_d , \f'''''''''_f'''''''''_Bool_5_argbuf_d );
  assign {\f'''''''''_f'''''''''_Bool_8_argbuf_r ,
          \f'''''''''_f'''''''''_Bool_7_argbuf_r ,
          \f'''''''''_f'''''''''_Bool_6_argbuf_r ,
          \f'''''''''_f'''''''''_Bool_5_argbuf_r } = {4 {(es_4_1es_5_1es_6_1es_7_1QNode_Bool_r && es_4_1es_5_1es_6_1es_7_1QNode_Bool_d[0])}};
  
  /* demux (Ty C8,
       Ty Pointer_QTree_Bool) : (f'''''''''_f'''''''''_Bool_choice,C8) (lizzieLet53_4Lf'''''''''_f'''''''''_Boolsbos_1_merge_merge_fork_2,Pointer_QTree_Bool) > [(f'''''''''_f'''''''''_Bool_1,Pointer_QTree_Bool),
                                                                                                                                                                 (f'''''''''_f'''''''''_Bool_2,Pointer_QTree_Bool),
                                                                                                                                                                 (f'''''''''_f'''''''''_Bool_3,Pointer_QTree_Bool),
                                                                                                                                                                 (f'''''''''_f'''''''''_Bool_4,Pointer_QTree_Bool),
                                                                                                                                                                 (f'''''''''_f'''''''''_Bool_5,Pointer_QTree_Bool),
                                                                                                                                                                 (f'''''''''_f'''''''''_Bool_6,Pointer_QTree_Bool),
                                                                                                                                                                 (f'''''''''_f'''''''''_Bool_7,Pointer_QTree_Bool),
                                                                                                                                                                 (f'''''''''_f'''''''''_Bool_8,Pointer_QTree_Bool)] */
  logic [7:0] \lizzieLet53_4Lf'''''''''_f'''''''''_Boolsbos_1_merge_merge_fork_2_onehotd ;
  always_comb
    if ((\f'''''''''_f'''''''''_Bool_choice_d [0] && \lizzieLet53_4Lf'''''''''_f'''''''''_Boolsbos_1_merge_merge_fork_2_d [0]))
      unique case (\f'''''''''_f'''''''''_Bool_choice_d [3:1])
        3'd0:
          \lizzieLet53_4Lf'''''''''_f'''''''''_Boolsbos_1_merge_merge_fork_2_onehotd  = 8'd1;
        3'd1:
          \lizzieLet53_4Lf'''''''''_f'''''''''_Boolsbos_1_merge_merge_fork_2_onehotd  = 8'd2;
        3'd2:
          \lizzieLet53_4Lf'''''''''_f'''''''''_Boolsbos_1_merge_merge_fork_2_onehotd  = 8'd4;
        3'd3:
          \lizzieLet53_4Lf'''''''''_f'''''''''_Boolsbos_1_merge_merge_fork_2_onehotd  = 8'd8;
        3'd4:
          \lizzieLet53_4Lf'''''''''_f'''''''''_Boolsbos_1_merge_merge_fork_2_onehotd  = 8'd16;
        3'd5:
          \lizzieLet53_4Lf'''''''''_f'''''''''_Boolsbos_1_merge_merge_fork_2_onehotd  = 8'd32;
        3'd6:
          \lizzieLet53_4Lf'''''''''_f'''''''''_Boolsbos_1_merge_merge_fork_2_onehotd  = 8'd64;
        3'd7:
          \lizzieLet53_4Lf'''''''''_f'''''''''_Boolsbos_1_merge_merge_fork_2_onehotd  = 8'd128;
        default:
          \lizzieLet53_4Lf'''''''''_f'''''''''_Boolsbos_1_merge_merge_fork_2_onehotd  = 8'd0;
      endcase
    else
      \lizzieLet53_4Lf'''''''''_f'''''''''_Boolsbos_1_merge_merge_fork_2_onehotd  = 8'd0;
  assign \f'''''''''_f'''''''''_Bool_1_d  = {\lizzieLet53_4Lf'''''''''_f'''''''''_Boolsbos_1_merge_merge_fork_2_d [16:1],
                                             \lizzieLet53_4Lf'''''''''_f'''''''''_Boolsbos_1_merge_merge_fork_2_onehotd [0]};
  assign \f'''''''''_f'''''''''_Bool_2_d  = {\lizzieLet53_4Lf'''''''''_f'''''''''_Boolsbos_1_merge_merge_fork_2_d [16:1],
                                             \lizzieLet53_4Lf'''''''''_f'''''''''_Boolsbos_1_merge_merge_fork_2_onehotd [1]};
  assign \f'''''''''_f'''''''''_Bool_3_d  = {\lizzieLet53_4Lf'''''''''_f'''''''''_Boolsbos_1_merge_merge_fork_2_d [16:1],
                                             \lizzieLet53_4Lf'''''''''_f'''''''''_Boolsbos_1_merge_merge_fork_2_onehotd [2]};
  assign \f'''''''''_f'''''''''_Bool_4_d  = {\lizzieLet53_4Lf'''''''''_f'''''''''_Boolsbos_1_merge_merge_fork_2_d [16:1],
                                             \lizzieLet53_4Lf'''''''''_f'''''''''_Boolsbos_1_merge_merge_fork_2_onehotd [3]};
  assign \f'''''''''_f'''''''''_Bool_5_d  = {\lizzieLet53_4Lf'''''''''_f'''''''''_Boolsbos_1_merge_merge_fork_2_d [16:1],
                                             \lizzieLet53_4Lf'''''''''_f'''''''''_Boolsbos_1_merge_merge_fork_2_onehotd [4]};
  assign \f'''''''''_f'''''''''_Bool_6_d  = {\lizzieLet53_4Lf'''''''''_f'''''''''_Boolsbos_1_merge_merge_fork_2_d [16:1],
                                             \lizzieLet53_4Lf'''''''''_f'''''''''_Boolsbos_1_merge_merge_fork_2_onehotd [5]};
  assign \f'''''''''_f'''''''''_Bool_7_d  = {\lizzieLet53_4Lf'''''''''_f'''''''''_Boolsbos_1_merge_merge_fork_2_d [16:1],
                                             \lizzieLet53_4Lf'''''''''_f'''''''''_Boolsbos_1_merge_merge_fork_2_onehotd [6]};
  assign \f'''''''''_f'''''''''_Bool_8_d  = {\lizzieLet53_4Lf'''''''''_f'''''''''_Boolsbos_1_merge_merge_fork_2_d [16:1],
                                             \lizzieLet53_4Lf'''''''''_f'''''''''_Boolsbos_1_merge_merge_fork_2_onehotd [7]};
  assign \lizzieLet53_4Lf'''''''''_f'''''''''_Boolsbos_1_merge_merge_fork_2_r  = (| (\lizzieLet53_4Lf'''''''''_f'''''''''_Boolsbos_1_merge_merge_fork_2_onehotd  & {\f'''''''''_f'''''''''_Bool_8_r ,
                                                                                                                                                                    \f'''''''''_f'''''''''_Bool_7_r ,
                                                                                                                                                                    \f'''''''''_f'''''''''_Bool_6_r ,
                                                                                                                                                                    \f'''''''''_f'''''''''_Bool_5_r ,
                                                                                                                                                                    \f'''''''''_f'''''''''_Bool_4_r ,
                                                                                                                                                                    \f'''''''''_f'''''''''_Bool_3_r ,
                                                                                                                                                                    \f'''''''''_f'''''''''_Bool_2_r ,
                                                                                                                                                                    \f'''''''''_f'''''''''_Bool_1_r }));
  assign \f'''''''''_f'''''''''_Bool_choice_r  = \lizzieLet53_4Lf'''''''''_f'''''''''_Boolsbos_1_merge_merge_fork_2_r ;
  
  /* destruct (Ty TupGo___Pointer_MaskQTree___Pointer_QTree_Bool,
          Dcon TupGo___Pointer_MaskQTree___Pointer_QTree_Bool) : (f'''''''''_f'''''''''_Bool_data,TupGo___Pointer_MaskQTree___Pointer_QTree_Bool) > [(f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Boolgo_7,Go),
                                                                                                                                                     (f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Boolq4a8w_1,Pointer_MaskQTree),
                                                                                                                                                     (f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Boolq4'a8x_1,Pointer_QTree_Bool)] */
  logic [2:0] \f'''''''''_f'''''''''_Bool_data_emitted ;
  logic [2:0] \f'''''''''_f'''''''''_Bool_data_done ;
  assign \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Boolgo_7_d  = (\f'''''''''_f'''''''''_Bool_data_d [0] && (! \f'''''''''_f'''''''''_Bool_data_emitted [0]));
  assign \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Boolq4a8w_1_d  = {\f'''''''''_f'''''''''_Bool_data_d [16:1],
                                                                                                (\f'''''''''_f'''''''''_Bool_data_d [0] && (! \f'''''''''_f'''''''''_Bool_data_emitted [1]))};
  assign \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Boolq4'a8x_1_d  = {\f'''''''''_f'''''''''_Bool_data_d [32:17],
                                                                                                 (\f'''''''''_f'''''''''_Bool_data_d [0] && (! \f'''''''''_f'''''''''_Bool_data_emitted [2]))};
  assign \f'''''''''_f'''''''''_Bool_data_done  = (\f'''''''''_f'''''''''_Bool_data_emitted  | ({\f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Boolq4'a8x_1_d [0],
                                                                                                 \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Boolq4a8w_1_d [0],
                                                                                                 \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Boolgo_7_d [0]} & {\f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Boolq4'a8x_1_r ,
                                                                                                                                                                                         \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Boolq4a8w_1_r ,
                                                                                                                                                                                         \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Boolgo_7_r }));
  assign \f'''''''''_f'''''''''_Bool_data_r  = (& \f'''''''''_f'''''''''_Bool_data_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f'''''''''_f'''''''''_Bool_data_emitted  <= 3'd0;
    else
      \f'''''''''_f'''''''''_Bool_data_emitted  <= (\f'''''''''_f'''''''''_Bool_data_r  ? 3'd0 :
                                                    \f'''''''''_f'''''''''_Bool_data_done );
  
  /* destruct (Ty TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool,
          Dcon TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool) : (f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_1,TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool) > [(f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolgo_6,Go),
                                                                                                                                                                           (f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolm2a8H_1,Pointer_QTree_Bool),
                                                                                                                                                                           (f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolm3a8I_1,Pointer_QTree_Bool)] */
  logic [2:0] \f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_1_emitted ;
  logic [2:0] \f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_1_done ;
  assign \f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolgo_6_d  = (\f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_1_d [0] && (! \f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_1_emitted [0]));
  assign \f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolm2a8H_1_d  = {\f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_1_d [16:1],
                                                                         (\f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_1_d [0] && (! \f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_1_emitted [1]))};
  assign \f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolm3a8I_1_d  = {\f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_1_d [32:17],
                                                                         (\f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_1_d [0] && (! \f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_1_emitted [2]))};
  assign \f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_1_done  = (\f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_1_emitted  | ({\f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolm3a8I_1_d [0],
                                                                                                                                         \f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolm2a8H_1_d [0],
                                                                                                                                         \f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolgo_6_d [0]} & {\f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolm3a8I_1_r ,
                                                                                                                                                                                                          \f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolm2a8H_1_r ,
                                                                                                                                                                                                          \f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolgo_6_r }));
  assign \f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_1_r  = (& \f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_1_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_1_emitted  <= 3'd0;
    else
      \f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_1_emitted  <= (\f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_1_r  ? 3'd0 :
                                                                        \f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_1_done );
  
  /* fork (Ty Go) : (f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolgo_6,Go) > [(go_6_1,Go),
                                                                             (go_6_2,Go)] */
  logic [1:0] \f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolgo_6_emitted ;
  logic [1:0] \f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolgo_6_done ;
  assign go_6_1_d = (\f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolgo_6_d [0] && (! \f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolgo_6_emitted [0]));
  assign go_6_2_d = (\f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolgo_6_d [0] && (! \f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolgo_6_emitted [1]));
  assign \f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolgo_6_done  = (\f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolgo_6_emitted  | ({go_6_2_d[0],
                                                                                                                                             go_6_1_d[0]} & {go_6_2_r,
                                                                                                                                                             go_6_1_r}));
  assign \f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolgo_6_r  = (& \f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolgo_6_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolgo_6_emitted  <= 2'd0;
    else
      \f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolgo_6_emitted  <= (\f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolgo_6_r  ? 2'd0 :
                                                                          \f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolgo_6_done );
  
  /* buf (Ty Pointer_QTree_Bool) : (f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolm2a8H_1,Pointer_QTree_Bool) > (m2a8H_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t \f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolm2a8H_1_bufchan_d ;
  logic \f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolm2a8H_1_bufchan_r ;
  assign \f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolm2a8H_1_r  = ((! \f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolm2a8H_1_bufchan_d [0]) || \f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolm2a8H_1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolm2a8H_1_bufchan_d  <= {16'd0,
                                                                               1'd0};
    else
      if (\f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolm2a8H_1_r )
        \f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolm2a8H_1_bufchan_d  <= \f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolm2a8H_1_d ;
  Pointer_QTree_Bool_t \f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolm2a8H_1_bufchan_buf ;
  assign \f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolm2a8H_1_bufchan_r  = (! \f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolm2a8H_1_bufchan_buf [0]);
  assign m2a8H_1_1_argbuf_d = (\f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolm2a8H_1_bufchan_buf [0] ? \f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolm2a8H_1_bufchan_buf  :
                               \f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolm2a8H_1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolm2a8H_1_bufchan_buf  <= {16'd0,
                                                                                 1'd0};
    else
      if ((m2a8H_1_1_argbuf_r && \f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolm2a8H_1_bufchan_buf [0]))
        \f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolm2a8H_1_bufchan_buf  <= {16'd0,
                                                                                   1'd0};
      else if (((! m2a8H_1_1_argbuf_r) && (! \f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolm2a8H_1_bufchan_buf [0])))
        \f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolm2a8H_1_bufchan_buf  <= \f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolm2a8H_1_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Bool) : (f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolm3a8I_1,Pointer_QTree_Bool) > (m3a8I_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t \f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolm3a8I_1_bufchan_d ;
  logic \f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolm3a8I_1_bufchan_r ;
  assign \f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolm3a8I_1_r  = ((! \f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolm3a8I_1_bufchan_d [0]) || \f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolm3a8I_1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolm3a8I_1_bufchan_d  <= {16'd0,
                                                                               1'd0};
    else
      if (\f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolm3a8I_1_r )
        \f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolm3a8I_1_bufchan_d  <= \f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolm3a8I_1_d ;
  Pointer_QTree_Bool_t \f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolm3a8I_1_bufchan_buf ;
  assign \f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolm3a8I_1_bufchan_r  = (! \f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolm3a8I_1_bufchan_buf [0]);
  assign m3a8I_1_1_argbuf_d = (\f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolm3a8I_1_bufchan_buf [0] ? \f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolm3a8I_1_bufchan_buf  :
                               \f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolm3a8I_1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolm3a8I_1_bufchan_buf  <= {16'd0,
                                                                                 1'd0};
    else
      if ((m3a8I_1_1_argbuf_r && \f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolm3a8I_1_bufchan_buf [0]))
        \f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolm3a8I_1_bufchan_buf  <= {16'd0,
                                                                                   1'd0};
      else if (((! m3a8I_1_1_argbuf_r) && (! \f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolm3a8I_1_bufchan_buf [0])))
        \f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolm3a8I_1_bufchan_buf  <= \f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Boolm3a8I_1_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Bool) : (f'_resbuf,Pointer_QTree_Bool) > (lizzieLet14_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t \f'_resbuf_bufchan_d ;
  logic \f'_resbuf_bufchan_r ;
  assign \f'_resbuf_r  = ((! \f'_resbuf_bufchan_d [0]) || \f'_resbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \f'_resbuf_bufchan_d  <= {16'd0, 1'd0};
    else if (\f'_resbuf_r ) \f'_resbuf_bufchan_d  <= \f'_resbuf_d ;
  Pointer_QTree_Bool_t \f'_resbuf_bufchan_buf ;
  assign \f'_resbuf_bufchan_r  = (! \f'_resbuf_bufchan_buf [0]);
  assign lizzieLet14_1_argbuf_d = (\f'_resbuf_bufchan_buf [0] ? \f'_resbuf_bufchan_buf  :
                                   \f'_resbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \f'_resbuf_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((lizzieLet14_1_argbuf_r && \f'_resbuf_bufchan_buf [0]))
        \f'_resbuf_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! lizzieLet14_1_argbuf_r) && (! \f'_resbuf_bufchan_buf [0])))
        \f'_resbuf_bufchan_buf  <= \f'_resbuf_bufchan_d ;
  
  /* destruct (Ty TupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool,
          Dcon TupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool) : (fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool_1,TupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool) > [(fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Boolgo_5,Go),
                                                                                                                                                                                                                                      (fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Boolm1a85_1,Pointer_MaskQTree),
                                                                                                                                                                                                                                      (fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Boolm2a86_1,Pointer_QTree_Bool),
                                                                                                                                                                                                                                      (fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Boolm3a87_1,Pointer_QTree_Bool)] */
  logic [3:0] fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool_1_emitted;
  logic [3:0] fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool_1_done;
  assign fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Boolgo_5_d = (fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool_1_d[0] && (! fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool_1_emitted[0]));
  assign fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Boolm1a85_1_d = {fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool_1_d[16:1],
                                                                                          (fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool_1_d[0] && (! fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool_1_emitted[1]))};
  assign fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Boolm2a86_1_d = {fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool_1_d[32:17],
                                                                                          (fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool_1_d[0] && (! fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool_1_emitted[2]))};
  assign fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Boolm3a87_1_d = {fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool_1_d[48:33],
                                                                                          (fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool_1_d[0] && (! fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool_1_emitted[3]))};
  assign fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool_1_done = (fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool_1_emitted | ({fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Boolm3a87_1_d[0],
                                                                                                                                                                           fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Boolm2a86_1_d[0],
                                                                                                                                                                           fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Boolm1a85_1_d[0],
                                                                                                                                                                           fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Boolgo_5_d[0]} & {fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Boolm3a87_1_r,
                                                                                                                                                                                                                                                             fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Boolm2a86_1_r,
                                                                                                                                                                                                                                                             fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Boolm1a85_1_r,
                                                                                                                                                                                                                                                             fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Boolgo_5_r}));
  assign fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool_1_r = (& fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool_1_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool_1_emitted <= 4'd0;
    else
      fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool_1_emitted <= (fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool_1_r ? 4'd0 :
                                                                                         fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool_1_done);
  
  /* fork (Ty Go) : (fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Boolgo_5,Go) > [(go_5_1,Go),
                                                                                                (go_5_2,Go)] */
  logic [1:0] fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Boolgo_5_emitted;
  logic [1:0] fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Boolgo_5_done;
  assign go_5_1_d = (fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Boolgo_5_d[0] && (! fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Boolgo_5_emitted[0]));
  assign go_5_2_d = (fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Boolgo_5_d[0] && (! fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Boolgo_5_emitted[1]));
  assign fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Boolgo_5_done = (fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Boolgo_5_emitted | ({go_5_2_d[0],
                                                                                                                                                                               go_5_1_d[0]} & {go_5_2_r,
                                                                                                                                                                                               go_5_1_r}));
  assign fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Boolgo_5_r = (& fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Boolgo_5_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Boolgo_5_emitted <= 2'd0;
    else
      fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Boolgo_5_emitted <= (fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Boolgo_5_r ? 2'd0 :
                                                                                           fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Boolgo_5_done);
  
  /* buf (Ty Pointer_MaskQTree) : (fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Boolm1a85_1,Pointer_MaskQTree) > (m1a85_1_1_argbuf,Pointer_MaskQTree) */
  Pointer_MaskQTree_t fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Boolm1a85_1_bufchan_d;
  logic fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Boolm1a85_1_bufchan_r;
  assign fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Boolm1a85_1_r = ((! fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Boolm1a85_1_bufchan_d[0]) || fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Boolm1a85_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Boolm1a85_1_bufchan_d <= {16'd0,
                                                                                                1'd0};
    else
      if (fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Boolm1a85_1_r)
        fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Boolm1a85_1_bufchan_d <= fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Boolm1a85_1_d;
  Pointer_MaskQTree_t fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Boolm1a85_1_bufchan_buf;
  assign fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Boolm1a85_1_bufchan_r = (! fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Boolm1a85_1_bufchan_buf[0]);
  assign m1a85_1_1_argbuf_d = (fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Boolm1a85_1_bufchan_buf[0] ? fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Boolm1a85_1_bufchan_buf :
                               fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Boolm1a85_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Boolm1a85_1_bufchan_buf <= {16'd0,
                                                                                                  1'd0};
    else
      if ((m1a85_1_1_argbuf_r && fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Boolm1a85_1_bufchan_buf[0]))
        fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Boolm1a85_1_bufchan_buf <= {16'd0,
                                                                                                    1'd0};
      else if (((! m1a85_1_1_argbuf_r) && (! fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Boolm1a85_1_bufchan_buf[0])))
        fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Boolm1a85_1_bufchan_buf <= fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Boolm1a85_1_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Boolm2a86_1,Pointer_QTree_Bool) > (m2a86_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Boolm2a86_1_bufchan_d;
  logic fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Boolm2a86_1_bufchan_r;
  assign fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Boolm2a86_1_r = ((! fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Boolm2a86_1_bufchan_d[0]) || fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Boolm2a86_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Boolm2a86_1_bufchan_d <= {16'd0,
                                                                                                1'd0};
    else
      if (fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Boolm2a86_1_r)
        fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Boolm2a86_1_bufchan_d <= fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Boolm2a86_1_d;
  Pointer_QTree_Bool_t fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Boolm2a86_1_bufchan_buf;
  assign fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Boolm2a86_1_bufchan_r = (! fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Boolm2a86_1_bufchan_buf[0]);
  assign m2a86_1_1_argbuf_d = (fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Boolm2a86_1_bufchan_buf[0] ? fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Boolm2a86_1_bufchan_buf :
                               fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Boolm2a86_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Boolm2a86_1_bufchan_buf <= {16'd0,
                                                                                                  1'd0};
    else
      if ((m2a86_1_1_argbuf_r && fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Boolm2a86_1_bufchan_buf[0]))
        fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Boolm2a86_1_bufchan_buf <= {16'd0,
                                                                                                    1'd0};
      else if (((! m2a86_1_1_argbuf_r) && (! fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Boolm2a86_1_bufchan_buf[0])))
        fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Boolm2a86_1_bufchan_buf <= fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Boolm2a86_1_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Boolm3a87_1,Pointer_QTree_Bool) > (m3a87_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Boolm3a87_1_bufchan_d;
  logic fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Boolm3a87_1_bufchan_r;
  assign fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Boolm3a87_1_r = ((! fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Boolm3a87_1_bufchan_d[0]) || fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Boolm3a87_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Boolm3a87_1_bufchan_d <= {16'd0,
                                                                                                1'd0};
    else
      if (fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Boolm3a87_1_r)
        fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Boolm3a87_1_bufchan_d <= fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Boolm3a87_1_d;
  Pointer_QTree_Bool_t fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Boolm3a87_1_bufchan_buf;
  assign fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Boolm3a87_1_bufchan_r = (! fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Boolm3a87_1_bufchan_buf[0]);
  assign m3a87_1_1_argbuf_d = (fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Boolm3a87_1_bufchan_buf[0] ? fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Boolm3a87_1_bufchan_buf :
                               fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Boolm3a87_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Boolm3a87_1_bufchan_buf <= {16'd0,
                                                                                                  1'd0};
    else
      if ((m3a87_1_1_argbuf_r && fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Boolm3a87_1_bufchan_buf[0]))
        fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Boolm3a87_1_bufchan_buf <= {16'd0,
                                                                                                    1'd0};
      else if (((! m3a87_1_1_argbuf_r) && (! fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Boolm3a87_1_bufchan_buf[0])))
        fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Boolm3a87_1_bufchan_buf <= fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Boolm3a87_1_bufchan_d;
  
  /* sink (Ty Pointer_QTree_Bool) : (f_resbuf,Pointer_QTree_Bool) > */
  assign {f_resbuf_r, f_resbuf_dout} = {f_resbuf_rout, f_resbuf_d};
  
  /* fork (Ty C12) : (go_10_goMux_choice,C12) > [(go_10_goMux_choice_1,C12),
                                            (go_10_goMux_choice_2,C12)] */
  logic [1:0] go_10_goMux_choice_emitted;
  logic [1:0] go_10_goMux_choice_done;
  assign go_10_goMux_choice_1_d = {go_10_goMux_choice_d[4:1],
                                   (go_10_goMux_choice_d[0] && (! go_10_goMux_choice_emitted[0]))};
  assign go_10_goMux_choice_2_d = {go_10_goMux_choice_d[4:1],
                                   (go_10_goMux_choice_d[0] && (! go_10_goMux_choice_emitted[1]))};
  assign go_10_goMux_choice_done = (go_10_goMux_choice_emitted | ({go_10_goMux_choice_2_d[0],
                                                                   go_10_goMux_choice_1_d[0]} & {go_10_goMux_choice_2_r,
                                                                                                 go_10_goMux_choice_1_r}));
  assign go_10_goMux_choice_r = (& go_10_goMux_choice_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_10_goMux_choice_emitted <= 2'd0;
    else
      go_10_goMux_choice_emitted <= (go_10_goMux_choice_r ? 2'd0 :
                                     go_10_goMux_choice_done);
  
  /* mux (Ty C12,
     Ty Pointer_QTree_Bool) : (go_10_goMux_choice_1,C12) [(lizzieLet20_1_6QNone_Bool_1_argbuf,Pointer_QTree_Bool),
                                                          (contRet_0_1_1_argbuf,Pointer_QTree_Bool),
                                                          (lizzieLet20_1_4QVal_Bool_4QNone_Bool_1_argbuf,Pointer_QTree_Bool),
                                                          (lizzieLet6_1_1_argbuf,Pointer_QTree_Bool),
                                                          (lizzieLet23_1_1_argbuf,Pointer_QTree_Bool),
                                                          (lizzieLet24_1_1_argbuf,Pointer_QTree_Bool),
                                                          (lizzieLet7_1_1_argbuf,Pointer_QTree_Bool),
                                                          (lizzieLet8_1_argbuf,Pointer_QTree_Bool),
                                                          (lizzieLet20_1_4QNode_Bool_4QNone_Bool_1_argbuf,Pointer_QTree_Bool),
                                                          (lizzieLet9_2_1_argbuf,Pointer_QTree_Bool),
                                                          (lizzieLet10_1_1_argbuf,Pointer_QTree_Bool),
                                                          (lizzieLet11_1_1_argbuf,Pointer_QTree_Bool)] > (srtarg_0_1_goMux_mux,Pointer_QTree_Bool) */
  logic [16:0] srtarg_0_1_goMux_mux_mux;
  logic [11:0] srtarg_0_1_goMux_mux_onehot;
  always_comb
    unique case (go_10_goMux_choice_1_d[4:1])
      4'd0:
        {srtarg_0_1_goMux_mux_onehot, srtarg_0_1_goMux_mux_mux} = {12'd1,
                                                                   lizzieLet20_1_6QNone_Bool_1_argbuf_d};
      4'd1:
        {srtarg_0_1_goMux_mux_onehot, srtarg_0_1_goMux_mux_mux} = {12'd2,
                                                                   contRet_0_1_1_argbuf_d};
      4'd2:
        {srtarg_0_1_goMux_mux_onehot, srtarg_0_1_goMux_mux_mux} = {12'd4,
                                                                   lizzieLet20_1_4QVal_Bool_4QNone_Bool_1_argbuf_d};
      4'd3:
        {srtarg_0_1_goMux_mux_onehot, srtarg_0_1_goMux_mux_mux} = {12'd8,
                                                                   lizzieLet6_1_1_argbuf_d};
      4'd4:
        {srtarg_0_1_goMux_mux_onehot, srtarg_0_1_goMux_mux_mux} = {12'd16,
                                                                   lizzieLet23_1_1_argbuf_d};
      4'd5:
        {srtarg_0_1_goMux_mux_onehot, srtarg_0_1_goMux_mux_mux} = {12'd32,
                                                                   lizzieLet24_1_1_argbuf_d};
      4'd6:
        {srtarg_0_1_goMux_mux_onehot, srtarg_0_1_goMux_mux_mux} = {12'd64,
                                                                   lizzieLet7_1_1_argbuf_d};
      4'd7:
        {srtarg_0_1_goMux_mux_onehot, srtarg_0_1_goMux_mux_mux} = {12'd128,
                                                                   lizzieLet8_1_argbuf_d};
      4'd8:
        {srtarg_0_1_goMux_mux_onehot, srtarg_0_1_goMux_mux_mux} = {12'd256,
                                                                   lizzieLet20_1_4QNode_Bool_4QNone_Bool_1_argbuf_d};
      4'd9:
        {srtarg_0_1_goMux_mux_onehot, srtarg_0_1_goMux_mux_mux} = {12'd512,
                                                                   lizzieLet9_2_1_argbuf_d};
      4'd10:
        {srtarg_0_1_goMux_mux_onehot,
         srtarg_0_1_goMux_mux_mux} = {12'd1024, lizzieLet10_1_1_argbuf_d};
      4'd11:
        {srtarg_0_1_goMux_mux_onehot,
         srtarg_0_1_goMux_mux_mux} = {12'd2048, lizzieLet11_1_1_argbuf_d};
      default:
        {srtarg_0_1_goMux_mux_onehot, srtarg_0_1_goMux_mux_mux} = {12'd0,
                                                                   {16'd0, 1'd0}};
    endcase
  assign srtarg_0_1_goMux_mux_d = {srtarg_0_1_goMux_mux_mux[16:1],
                                   (srtarg_0_1_goMux_mux_mux[0] && go_10_goMux_choice_1_d[0])};
  assign go_10_goMux_choice_1_r = (srtarg_0_1_goMux_mux_d[0] && srtarg_0_1_goMux_mux_r);
  assign {lizzieLet11_1_1_argbuf_r,
          lizzieLet10_1_1_argbuf_r,
          lizzieLet9_2_1_argbuf_r,
          lizzieLet20_1_4QNode_Bool_4QNone_Bool_1_argbuf_r,
          lizzieLet8_1_argbuf_r,
          lizzieLet7_1_1_argbuf_r,
          lizzieLet24_1_1_argbuf_r,
          lizzieLet23_1_1_argbuf_r,
          lizzieLet6_1_1_argbuf_r,
          lizzieLet20_1_4QVal_Bool_4QNone_Bool_1_argbuf_r,
          contRet_0_1_1_argbuf_r,
          lizzieLet20_1_6QNone_Bool_1_argbuf_r} = (go_10_goMux_choice_1_r ? srtarg_0_1_goMux_mux_onehot :
                                                   12'd0);
  
  /* mux (Ty C12,
     Ty Pointer_CTf') : (go_10_goMux_choice_2,C12) [(lizzieLet20_1_7QNone_Bool_1_argbuf,Pointer_CTf'),
                                                    (sc_0_10_1_argbuf,Pointer_CTf'),
                                                    (lizzieLet20_1_4QVal_Bool_5QNone_Bool_1_argbuf,Pointer_CTf'),
                                                    (lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_2MyFalse_1_argbuf,Pointer_CTf'),
                                                    (lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_2MyTrue_1_argbuf,Pointer_CTf'),
                                                    (lizzieLet20_1_4QVal_Bool_6QVal_Bool_2MyTrue_1_argbuf,Pointer_CTf'),
                                                    (lizzieLet20_1_4QVal_Bool_5QNode_Bool_1_argbuf,Pointer_CTf'),
                                                    (lizzieLet20_1_4QVal_Bool_5QError_Bool_1_argbuf,Pointer_CTf'),
                                                    (lizzieLet20_1_4QNode_Bool_5QNone_Bool_1_argbuf,Pointer_CTf'),
                                                    (lizzieLet20_1_4QNode_Bool_5QVal_Bool_1_argbuf,Pointer_CTf'),
                                                    (lizzieLet20_1_4QNode_Bool_5QError_Bool_1_argbuf,Pointer_CTf'),
                                                    (lizzieLet20_1_7QError_Bool_1_argbuf,Pointer_CTf')] > (scfarg_0_1_goMux_mux,Pointer_CTf') */
  logic [16:0] scfarg_0_1_goMux_mux_mux;
  logic [11:0] scfarg_0_1_goMux_mux_onehot;
  always_comb
    unique case (go_10_goMux_choice_2_d[4:1])
      4'd0:
        {scfarg_0_1_goMux_mux_onehot, scfarg_0_1_goMux_mux_mux} = {12'd1,
                                                                   lizzieLet20_1_7QNone_Bool_1_argbuf_d};
      4'd1:
        {scfarg_0_1_goMux_mux_onehot, scfarg_0_1_goMux_mux_mux} = {12'd2,
                                                                   sc_0_10_1_argbuf_d};
      4'd2:
        {scfarg_0_1_goMux_mux_onehot, scfarg_0_1_goMux_mux_mux} = {12'd4,
                                                                   lizzieLet20_1_4QVal_Bool_5QNone_Bool_1_argbuf_d};
      4'd3:
        {scfarg_0_1_goMux_mux_onehot, scfarg_0_1_goMux_mux_mux} = {12'd8,
                                                                   lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_2MyFalse_1_argbuf_d};
      4'd4:
        {scfarg_0_1_goMux_mux_onehot, scfarg_0_1_goMux_mux_mux} = {12'd16,
                                                                   lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_2MyTrue_1_argbuf_d};
      4'd5:
        {scfarg_0_1_goMux_mux_onehot, scfarg_0_1_goMux_mux_mux} = {12'd32,
                                                                   lizzieLet20_1_4QVal_Bool_6QVal_Bool_2MyTrue_1_argbuf_d};
      4'd6:
        {scfarg_0_1_goMux_mux_onehot, scfarg_0_1_goMux_mux_mux} = {12'd64,
                                                                   lizzieLet20_1_4QVal_Bool_5QNode_Bool_1_argbuf_d};
      4'd7:
        {scfarg_0_1_goMux_mux_onehot, scfarg_0_1_goMux_mux_mux} = {12'd128,
                                                                   lizzieLet20_1_4QVal_Bool_5QError_Bool_1_argbuf_d};
      4'd8:
        {scfarg_0_1_goMux_mux_onehot, scfarg_0_1_goMux_mux_mux} = {12'd256,
                                                                   lizzieLet20_1_4QNode_Bool_5QNone_Bool_1_argbuf_d};
      4'd9:
        {scfarg_0_1_goMux_mux_onehot, scfarg_0_1_goMux_mux_mux} = {12'd512,
                                                                   lizzieLet20_1_4QNode_Bool_5QVal_Bool_1_argbuf_d};
      4'd10:
        {scfarg_0_1_goMux_mux_onehot,
         scfarg_0_1_goMux_mux_mux} = {12'd1024,
                                      lizzieLet20_1_4QNode_Bool_5QError_Bool_1_argbuf_d};
      4'd11:
        {scfarg_0_1_goMux_mux_onehot,
         scfarg_0_1_goMux_mux_mux} = {12'd2048,
                                      lizzieLet20_1_7QError_Bool_1_argbuf_d};
      default:
        {scfarg_0_1_goMux_mux_onehot, scfarg_0_1_goMux_mux_mux} = {12'd0,
                                                                   {16'd0, 1'd0}};
    endcase
  assign scfarg_0_1_goMux_mux_d = {scfarg_0_1_goMux_mux_mux[16:1],
                                   (scfarg_0_1_goMux_mux_mux[0] && go_10_goMux_choice_2_d[0])};
  assign go_10_goMux_choice_2_r = (scfarg_0_1_goMux_mux_d[0] && scfarg_0_1_goMux_mux_r);
  assign {lizzieLet20_1_7QError_Bool_1_argbuf_r,
          lizzieLet20_1_4QNode_Bool_5QError_Bool_1_argbuf_r,
          lizzieLet20_1_4QNode_Bool_5QVal_Bool_1_argbuf_r,
          lizzieLet20_1_4QNode_Bool_5QNone_Bool_1_argbuf_r,
          lizzieLet20_1_4QVal_Bool_5QError_Bool_1_argbuf_r,
          lizzieLet20_1_4QVal_Bool_5QNode_Bool_1_argbuf_r,
          lizzieLet20_1_4QVal_Bool_6QVal_Bool_2MyTrue_1_argbuf_r,
          lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_2MyTrue_1_argbuf_r,
          lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_2MyFalse_1_argbuf_r,
          lizzieLet20_1_4QVal_Bool_5QNone_Bool_1_argbuf_r,
          sc_0_10_1_argbuf_r,
          lizzieLet20_1_7QNone_Bool_1_argbuf_r} = (go_10_goMux_choice_2_r ? scfarg_0_1_goMux_mux_onehot :
                                                   12'd0);
  
  /* fork (Ty C6) : (go_11_goMux_choice,C6) > [(go_11_goMux_choice_1,C6),
                                          (go_11_goMux_choice_2,C6)] */
  logic [1:0] go_11_goMux_choice_emitted;
  logic [1:0] go_11_goMux_choice_done;
  assign go_11_goMux_choice_1_d = {go_11_goMux_choice_d[3:1],
                                   (go_11_goMux_choice_d[0] && (! go_11_goMux_choice_emitted[0]))};
  assign go_11_goMux_choice_2_d = {go_11_goMux_choice_d[3:1],
                                   (go_11_goMux_choice_d[0] && (! go_11_goMux_choice_emitted[1]))};
  assign go_11_goMux_choice_done = (go_11_goMux_choice_emitted | ({go_11_goMux_choice_2_d[0],
                                                                   go_11_goMux_choice_1_d[0]} & {go_11_goMux_choice_2_r,
                                                                                                 go_11_goMux_choice_1_r}));
  assign go_11_goMux_choice_r = (& go_11_goMux_choice_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_11_goMux_choice_emitted <= 2'd0;
    else
      go_11_goMux_choice_emitted <= (go_11_goMux_choice_r ? 2'd0 :
                                     go_11_goMux_choice_done);
  
  /* mux (Ty C6,
     Ty Pointer_QTree_Bool) : (go_11_goMux_choice_1,C6) [(lizzieLet1_1_1_argbuf,Pointer_QTree_Bool),
                                                         (contRet_0_2_1_argbuf,Pointer_QTree_Bool),
                                                         (lizzieLet32_5MQVal_1_argbuf,Pointer_QTree_Bool),
                                                         (lizzieLet2_1_1_argbuf,Pointer_QTree_Bool),
                                                         (lizzieLet3_1_1_argbuf,Pointer_QTree_Bool),
                                                         (lizzieLet4_1_1_argbuf,Pointer_QTree_Bool)] > (srtarg_0_2_goMux_mux,Pointer_QTree_Bool) */
  logic [16:0] srtarg_0_2_goMux_mux_mux;
  logic [5:0] srtarg_0_2_goMux_mux_onehot;
  always_comb
    unique case (go_11_goMux_choice_1_d[3:1])
      3'd0:
        {srtarg_0_2_goMux_mux_onehot, srtarg_0_2_goMux_mux_mux} = {6'd1,
                                                                   lizzieLet1_1_1_argbuf_d};
      3'd1:
        {srtarg_0_2_goMux_mux_onehot, srtarg_0_2_goMux_mux_mux} = {6'd2,
                                                                   contRet_0_2_1_argbuf_d};
      3'd2:
        {srtarg_0_2_goMux_mux_onehot, srtarg_0_2_goMux_mux_mux} = {6'd4,
                                                                   lizzieLet32_5MQVal_1_argbuf_d};
      3'd3:
        {srtarg_0_2_goMux_mux_onehot, srtarg_0_2_goMux_mux_mux} = {6'd8,
                                                                   lizzieLet2_1_1_argbuf_d};
      3'd4:
        {srtarg_0_2_goMux_mux_onehot, srtarg_0_2_goMux_mux_mux} = {6'd16,
                                                                   lizzieLet3_1_1_argbuf_d};
      3'd5:
        {srtarg_0_2_goMux_mux_onehot, srtarg_0_2_goMux_mux_mux} = {6'd32,
                                                                   lizzieLet4_1_1_argbuf_d};
      default:
        {srtarg_0_2_goMux_mux_onehot, srtarg_0_2_goMux_mux_mux} = {6'd0,
                                                                   {16'd0, 1'd0}};
    endcase
  assign srtarg_0_2_goMux_mux_d = {srtarg_0_2_goMux_mux_mux[16:1],
                                   (srtarg_0_2_goMux_mux_mux[0] && go_11_goMux_choice_1_d[0])};
  assign go_11_goMux_choice_1_r = (srtarg_0_2_goMux_mux_d[0] && srtarg_0_2_goMux_mux_r);
  assign {lizzieLet4_1_1_argbuf_r,
          lizzieLet3_1_1_argbuf_r,
          lizzieLet2_1_1_argbuf_r,
          lizzieLet32_5MQVal_1_argbuf_r,
          contRet_0_2_1_argbuf_r,
          lizzieLet1_1_1_argbuf_r} = (go_11_goMux_choice_1_r ? srtarg_0_2_goMux_mux_onehot :
                                      6'd0);
  
  /* mux (Ty C6,
     Ty Pointer_CTf'''''''''_f'''''''''_Bool) : (go_11_goMux_choice_2,C6) [(lizzieLet32_6MQNone_1_argbuf,Pointer_CTf'''''''''_f'''''''''_Bool),
                                                                           (sc_0_14_1_argbuf,Pointer_CTf'''''''''_f'''''''''_Bool),
                                                                           (lizzieLet32_6MQVal_1_argbuf,Pointer_CTf'''''''''_f'''''''''_Bool),
                                                                           (lizzieLet32_4MQNode_4QNone_Bool_1_argbuf,Pointer_CTf'''''''''_f'''''''''_Bool),
                                                                           (lizzieLet32_4MQNode_4QVal_Bool_1_argbuf,Pointer_CTf'''''''''_f'''''''''_Bool),
                                                                           (lizzieLet32_4MQNode_4QError_Bool_1_argbuf,Pointer_CTf'''''''''_f'''''''''_Bool)] > (scfarg_0_2_goMux_mux,Pointer_CTf'''''''''_f'''''''''_Bool) */
  logic [16:0] scfarg_0_2_goMux_mux_mux;
  logic [5:0] scfarg_0_2_goMux_mux_onehot;
  always_comb
    unique case (go_11_goMux_choice_2_d[3:1])
      3'd0:
        {scfarg_0_2_goMux_mux_onehot, scfarg_0_2_goMux_mux_mux} = {6'd1,
                                                                   lizzieLet32_6MQNone_1_argbuf_d};
      3'd1:
        {scfarg_0_2_goMux_mux_onehot, scfarg_0_2_goMux_mux_mux} = {6'd2,
                                                                   sc_0_14_1_argbuf_d};
      3'd2:
        {scfarg_0_2_goMux_mux_onehot, scfarg_0_2_goMux_mux_mux} = {6'd4,
                                                                   lizzieLet32_6MQVal_1_argbuf_d};
      3'd3:
        {scfarg_0_2_goMux_mux_onehot, scfarg_0_2_goMux_mux_mux} = {6'd8,
                                                                   lizzieLet32_4MQNode_4QNone_Bool_1_argbuf_d};
      3'd4:
        {scfarg_0_2_goMux_mux_onehot, scfarg_0_2_goMux_mux_mux} = {6'd16,
                                                                   lizzieLet32_4MQNode_4QVal_Bool_1_argbuf_d};
      3'd5:
        {scfarg_0_2_goMux_mux_onehot, scfarg_0_2_goMux_mux_mux} = {6'd32,
                                                                   lizzieLet32_4MQNode_4QError_Bool_1_argbuf_d};
      default:
        {scfarg_0_2_goMux_mux_onehot, scfarg_0_2_goMux_mux_mux} = {6'd0,
                                                                   {16'd0, 1'd0}};
    endcase
  assign scfarg_0_2_goMux_mux_d = {scfarg_0_2_goMux_mux_mux[16:1],
                                   (scfarg_0_2_goMux_mux_mux[0] && go_11_goMux_choice_2_d[0])};
  assign go_11_goMux_choice_2_r = (scfarg_0_2_goMux_mux_d[0] && scfarg_0_2_goMux_mux_r);
  assign {lizzieLet32_4MQNode_4QError_Bool_1_argbuf_r,
          lizzieLet32_4MQNode_4QVal_Bool_1_argbuf_r,
          lizzieLet32_4MQNode_4QNone_Bool_1_argbuf_r,
          lizzieLet32_6MQVal_1_argbuf_r,
          sc_0_14_1_argbuf_r,
          lizzieLet32_6MQNone_1_argbuf_r} = (go_11_goMux_choice_2_r ? scfarg_0_2_goMux_mux_onehot :
                                             6'd0);
  
  /* dcon (Ty TupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool,
      Dcon TupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool) : [(go_1_argbuf,Go),
                                                                                   (m1a82_0,Pointer_MaskQTree),
                                                                                   (m2a83_1,Pointer_QTree_Bool),
                                                                                   (m3a84_2,Pointer_QTree_Bool)] > (fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool_1,TupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool) */
  assign fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool_1_d = TupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool_dc((& {go_1_argbuf_d[0],
                                                                                                                                                               m1a82_0_d[0],
                                                                                                                                                               m2a83_1_d[0],
                                                                                                                                                               m3a84_2_d[0]}), go_1_argbuf_d, m1a82_0_d, m2a83_1_d, m3a84_2_d);
  assign {go_1_argbuf_r,
          m1a82_0_r,
          m2a83_1_r,
          m3a84_2_r} = {4 {(fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool_1_r && fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool_1_d[0])}};
  
  /* fork (Ty C5) : (go_2_goMux_choice,C5) > [(go_2_goMux_choice_1,C5),
                                         (go_2_goMux_choice_2,C5),
                                         (go_2_goMux_choice_3,C5),
                                         (go_2_goMux_choice_4,C5)] */
  logic [3:0] go_2_goMux_choice_emitted;
  logic [3:0] go_2_goMux_choice_done;
  assign go_2_goMux_choice_1_d = {go_2_goMux_choice_d[3:1],
                                  (go_2_goMux_choice_d[0] && (! go_2_goMux_choice_emitted[0]))};
  assign go_2_goMux_choice_2_d = {go_2_goMux_choice_d[3:1],
                                  (go_2_goMux_choice_d[0] && (! go_2_goMux_choice_emitted[1]))};
  assign go_2_goMux_choice_3_d = {go_2_goMux_choice_d[3:1],
                                  (go_2_goMux_choice_d[0] && (! go_2_goMux_choice_emitted[2]))};
  assign go_2_goMux_choice_4_d = {go_2_goMux_choice_d[3:1],
                                  (go_2_goMux_choice_d[0] && (! go_2_goMux_choice_emitted[3]))};
  assign go_2_goMux_choice_done = (go_2_goMux_choice_emitted | ({go_2_goMux_choice_4_d[0],
                                                                 go_2_goMux_choice_3_d[0],
                                                                 go_2_goMux_choice_2_d[0],
                                                                 go_2_goMux_choice_1_d[0]} & {go_2_goMux_choice_4_r,
                                                                                              go_2_goMux_choice_3_r,
                                                                                              go_2_goMux_choice_2_r,
                                                                                              go_2_goMux_choice_1_r}));
  assign go_2_goMux_choice_r = (& go_2_goMux_choice_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_2_goMux_choice_emitted <= 4'd0;
    else
      go_2_goMux_choice_emitted <= (go_2_goMux_choice_r ? 4'd0 :
                                    go_2_goMux_choice_done);
  
  /* mux (Ty C5,
     Ty Pointer_MaskQTree) : (go_2_goMux_choice_1,C5) [(call_f_goMux2,Pointer_MaskQTree),
                                                       (q3a8a_1_1_argbuf,Pointer_MaskQTree),
                                                       (q2a89_2_1_argbuf,Pointer_MaskQTree),
                                                       (q1a88_3_1_argbuf,Pointer_MaskQTree),
                                                       (lizzieLet0_4MQNode_4QNode_Bool_8QNode_Bool_1_argbuf,Pointer_MaskQTree)] > (m1a85_goMux_mux,Pointer_MaskQTree) */
  logic [16:0] m1a85_goMux_mux_mux;
  logic [4:0] m1a85_goMux_mux_onehot;
  always_comb
    unique case (go_2_goMux_choice_1_d[3:1])
      3'd0:
        {m1a85_goMux_mux_onehot, m1a85_goMux_mux_mux} = {5'd1,
                                                         call_f_goMux2_d};
      3'd1:
        {m1a85_goMux_mux_onehot, m1a85_goMux_mux_mux} = {5'd2,
                                                         q3a8a_1_1_argbuf_d};
      3'd2:
        {m1a85_goMux_mux_onehot, m1a85_goMux_mux_mux} = {5'd4,
                                                         q2a89_2_1_argbuf_d};
      3'd3:
        {m1a85_goMux_mux_onehot, m1a85_goMux_mux_mux} = {5'd8,
                                                         q1a88_3_1_argbuf_d};
      3'd4:
        {m1a85_goMux_mux_onehot, m1a85_goMux_mux_mux} = {5'd16,
                                                         lizzieLet0_4MQNode_4QNode_Bool_8QNode_Bool_1_argbuf_d};
      default:
        {m1a85_goMux_mux_onehot, m1a85_goMux_mux_mux} = {5'd0,
                                                         {16'd0, 1'd0}};
    endcase
  assign m1a85_goMux_mux_d = {m1a85_goMux_mux_mux[16:1],
                              (m1a85_goMux_mux_mux[0] && go_2_goMux_choice_1_d[0])};
  assign go_2_goMux_choice_1_r = (m1a85_goMux_mux_d[0] && m1a85_goMux_mux_r);
  assign {lizzieLet0_4MQNode_4QNode_Bool_8QNode_Bool_1_argbuf_r,
          q1a88_3_1_argbuf_r,
          q2a89_2_1_argbuf_r,
          q3a8a_1_1_argbuf_r,
          call_f_goMux2_r} = (go_2_goMux_choice_1_r ? m1a85_goMux_mux_onehot :
                              5'd0);
  
  /* mux (Ty C5,
     Ty Pointer_QTree_Bool) : (go_2_goMux_choice_2,C5) [(call_f_goMux3,Pointer_QTree_Bool),
                                                        (q3'a8p_1_1_argbuf,Pointer_QTree_Bool),
                                                        (q2'a8o_2_1_argbuf,Pointer_QTree_Bool),
                                                        (q1'a8n_3_1_argbuf,Pointer_QTree_Bool),
                                                        (lizzieLet0_4MQNode_4QNode_Bool_12QNode_Bool_1_argbuf,Pointer_QTree_Bool)] > (m2a86_goMux_mux,Pointer_QTree_Bool) */
  logic [16:0] m2a86_goMux_mux_mux;
  logic [4:0] m2a86_goMux_mux_onehot;
  always_comb
    unique case (go_2_goMux_choice_2_d[3:1])
      3'd0:
        {m2a86_goMux_mux_onehot, m2a86_goMux_mux_mux} = {5'd1,
                                                         call_f_goMux3_d};
      3'd1:
        {m2a86_goMux_mux_onehot, m2a86_goMux_mux_mux} = {5'd2,
                                                         \q3'a8p_1_1_argbuf_d };
      3'd2:
        {m2a86_goMux_mux_onehot, m2a86_goMux_mux_mux} = {5'd4,
                                                         \q2'a8o_2_1_argbuf_d };
      3'd3:
        {m2a86_goMux_mux_onehot, m2a86_goMux_mux_mux} = {5'd8,
                                                         \q1'a8n_3_1_argbuf_d };
      3'd4:
        {m2a86_goMux_mux_onehot, m2a86_goMux_mux_mux} = {5'd16,
                                                         lizzieLet0_4MQNode_4QNode_Bool_12QNode_Bool_1_argbuf_d};
      default:
        {m2a86_goMux_mux_onehot, m2a86_goMux_mux_mux} = {5'd0,
                                                         {16'd0, 1'd0}};
    endcase
  assign m2a86_goMux_mux_d = {m2a86_goMux_mux_mux[16:1],
                              (m2a86_goMux_mux_mux[0] && go_2_goMux_choice_2_d[0])};
  assign go_2_goMux_choice_2_r = (m2a86_goMux_mux_d[0] && m2a86_goMux_mux_r);
  assign {lizzieLet0_4MQNode_4QNode_Bool_12QNode_Bool_1_argbuf_r,
          \q1'a8n_3_1_argbuf_r ,
          \q2'a8o_2_1_argbuf_r ,
          \q3'a8p_1_1_argbuf_r ,
          call_f_goMux3_r} = (go_2_goMux_choice_2_r ? m2a86_goMux_mux_onehot :
                              5'd0);
  
  /* mux (Ty C5,
     Ty Pointer_QTree_Bool) : (go_2_goMux_choice_3,C5) [(call_f_goMux4,Pointer_QTree_Bool),
                                                        (t3a8u_1_1_argbuf,Pointer_QTree_Bool),
                                                        (t2a8t_2_1_argbuf,Pointer_QTree_Bool),
                                                        (t1a8s_3_1_argbuf,Pointer_QTree_Bool),
                                                        (t4a8v_1_argbuf,Pointer_QTree_Bool)] > (m3a87_goMux_mux,Pointer_QTree_Bool) */
  logic [16:0] m3a87_goMux_mux_mux;
  logic [4:0] m3a87_goMux_mux_onehot;
  always_comb
    unique case (go_2_goMux_choice_3_d[3:1])
      3'd0:
        {m3a87_goMux_mux_onehot, m3a87_goMux_mux_mux} = {5'd1,
                                                         call_f_goMux4_d};
      3'd1:
        {m3a87_goMux_mux_onehot, m3a87_goMux_mux_mux} = {5'd2,
                                                         t3a8u_1_1_argbuf_d};
      3'd2:
        {m3a87_goMux_mux_onehot, m3a87_goMux_mux_mux} = {5'd4,
                                                         t2a8t_2_1_argbuf_d};
      3'd3:
        {m3a87_goMux_mux_onehot, m3a87_goMux_mux_mux} = {5'd8,
                                                         t1a8s_3_1_argbuf_d};
      3'd4:
        {m3a87_goMux_mux_onehot, m3a87_goMux_mux_mux} = {5'd16,
                                                         t4a8v_1_argbuf_d};
      default:
        {m3a87_goMux_mux_onehot, m3a87_goMux_mux_mux} = {5'd0,
                                                         {16'd0, 1'd0}};
    endcase
  assign m3a87_goMux_mux_d = {m3a87_goMux_mux_mux[16:1],
                              (m3a87_goMux_mux_mux[0] && go_2_goMux_choice_3_d[0])};
  assign go_2_goMux_choice_3_r = (m3a87_goMux_mux_d[0] && m3a87_goMux_mux_r);
  assign {t4a8v_1_argbuf_r,
          t1a8s_3_1_argbuf_r,
          t2a8t_2_1_argbuf_r,
          t3a8u_1_1_argbuf_r,
          call_f_goMux4_r} = (go_2_goMux_choice_3_r ? m3a87_goMux_mux_onehot :
                              5'd0);
  
  /* mux (Ty C5,
     Ty Pointer_CTf) : (go_2_goMux_choice_4,C5) [(call_f_goMux5,Pointer_CTf),
                                                 (sca2_1_argbuf,Pointer_CTf),
                                                 (sca1_1_argbuf,Pointer_CTf),
                                                 (sca0_1_argbuf,Pointer_CTf),
                                                 (sca3_1_argbuf,Pointer_CTf)] > (sc_0_goMux_mux,Pointer_CTf) */
  logic [16:0] sc_0_goMux_mux_mux;
  logic [4:0] sc_0_goMux_mux_onehot;
  always_comb
    unique case (go_2_goMux_choice_4_d[3:1])
      3'd0:
        {sc_0_goMux_mux_onehot, sc_0_goMux_mux_mux} = {5'd1,
                                                       call_f_goMux5_d};
      3'd1:
        {sc_0_goMux_mux_onehot, sc_0_goMux_mux_mux} = {5'd2,
                                                       sca2_1_argbuf_d};
      3'd2:
        {sc_0_goMux_mux_onehot, sc_0_goMux_mux_mux} = {5'd4,
                                                       sca1_1_argbuf_d};
      3'd3:
        {sc_0_goMux_mux_onehot, sc_0_goMux_mux_mux} = {5'd8,
                                                       sca0_1_argbuf_d};
      3'd4:
        {sc_0_goMux_mux_onehot, sc_0_goMux_mux_mux} = {5'd16,
                                                       sca3_1_argbuf_d};
      default:
        {sc_0_goMux_mux_onehot, sc_0_goMux_mux_mux} = {5'd0,
                                                       {16'd0, 1'd0}};
    endcase
  assign sc_0_goMux_mux_d = {sc_0_goMux_mux_mux[16:1],
                             (sc_0_goMux_mux_mux[0] && go_2_goMux_choice_4_d[0])};
  assign go_2_goMux_choice_4_r = (sc_0_goMux_mux_d[0] && sc_0_goMux_mux_r);
  assign {sca3_1_argbuf_r,
          sca0_1_argbuf_r,
          sca1_1_argbuf_r,
          sca2_1_argbuf_r,
          call_f_goMux5_r} = (go_2_goMux_choice_4_r ? sc_0_goMux_mux_onehot :
                              5'd0);
  
  /* fork (Ty C5) : (go_3_goMux_choice,C5) > [(go_3_goMux_choice_1,C5),
                                         (go_3_goMux_choice_2,C5),
                                         (go_3_goMux_choice_3,C5)] */
  logic [2:0] go_3_goMux_choice_emitted;
  logic [2:0] go_3_goMux_choice_done;
  assign go_3_goMux_choice_1_d = {go_3_goMux_choice_d[3:1],
                                  (go_3_goMux_choice_d[0] && (! go_3_goMux_choice_emitted[0]))};
  assign go_3_goMux_choice_2_d = {go_3_goMux_choice_d[3:1],
                                  (go_3_goMux_choice_d[0] && (! go_3_goMux_choice_emitted[1]))};
  assign go_3_goMux_choice_3_d = {go_3_goMux_choice_d[3:1],
                                  (go_3_goMux_choice_d[0] && (! go_3_goMux_choice_emitted[2]))};
  assign go_3_goMux_choice_done = (go_3_goMux_choice_emitted | ({go_3_goMux_choice_3_d[0],
                                                                 go_3_goMux_choice_2_d[0],
                                                                 go_3_goMux_choice_1_d[0]} & {go_3_goMux_choice_3_r,
                                                                                              go_3_goMux_choice_2_r,
                                                                                              go_3_goMux_choice_1_r}));
  assign go_3_goMux_choice_r = (& go_3_goMux_choice_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_3_goMux_choice_emitted <= 3'd0;
    else
      go_3_goMux_choice_emitted <= (go_3_goMux_choice_r ? 3'd0 :
                                    go_3_goMux_choice_done);
  
  /* mux (Ty C5,
     Ty Pointer_QTree_Bool) : (go_3_goMux_choice_1,C5) [(call_f'_goMux2,Pointer_QTree_Bool),
                                                        (q3a8R_1_1_argbuf,Pointer_QTree_Bool),
                                                        (q2a8Q_2_1_argbuf,Pointer_QTree_Bool),
                                                        (q1a8P_3_1_argbuf,Pointer_QTree_Bool),
                                                        (lizzieLet20_1_4QNode_Bool_9QNode_Bool_1_argbuf,Pointer_QTree_Bool)] > (m2a8H_goMux_mux,Pointer_QTree_Bool) */
  logic [16:0] m2a8H_goMux_mux_mux;
  logic [4:0] m2a8H_goMux_mux_onehot;
  always_comb
    unique case (go_3_goMux_choice_1_d[3:1])
      3'd0:
        {m2a8H_goMux_mux_onehot, m2a8H_goMux_mux_mux} = {5'd1,
                                                         \call_f'_goMux2_d };
      3'd1:
        {m2a8H_goMux_mux_onehot, m2a8H_goMux_mux_mux} = {5'd2,
                                                         q3a8R_1_1_argbuf_d};
      3'd2:
        {m2a8H_goMux_mux_onehot, m2a8H_goMux_mux_mux} = {5'd4,
                                                         q2a8Q_2_1_argbuf_d};
      3'd3:
        {m2a8H_goMux_mux_onehot, m2a8H_goMux_mux_mux} = {5'd8,
                                                         q1a8P_3_1_argbuf_d};
      3'd4:
        {m2a8H_goMux_mux_onehot, m2a8H_goMux_mux_mux} = {5'd16,
                                                         lizzieLet20_1_4QNode_Bool_9QNode_Bool_1_argbuf_d};
      default:
        {m2a8H_goMux_mux_onehot, m2a8H_goMux_mux_mux} = {5'd0,
                                                         {16'd0, 1'd0}};
    endcase
  assign m2a8H_goMux_mux_d = {m2a8H_goMux_mux_mux[16:1],
                              (m2a8H_goMux_mux_mux[0] && go_3_goMux_choice_1_d[0])};
  assign go_3_goMux_choice_1_r = (m2a8H_goMux_mux_d[0] && m2a8H_goMux_mux_r);
  assign {lizzieLet20_1_4QNode_Bool_9QNode_Bool_1_argbuf_r,
          q1a8P_3_1_argbuf_r,
          q2a8Q_2_1_argbuf_r,
          q3a8R_1_1_argbuf_r,
          \call_f'_goMux2_r } = (go_3_goMux_choice_1_r ? m2a8H_goMux_mux_onehot :
                                 5'd0);
  
  /* mux (Ty C5,
     Ty Pointer_QTree_Bool) : (go_3_goMux_choice_2,C5) [(call_f'_goMux3,Pointer_QTree_Bool),
                                                        (t3a8W_1_1_argbuf,Pointer_QTree_Bool),
                                                        (t2a8V_2_1_argbuf,Pointer_QTree_Bool),
                                                        (t1a8U_3_1_argbuf,Pointer_QTree_Bool),
                                                        (t4a8X_1_argbuf,Pointer_QTree_Bool)] > (m3a8I_goMux_mux,Pointer_QTree_Bool) */
  logic [16:0] m3a8I_goMux_mux_mux;
  logic [4:0] m3a8I_goMux_mux_onehot;
  always_comb
    unique case (go_3_goMux_choice_2_d[3:1])
      3'd0:
        {m3a8I_goMux_mux_onehot, m3a8I_goMux_mux_mux} = {5'd1,
                                                         \call_f'_goMux3_d };
      3'd1:
        {m3a8I_goMux_mux_onehot, m3a8I_goMux_mux_mux} = {5'd2,
                                                         t3a8W_1_1_argbuf_d};
      3'd2:
        {m3a8I_goMux_mux_onehot, m3a8I_goMux_mux_mux} = {5'd4,
                                                         t2a8V_2_1_argbuf_d};
      3'd3:
        {m3a8I_goMux_mux_onehot, m3a8I_goMux_mux_mux} = {5'd8,
                                                         t1a8U_3_1_argbuf_d};
      3'd4:
        {m3a8I_goMux_mux_onehot, m3a8I_goMux_mux_mux} = {5'd16,
                                                         t4a8X_1_argbuf_d};
      default:
        {m3a8I_goMux_mux_onehot, m3a8I_goMux_mux_mux} = {5'd0,
                                                         {16'd0, 1'd0}};
    endcase
  assign m3a8I_goMux_mux_d = {m3a8I_goMux_mux_mux[16:1],
                              (m3a8I_goMux_mux_mux[0] && go_3_goMux_choice_2_d[0])};
  assign go_3_goMux_choice_2_r = (m3a8I_goMux_mux_d[0] && m3a8I_goMux_mux_r);
  assign {t4a8X_1_argbuf_r,
          t1a8U_3_1_argbuf_r,
          t2a8V_2_1_argbuf_r,
          t3a8W_1_1_argbuf_r,
          \call_f'_goMux3_r } = (go_3_goMux_choice_2_r ? m3a8I_goMux_mux_onehot :
                                 5'd0);
  
  /* mux (Ty C5,
     Ty Pointer_CTf') : (go_3_goMux_choice_3,C5) [(call_f'_goMux4,Pointer_CTf'),
                                                  (sca2_1_1_argbuf,Pointer_CTf'),
                                                  (sca1_1_1_argbuf,Pointer_CTf'),
                                                  (sca0_1_1_argbuf,Pointer_CTf'),
                                                  (sca3_1_1_argbuf,Pointer_CTf')] > (sc_0_1_goMux_mux,Pointer_CTf') */
  logic [16:0] sc_0_1_goMux_mux_mux;
  logic [4:0] sc_0_1_goMux_mux_onehot;
  always_comb
    unique case (go_3_goMux_choice_3_d[3:1])
      3'd0:
        {sc_0_1_goMux_mux_onehot, sc_0_1_goMux_mux_mux} = {5'd1,
                                                           \call_f'_goMux4_d };
      3'd1:
        {sc_0_1_goMux_mux_onehot, sc_0_1_goMux_mux_mux} = {5'd2,
                                                           sca2_1_1_argbuf_d};
      3'd2:
        {sc_0_1_goMux_mux_onehot, sc_0_1_goMux_mux_mux} = {5'd4,
                                                           sca1_1_1_argbuf_d};
      3'd3:
        {sc_0_1_goMux_mux_onehot, sc_0_1_goMux_mux_mux} = {5'd8,
                                                           sca0_1_1_argbuf_d};
      3'd4:
        {sc_0_1_goMux_mux_onehot, sc_0_1_goMux_mux_mux} = {5'd16,
                                                           sca3_1_1_argbuf_d};
      default:
        {sc_0_1_goMux_mux_onehot, sc_0_1_goMux_mux_mux} = {5'd0,
                                                           {16'd0, 1'd0}};
    endcase
  assign sc_0_1_goMux_mux_d = {sc_0_1_goMux_mux_mux[16:1],
                               (sc_0_1_goMux_mux_mux[0] && go_3_goMux_choice_3_d[0])};
  assign go_3_goMux_choice_3_r = (sc_0_1_goMux_mux_d[0] && sc_0_1_goMux_mux_r);
  assign {sca3_1_1_argbuf_r,
          sca0_1_1_argbuf_r,
          sca1_1_1_argbuf_r,
          sca2_1_1_argbuf_r,
          \call_f'_goMux4_r } = (go_3_goMux_choice_3_r ? sc_0_1_goMux_mux_onehot :
                                 5'd0);
  
  /* fork (Ty C5) : (go_4_goMux_choice,C5) > [(go_4_goMux_choice_1,C5),
                                         (go_4_goMux_choice_2,C5),
                                         (go_4_goMux_choice_3,C5)] */
  logic [2:0] go_4_goMux_choice_emitted;
  logic [2:0] go_4_goMux_choice_done;
  assign go_4_goMux_choice_1_d = {go_4_goMux_choice_d[3:1],
                                  (go_4_goMux_choice_d[0] && (! go_4_goMux_choice_emitted[0]))};
  assign go_4_goMux_choice_2_d = {go_4_goMux_choice_d[3:1],
                                  (go_4_goMux_choice_d[0] && (! go_4_goMux_choice_emitted[1]))};
  assign go_4_goMux_choice_3_d = {go_4_goMux_choice_d[3:1],
                                  (go_4_goMux_choice_d[0] && (! go_4_goMux_choice_emitted[2]))};
  assign go_4_goMux_choice_done = (go_4_goMux_choice_emitted | ({go_4_goMux_choice_3_d[0],
                                                                 go_4_goMux_choice_2_d[0],
                                                                 go_4_goMux_choice_1_d[0]} & {go_4_goMux_choice_3_r,
                                                                                              go_4_goMux_choice_2_r,
                                                                                              go_4_goMux_choice_1_r}));
  assign go_4_goMux_choice_r = (& go_4_goMux_choice_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_4_goMux_choice_emitted <= 3'd0;
    else
      go_4_goMux_choice_emitted <= (go_4_goMux_choice_r ? 3'd0 :
                                    go_4_goMux_choice_done);
  
  /* mux (Ty C5,
     Ty Pointer_MaskQTree) : (go_4_goMux_choice_1,C5) [(call_f'''''''''_f'''''''''_Bool_goMux2,Pointer_MaskQTree),
                                                       (q3a8A_1_1_argbuf,Pointer_MaskQTree),
                                                       (q2a8z_2_1_argbuf,Pointer_MaskQTree),
                                                       (q1a8y_3_1_argbuf,Pointer_MaskQTree),
                                                       (lizzieLet32_4MQNode_8QNode_Bool_1_argbuf,Pointer_MaskQTree)] > (q4a8w_goMux_mux,Pointer_MaskQTree) */
  logic [16:0] q4a8w_goMux_mux_mux;
  logic [4:0] q4a8w_goMux_mux_onehot;
  always_comb
    unique case (go_4_goMux_choice_1_d[3:1])
      3'd0:
        {q4a8w_goMux_mux_onehot, q4a8w_goMux_mux_mux} = {5'd1,
                                                         \call_f'''''''''_f'''''''''_Bool_goMux2_d };
      3'd1:
        {q4a8w_goMux_mux_onehot, q4a8w_goMux_mux_mux} = {5'd2,
                                                         q3a8A_1_1_argbuf_d};
      3'd2:
        {q4a8w_goMux_mux_onehot, q4a8w_goMux_mux_mux} = {5'd4,
                                                         q2a8z_2_1_argbuf_d};
      3'd3:
        {q4a8w_goMux_mux_onehot, q4a8w_goMux_mux_mux} = {5'd8,
                                                         q1a8y_3_1_argbuf_d};
      3'd4:
        {q4a8w_goMux_mux_onehot, q4a8w_goMux_mux_mux} = {5'd16,
                                                         lizzieLet32_4MQNode_8QNode_Bool_1_argbuf_d};
      default:
        {q4a8w_goMux_mux_onehot, q4a8w_goMux_mux_mux} = {5'd0,
                                                         {16'd0, 1'd0}};
    endcase
  assign q4a8w_goMux_mux_d = {q4a8w_goMux_mux_mux[16:1],
                              (q4a8w_goMux_mux_mux[0] && go_4_goMux_choice_1_d[0])};
  assign go_4_goMux_choice_1_r = (q4a8w_goMux_mux_d[0] && q4a8w_goMux_mux_r);
  assign {lizzieLet32_4MQNode_8QNode_Bool_1_argbuf_r,
          q1a8y_3_1_argbuf_r,
          q2a8z_2_1_argbuf_r,
          q3a8A_1_1_argbuf_r,
          \call_f'''''''''_f'''''''''_Bool_goMux2_r } = (go_4_goMux_choice_1_r ? q4a8w_goMux_mux_onehot :
                                                         5'd0);
  
  /* mux (Ty C5,
     Ty Pointer_QTree_Bool) : (go_4_goMux_choice_2,C5) [(call_f'''''''''_f'''''''''_Bool_goMux3,Pointer_QTree_Bool),
                                                        (t3a8F_1_1_argbuf,Pointer_QTree_Bool),
                                                        (t2a8E_2_1_argbuf,Pointer_QTree_Bool),
                                                        (t1a8D_3_1_argbuf,Pointer_QTree_Bool),
                                                        (t4a8G_1_argbuf,Pointer_QTree_Bool)] > (q4'a8x_goMux_mux,Pointer_QTree_Bool) */
  logic [16:0] \q4'a8x_goMux_mux_mux ;
  logic [4:0] \q4'a8x_goMux_mux_onehot ;
  always_comb
    unique case (go_4_goMux_choice_2_d[3:1])
      3'd0:
        {\q4'a8x_goMux_mux_onehot , \q4'a8x_goMux_mux_mux } = {5'd1,
                                                               \call_f'''''''''_f'''''''''_Bool_goMux3_d };
      3'd1:
        {\q4'a8x_goMux_mux_onehot , \q4'a8x_goMux_mux_mux } = {5'd2,
                                                               t3a8F_1_1_argbuf_d};
      3'd2:
        {\q4'a8x_goMux_mux_onehot , \q4'a8x_goMux_mux_mux } = {5'd4,
                                                               t2a8E_2_1_argbuf_d};
      3'd3:
        {\q4'a8x_goMux_mux_onehot , \q4'a8x_goMux_mux_mux } = {5'd8,
                                                               t1a8D_3_1_argbuf_d};
      3'd4:
        {\q4'a8x_goMux_mux_onehot , \q4'a8x_goMux_mux_mux } = {5'd16,
                                                               t4a8G_1_argbuf_d};
      default:
        {\q4'a8x_goMux_mux_onehot , \q4'a8x_goMux_mux_mux } = {5'd0,
                                                               {16'd0, 1'd0}};
    endcase
  assign \q4'a8x_goMux_mux_d  = {\q4'a8x_goMux_mux_mux [16:1],
                                 (\q4'a8x_goMux_mux_mux [0] && go_4_goMux_choice_2_d[0])};
  assign go_4_goMux_choice_2_r = (\q4'a8x_goMux_mux_d [0] && \q4'a8x_goMux_mux_r );
  assign {t4a8G_1_argbuf_r,
          t1a8D_3_1_argbuf_r,
          t2a8E_2_1_argbuf_r,
          t3a8F_1_1_argbuf_r,
          \call_f'''''''''_f'''''''''_Bool_goMux3_r } = (go_4_goMux_choice_2_r ? \q4'a8x_goMux_mux_onehot  :
                                                         5'd0);
  
  /* mux (Ty C5,
     Ty Pointer_CTf'''''''''_f'''''''''_Bool) : (go_4_goMux_choice_3,C5) [(call_f'''''''''_f'''''''''_Bool_goMux4,Pointer_CTf'''''''''_f'''''''''_Bool),
                                                                          (sca2_2_1_argbuf,Pointer_CTf'''''''''_f'''''''''_Bool),
                                                                          (sca1_2_1_argbuf,Pointer_CTf'''''''''_f'''''''''_Bool),
                                                                          (sca0_2_1_argbuf,Pointer_CTf'''''''''_f'''''''''_Bool),
                                                                          (sca3_2_1_argbuf,Pointer_CTf'''''''''_f'''''''''_Bool)] > (sc_0_2_goMux_mux,Pointer_CTf'''''''''_f'''''''''_Bool) */
  logic [16:0] sc_0_2_goMux_mux_mux;
  logic [4:0] sc_0_2_goMux_mux_onehot;
  always_comb
    unique case (go_4_goMux_choice_3_d[3:1])
      3'd0:
        {sc_0_2_goMux_mux_onehot, sc_0_2_goMux_mux_mux} = {5'd1,
                                                           \call_f'''''''''_f'''''''''_Bool_goMux4_d };
      3'd1:
        {sc_0_2_goMux_mux_onehot, sc_0_2_goMux_mux_mux} = {5'd2,
                                                           sca2_2_1_argbuf_d};
      3'd2:
        {sc_0_2_goMux_mux_onehot, sc_0_2_goMux_mux_mux} = {5'd4,
                                                           sca1_2_1_argbuf_d};
      3'd3:
        {sc_0_2_goMux_mux_onehot, sc_0_2_goMux_mux_mux} = {5'd8,
                                                           sca0_2_1_argbuf_d};
      3'd4:
        {sc_0_2_goMux_mux_onehot, sc_0_2_goMux_mux_mux} = {5'd16,
                                                           sca3_2_1_argbuf_d};
      default:
        {sc_0_2_goMux_mux_onehot, sc_0_2_goMux_mux_mux} = {5'd0,
                                                           {16'd0, 1'd0}};
    endcase
  assign sc_0_2_goMux_mux_d = {sc_0_2_goMux_mux_mux[16:1],
                               (sc_0_2_goMux_mux_mux[0] && go_4_goMux_choice_3_d[0])};
  assign go_4_goMux_choice_3_r = (sc_0_2_goMux_mux_d[0] && sc_0_2_goMux_mux_r);
  assign {sca3_2_1_argbuf_r,
          sca0_2_1_argbuf_r,
          sca1_2_1_argbuf_r,
          sca2_2_1_argbuf_r,
          \call_f'''''''''_f'''''''''_Bool_goMux4_r } = (go_4_goMux_choice_3_r ? sc_0_2_goMux_mux_onehot :
                                                         5'd0);
  
  /* dcon (Ty CTf,Dcon Lfsbos) : [(go_5_1,Go)] > (go_5_1Lfsbos,CTf) */
  assign go_5_1Lfsbos_d = Lfsbos_dc((& {go_5_1_d[0]}), go_5_1_d);
  assign {go_5_1_r} = {1 {(go_5_1Lfsbos_r && go_5_1Lfsbos_d[0])}};
  
  /* buf (Ty CTf) : (go_5_1Lfsbos,CTf) > (lizzieLet39_1_argbuf,CTf) */
  CTf_t go_5_1Lfsbos_bufchan_d;
  logic go_5_1Lfsbos_bufchan_r;
  assign go_5_1Lfsbos_r = ((! go_5_1Lfsbos_bufchan_d[0]) || go_5_1Lfsbos_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_5_1Lfsbos_bufchan_d <= {163'd0, 1'd0};
    else if (go_5_1Lfsbos_r) go_5_1Lfsbos_bufchan_d <= go_5_1Lfsbos_d;
  CTf_t go_5_1Lfsbos_bufchan_buf;
  assign go_5_1Lfsbos_bufchan_r = (! go_5_1Lfsbos_bufchan_buf[0]);
  assign lizzieLet39_1_argbuf_d = (go_5_1Lfsbos_bufchan_buf[0] ? go_5_1Lfsbos_bufchan_buf :
                                   go_5_1Lfsbos_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_5_1Lfsbos_bufchan_buf <= {163'd0, 1'd0};
    else
      if ((lizzieLet39_1_argbuf_r && go_5_1Lfsbos_bufchan_buf[0]))
        go_5_1Lfsbos_bufchan_buf <= {163'd0, 1'd0};
      else if (((! lizzieLet39_1_argbuf_r) && (! go_5_1Lfsbos_bufchan_buf[0])))
        go_5_1Lfsbos_bufchan_buf <= go_5_1Lfsbos_bufchan_d;
  
  /* buf (Ty Go) : (go_5_2,Go) > (go_5_2_argbuf,Go) */
  Go_t go_5_2_bufchan_d;
  logic go_5_2_bufchan_r;
  assign go_5_2_r = ((! go_5_2_bufchan_d[0]) || go_5_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_5_2_bufchan_d <= 1'd0;
    else if (go_5_2_r) go_5_2_bufchan_d <= go_5_2_d;
  Go_t go_5_2_bufchan_buf;
  assign go_5_2_bufchan_r = (! go_5_2_bufchan_buf[0]);
  assign go_5_2_argbuf_d = (go_5_2_bufchan_buf[0] ? go_5_2_bufchan_buf :
                            go_5_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_5_2_bufchan_buf <= 1'd0;
    else
      if ((go_5_2_argbuf_r && go_5_2_bufchan_buf[0]))
        go_5_2_bufchan_buf <= 1'd0;
      else if (((! go_5_2_argbuf_r) && (! go_5_2_bufchan_buf[0])))
        go_5_2_bufchan_buf <= go_5_2_bufchan_d;
  
  /* dcon (Ty TupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf,
      Dcon TupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf) : [(go_5_2_argbuf,Go),
                                                                                                 (m1a85_1_1_argbuf,Pointer_MaskQTree),
                                                                                                 (m2a86_1_1_argbuf,Pointer_QTree_Bool),
                                                                                                 (m3a87_1_1_argbuf,Pointer_QTree_Bool),
                                                                                                 (lizzieLet28_1_1_argbuf,Pointer_CTf)] > (call_fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf_1,TupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf) */
  assign call_fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf_1_d = TupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf_dc((& {go_5_2_argbuf_d[0],
                                                                                                                                                                                                m1a85_1_1_argbuf_d[0],
                                                                                                                                                                                                m2a86_1_1_argbuf_d[0],
                                                                                                                                                                                                m3a87_1_1_argbuf_d[0],
                                                                                                                                                                                                lizzieLet28_1_1_argbuf_d[0]}), go_5_2_argbuf_d, m1a85_1_1_argbuf_d, m2a86_1_1_argbuf_d, m3a87_1_1_argbuf_d, lizzieLet28_1_1_argbuf_d);
  assign {go_5_2_argbuf_r,
          m1a85_1_1_argbuf_r,
          m2a86_1_1_argbuf_r,
          m3a87_1_1_argbuf_r,
          lizzieLet28_1_1_argbuf_r} = {5 {(call_fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf_1_r && call_fTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf_1_d[0])}};
  
  /* dcon (Ty CTf',Dcon Lf'sbos) : [(go_6_1,Go)] > (go_6_1Lf'sbos,CTf') */
  assign \go_6_1Lf'sbos_d  = \Lf'sbos_dc ((& {go_6_1_d[0]}), go_6_1_d);
  assign {go_6_1_r} = {1 {(\go_6_1Lf'sbos_r  && \go_6_1Lf'sbos_d [0])}};
  
  /* buf (Ty CTf') : (go_6_1Lf'sbos,CTf') > (lizzieLet40_1_argbuf,CTf') */
  \CTf'_t  \go_6_1Lf'sbos_bufchan_d ;
  logic \go_6_1Lf'sbos_bufchan_r ;
  assign \go_6_1Lf'sbos_r  = ((! \go_6_1Lf'sbos_bufchan_d [0]) || \go_6_1Lf'sbos_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \go_6_1Lf'sbos_bufchan_d  <= {115'd0, 1'd0};
    else
      if (\go_6_1Lf'sbos_r )
        \go_6_1Lf'sbos_bufchan_d  <= \go_6_1Lf'sbos_d ;
  \CTf'_t  \go_6_1Lf'sbos_bufchan_buf ;
  assign \go_6_1Lf'sbos_bufchan_r  = (! \go_6_1Lf'sbos_bufchan_buf [0]);
  assign lizzieLet40_1_argbuf_d = (\go_6_1Lf'sbos_bufchan_buf [0] ? \go_6_1Lf'sbos_bufchan_buf  :
                                   \go_6_1Lf'sbos_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \go_6_1Lf'sbos_bufchan_buf  <= {115'd0, 1'd0};
    else
      if ((lizzieLet40_1_argbuf_r && \go_6_1Lf'sbos_bufchan_buf [0]))
        \go_6_1Lf'sbos_bufchan_buf  <= {115'd0, 1'd0};
      else if (((! lizzieLet40_1_argbuf_r) && (! \go_6_1Lf'sbos_bufchan_buf [0])))
        \go_6_1Lf'sbos_bufchan_buf  <= \go_6_1Lf'sbos_bufchan_d ;
  
  /* buf (Ty Go) : (go_6_2,Go) > (go_6_2_argbuf,Go) */
  Go_t go_6_2_bufchan_d;
  logic go_6_2_bufchan_r;
  assign go_6_2_r = ((! go_6_2_bufchan_d[0]) || go_6_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_6_2_bufchan_d <= 1'd0;
    else if (go_6_2_r) go_6_2_bufchan_d <= go_6_2_d;
  Go_t go_6_2_bufchan_buf;
  assign go_6_2_bufchan_r = (! go_6_2_bufchan_buf[0]);
  assign go_6_2_argbuf_d = (go_6_2_bufchan_buf[0] ? go_6_2_bufchan_buf :
                            go_6_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_6_2_bufchan_buf <= 1'd0;
    else
      if ((go_6_2_argbuf_r && go_6_2_bufchan_buf[0]))
        go_6_2_bufchan_buf <= 1'd0;
      else if (((! go_6_2_argbuf_r) && (! go_6_2_bufchan_buf[0])))
        go_6_2_bufchan_buf <= go_6_2_bufchan_d;
  
  /* dcon (Ty TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf',
      Dcon TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf') : [(go_6_2_argbuf,Go),
                                                                              (m2a8H_1_1_argbuf,Pointer_QTree_Bool),
                                                                              (m3a8I_1_1_argbuf,Pointer_QTree_Bool),
                                                                              (lizzieLet12_1_1_argbuf,Pointer_CTf')] > (call_f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf'_1,TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf') */
  assign \call_f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf'_1_d  = \TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf'_dc ((& {go_6_2_argbuf_d[0],
                                                                                                                                                               m2a8H_1_1_argbuf_d[0],
                                                                                                                                                               m3a8I_1_1_argbuf_d[0],
                                                                                                                                                               lizzieLet12_1_1_argbuf_d[0]}), go_6_2_argbuf_d, m2a8H_1_1_argbuf_d, m3a8I_1_1_argbuf_d, lizzieLet12_1_1_argbuf_d);
  assign {go_6_2_argbuf_r,
          m2a8H_1_1_argbuf_r,
          m3a8I_1_1_argbuf_r,
          lizzieLet12_1_1_argbuf_r} = {4 {(\call_f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf'_1_r  && \call_f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf'_1_d [0])}};
  
  /* dcon (Ty CTf'''''''''_f'''''''''_Bool,
      Dcon Lf'''''''''_f'''''''''_Boolsbos) : [(go_7_1,Go)] > (go_7_1Lf'''''''''_f'''''''''_Boolsbos,CTf'''''''''_f'''''''''_Bool) */
  assign \go_7_1Lf'''''''''_f'''''''''_Boolsbos_d  = \Lf'''''''''_f'''''''''_Boolsbos_dc ((& {go_7_1_d[0]}), go_7_1_d);
  assign {go_7_1_r} = {1 {(\go_7_1Lf'''''''''_f'''''''''_Boolsbos_r  && \go_7_1Lf'''''''''_f'''''''''_Boolsbos_d [0])}};
  
  /* buf (Ty CTf'''''''''_f'''''''''_Bool) : (go_7_1Lf'''''''''_f'''''''''_Boolsbos,CTf'''''''''_f'''''''''_Bool) > (lizzieLet41_1_argbuf,CTf'''''''''_f'''''''''_Bool) */
  \CTf'''''''''_f'''''''''_Bool_t  \go_7_1Lf'''''''''_f'''''''''_Boolsbos_bufchan_d ;
  logic \go_7_1Lf'''''''''_f'''''''''_Boolsbos_bufchan_r ;
  assign \go_7_1Lf'''''''''_f'''''''''_Boolsbos_r  = ((! \go_7_1Lf'''''''''_f'''''''''_Boolsbos_bufchan_d [0]) || \go_7_1Lf'''''''''_f'''''''''_Boolsbos_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \go_7_1Lf'''''''''_f'''''''''_Boolsbos_bufchan_d  <= {115'd0,
                                                            1'd0};
    else
      if (\go_7_1Lf'''''''''_f'''''''''_Boolsbos_r )
        \go_7_1Lf'''''''''_f'''''''''_Boolsbos_bufchan_d  <= \go_7_1Lf'''''''''_f'''''''''_Boolsbos_d ;
  \CTf'''''''''_f'''''''''_Bool_t  \go_7_1Lf'''''''''_f'''''''''_Boolsbos_bufchan_buf ;
  assign \go_7_1Lf'''''''''_f'''''''''_Boolsbos_bufchan_r  = (! \go_7_1Lf'''''''''_f'''''''''_Boolsbos_bufchan_buf [0]);
  assign lizzieLet41_1_argbuf_d = (\go_7_1Lf'''''''''_f'''''''''_Boolsbos_bufchan_buf [0] ? \go_7_1Lf'''''''''_f'''''''''_Boolsbos_bufchan_buf  :
                                   \go_7_1Lf'''''''''_f'''''''''_Boolsbos_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \go_7_1Lf'''''''''_f'''''''''_Boolsbos_bufchan_buf  <= {115'd0,
                                                              1'd0};
    else
      if ((lizzieLet41_1_argbuf_r && \go_7_1Lf'''''''''_f'''''''''_Boolsbos_bufchan_buf [0]))
        \go_7_1Lf'''''''''_f'''''''''_Boolsbos_bufchan_buf  <= {115'd0,
                                                                1'd0};
      else if (((! lizzieLet41_1_argbuf_r) && (! \go_7_1Lf'''''''''_f'''''''''_Boolsbos_bufchan_buf [0])))
        \go_7_1Lf'''''''''_f'''''''''_Boolsbos_bufchan_buf  <= \go_7_1Lf'''''''''_f'''''''''_Boolsbos_bufchan_d ;
  
  /* buf (Ty Go) : (go_7_2,Go) > (go_7_2_argbuf,Go) */
  Go_t go_7_2_bufchan_d;
  logic go_7_2_bufchan_r;
  assign go_7_2_r = ((! go_7_2_bufchan_d[0]) || go_7_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_7_2_bufchan_d <= 1'd0;
    else if (go_7_2_r) go_7_2_bufchan_d <= go_7_2_d;
  Go_t go_7_2_bufchan_buf;
  assign go_7_2_bufchan_r = (! go_7_2_bufchan_buf[0]);
  assign go_7_2_argbuf_d = (go_7_2_bufchan_buf[0] ? go_7_2_bufchan_buf :
                            go_7_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_7_2_bufchan_buf <= 1'd0;
    else
      if ((go_7_2_argbuf_r && go_7_2_bufchan_buf[0]))
        go_7_2_bufchan_buf <= 1'd0;
      else if (((! go_7_2_argbuf_r) && (! go_7_2_bufchan_buf[0])))
        go_7_2_bufchan_buf <= go_7_2_bufchan_d;
  
  /* dcon (Ty TupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_CTf'''''''''_f'''''''''_Bool,
      Dcon TupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_CTf'''''''''_f'''''''''_Bool) : [(go_7_2_argbuf,Go),
                                                                                                     (q4a8w_1_1_argbuf,Pointer_MaskQTree),
                                                                                                     (q4'a8x_1_1_argbuf,Pointer_QTree_Bool),
                                                                                                     (lizzieLet5_1_1_argbuf,Pointer_CTf'''''''''_f'''''''''_Bool)] > (call_f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_CTf'''''''''_f'''''''''_Bool_1,TupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_CTf'''''''''_f'''''''''_Bool) */
  assign \call_f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_CTf'''''''''_f'''''''''_Bool_1_d  = \TupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_CTf'''''''''_f'''''''''_Bool_dc ((& {go_7_2_argbuf_d[0],
                                                                                                                                                                                                                                     q4a8w_1_1_argbuf_d[0],
                                                                                                                                                                                                                                     \q4'a8x_1_1_argbuf_d [0],
                                                                                                                                                                                                                                     lizzieLet5_1_1_argbuf_d[0]}), go_7_2_argbuf_d, q4a8w_1_1_argbuf_d, \q4'a8x_1_1_argbuf_d , lizzieLet5_1_1_argbuf_d);
  assign {go_7_2_argbuf_r,
          q4a8w_1_1_argbuf_r,
          \q4'a8x_1_1_argbuf_r ,
          lizzieLet5_1_1_argbuf_r} = {4 {(\call_f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_CTf'''''''''_f'''''''''_Bool_1_r  && \call_f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_CTf'''''''''_f'''''''''_Bool_1_d [0])}};
  
  /* dcon (Ty QTree_Bool,
      Dcon QVal_Bool) : [(go_8_1MyTrue,MyBool)] > (lizzieLet0_1_1QVal_Bool,QTree_Bool) */
  assign lizzieLet0_1_1QVal_Bool_d = QVal_Bool_dc((& {go_8_1MyTrue_d[0]}), go_8_1MyTrue_d);
  assign {go_8_1MyTrue_r} = {1 {(lizzieLet0_1_1QVal_Bool_r && lizzieLet0_1_1QVal_Bool_d[0])}};
  
  /* fork (Ty C17) : (go_9_goMux_choice,C17) > [(go_9_goMux_choice_1,C17),
                                           (go_9_goMux_choice_2,C17)] */
  logic [1:0] go_9_goMux_choice_emitted;
  logic [1:0] go_9_goMux_choice_done;
  assign go_9_goMux_choice_1_d = {go_9_goMux_choice_d[5:1],
                                  (go_9_goMux_choice_d[0] && (! go_9_goMux_choice_emitted[0]))};
  assign go_9_goMux_choice_2_d = {go_9_goMux_choice_d[5:1],
                                  (go_9_goMux_choice_d[0] && (! go_9_goMux_choice_emitted[1]))};
  assign go_9_goMux_choice_done = (go_9_goMux_choice_emitted | ({go_9_goMux_choice_2_d[0],
                                                                 go_9_goMux_choice_1_d[0]} & {go_9_goMux_choice_2_r,
                                                                                              go_9_goMux_choice_1_r}));
  assign go_9_goMux_choice_r = (& go_9_goMux_choice_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_9_goMux_choice_emitted <= 2'd0;
    else
      go_9_goMux_choice_emitted <= (go_9_goMux_choice_r ? 2'd0 :
                                    go_9_goMux_choice_done);
  
  /* mux (Ty C17,
     Ty Pointer_QTree_Bool) : (go_9_goMux_choice_1,C17) [(lizzieLet13_1_argbuf,Pointer_QTree_Bool),
                                                         (contRet_0_1_argbuf,Pointer_QTree_Bool),
                                                         (lizzieLet14_1_argbuf,Pointer_QTree_Bool),
                                                         (lizzieLet15_1_argbuf,Pointer_QTree_Bool),
                                                         (lizzieLet16_1_argbuf,Pointer_QTree_Bool),
                                                         (lizzieLet17_1_argbuf,Pointer_QTree_Bool),
                                                         (lizzieLet18_1_argbuf,Pointer_QTree_Bool),
                                                         (lizzieLet19_1_argbuf,Pointer_QTree_Bool),
                                                         (lizzieLet20_1_argbuf,Pointer_QTree_Bool),
                                                         (lizzieLet21_1_argbuf,Pointer_QTree_Bool),
                                                         (lizzieLet22_1_argbuf,Pointer_QTree_Bool),
                                                         (lizzieLet23_1_argbuf,Pointer_QTree_Bool),
                                                         (lizzieLet19_1_1_argbuf,Pointer_QTree_Bool),
                                                         (lizzieLet24_1_argbuf,Pointer_QTree_Bool),
                                                         (lizzieLet25_1_argbuf,Pointer_QTree_Bool),
                                                         (lizzieLet26_1_argbuf,Pointer_QTree_Bool),
                                                         (lizzieLet27_1_argbuf,Pointer_QTree_Bool)] > (srtarg_0_goMux_mux,Pointer_QTree_Bool) */
  logic [16:0] srtarg_0_goMux_mux_mux;
  logic [16:0] srtarg_0_goMux_mux_onehot;
  always_comb
    unique case (go_9_goMux_choice_1_d[5:1])
      5'd0:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {17'd1,
                                                               lizzieLet13_1_argbuf_d};
      5'd1:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {17'd2,
                                                               contRet_0_1_argbuf_d};
      5'd2:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {17'd4,
                                                               lizzieLet14_1_argbuf_d};
      5'd3:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {17'd8,
                                                               lizzieLet15_1_argbuf_d};
      5'd4:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {17'd16,
                                                               lizzieLet16_1_argbuf_d};
      5'd5:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {17'd32,
                                                               lizzieLet17_1_argbuf_d};
      5'd6:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {17'd64,
                                                               lizzieLet18_1_argbuf_d};
      5'd7:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {17'd128,
                                                               lizzieLet19_1_argbuf_d};
      5'd8:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {17'd256,
                                                               lizzieLet20_1_argbuf_d};
      5'd9:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {17'd512,
                                                               lizzieLet21_1_argbuf_d};
      5'd10:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {17'd1024,
                                                               lizzieLet22_1_argbuf_d};
      5'd11:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {17'd2048,
                                                               lizzieLet23_1_argbuf_d};
      5'd12:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {17'd4096,
                                                               lizzieLet19_1_1_argbuf_d};
      5'd13:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {17'd8192,
                                                               lizzieLet24_1_argbuf_d};
      5'd14:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {17'd16384,
                                                               lizzieLet25_1_argbuf_d};
      5'd15:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {17'd32768,
                                                               lizzieLet26_1_argbuf_d};
      5'd16:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {17'd65536,
                                                               lizzieLet27_1_argbuf_d};
      default:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {17'd0,
                                                               {16'd0, 1'd0}};
    endcase
  assign srtarg_0_goMux_mux_d = {srtarg_0_goMux_mux_mux[16:1],
                                 (srtarg_0_goMux_mux_mux[0] && go_9_goMux_choice_1_d[0])};
  assign go_9_goMux_choice_1_r = (srtarg_0_goMux_mux_d[0] && srtarg_0_goMux_mux_r);
  assign {lizzieLet27_1_argbuf_r,
          lizzieLet26_1_argbuf_r,
          lizzieLet25_1_argbuf_r,
          lizzieLet24_1_argbuf_r,
          lizzieLet19_1_1_argbuf_r,
          lizzieLet23_1_argbuf_r,
          lizzieLet22_1_argbuf_r,
          lizzieLet21_1_argbuf_r,
          lizzieLet20_1_argbuf_r,
          lizzieLet19_1_argbuf_r,
          lizzieLet18_1_argbuf_r,
          lizzieLet17_1_argbuf_r,
          lizzieLet16_1_argbuf_r,
          lizzieLet15_1_argbuf_r,
          lizzieLet14_1_argbuf_r,
          contRet_0_1_argbuf_r,
          lizzieLet13_1_argbuf_r} = (go_9_goMux_choice_1_r ? srtarg_0_goMux_mux_onehot :
                                     17'd0);
  
  /* mux (Ty C17,
     Ty Pointer_CTf) : (go_9_goMux_choice_2,C17) [(lizzieLet0_8MQNone_1_argbuf,Pointer_CTf),
                                                  (sc_0_6_1_argbuf,Pointer_CTf),
                                                  (lizzieLet0_8MQVal_1_argbuf,Pointer_CTf),
                                                  (lizzieLet0_4MQNode_4QNone_Bool_4QNone_Bool_1_argbuf,Pointer_CTf),
                                                  (lizzieLet0_4MQNode_4QNone_Bool_4QVal_Bool_1_argbuf,Pointer_CTf),
                                                  (lizzieLet0_4MQNode_4QNone_Bool_4QNode_Bool_1_argbuf,Pointer_CTf),
                                                  (lizzieLet0_4MQNode_4QNone_Bool_4QError_Bool_1_argbuf,Pointer_CTf),
                                                  (lizzieLet0_4MQNode_4QVal_Bool_4QNone_Bool_1_argbuf,Pointer_CTf),
                                                  (lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_2MyFalse_1_argbuf,Pointer_CTf),
                                                  (lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_2MyTrue_1_argbuf,Pointer_CTf),
                                                  (lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_2MyTrue_1_argbuf,Pointer_CTf),
                                                  (lizzieLet0_4MQNode_4QVal_Bool_4QNode_Bool_1_argbuf,Pointer_CTf),
                                                  (lizzieLet0_4MQNode_4QVal_Bool_4QError_Bool_1_argbuf,Pointer_CTf),
                                                  (lizzieLet0_4MQNode_4QNode_Bool_4QNone_Bool_1_argbuf,Pointer_CTf),
                                                  (lizzieLet0_4MQNode_4QNode_Bool_4QVal_Bool_1_argbuf,Pointer_CTf),
                                                  (lizzieLet0_4MQNode_4QNode_Bool_4QError_Bool_1_argbuf,Pointer_CTf),
                                                  (lizzieLet0_4MQNode_5QError_Bool_1_argbuf,Pointer_CTf)] > (scfarg_0_goMux_mux,Pointer_CTf) */
  logic [16:0] scfarg_0_goMux_mux_mux;
  logic [16:0] scfarg_0_goMux_mux_onehot;
  always_comb
    unique case (go_9_goMux_choice_2_d[5:1])
      5'd0:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {17'd1,
                                                               lizzieLet0_8MQNone_1_argbuf_d};
      5'd1:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {17'd2,
                                                               sc_0_6_1_argbuf_d};
      5'd2:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {17'd4,
                                                               lizzieLet0_8MQVal_1_argbuf_d};
      5'd3:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {17'd8,
                                                               lizzieLet0_4MQNode_4QNone_Bool_4QNone_Bool_1_argbuf_d};
      5'd4:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {17'd16,
                                                               lizzieLet0_4MQNode_4QNone_Bool_4QVal_Bool_1_argbuf_d};
      5'd5:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {17'd32,
                                                               lizzieLet0_4MQNode_4QNone_Bool_4QNode_Bool_1_argbuf_d};
      5'd6:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {17'd64,
                                                               lizzieLet0_4MQNode_4QNone_Bool_4QError_Bool_1_argbuf_d};
      5'd7:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {17'd128,
                                                               lizzieLet0_4MQNode_4QVal_Bool_4QNone_Bool_1_argbuf_d};
      5'd8:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {17'd256,
                                                               lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_2MyFalse_1_argbuf_d};
      5'd9:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {17'd512,
                                                               lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_2MyTrue_1_argbuf_d};
      5'd10:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {17'd1024,
                                                               lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_2MyTrue_1_argbuf_d};
      5'd11:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {17'd2048,
                                                               lizzieLet0_4MQNode_4QVal_Bool_4QNode_Bool_1_argbuf_d};
      5'd12:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {17'd4096,
                                                               lizzieLet0_4MQNode_4QVal_Bool_4QError_Bool_1_argbuf_d};
      5'd13:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {17'd8192,
                                                               lizzieLet0_4MQNode_4QNode_Bool_4QNone_Bool_1_argbuf_d};
      5'd14:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {17'd16384,
                                                               lizzieLet0_4MQNode_4QNode_Bool_4QVal_Bool_1_argbuf_d};
      5'd15:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {17'd32768,
                                                               lizzieLet0_4MQNode_4QNode_Bool_4QError_Bool_1_argbuf_d};
      5'd16:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {17'd65536,
                                                               lizzieLet0_4MQNode_5QError_Bool_1_argbuf_d};
      default:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {17'd0,
                                                               {16'd0, 1'd0}};
    endcase
  assign scfarg_0_goMux_mux_d = {scfarg_0_goMux_mux_mux[16:1],
                                 (scfarg_0_goMux_mux_mux[0] && go_9_goMux_choice_2_d[0])};
  assign go_9_goMux_choice_2_r = (scfarg_0_goMux_mux_d[0] && scfarg_0_goMux_mux_r);
  assign {lizzieLet0_4MQNode_5QError_Bool_1_argbuf_r,
          lizzieLet0_4MQNode_4QNode_Bool_4QError_Bool_1_argbuf_r,
          lizzieLet0_4MQNode_4QNode_Bool_4QVal_Bool_1_argbuf_r,
          lizzieLet0_4MQNode_4QNode_Bool_4QNone_Bool_1_argbuf_r,
          lizzieLet0_4MQNode_4QVal_Bool_4QError_Bool_1_argbuf_r,
          lizzieLet0_4MQNode_4QVal_Bool_4QNode_Bool_1_argbuf_r,
          lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_2MyTrue_1_argbuf_r,
          lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_2MyTrue_1_argbuf_r,
          lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_2MyFalse_1_argbuf_r,
          lizzieLet0_4MQNode_4QVal_Bool_4QNone_Bool_1_argbuf_r,
          lizzieLet0_4MQNode_4QNone_Bool_4QError_Bool_1_argbuf_r,
          lizzieLet0_4MQNode_4QNone_Bool_4QNode_Bool_1_argbuf_r,
          lizzieLet0_4MQNode_4QNone_Bool_4QVal_Bool_1_argbuf_r,
          lizzieLet0_4MQNode_4QNone_Bool_4QNone_Bool_1_argbuf_r,
          lizzieLet0_8MQVal_1_argbuf_r,
          sc_0_6_1_argbuf_r,
          lizzieLet0_8MQNone_1_argbuf_r} = (go_9_goMux_choice_2_r ? scfarg_0_goMux_mux_onehot :
                                            17'd0);
  
  /* destruct (Ty MaskQTree,
          Dcon MQNode) : (lizzieLet0_1MQNode,MaskQTree) > [(q1a88_destruct,Pointer_MaskQTree),
                                                           (q2a89_destruct,Pointer_MaskQTree),
                                                           (q3a8a_destruct,Pointer_MaskQTree),
                                                           (q4a8b_destruct,Pointer_MaskQTree)] */
  logic [3:0] lizzieLet0_1MQNode_emitted;
  logic [3:0] lizzieLet0_1MQNode_done;
  assign q1a88_destruct_d = {lizzieLet0_1MQNode_d[18:3],
                             (lizzieLet0_1MQNode_d[0] && (! lizzieLet0_1MQNode_emitted[0]))};
  assign q2a89_destruct_d = {lizzieLet0_1MQNode_d[34:19],
                             (lizzieLet0_1MQNode_d[0] && (! lizzieLet0_1MQNode_emitted[1]))};
  assign q3a8a_destruct_d = {lizzieLet0_1MQNode_d[50:35],
                             (lizzieLet0_1MQNode_d[0] && (! lizzieLet0_1MQNode_emitted[2]))};
  assign q4a8b_destruct_d = {lizzieLet0_1MQNode_d[66:51],
                             (lizzieLet0_1MQNode_d[0] && (! lizzieLet0_1MQNode_emitted[3]))};
  assign lizzieLet0_1MQNode_done = (lizzieLet0_1MQNode_emitted | ({q4a8b_destruct_d[0],
                                                                   q3a8a_destruct_d[0],
                                                                   q2a89_destruct_d[0],
                                                                   q1a88_destruct_d[0]} & {q4a8b_destruct_r,
                                                                                           q3a8a_destruct_r,
                                                                                           q2a89_destruct_r,
                                                                                           q1a88_destruct_r}));
  assign lizzieLet0_1MQNode_r = (& lizzieLet0_1MQNode_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet0_1MQNode_emitted <= 4'd0;
    else
      lizzieLet0_1MQNode_emitted <= (lizzieLet0_1MQNode_r ? 4'd0 :
                                     lizzieLet0_1MQNode_done);
  
  /* buf (Ty QTree_Bool) : (lizzieLet0_1_1QVal_Bool,QTree_Bool) > (lizzieLet42_1_argbuf,QTree_Bool) */
  QTree_Bool_t lizzieLet0_1_1QVal_Bool_bufchan_d;
  logic lizzieLet0_1_1QVal_Bool_bufchan_r;
  assign lizzieLet0_1_1QVal_Bool_r = ((! lizzieLet0_1_1QVal_Bool_bufchan_d[0]) || lizzieLet0_1_1QVal_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_1_1QVal_Bool_bufchan_d <= {66'd0, 1'd0};
    else
      if (lizzieLet0_1_1QVal_Bool_r)
        lizzieLet0_1_1QVal_Bool_bufchan_d <= lizzieLet0_1_1QVal_Bool_d;
  QTree_Bool_t lizzieLet0_1_1QVal_Bool_bufchan_buf;
  assign lizzieLet0_1_1QVal_Bool_bufchan_r = (! lizzieLet0_1_1QVal_Bool_bufchan_buf[0]);
  assign lizzieLet42_1_argbuf_d = (lizzieLet0_1_1QVal_Bool_bufchan_buf[0] ? lizzieLet0_1_1QVal_Bool_bufchan_buf :
                                   lizzieLet0_1_1QVal_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_1_1QVal_Bool_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((lizzieLet42_1_argbuf_r && lizzieLet0_1_1QVal_Bool_bufchan_buf[0]))
        lizzieLet0_1_1QVal_Bool_bufchan_buf <= {66'd0, 1'd0};
      else if (((! lizzieLet42_1_argbuf_r) && (! lizzieLet0_1_1QVal_Bool_bufchan_buf[0])))
        lizzieLet0_1_1QVal_Bool_bufchan_buf <= lizzieLet0_1_1QVal_Bool_bufchan_d;
  
  /* demux (Ty MaskQTree,
       Ty MaskQTree) : (lizzieLet0_2,MaskQTree) (lizzieLet0_1,MaskQTree) > [(_125,MaskQTree),
                                                                            (_124,MaskQTree),
                                                                            (lizzieLet0_1MQNode,MaskQTree)] */
  logic [2:0] lizzieLet0_1_onehotd;
  always_comb
    if ((lizzieLet0_2_d[0] && lizzieLet0_1_d[0]))
      unique case (lizzieLet0_2_d[2:1])
        2'd0: lizzieLet0_1_onehotd = 3'd1;
        2'd1: lizzieLet0_1_onehotd = 3'd2;
        2'd2: lizzieLet0_1_onehotd = 3'd4;
        default: lizzieLet0_1_onehotd = 3'd0;
      endcase
    else lizzieLet0_1_onehotd = 3'd0;
  assign _125_d = {lizzieLet0_1_d[66:1], lizzieLet0_1_onehotd[0]};
  assign _124_d = {lizzieLet0_1_d[66:1], lizzieLet0_1_onehotd[1]};
  assign lizzieLet0_1MQNode_d = {lizzieLet0_1_d[66:1],
                                 lizzieLet0_1_onehotd[2]};
  assign lizzieLet0_1_r = (| (lizzieLet0_1_onehotd & {lizzieLet0_1MQNode_r,
                                                      _124_r,
                                                      _125_r}));
  assign lizzieLet0_2_r = lizzieLet0_1_r;
  
  /* demux (Ty MaskQTree,
       Ty Go) : (lizzieLet0_3,MaskQTree) (go_2_goMux_data,Go) > [(lizzieLet0_3MQNone,Go),
                                                                 (lizzieLet0_3MQVal,Go),
                                                                 (lizzieLet0_3MQNode,Go)] */
  logic [2:0] go_2_goMux_data_onehotd;
  always_comb
    if ((lizzieLet0_3_d[0] && go_2_goMux_data_d[0]))
      unique case (lizzieLet0_3_d[2:1])
        2'd0: go_2_goMux_data_onehotd = 3'd1;
        2'd1: go_2_goMux_data_onehotd = 3'd2;
        2'd2: go_2_goMux_data_onehotd = 3'd4;
        default: go_2_goMux_data_onehotd = 3'd0;
      endcase
    else go_2_goMux_data_onehotd = 3'd0;
  assign lizzieLet0_3MQNone_d = go_2_goMux_data_onehotd[0];
  assign lizzieLet0_3MQVal_d = go_2_goMux_data_onehotd[1];
  assign lizzieLet0_3MQNode_d = go_2_goMux_data_onehotd[2];
  assign go_2_goMux_data_r = (| (go_2_goMux_data_onehotd & {lizzieLet0_3MQNode_r,
                                                            lizzieLet0_3MQVal_r,
                                                            lizzieLet0_3MQNone_r}));
  assign lizzieLet0_3_r = go_2_goMux_data_r;
  
  /* fork (Ty Go) : (lizzieLet0_3MQNone,Go) > [(lizzieLet0_3MQNone_1,Go),
                                          (lizzieLet0_3MQNone_2,Go)] */
  logic [1:0] lizzieLet0_3MQNone_emitted;
  logic [1:0] lizzieLet0_3MQNone_done;
  assign lizzieLet0_3MQNone_1_d = (lizzieLet0_3MQNone_d[0] && (! lizzieLet0_3MQNone_emitted[0]));
  assign lizzieLet0_3MQNone_2_d = (lizzieLet0_3MQNone_d[0] && (! lizzieLet0_3MQNone_emitted[1]));
  assign lizzieLet0_3MQNone_done = (lizzieLet0_3MQNone_emitted | ({lizzieLet0_3MQNone_2_d[0],
                                                                   lizzieLet0_3MQNone_1_d[0]} & {lizzieLet0_3MQNone_2_r,
                                                                                                 lizzieLet0_3MQNone_1_r}));
  assign lizzieLet0_3MQNone_r = (& lizzieLet0_3MQNone_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet0_3MQNone_emitted <= 2'd0;
    else
      lizzieLet0_3MQNone_emitted <= (lizzieLet0_3MQNone_r ? 2'd0 :
                                     lizzieLet0_3MQNone_done);
  
  /* dcon (Ty QTree_Bool,
      Dcon QNone_Bool) : [(lizzieLet0_3MQNone_1,Go)] > (lizzieLet0_3MQNone_1QNone_Bool,QTree_Bool) */
  assign lizzieLet0_3MQNone_1QNone_Bool_d = QNone_Bool_dc((& {lizzieLet0_3MQNone_1_d[0]}), lizzieLet0_3MQNone_1_d);
  assign {lizzieLet0_3MQNone_1_r} = {1 {(lizzieLet0_3MQNone_1QNone_Bool_r && lizzieLet0_3MQNone_1QNone_Bool_d[0])}};
  
  /* buf (Ty QTree_Bool) : (lizzieLet0_3MQNone_1QNone_Bool,QTree_Bool) > (lizzieLet1_1_argbuf,QTree_Bool) */
  QTree_Bool_t lizzieLet0_3MQNone_1QNone_Bool_bufchan_d;
  logic lizzieLet0_3MQNone_1QNone_Bool_bufchan_r;
  assign lizzieLet0_3MQNone_1QNone_Bool_r = ((! lizzieLet0_3MQNone_1QNone_Bool_bufchan_d[0]) || lizzieLet0_3MQNone_1QNone_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_3MQNone_1QNone_Bool_bufchan_d <= {66'd0, 1'd0};
    else
      if (lizzieLet0_3MQNone_1QNone_Bool_r)
        lizzieLet0_3MQNone_1QNone_Bool_bufchan_d <= lizzieLet0_3MQNone_1QNone_Bool_d;
  QTree_Bool_t lizzieLet0_3MQNone_1QNone_Bool_bufchan_buf;
  assign lizzieLet0_3MQNone_1QNone_Bool_bufchan_r = (! lizzieLet0_3MQNone_1QNone_Bool_bufchan_buf[0]);
  assign lizzieLet1_1_argbuf_d = (lizzieLet0_3MQNone_1QNone_Bool_bufchan_buf[0] ? lizzieLet0_3MQNone_1QNone_Bool_bufchan_buf :
                                  lizzieLet0_3MQNone_1QNone_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_3MQNone_1QNone_Bool_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((lizzieLet1_1_argbuf_r && lizzieLet0_3MQNone_1QNone_Bool_bufchan_buf[0]))
        lizzieLet0_3MQNone_1QNone_Bool_bufchan_buf <= {66'd0, 1'd0};
      else if (((! lizzieLet1_1_argbuf_r) && (! lizzieLet0_3MQNone_1QNone_Bool_bufchan_buf[0])))
        lizzieLet0_3MQNone_1QNone_Bool_bufchan_buf <= lizzieLet0_3MQNone_1QNone_Bool_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet0_3MQNone_2,Go) > (lizzieLet0_3MQNone_2_argbuf,Go) */
  Go_t lizzieLet0_3MQNone_2_bufchan_d;
  logic lizzieLet0_3MQNone_2_bufchan_r;
  assign lizzieLet0_3MQNone_2_r = ((! lizzieLet0_3MQNone_2_bufchan_d[0]) || lizzieLet0_3MQNone_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet0_3MQNone_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet0_3MQNone_2_r)
        lizzieLet0_3MQNone_2_bufchan_d <= lizzieLet0_3MQNone_2_d;
  Go_t lizzieLet0_3MQNone_2_bufchan_buf;
  assign lizzieLet0_3MQNone_2_bufchan_r = (! lizzieLet0_3MQNone_2_bufchan_buf[0]);
  assign lizzieLet0_3MQNone_2_argbuf_d = (lizzieLet0_3MQNone_2_bufchan_buf[0] ? lizzieLet0_3MQNone_2_bufchan_buf :
                                          lizzieLet0_3MQNone_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet0_3MQNone_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet0_3MQNone_2_argbuf_r && lizzieLet0_3MQNone_2_bufchan_buf[0]))
        lizzieLet0_3MQNone_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet0_3MQNone_2_argbuf_r) && (! lizzieLet0_3MQNone_2_bufchan_buf[0])))
        lizzieLet0_3MQNone_2_bufchan_buf <= lizzieLet0_3MQNone_2_bufchan_d;
  
  /* mergectrl (Ty C17,Ty Go) : [(lizzieLet0_3MQNone_2_argbuf,Go),
                            (lizzieLet43_3Lcall_f0_1_argbuf,Go),
                            (lizzieLet0_3MQVal_2_argbuf,Go),
                            (lizzieLet0_4MQNode_4QNone_Bool_3QNone_Bool_2_argbuf,Go),
                            (lizzieLet0_4MQNode_4QNone_Bool_3QVal_Bool_2_argbuf,Go),
                            (lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_5_argbuf,Go),
                            (lizzieLet0_4MQNode_4QNone_Bool_3QError_Bool_2_argbuf,Go),
                            (lizzieLet0_4MQNode_4QVal_Bool_3QNone_Bool_2_argbuf,Go),
                            (lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyFalse_2_argbuf,Go),
                            (lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyTrue_2_argbuf,Go),
                            (lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyTrue_2_argbuf,Go),
                            (lizzieLet0_4MQNode_4QVal_Bool_3QNode_Bool_2_argbuf,Go),
                            (lizzieLet0_4MQNode_4QVal_Bool_3QError_Bool_2_argbuf,Go),
                            (lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_5_argbuf,Go),
                            (lizzieLet0_4MQNode_4QNode_Bool_3QVal_Bool_2_argbuf,Go),
                            (lizzieLet0_4MQNode_4QNode_Bool_3QError_Bool_2_argbuf,Go),
                            (lizzieLet0_4MQNode_3QError_Bool_2_argbuf,Go)] > (go_9_goMux_choice,C17) (go_9_goMux_data,Go) */
  logic [16:0] lizzieLet0_3MQNone_2_argbuf_select_d;
  assign lizzieLet0_3MQNone_2_argbuf_select_d = ((| lizzieLet0_3MQNone_2_argbuf_select_q) ? lizzieLet0_3MQNone_2_argbuf_select_q :
                                                 (lizzieLet0_3MQNone_2_argbuf_d[0] ? 17'd1 :
                                                  (lizzieLet43_3Lcall_f0_1_argbuf_d[0] ? 17'd2 :
                                                   (lizzieLet0_3MQVal_2_argbuf_d[0] ? 17'd4 :
                                                    (lizzieLet0_4MQNode_4QNone_Bool_3QNone_Bool_2_argbuf_d[0] ? 17'd8 :
                                                     (lizzieLet0_4MQNode_4QNone_Bool_3QVal_Bool_2_argbuf_d[0] ? 17'd16 :
                                                      (lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_5_argbuf_d[0] ? 17'd32 :
                                                       (lizzieLet0_4MQNode_4QNone_Bool_3QError_Bool_2_argbuf_d[0] ? 17'd64 :
                                                        (lizzieLet0_4MQNode_4QVal_Bool_3QNone_Bool_2_argbuf_d[0] ? 17'd128 :
                                                         (lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyFalse_2_argbuf_d[0] ? 17'd256 :
                                                          (lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyTrue_2_argbuf_d[0] ? 17'd512 :
                                                           (lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyTrue_2_argbuf_d[0] ? 17'd1024 :
                                                            (lizzieLet0_4MQNode_4QVal_Bool_3QNode_Bool_2_argbuf_d[0] ? 17'd2048 :
                                                             (lizzieLet0_4MQNode_4QVal_Bool_3QError_Bool_2_argbuf_d[0] ? 17'd4096 :
                                                              (lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_5_argbuf_d[0] ? 17'd8192 :
                                                               (lizzieLet0_4MQNode_4QNode_Bool_3QVal_Bool_2_argbuf_d[0] ? 17'd16384 :
                                                                (lizzieLet0_4MQNode_4QNode_Bool_3QError_Bool_2_argbuf_d[0] ? 17'd32768 :
                                                                 (lizzieLet0_4MQNode_3QError_Bool_2_argbuf_d[0] ? 17'd65536 :
                                                                  17'd0))))))))))))))))));
  logic [16:0] lizzieLet0_3MQNone_2_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet0_3MQNone_2_argbuf_select_q <= 17'd0;
    else
      lizzieLet0_3MQNone_2_argbuf_select_q <= (lizzieLet0_3MQNone_2_argbuf_done ? 17'd0 :
                                               lizzieLet0_3MQNone_2_argbuf_select_d);
  logic [1:0] lizzieLet0_3MQNone_2_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet0_3MQNone_2_argbuf_emit_q <= 2'd0;
    else
      lizzieLet0_3MQNone_2_argbuf_emit_q <= (lizzieLet0_3MQNone_2_argbuf_done ? 2'd0 :
                                             lizzieLet0_3MQNone_2_argbuf_emit_d);
  logic [1:0] lizzieLet0_3MQNone_2_argbuf_emit_d;
  assign lizzieLet0_3MQNone_2_argbuf_emit_d = (lizzieLet0_3MQNone_2_argbuf_emit_q | ({go_9_goMux_choice_d[0],
                                                                                      go_9_goMux_data_d[0]} & {go_9_goMux_choice_r,
                                                                                                               go_9_goMux_data_r}));
  logic lizzieLet0_3MQNone_2_argbuf_done;
  assign lizzieLet0_3MQNone_2_argbuf_done = (& lizzieLet0_3MQNone_2_argbuf_emit_d);
  assign {lizzieLet0_4MQNode_3QError_Bool_2_argbuf_r,
          lizzieLet0_4MQNode_4QNode_Bool_3QError_Bool_2_argbuf_r,
          lizzieLet0_4MQNode_4QNode_Bool_3QVal_Bool_2_argbuf_r,
          lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_5_argbuf_r,
          lizzieLet0_4MQNode_4QVal_Bool_3QError_Bool_2_argbuf_r,
          lizzieLet0_4MQNode_4QVal_Bool_3QNode_Bool_2_argbuf_r,
          lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyTrue_2_argbuf_r,
          lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyTrue_2_argbuf_r,
          lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyFalse_2_argbuf_r,
          lizzieLet0_4MQNode_4QVal_Bool_3QNone_Bool_2_argbuf_r,
          lizzieLet0_4MQNode_4QNone_Bool_3QError_Bool_2_argbuf_r,
          lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_5_argbuf_r,
          lizzieLet0_4MQNode_4QNone_Bool_3QVal_Bool_2_argbuf_r,
          lizzieLet0_4MQNode_4QNone_Bool_3QNone_Bool_2_argbuf_r,
          lizzieLet0_3MQVal_2_argbuf_r,
          lizzieLet43_3Lcall_f0_1_argbuf_r,
          lizzieLet0_3MQNone_2_argbuf_r} = (lizzieLet0_3MQNone_2_argbuf_done ? lizzieLet0_3MQNone_2_argbuf_select_d :
                                            17'd0);
  assign go_9_goMux_data_d = ((lizzieLet0_3MQNone_2_argbuf_select_d[0] && (! lizzieLet0_3MQNone_2_argbuf_emit_q[0])) ? lizzieLet0_3MQNone_2_argbuf_d :
                              ((lizzieLet0_3MQNone_2_argbuf_select_d[1] && (! lizzieLet0_3MQNone_2_argbuf_emit_q[0])) ? lizzieLet43_3Lcall_f0_1_argbuf_d :
                               ((lizzieLet0_3MQNone_2_argbuf_select_d[2] && (! lizzieLet0_3MQNone_2_argbuf_emit_q[0])) ? lizzieLet0_3MQVal_2_argbuf_d :
                                ((lizzieLet0_3MQNone_2_argbuf_select_d[3] && (! lizzieLet0_3MQNone_2_argbuf_emit_q[0])) ? lizzieLet0_4MQNode_4QNone_Bool_3QNone_Bool_2_argbuf_d :
                                 ((lizzieLet0_3MQNone_2_argbuf_select_d[4] && (! lizzieLet0_3MQNone_2_argbuf_emit_q[0])) ? lizzieLet0_4MQNode_4QNone_Bool_3QVal_Bool_2_argbuf_d :
                                  ((lizzieLet0_3MQNone_2_argbuf_select_d[5] && (! lizzieLet0_3MQNone_2_argbuf_emit_q[0])) ? lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_5_argbuf_d :
                                   ((lizzieLet0_3MQNone_2_argbuf_select_d[6] && (! lizzieLet0_3MQNone_2_argbuf_emit_q[0])) ? lizzieLet0_4MQNode_4QNone_Bool_3QError_Bool_2_argbuf_d :
                                    ((lizzieLet0_3MQNone_2_argbuf_select_d[7] && (! lizzieLet0_3MQNone_2_argbuf_emit_q[0])) ? lizzieLet0_4MQNode_4QVal_Bool_3QNone_Bool_2_argbuf_d :
                                     ((lizzieLet0_3MQNone_2_argbuf_select_d[8] && (! lizzieLet0_3MQNone_2_argbuf_emit_q[0])) ? lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyFalse_2_argbuf_d :
                                      ((lizzieLet0_3MQNone_2_argbuf_select_d[9] && (! lizzieLet0_3MQNone_2_argbuf_emit_q[0])) ? lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyTrue_2_argbuf_d :
                                       ((lizzieLet0_3MQNone_2_argbuf_select_d[10] && (! lizzieLet0_3MQNone_2_argbuf_emit_q[0])) ? lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyTrue_2_argbuf_d :
                                        ((lizzieLet0_3MQNone_2_argbuf_select_d[11] && (! lizzieLet0_3MQNone_2_argbuf_emit_q[0])) ? lizzieLet0_4MQNode_4QVal_Bool_3QNode_Bool_2_argbuf_d :
                                         ((lizzieLet0_3MQNone_2_argbuf_select_d[12] && (! lizzieLet0_3MQNone_2_argbuf_emit_q[0])) ? lizzieLet0_4MQNode_4QVal_Bool_3QError_Bool_2_argbuf_d :
                                          ((lizzieLet0_3MQNone_2_argbuf_select_d[13] && (! lizzieLet0_3MQNone_2_argbuf_emit_q[0])) ? lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_5_argbuf_d :
                                           ((lizzieLet0_3MQNone_2_argbuf_select_d[14] && (! lizzieLet0_3MQNone_2_argbuf_emit_q[0])) ? lizzieLet0_4MQNode_4QNode_Bool_3QVal_Bool_2_argbuf_d :
                                            ((lizzieLet0_3MQNone_2_argbuf_select_d[15] && (! lizzieLet0_3MQNone_2_argbuf_emit_q[0])) ? lizzieLet0_4MQNode_4QNode_Bool_3QError_Bool_2_argbuf_d :
                                             ((lizzieLet0_3MQNone_2_argbuf_select_d[16] && (! lizzieLet0_3MQNone_2_argbuf_emit_q[0])) ? lizzieLet0_4MQNode_3QError_Bool_2_argbuf_d :
                                              1'd0)))))))))))))))));
  assign go_9_goMux_choice_d = ((lizzieLet0_3MQNone_2_argbuf_select_d[0] && (! lizzieLet0_3MQNone_2_argbuf_emit_q[1])) ? C1_17_dc(1'd1) :
                                ((lizzieLet0_3MQNone_2_argbuf_select_d[1] && (! lizzieLet0_3MQNone_2_argbuf_emit_q[1])) ? C2_17_dc(1'd1) :
                                 ((lizzieLet0_3MQNone_2_argbuf_select_d[2] && (! lizzieLet0_3MQNone_2_argbuf_emit_q[1])) ? C3_17_dc(1'd1) :
                                  ((lizzieLet0_3MQNone_2_argbuf_select_d[3] && (! lizzieLet0_3MQNone_2_argbuf_emit_q[1])) ? C4_17_dc(1'd1) :
                                   ((lizzieLet0_3MQNone_2_argbuf_select_d[4] && (! lizzieLet0_3MQNone_2_argbuf_emit_q[1])) ? C5_17_dc(1'd1) :
                                    ((lizzieLet0_3MQNone_2_argbuf_select_d[5] && (! lizzieLet0_3MQNone_2_argbuf_emit_q[1])) ? C6_17_dc(1'd1) :
                                     ((lizzieLet0_3MQNone_2_argbuf_select_d[6] && (! lizzieLet0_3MQNone_2_argbuf_emit_q[1])) ? C7_17_dc(1'd1) :
                                      ((lizzieLet0_3MQNone_2_argbuf_select_d[7] && (! lizzieLet0_3MQNone_2_argbuf_emit_q[1])) ? C8_17_dc(1'd1) :
                                       ((lizzieLet0_3MQNone_2_argbuf_select_d[8] && (! lizzieLet0_3MQNone_2_argbuf_emit_q[1])) ? C9_17_dc(1'd1) :
                                        ((lizzieLet0_3MQNone_2_argbuf_select_d[9] && (! lizzieLet0_3MQNone_2_argbuf_emit_q[1])) ? C10_17_dc(1'd1) :
                                         ((lizzieLet0_3MQNone_2_argbuf_select_d[10] && (! lizzieLet0_3MQNone_2_argbuf_emit_q[1])) ? C11_17_dc(1'd1) :
                                          ((lizzieLet0_3MQNone_2_argbuf_select_d[11] && (! lizzieLet0_3MQNone_2_argbuf_emit_q[1])) ? C12_17_dc(1'd1) :
                                           ((lizzieLet0_3MQNone_2_argbuf_select_d[12] && (! lizzieLet0_3MQNone_2_argbuf_emit_q[1])) ? C13_17_dc(1'd1) :
                                            ((lizzieLet0_3MQNone_2_argbuf_select_d[13] && (! lizzieLet0_3MQNone_2_argbuf_emit_q[1])) ? C14_17_dc(1'd1) :
                                             ((lizzieLet0_3MQNone_2_argbuf_select_d[14] && (! lizzieLet0_3MQNone_2_argbuf_emit_q[1])) ? C15_17_dc(1'd1) :
                                              ((lizzieLet0_3MQNone_2_argbuf_select_d[15] && (! lizzieLet0_3MQNone_2_argbuf_emit_q[1])) ? C16_17_dc(1'd1) :
                                               ((lizzieLet0_3MQNone_2_argbuf_select_d[16] && (! lizzieLet0_3MQNone_2_argbuf_emit_q[1])) ? C17_17_dc(1'd1) :
                                                {5'd0, 1'd0})))))))))))))))));
  
  /* fork (Ty Go) : (lizzieLet0_3MQVal,Go) > [(lizzieLet0_3MQVal_1,Go),
                                         (lizzieLet0_3MQVal_2,Go)] */
  logic [1:0] lizzieLet0_3MQVal_emitted;
  logic [1:0] lizzieLet0_3MQVal_done;
  assign lizzieLet0_3MQVal_1_d = (lizzieLet0_3MQVal_d[0] && (! lizzieLet0_3MQVal_emitted[0]));
  assign lizzieLet0_3MQVal_2_d = (lizzieLet0_3MQVal_d[0] && (! lizzieLet0_3MQVal_emitted[1]));
  assign lizzieLet0_3MQVal_done = (lizzieLet0_3MQVal_emitted | ({lizzieLet0_3MQVal_2_d[0],
                                                                 lizzieLet0_3MQVal_1_d[0]} & {lizzieLet0_3MQVal_2_r,
                                                                                              lizzieLet0_3MQVal_1_r}));
  assign lizzieLet0_3MQVal_r = (& lizzieLet0_3MQVal_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet0_3MQVal_emitted <= 2'd0;
    else
      lizzieLet0_3MQVal_emitted <= (lizzieLet0_3MQVal_r ? 2'd0 :
                                    lizzieLet0_3MQVal_done);
  
  /* buf (Ty Go) : (lizzieLet0_3MQVal_1,Go) > (lizzieLet0_3MQVal_1_argbuf,Go) */
  Go_t lizzieLet0_3MQVal_1_bufchan_d;
  logic lizzieLet0_3MQVal_1_bufchan_r;
  assign lizzieLet0_3MQVal_1_r = ((! lizzieLet0_3MQVal_1_bufchan_d[0]) || lizzieLet0_3MQVal_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet0_3MQVal_1_bufchan_d <= 1'd0;
    else
      if (lizzieLet0_3MQVal_1_r)
        lizzieLet0_3MQVal_1_bufchan_d <= lizzieLet0_3MQVal_1_d;
  Go_t lizzieLet0_3MQVal_1_bufchan_buf;
  assign lizzieLet0_3MQVal_1_bufchan_r = (! lizzieLet0_3MQVal_1_bufchan_buf[0]);
  assign lizzieLet0_3MQVal_1_argbuf_d = (lizzieLet0_3MQVal_1_bufchan_buf[0] ? lizzieLet0_3MQVal_1_bufchan_buf :
                                         lizzieLet0_3MQVal_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet0_3MQVal_1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet0_3MQVal_1_argbuf_r && lizzieLet0_3MQVal_1_bufchan_buf[0]))
        lizzieLet0_3MQVal_1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet0_3MQVal_1_argbuf_r) && (! lizzieLet0_3MQVal_1_bufchan_buf[0])))
        lizzieLet0_3MQVal_1_bufchan_buf <= lizzieLet0_3MQVal_1_bufchan_d;
  
  /* dcon (Ty TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool,
      Dcon TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool) : [(lizzieLet0_3MQVal_1_argbuf,Go),
                                                               (lizzieLet0_6MQVal_1_argbuf,Pointer_QTree_Bool),
                                                               (lizzieLet0_7MQVal_1_argbuf,Pointer_QTree_Bool)] > (f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_1,TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool) */
  assign \f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_1_d  = TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_dc((& {lizzieLet0_3MQVal_1_argbuf_d[0],
                                                                                                                          lizzieLet0_6MQVal_1_argbuf_d[0],
                                                                                                                          lizzieLet0_7MQVal_1_argbuf_d[0]}), lizzieLet0_3MQVal_1_argbuf_d, lizzieLet0_6MQVal_1_argbuf_d, lizzieLet0_7MQVal_1_argbuf_d);
  assign {lizzieLet0_3MQVal_1_argbuf_r,
          lizzieLet0_6MQVal_1_argbuf_r,
          lizzieLet0_7MQVal_1_argbuf_r} = {3 {(\f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_1_r  && \f'TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_1_d [0])}};
  
  /* buf (Ty Go) : (lizzieLet0_3MQVal_2,Go) > (lizzieLet0_3MQVal_2_argbuf,Go) */
  Go_t lizzieLet0_3MQVal_2_bufchan_d;
  logic lizzieLet0_3MQVal_2_bufchan_r;
  assign lizzieLet0_3MQVal_2_r = ((! lizzieLet0_3MQVal_2_bufchan_d[0]) || lizzieLet0_3MQVal_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet0_3MQVal_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet0_3MQVal_2_r)
        lizzieLet0_3MQVal_2_bufchan_d <= lizzieLet0_3MQVal_2_d;
  Go_t lizzieLet0_3MQVal_2_bufchan_buf;
  assign lizzieLet0_3MQVal_2_bufchan_r = (! lizzieLet0_3MQVal_2_bufchan_buf[0]);
  assign lizzieLet0_3MQVal_2_argbuf_d = (lizzieLet0_3MQVal_2_bufchan_buf[0] ? lizzieLet0_3MQVal_2_bufchan_buf :
                                         lizzieLet0_3MQVal_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet0_3MQVal_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet0_3MQVal_2_argbuf_r && lizzieLet0_3MQVal_2_bufchan_buf[0]))
        lizzieLet0_3MQVal_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet0_3MQVal_2_argbuf_r) && (! lizzieLet0_3MQVal_2_bufchan_buf[0])))
        lizzieLet0_3MQVal_2_bufchan_buf <= lizzieLet0_3MQVal_2_bufchan_d;
  
  /* demux (Ty MaskQTree,
       Ty QTree_Bool) : (lizzieLet0_4,MaskQTree) (readPointer_QTree_Boolm2a86_1_argbuf_rwb,QTree_Bool) > [(_123,QTree_Bool),
                                                                                                          (_122,QTree_Bool),
                                                                                                          (lizzieLet0_4MQNode,QTree_Bool)] */
  logic [2:0] readPointer_QTree_Boolm2a86_1_argbuf_rwb_onehotd;
  always_comb
    if ((lizzieLet0_4_d[0] && readPointer_QTree_Boolm2a86_1_argbuf_rwb_d[0]))
      unique case (lizzieLet0_4_d[2:1])
        2'd0: readPointer_QTree_Boolm2a86_1_argbuf_rwb_onehotd = 3'd1;
        2'd1: readPointer_QTree_Boolm2a86_1_argbuf_rwb_onehotd = 3'd2;
        2'd2: readPointer_QTree_Boolm2a86_1_argbuf_rwb_onehotd = 3'd4;
        default: readPointer_QTree_Boolm2a86_1_argbuf_rwb_onehotd = 3'd0;
      endcase
    else readPointer_QTree_Boolm2a86_1_argbuf_rwb_onehotd = 3'd0;
  assign _123_d = {readPointer_QTree_Boolm2a86_1_argbuf_rwb_d[66:1],
                   readPointer_QTree_Boolm2a86_1_argbuf_rwb_onehotd[0]};
  assign _122_d = {readPointer_QTree_Boolm2a86_1_argbuf_rwb_d[66:1],
                   readPointer_QTree_Boolm2a86_1_argbuf_rwb_onehotd[1]};
  assign lizzieLet0_4MQNode_d = {readPointer_QTree_Boolm2a86_1_argbuf_rwb_d[66:1],
                                 readPointer_QTree_Boolm2a86_1_argbuf_rwb_onehotd[2]};
  assign readPointer_QTree_Boolm2a86_1_argbuf_rwb_r = (| (readPointer_QTree_Boolm2a86_1_argbuf_rwb_onehotd & {lizzieLet0_4MQNode_r,
                                                                                                              _122_r,
                                                                                                              _123_r}));
  assign lizzieLet0_4_r = readPointer_QTree_Boolm2a86_1_argbuf_rwb_r;
  
  /* fork (Ty QTree_Bool) : (lizzieLet0_4MQNode,QTree_Bool) > [(lizzieLet0_4MQNode_1,QTree_Bool),
                                                          (lizzieLet0_4MQNode_2,QTree_Bool),
                                                          (lizzieLet0_4MQNode_3,QTree_Bool),
                                                          (lizzieLet0_4MQNode_4,QTree_Bool),
                                                          (lizzieLet0_4MQNode_5,QTree_Bool),
                                                          (lizzieLet0_4MQNode_6,QTree_Bool),
                                                          (lizzieLet0_4MQNode_7,QTree_Bool),
                                                          (lizzieLet0_4MQNode_8,QTree_Bool),
                                                          (lizzieLet0_4MQNode_9,QTree_Bool)] */
  logic [8:0] lizzieLet0_4MQNode_emitted;
  logic [8:0] lizzieLet0_4MQNode_done;
  assign lizzieLet0_4MQNode_1_d = {lizzieLet0_4MQNode_d[66:1],
                                   (lizzieLet0_4MQNode_d[0] && (! lizzieLet0_4MQNode_emitted[0]))};
  assign lizzieLet0_4MQNode_2_d = {lizzieLet0_4MQNode_d[66:1],
                                   (lizzieLet0_4MQNode_d[0] && (! lizzieLet0_4MQNode_emitted[1]))};
  assign lizzieLet0_4MQNode_3_d = {lizzieLet0_4MQNode_d[66:1],
                                   (lizzieLet0_4MQNode_d[0] && (! lizzieLet0_4MQNode_emitted[2]))};
  assign lizzieLet0_4MQNode_4_d = {lizzieLet0_4MQNode_d[66:1],
                                   (lizzieLet0_4MQNode_d[0] && (! lizzieLet0_4MQNode_emitted[3]))};
  assign lizzieLet0_4MQNode_5_d = {lizzieLet0_4MQNode_d[66:1],
                                   (lizzieLet0_4MQNode_d[0] && (! lizzieLet0_4MQNode_emitted[4]))};
  assign lizzieLet0_4MQNode_6_d = {lizzieLet0_4MQNode_d[66:1],
                                   (lizzieLet0_4MQNode_d[0] && (! lizzieLet0_4MQNode_emitted[5]))};
  assign lizzieLet0_4MQNode_7_d = {lizzieLet0_4MQNode_d[66:1],
                                   (lizzieLet0_4MQNode_d[0] && (! lizzieLet0_4MQNode_emitted[6]))};
  assign lizzieLet0_4MQNode_8_d = {lizzieLet0_4MQNode_d[66:1],
                                   (lizzieLet0_4MQNode_d[0] && (! lizzieLet0_4MQNode_emitted[7]))};
  assign lizzieLet0_4MQNode_9_d = {lizzieLet0_4MQNode_d[66:1],
                                   (lizzieLet0_4MQNode_d[0] && (! lizzieLet0_4MQNode_emitted[8]))};
  assign lizzieLet0_4MQNode_done = (lizzieLet0_4MQNode_emitted | ({lizzieLet0_4MQNode_9_d[0],
                                                                   lizzieLet0_4MQNode_8_d[0],
                                                                   lizzieLet0_4MQNode_7_d[0],
                                                                   lizzieLet0_4MQNode_6_d[0],
                                                                   lizzieLet0_4MQNode_5_d[0],
                                                                   lizzieLet0_4MQNode_4_d[0],
                                                                   lizzieLet0_4MQNode_3_d[0],
                                                                   lizzieLet0_4MQNode_2_d[0],
                                                                   lizzieLet0_4MQNode_1_d[0]} & {lizzieLet0_4MQNode_9_r,
                                                                                                 lizzieLet0_4MQNode_8_r,
                                                                                                 lizzieLet0_4MQNode_7_r,
                                                                                                 lizzieLet0_4MQNode_6_r,
                                                                                                 lizzieLet0_4MQNode_5_r,
                                                                                                 lizzieLet0_4MQNode_4_r,
                                                                                                 lizzieLet0_4MQNode_3_r,
                                                                                                 lizzieLet0_4MQNode_2_r,
                                                                                                 lizzieLet0_4MQNode_1_r}));
  assign lizzieLet0_4MQNode_r = (& lizzieLet0_4MQNode_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet0_4MQNode_emitted <= 9'd0;
    else
      lizzieLet0_4MQNode_emitted <= (lizzieLet0_4MQNode_r ? 9'd0 :
                                     lizzieLet0_4MQNode_done);
  
  /* destruct (Ty QTree_Bool,
          Dcon QNode_Bool) : (lizzieLet0_4MQNode_1QNode_Bool,QTree_Bool) > [(q1'a8n_destruct,Pointer_QTree_Bool),
                                                                            (q2'a8o_destruct,Pointer_QTree_Bool),
                                                                            (q3'a8p_destruct,Pointer_QTree_Bool),
                                                                            (q4'a8q_destruct,Pointer_QTree_Bool)] */
  logic [3:0] lizzieLet0_4MQNode_1QNode_Bool_emitted;
  logic [3:0] lizzieLet0_4MQNode_1QNode_Bool_done;
  assign \q1'a8n_destruct_d  = {lizzieLet0_4MQNode_1QNode_Bool_d[18:3],
                                (lizzieLet0_4MQNode_1QNode_Bool_d[0] && (! lizzieLet0_4MQNode_1QNode_Bool_emitted[0]))};
  assign \q2'a8o_destruct_d  = {lizzieLet0_4MQNode_1QNode_Bool_d[34:19],
                                (lizzieLet0_4MQNode_1QNode_Bool_d[0] && (! lizzieLet0_4MQNode_1QNode_Bool_emitted[1]))};
  assign \q3'a8p_destruct_d  = {lizzieLet0_4MQNode_1QNode_Bool_d[50:35],
                                (lizzieLet0_4MQNode_1QNode_Bool_d[0] && (! lizzieLet0_4MQNode_1QNode_Bool_emitted[2]))};
  assign \q4'a8q_destruct_d  = {lizzieLet0_4MQNode_1QNode_Bool_d[66:51],
                                (lizzieLet0_4MQNode_1QNode_Bool_d[0] && (! lizzieLet0_4MQNode_1QNode_Bool_emitted[3]))};
  assign lizzieLet0_4MQNode_1QNode_Bool_done = (lizzieLet0_4MQNode_1QNode_Bool_emitted | ({\q4'a8q_destruct_d [0],
                                                                                           \q3'a8p_destruct_d [0],
                                                                                           \q2'a8o_destruct_d [0],
                                                                                           \q1'a8n_destruct_d [0]} & {\q4'a8q_destruct_r ,
                                                                                                                      \q3'a8p_destruct_r ,
                                                                                                                      \q2'a8o_destruct_r ,
                                                                                                                      \q1'a8n_destruct_r }));
  assign lizzieLet0_4MQNode_1QNode_Bool_r = (& lizzieLet0_4MQNode_1QNode_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_1QNode_Bool_emitted <= 4'd0;
    else
      lizzieLet0_4MQNode_1QNode_Bool_emitted <= (lizzieLet0_4MQNode_1QNode_Bool_r ? 4'd0 :
                                                 lizzieLet0_4MQNode_1QNode_Bool_done);
  
  /* destruct (Ty QTree_Bool,
          Dcon QVal_Bool) : (lizzieLet0_4MQNode_1QVal_Bool,QTree_Bool) > [(v1a8h_destruct,MyBool)] */
  assign v1a8h_destruct_d = {lizzieLet0_4MQNode_1QVal_Bool_d[3:3],
                             lizzieLet0_4MQNode_1QVal_Bool_d[0]};
  assign lizzieLet0_4MQNode_1QVal_Bool_r = v1a8h_destruct_r;
  
  /* demux (Ty QTree_Bool,
       Ty QTree_Bool) : (lizzieLet0_4MQNode_2,QTree_Bool) (lizzieLet0_4MQNode_1,QTree_Bool) > [(_121,QTree_Bool),
                                                                                               (lizzieLet0_4MQNode_1QVal_Bool,QTree_Bool),
                                                                                               (lizzieLet0_4MQNode_1QNode_Bool,QTree_Bool),
                                                                                               (_120,QTree_Bool)] */
  logic [3:0] lizzieLet0_4MQNode_1_onehotd;
  always_comb
    if ((lizzieLet0_4MQNode_2_d[0] && lizzieLet0_4MQNode_1_d[0]))
      unique case (lizzieLet0_4MQNode_2_d[2:1])
        2'd0: lizzieLet0_4MQNode_1_onehotd = 4'd1;
        2'd1: lizzieLet0_4MQNode_1_onehotd = 4'd2;
        2'd2: lizzieLet0_4MQNode_1_onehotd = 4'd4;
        2'd3: lizzieLet0_4MQNode_1_onehotd = 4'd8;
        default: lizzieLet0_4MQNode_1_onehotd = 4'd0;
      endcase
    else lizzieLet0_4MQNode_1_onehotd = 4'd0;
  assign _121_d = {lizzieLet0_4MQNode_1_d[66:1],
                   lizzieLet0_4MQNode_1_onehotd[0]};
  assign lizzieLet0_4MQNode_1QVal_Bool_d = {lizzieLet0_4MQNode_1_d[66:1],
                                            lizzieLet0_4MQNode_1_onehotd[1]};
  assign lizzieLet0_4MQNode_1QNode_Bool_d = {lizzieLet0_4MQNode_1_d[66:1],
                                             lizzieLet0_4MQNode_1_onehotd[2]};
  assign _120_d = {lizzieLet0_4MQNode_1_d[66:1],
                   lizzieLet0_4MQNode_1_onehotd[3]};
  assign lizzieLet0_4MQNode_1_r = (| (lizzieLet0_4MQNode_1_onehotd & {_120_r,
                                                                      lizzieLet0_4MQNode_1QNode_Bool_r,
                                                                      lizzieLet0_4MQNode_1QVal_Bool_r,
                                                                      _121_r}));
  assign lizzieLet0_4MQNode_2_r = lizzieLet0_4MQNode_1_r;
  
  /* demux (Ty QTree_Bool,
       Ty Go) : (lizzieLet0_4MQNode_3,QTree_Bool) (lizzieLet0_3MQNode,Go) > [(lizzieLet0_4MQNode_3QNone_Bool,Go),
                                                                             (lizzieLet0_4MQNode_3QVal_Bool,Go),
                                                                             (lizzieLet0_4MQNode_3QNode_Bool,Go),
                                                                             (lizzieLet0_4MQNode_3QError_Bool,Go)] */
  logic [3:0] lizzieLet0_3MQNode_onehotd;
  always_comb
    if ((lizzieLet0_4MQNode_3_d[0] && lizzieLet0_3MQNode_d[0]))
      unique case (lizzieLet0_4MQNode_3_d[2:1])
        2'd0: lizzieLet0_3MQNode_onehotd = 4'd1;
        2'd1: lizzieLet0_3MQNode_onehotd = 4'd2;
        2'd2: lizzieLet0_3MQNode_onehotd = 4'd4;
        2'd3: lizzieLet0_3MQNode_onehotd = 4'd8;
        default: lizzieLet0_3MQNode_onehotd = 4'd0;
      endcase
    else lizzieLet0_3MQNode_onehotd = 4'd0;
  assign lizzieLet0_4MQNode_3QNone_Bool_d = lizzieLet0_3MQNode_onehotd[0];
  assign lizzieLet0_4MQNode_3QVal_Bool_d = lizzieLet0_3MQNode_onehotd[1];
  assign lizzieLet0_4MQNode_3QNode_Bool_d = lizzieLet0_3MQNode_onehotd[2];
  assign lizzieLet0_4MQNode_3QError_Bool_d = lizzieLet0_3MQNode_onehotd[3];
  assign lizzieLet0_3MQNode_r = (| (lizzieLet0_3MQNode_onehotd & {lizzieLet0_4MQNode_3QError_Bool_r,
                                                                  lizzieLet0_4MQNode_3QNode_Bool_r,
                                                                  lizzieLet0_4MQNode_3QVal_Bool_r,
                                                                  lizzieLet0_4MQNode_3QNone_Bool_r}));
  assign lizzieLet0_4MQNode_3_r = lizzieLet0_3MQNode_r;
  
  /* fork (Ty Go) : (lizzieLet0_4MQNode_3QError_Bool,Go) > [(lizzieLet0_4MQNode_3QError_Bool_1,Go),
                                                       (lizzieLet0_4MQNode_3QError_Bool_2,Go)] */
  logic [1:0] lizzieLet0_4MQNode_3QError_Bool_emitted;
  logic [1:0] lizzieLet0_4MQNode_3QError_Bool_done;
  assign lizzieLet0_4MQNode_3QError_Bool_1_d = (lizzieLet0_4MQNode_3QError_Bool_d[0] && (! lizzieLet0_4MQNode_3QError_Bool_emitted[0]));
  assign lizzieLet0_4MQNode_3QError_Bool_2_d = (lizzieLet0_4MQNode_3QError_Bool_d[0] && (! lizzieLet0_4MQNode_3QError_Bool_emitted[1]));
  assign lizzieLet0_4MQNode_3QError_Bool_done = (lizzieLet0_4MQNode_3QError_Bool_emitted | ({lizzieLet0_4MQNode_3QError_Bool_2_d[0],
                                                                                             lizzieLet0_4MQNode_3QError_Bool_1_d[0]} & {lizzieLet0_4MQNode_3QError_Bool_2_r,
                                                                                                                                        lizzieLet0_4MQNode_3QError_Bool_1_r}));
  assign lizzieLet0_4MQNode_3QError_Bool_r = (& lizzieLet0_4MQNode_3QError_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_3QError_Bool_emitted <= 2'd0;
    else
      lizzieLet0_4MQNode_3QError_Bool_emitted <= (lizzieLet0_4MQNode_3QError_Bool_r ? 2'd0 :
                                                  lizzieLet0_4MQNode_3QError_Bool_done);
  
  /* dcon (Ty QTree_Bool,
      Dcon QError_Bool) : [(lizzieLet0_4MQNode_3QError_Bool_1,Go)] > (lizzieLet0_4MQNode_3QError_Bool_1QError_Bool,QTree_Bool) */
  assign lizzieLet0_4MQNode_3QError_Bool_1QError_Bool_d = QError_Bool_dc((& {lizzieLet0_4MQNode_3QError_Bool_1_d[0]}), lizzieLet0_4MQNode_3QError_Bool_1_d);
  assign {lizzieLet0_4MQNode_3QError_Bool_1_r} = {1 {(lizzieLet0_4MQNode_3QError_Bool_1QError_Bool_r && lizzieLet0_4MQNode_3QError_Bool_1QError_Bool_d[0])}};
  
  /* buf (Ty QTree_Bool) : (lizzieLet0_4MQNode_3QError_Bool_1QError_Bool,QTree_Bool) > (lizzieLet19_2_1_argbuf,QTree_Bool) */
  QTree_Bool_t lizzieLet0_4MQNode_3QError_Bool_1QError_Bool_bufchan_d;
  logic lizzieLet0_4MQNode_3QError_Bool_1QError_Bool_bufchan_r;
  assign lizzieLet0_4MQNode_3QError_Bool_1QError_Bool_r = ((! lizzieLet0_4MQNode_3QError_Bool_1QError_Bool_bufchan_d[0]) || lizzieLet0_4MQNode_3QError_Bool_1QError_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_3QError_Bool_1QError_Bool_bufchan_d <= {66'd0,
                                                                 1'd0};
    else
      if (lizzieLet0_4MQNode_3QError_Bool_1QError_Bool_r)
        lizzieLet0_4MQNode_3QError_Bool_1QError_Bool_bufchan_d <= lizzieLet0_4MQNode_3QError_Bool_1QError_Bool_d;
  QTree_Bool_t lizzieLet0_4MQNode_3QError_Bool_1QError_Bool_bufchan_buf;
  assign lizzieLet0_4MQNode_3QError_Bool_1QError_Bool_bufchan_r = (! lizzieLet0_4MQNode_3QError_Bool_1QError_Bool_bufchan_buf[0]);
  assign lizzieLet19_2_1_argbuf_d = (lizzieLet0_4MQNode_3QError_Bool_1QError_Bool_bufchan_buf[0] ? lizzieLet0_4MQNode_3QError_Bool_1QError_Bool_bufchan_buf :
                                     lizzieLet0_4MQNode_3QError_Bool_1QError_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_3QError_Bool_1QError_Bool_bufchan_buf <= {66'd0,
                                                                   1'd0};
    else
      if ((lizzieLet19_2_1_argbuf_r && lizzieLet0_4MQNode_3QError_Bool_1QError_Bool_bufchan_buf[0]))
        lizzieLet0_4MQNode_3QError_Bool_1QError_Bool_bufchan_buf <= {66'd0,
                                                                     1'd0};
      else if (((! lizzieLet19_2_1_argbuf_r) && (! lizzieLet0_4MQNode_3QError_Bool_1QError_Bool_bufchan_buf[0])))
        lizzieLet0_4MQNode_3QError_Bool_1QError_Bool_bufchan_buf <= lizzieLet0_4MQNode_3QError_Bool_1QError_Bool_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet0_4MQNode_3QError_Bool_2,Go) > (lizzieLet0_4MQNode_3QError_Bool_2_argbuf,Go) */
  Go_t lizzieLet0_4MQNode_3QError_Bool_2_bufchan_d;
  logic lizzieLet0_4MQNode_3QError_Bool_2_bufchan_r;
  assign lizzieLet0_4MQNode_3QError_Bool_2_r = ((! lizzieLet0_4MQNode_3QError_Bool_2_bufchan_d[0]) || lizzieLet0_4MQNode_3QError_Bool_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_3QError_Bool_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet0_4MQNode_3QError_Bool_2_r)
        lizzieLet0_4MQNode_3QError_Bool_2_bufchan_d <= lizzieLet0_4MQNode_3QError_Bool_2_d;
  Go_t lizzieLet0_4MQNode_3QError_Bool_2_bufchan_buf;
  assign lizzieLet0_4MQNode_3QError_Bool_2_bufchan_r = (! lizzieLet0_4MQNode_3QError_Bool_2_bufchan_buf[0]);
  assign lizzieLet0_4MQNode_3QError_Bool_2_argbuf_d = (lizzieLet0_4MQNode_3QError_Bool_2_bufchan_buf[0] ? lizzieLet0_4MQNode_3QError_Bool_2_bufchan_buf :
                                                       lizzieLet0_4MQNode_3QError_Bool_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_3QError_Bool_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet0_4MQNode_3QError_Bool_2_argbuf_r && lizzieLet0_4MQNode_3QError_Bool_2_bufchan_buf[0]))
        lizzieLet0_4MQNode_3QError_Bool_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet0_4MQNode_3QError_Bool_2_argbuf_r) && (! lizzieLet0_4MQNode_3QError_Bool_2_bufchan_buf[0])))
        lizzieLet0_4MQNode_3QError_Bool_2_bufchan_buf <= lizzieLet0_4MQNode_3QError_Bool_2_bufchan_d;
  
  /* demux (Ty QTree_Bool,
       Ty QTree_Bool) : (lizzieLet0_4MQNode_4,QTree_Bool) (lizzieLet0_5MQNode,QTree_Bool) > [(lizzieLet0_4MQNode_4QNone_Bool,QTree_Bool),
                                                                                             (lizzieLet0_4MQNode_4QVal_Bool,QTree_Bool),
                                                                                             (lizzieLet0_4MQNode_4QNode_Bool,QTree_Bool),
                                                                                             (_119,QTree_Bool)] */
  logic [3:0] lizzieLet0_5MQNode_onehotd;
  always_comb
    if ((lizzieLet0_4MQNode_4_d[0] && lizzieLet0_5MQNode_d[0]))
      unique case (lizzieLet0_4MQNode_4_d[2:1])
        2'd0: lizzieLet0_5MQNode_onehotd = 4'd1;
        2'd1: lizzieLet0_5MQNode_onehotd = 4'd2;
        2'd2: lizzieLet0_5MQNode_onehotd = 4'd4;
        2'd3: lizzieLet0_5MQNode_onehotd = 4'd8;
        default: lizzieLet0_5MQNode_onehotd = 4'd0;
      endcase
    else lizzieLet0_5MQNode_onehotd = 4'd0;
  assign lizzieLet0_4MQNode_4QNone_Bool_d = {lizzieLet0_5MQNode_d[66:1],
                                             lizzieLet0_5MQNode_onehotd[0]};
  assign lizzieLet0_4MQNode_4QVal_Bool_d = {lizzieLet0_5MQNode_d[66:1],
                                            lizzieLet0_5MQNode_onehotd[1]};
  assign lizzieLet0_4MQNode_4QNode_Bool_d = {lizzieLet0_5MQNode_d[66:1],
                                             lizzieLet0_5MQNode_onehotd[2]};
  assign _119_d = {lizzieLet0_5MQNode_d[66:1],
                   lizzieLet0_5MQNode_onehotd[3]};
  assign lizzieLet0_5MQNode_r = (| (lizzieLet0_5MQNode_onehotd & {_119_r,
                                                                  lizzieLet0_4MQNode_4QNode_Bool_r,
                                                                  lizzieLet0_4MQNode_4QVal_Bool_r,
                                                                  lizzieLet0_4MQNode_4QNone_Bool_r}));
  assign lizzieLet0_4MQNode_4_r = lizzieLet0_5MQNode_r;
  
  /* fork (Ty QTree_Bool) : (lizzieLet0_4MQNode_4QNode_Bool,QTree_Bool) > [(lizzieLet0_4MQNode_4QNode_Bool_1,QTree_Bool),
                                                                      (lizzieLet0_4MQNode_4QNode_Bool_2,QTree_Bool),
                                                                      (lizzieLet0_4MQNode_4QNode_Bool_3,QTree_Bool),
                                                                      (lizzieLet0_4MQNode_4QNode_Bool_4,QTree_Bool),
                                                                      (lizzieLet0_4MQNode_4QNode_Bool_5,QTree_Bool),
                                                                      (lizzieLet0_4MQNode_4QNode_Bool_6,QTree_Bool),
                                                                      (lizzieLet0_4MQNode_4QNode_Bool_7,QTree_Bool),
                                                                      (lizzieLet0_4MQNode_4QNode_Bool_8,QTree_Bool),
                                                                      (lizzieLet0_4MQNode_4QNode_Bool_9,QTree_Bool),
                                                                      (lizzieLet0_4MQNode_4QNode_Bool_10,QTree_Bool),
                                                                      (lizzieLet0_4MQNode_4QNode_Bool_11,QTree_Bool),
                                                                      (lizzieLet0_4MQNode_4QNode_Bool_12,QTree_Bool)] */
  logic [11:0] lizzieLet0_4MQNode_4QNode_Bool_emitted;
  logic [11:0] lizzieLet0_4MQNode_4QNode_Bool_done;
  assign lizzieLet0_4MQNode_4QNode_Bool_1_d = {lizzieLet0_4MQNode_4QNode_Bool_d[66:1],
                                               (lizzieLet0_4MQNode_4QNode_Bool_d[0] && (! lizzieLet0_4MQNode_4QNode_Bool_emitted[0]))};
  assign lizzieLet0_4MQNode_4QNode_Bool_2_d = {lizzieLet0_4MQNode_4QNode_Bool_d[66:1],
                                               (lizzieLet0_4MQNode_4QNode_Bool_d[0] && (! lizzieLet0_4MQNode_4QNode_Bool_emitted[1]))};
  assign lizzieLet0_4MQNode_4QNode_Bool_3_d = {lizzieLet0_4MQNode_4QNode_Bool_d[66:1],
                                               (lizzieLet0_4MQNode_4QNode_Bool_d[0] && (! lizzieLet0_4MQNode_4QNode_Bool_emitted[2]))};
  assign lizzieLet0_4MQNode_4QNode_Bool_4_d = {lizzieLet0_4MQNode_4QNode_Bool_d[66:1],
                                               (lizzieLet0_4MQNode_4QNode_Bool_d[0] && (! lizzieLet0_4MQNode_4QNode_Bool_emitted[3]))};
  assign lizzieLet0_4MQNode_4QNode_Bool_5_d = {lizzieLet0_4MQNode_4QNode_Bool_d[66:1],
                                               (lizzieLet0_4MQNode_4QNode_Bool_d[0] && (! lizzieLet0_4MQNode_4QNode_Bool_emitted[4]))};
  assign lizzieLet0_4MQNode_4QNode_Bool_6_d = {lizzieLet0_4MQNode_4QNode_Bool_d[66:1],
                                               (lizzieLet0_4MQNode_4QNode_Bool_d[0] && (! lizzieLet0_4MQNode_4QNode_Bool_emitted[5]))};
  assign lizzieLet0_4MQNode_4QNode_Bool_7_d = {lizzieLet0_4MQNode_4QNode_Bool_d[66:1],
                                               (lizzieLet0_4MQNode_4QNode_Bool_d[0] && (! lizzieLet0_4MQNode_4QNode_Bool_emitted[6]))};
  assign lizzieLet0_4MQNode_4QNode_Bool_8_d = {lizzieLet0_4MQNode_4QNode_Bool_d[66:1],
                                               (lizzieLet0_4MQNode_4QNode_Bool_d[0] && (! lizzieLet0_4MQNode_4QNode_Bool_emitted[7]))};
  assign lizzieLet0_4MQNode_4QNode_Bool_9_d = {lizzieLet0_4MQNode_4QNode_Bool_d[66:1],
                                               (lizzieLet0_4MQNode_4QNode_Bool_d[0] && (! lizzieLet0_4MQNode_4QNode_Bool_emitted[8]))};
  assign lizzieLet0_4MQNode_4QNode_Bool_10_d = {lizzieLet0_4MQNode_4QNode_Bool_d[66:1],
                                                (lizzieLet0_4MQNode_4QNode_Bool_d[0] && (! lizzieLet0_4MQNode_4QNode_Bool_emitted[9]))};
  assign lizzieLet0_4MQNode_4QNode_Bool_11_d = {lizzieLet0_4MQNode_4QNode_Bool_d[66:1],
                                                (lizzieLet0_4MQNode_4QNode_Bool_d[0] && (! lizzieLet0_4MQNode_4QNode_Bool_emitted[10]))};
  assign lizzieLet0_4MQNode_4QNode_Bool_12_d = {lizzieLet0_4MQNode_4QNode_Bool_d[66:1],
                                                (lizzieLet0_4MQNode_4QNode_Bool_d[0] && (! lizzieLet0_4MQNode_4QNode_Bool_emitted[11]))};
  assign lizzieLet0_4MQNode_4QNode_Bool_done = (lizzieLet0_4MQNode_4QNode_Bool_emitted | ({lizzieLet0_4MQNode_4QNode_Bool_12_d[0],
                                                                                           lizzieLet0_4MQNode_4QNode_Bool_11_d[0],
                                                                                           lizzieLet0_4MQNode_4QNode_Bool_10_d[0],
                                                                                           lizzieLet0_4MQNode_4QNode_Bool_9_d[0],
                                                                                           lizzieLet0_4MQNode_4QNode_Bool_8_d[0],
                                                                                           lizzieLet0_4MQNode_4QNode_Bool_7_d[0],
                                                                                           lizzieLet0_4MQNode_4QNode_Bool_6_d[0],
                                                                                           lizzieLet0_4MQNode_4QNode_Bool_5_d[0],
                                                                                           lizzieLet0_4MQNode_4QNode_Bool_4_d[0],
                                                                                           lizzieLet0_4MQNode_4QNode_Bool_3_d[0],
                                                                                           lizzieLet0_4MQNode_4QNode_Bool_2_d[0],
                                                                                           lizzieLet0_4MQNode_4QNode_Bool_1_d[0]} & {lizzieLet0_4MQNode_4QNode_Bool_12_r,
                                                                                                                                     lizzieLet0_4MQNode_4QNode_Bool_11_r,
                                                                                                                                     lizzieLet0_4MQNode_4QNode_Bool_10_r,
                                                                                                                                     lizzieLet0_4MQNode_4QNode_Bool_9_r,
                                                                                                                                     lizzieLet0_4MQNode_4QNode_Bool_8_r,
                                                                                                                                     lizzieLet0_4MQNode_4QNode_Bool_7_r,
                                                                                                                                     lizzieLet0_4MQNode_4QNode_Bool_6_r,
                                                                                                                                     lizzieLet0_4MQNode_4QNode_Bool_5_r,
                                                                                                                                     lizzieLet0_4MQNode_4QNode_Bool_4_r,
                                                                                                                                     lizzieLet0_4MQNode_4QNode_Bool_3_r,
                                                                                                                                     lizzieLet0_4MQNode_4QNode_Bool_2_r,
                                                                                                                                     lizzieLet0_4MQNode_4QNode_Bool_1_r}));
  assign lizzieLet0_4MQNode_4QNode_Bool_r = (& lizzieLet0_4MQNode_4QNode_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QNode_Bool_emitted <= 12'd0;
    else
      lizzieLet0_4MQNode_4QNode_Bool_emitted <= (lizzieLet0_4MQNode_4QNode_Bool_r ? 12'd0 :
                                                 lizzieLet0_4MQNode_4QNode_Bool_done);
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_QTree_Bool) : (lizzieLet0_4MQNode_4QNode_Bool_10,QTree_Bool) (q2'a8o_destruct,Pointer_QTree_Bool) > [(lizzieLet0_4MQNode_4QNode_Bool_10QNone_Bool,Pointer_QTree_Bool),
                                                                                                                       (_118,Pointer_QTree_Bool),
                                                                                                                       (lizzieLet0_4MQNode_4QNode_Bool_10QNode_Bool,Pointer_QTree_Bool),
                                                                                                                       (_117,Pointer_QTree_Bool)] */
  logic [3:0] \q2'a8o_destruct_onehotd ;
  always_comb
    if ((lizzieLet0_4MQNode_4QNode_Bool_10_d[0] && \q2'a8o_destruct_d [0]))
      unique case (lizzieLet0_4MQNode_4QNode_Bool_10_d[2:1])
        2'd0: \q2'a8o_destruct_onehotd  = 4'd1;
        2'd1: \q2'a8o_destruct_onehotd  = 4'd2;
        2'd2: \q2'a8o_destruct_onehotd  = 4'd4;
        2'd3: \q2'a8o_destruct_onehotd  = 4'd8;
        default: \q2'a8o_destruct_onehotd  = 4'd0;
      endcase
    else \q2'a8o_destruct_onehotd  = 4'd0;
  assign lizzieLet0_4MQNode_4QNode_Bool_10QNone_Bool_d = {\q2'a8o_destruct_d [16:1],
                                                          \q2'a8o_destruct_onehotd [0]};
  assign _118_d = {\q2'a8o_destruct_d [16:1],
                   \q2'a8o_destruct_onehotd [1]};
  assign lizzieLet0_4MQNode_4QNode_Bool_10QNode_Bool_d = {\q2'a8o_destruct_d [16:1],
                                                          \q2'a8o_destruct_onehotd [2]};
  assign _117_d = {\q2'a8o_destruct_d [16:1],
                   \q2'a8o_destruct_onehotd [3]};
  assign \q2'a8o_destruct_r  = (| (\q2'a8o_destruct_onehotd  & {_117_r,
                                                                lizzieLet0_4MQNode_4QNode_Bool_10QNode_Bool_r,
                                                                _118_r,
                                                                lizzieLet0_4MQNode_4QNode_Bool_10QNone_Bool_r}));
  assign lizzieLet0_4MQNode_4QNode_Bool_10_r = \q2'a8o_destruct_r ;
  
  /* buf (Ty Pointer_QTree_Bool) : (lizzieLet0_4MQNode_4QNode_Bool_10QNone_Bool,Pointer_QTree_Bool) > (lizzieLet0_4MQNode_4QNode_Bool_10QNone_Bool_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t lizzieLet0_4MQNode_4QNode_Bool_10QNone_Bool_bufchan_d;
  logic lizzieLet0_4MQNode_4QNode_Bool_10QNone_Bool_bufchan_r;
  assign lizzieLet0_4MQNode_4QNode_Bool_10QNone_Bool_r = ((! lizzieLet0_4MQNode_4QNode_Bool_10QNone_Bool_bufchan_d[0]) || lizzieLet0_4MQNode_4QNode_Bool_10QNone_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QNode_Bool_10QNone_Bool_bufchan_d <= {16'd0,
                                                                1'd0};
    else
      if (lizzieLet0_4MQNode_4QNode_Bool_10QNone_Bool_r)
        lizzieLet0_4MQNode_4QNode_Bool_10QNone_Bool_bufchan_d <= lizzieLet0_4MQNode_4QNode_Bool_10QNone_Bool_d;
  Pointer_QTree_Bool_t lizzieLet0_4MQNode_4QNode_Bool_10QNone_Bool_bufchan_buf;
  assign lizzieLet0_4MQNode_4QNode_Bool_10QNone_Bool_bufchan_r = (! lizzieLet0_4MQNode_4QNode_Bool_10QNone_Bool_bufchan_buf[0]);
  assign lizzieLet0_4MQNode_4QNode_Bool_10QNone_Bool_1_argbuf_d = (lizzieLet0_4MQNode_4QNode_Bool_10QNone_Bool_bufchan_buf[0] ? lizzieLet0_4MQNode_4QNode_Bool_10QNone_Bool_bufchan_buf :
                                                                   lizzieLet0_4MQNode_4QNode_Bool_10QNone_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QNode_Bool_10QNone_Bool_bufchan_buf <= {16'd0,
                                                                  1'd0};
    else
      if ((lizzieLet0_4MQNode_4QNode_Bool_10QNone_Bool_1_argbuf_r && lizzieLet0_4MQNode_4QNode_Bool_10QNone_Bool_bufchan_buf[0]))
        lizzieLet0_4MQNode_4QNode_Bool_10QNone_Bool_bufchan_buf <= {16'd0,
                                                                    1'd0};
      else if (((! lizzieLet0_4MQNode_4QNode_Bool_10QNone_Bool_1_argbuf_r) && (! lizzieLet0_4MQNode_4QNode_Bool_10QNone_Bool_bufchan_buf[0])))
        lizzieLet0_4MQNode_4QNode_Bool_10QNone_Bool_bufchan_buf <= lizzieLet0_4MQNode_4QNode_Bool_10QNone_Bool_bufchan_d;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_QTree_Bool) : (lizzieLet0_4MQNode_4QNode_Bool_11,QTree_Bool) (q3'a8p_destruct,Pointer_QTree_Bool) > [(lizzieLet0_4MQNode_4QNode_Bool_11QNone_Bool,Pointer_QTree_Bool),
                                                                                                                       (_116,Pointer_QTree_Bool),
                                                                                                                       (lizzieLet0_4MQNode_4QNode_Bool_11QNode_Bool,Pointer_QTree_Bool),
                                                                                                                       (_115,Pointer_QTree_Bool)] */
  logic [3:0] \q3'a8p_destruct_onehotd ;
  always_comb
    if ((lizzieLet0_4MQNode_4QNode_Bool_11_d[0] && \q3'a8p_destruct_d [0]))
      unique case (lizzieLet0_4MQNode_4QNode_Bool_11_d[2:1])
        2'd0: \q3'a8p_destruct_onehotd  = 4'd1;
        2'd1: \q3'a8p_destruct_onehotd  = 4'd2;
        2'd2: \q3'a8p_destruct_onehotd  = 4'd4;
        2'd3: \q3'a8p_destruct_onehotd  = 4'd8;
        default: \q3'a8p_destruct_onehotd  = 4'd0;
      endcase
    else \q3'a8p_destruct_onehotd  = 4'd0;
  assign lizzieLet0_4MQNode_4QNode_Bool_11QNone_Bool_d = {\q3'a8p_destruct_d [16:1],
                                                          \q3'a8p_destruct_onehotd [0]};
  assign _116_d = {\q3'a8p_destruct_d [16:1],
                   \q3'a8p_destruct_onehotd [1]};
  assign lizzieLet0_4MQNode_4QNode_Bool_11QNode_Bool_d = {\q3'a8p_destruct_d [16:1],
                                                          \q3'a8p_destruct_onehotd [2]};
  assign _115_d = {\q3'a8p_destruct_d [16:1],
                   \q3'a8p_destruct_onehotd [3]};
  assign \q3'a8p_destruct_r  = (| (\q3'a8p_destruct_onehotd  & {_115_r,
                                                                lizzieLet0_4MQNode_4QNode_Bool_11QNode_Bool_r,
                                                                _116_r,
                                                                lizzieLet0_4MQNode_4QNode_Bool_11QNone_Bool_r}));
  assign lizzieLet0_4MQNode_4QNode_Bool_11_r = \q3'a8p_destruct_r ;
  
  /* buf (Ty Pointer_QTree_Bool) : (lizzieLet0_4MQNode_4QNode_Bool_11QNone_Bool,Pointer_QTree_Bool) > (lizzieLet0_4MQNode_4QNode_Bool_11QNone_Bool_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t lizzieLet0_4MQNode_4QNode_Bool_11QNone_Bool_bufchan_d;
  logic lizzieLet0_4MQNode_4QNode_Bool_11QNone_Bool_bufchan_r;
  assign lizzieLet0_4MQNode_4QNode_Bool_11QNone_Bool_r = ((! lizzieLet0_4MQNode_4QNode_Bool_11QNone_Bool_bufchan_d[0]) || lizzieLet0_4MQNode_4QNode_Bool_11QNone_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QNode_Bool_11QNone_Bool_bufchan_d <= {16'd0,
                                                                1'd0};
    else
      if (lizzieLet0_4MQNode_4QNode_Bool_11QNone_Bool_r)
        lizzieLet0_4MQNode_4QNode_Bool_11QNone_Bool_bufchan_d <= lizzieLet0_4MQNode_4QNode_Bool_11QNone_Bool_d;
  Pointer_QTree_Bool_t lizzieLet0_4MQNode_4QNode_Bool_11QNone_Bool_bufchan_buf;
  assign lizzieLet0_4MQNode_4QNode_Bool_11QNone_Bool_bufchan_r = (! lizzieLet0_4MQNode_4QNode_Bool_11QNone_Bool_bufchan_buf[0]);
  assign lizzieLet0_4MQNode_4QNode_Bool_11QNone_Bool_1_argbuf_d = (lizzieLet0_4MQNode_4QNode_Bool_11QNone_Bool_bufchan_buf[0] ? lizzieLet0_4MQNode_4QNode_Bool_11QNone_Bool_bufchan_buf :
                                                                   lizzieLet0_4MQNode_4QNode_Bool_11QNone_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QNode_Bool_11QNone_Bool_bufchan_buf <= {16'd0,
                                                                  1'd0};
    else
      if ((lizzieLet0_4MQNode_4QNode_Bool_11QNone_Bool_1_argbuf_r && lizzieLet0_4MQNode_4QNode_Bool_11QNone_Bool_bufchan_buf[0]))
        lizzieLet0_4MQNode_4QNode_Bool_11QNone_Bool_bufchan_buf <= {16'd0,
                                                                    1'd0};
      else if (((! lizzieLet0_4MQNode_4QNode_Bool_11QNone_Bool_1_argbuf_r) && (! lizzieLet0_4MQNode_4QNode_Bool_11QNone_Bool_bufchan_buf[0])))
        lizzieLet0_4MQNode_4QNode_Bool_11QNone_Bool_bufchan_buf <= lizzieLet0_4MQNode_4QNode_Bool_11QNone_Bool_bufchan_d;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_QTree_Bool) : (lizzieLet0_4MQNode_4QNode_Bool_12,QTree_Bool) (q4'a8q_destruct,Pointer_QTree_Bool) > [(lizzieLet0_4MQNode_4QNode_Bool_12QNone_Bool,Pointer_QTree_Bool),
                                                                                                                       (_114,Pointer_QTree_Bool),
                                                                                                                       (lizzieLet0_4MQNode_4QNode_Bool_12QNode_Bool,Pointer_QTree_Bool),
                                                                                                                       (_113,Pointer_QTree_Bool)] */
  logic [3:0] \q4'a8q_destruct_onehotd ;
  always_comb
    if ((lizzieLet0_4MQNode_4QNode_Bool_12_d[0] && \q4'a8q_destruct_d [0]))
      unique case (lizzieLet0_4MQNode_4QNode_Bool_12_d[2:1])
        2'd0: \q4'a8q_destruct_onehotd  = 4'd1;
        2'd1: \q4'a8q_destruct_onehotd  = 4'd2;
        2'd2: \q4'a8q_destruct_onehotd  = 4'd4;
        2'd3: \q4'a8q_destruct_onehotd  = 4'd8;
        default: \q4'a8q_destruct_onehotd  = 4'd0;
      endcase
    else \q4'a8q_destruct_onehotd  = 4'd0;
  assign lizzieLet0_4MQNode_4QNode_Bool_12QNone_Bool_d = {\q4'a8q_destruct_d [16:1],
                                                          \q4'a8q_destruct_onehotd [0]};
  assign _114_d = {\q4'a8q_destruct_d [16:1],
                   \q4'a8q_destruct_onehotd [1]};
  assign lizzieLet0_4MQNode_4QNode_Bool_12QNode_Bool_d = {\q4'a8q_destruct_d [16:1],
                                                          \q4'a8q_destruct_onehotd [2]};
  assign _113_d = {\q4'a8q_destruct_d [16:1],
                   \q4'a8q_destruct_onehotd [3]};
  assign \q4'a8q_destruct_r  = (| (\q4'a8q_destruct_onehotd  & {_113_r,
                                                                lizzieLet0_4MQNode_4QNode_Bool_12QNode_Bool_r,
                                                                _114_r,
                                                                lizzieLet0_4MQNode_4QNode_Bool_12QNone_Bool_r}));
  assign lizzieLet0_4MQNode_4QNode_Bool_12_r = \q4'a8q_destruct_r ;
  
  /* buf (Ty Pointer_QTree_Bool) : (lizzieLet0_4MQNode_4QNode_Bool_12QNode_Bool,Pointer_QTree_Bool) > (lizzieLet0_4MQNode_4QNode_Bool_12QNode_Bool_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t lizzieLet0_4MQNode_4QNode_Bool_12QNode_Bool_bufchan_d;
  logic lizzieLet0_4MQNode_4QNode_Bool_12QNode_Bool_bufchan_r;
  assign lizzieLet0_4MQNode_4QNode_Bool_12QNode_Bool_r = ((! lizzieLet0_4MQNode_4QNode_Bool_12QNode_Bool_bufchan_d[0]) || lizzieLet0_4MQNode_4QNode_Bool_12QNode_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QNode_Bool_12QNode_Bool_bufchan_d <= {16'd0,
                                                                1'd0};
    else
      if (lizzieLet0_4MQNode_4QNode_Bool_12QNode_Bool_r)
        lizzieLet0_4MQNode_4QNode_Bool_12QNode_Bool_bufchan_d <= lizzieLet0_4MQNode_4QNode_Bool_12QNode_Bool_d;
  Pointer_QTree_Bool_t lizzieLet0_4MQNode_4QNode_Bool_12QNode_Bool_bufchan_buf;
  assign lizzieLet0_4MQNode_4QNode_Bool_12QNode_Bool_bufchan_r = (! lizzieLet0_4MQNode_4QNode_Bool_12QNode_Bool_bufchan_buf[0]);
  assign lizzieLet0_4MQNode_4QNode_Bool_12QNode_Bool_1_argbuf_d = (lizzieLet0_4MQNode_4QNode_Bool_12QNode_Bool_bufchan_buf[0] ? lizzieLet0_4MQNode_4QNode_Bool_12QNode_Bool_bufchan_buf :
                                                                   lizzieLet0_4MQNode_4QNode_Bool_12QNode_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QNode_Bool_12QNode_Bool_bufchan_buf <= {16'd0,
                                                                  1'd0};
    else
      if ((lizzieLet0_4MQNode_4QNode_Bool_12QNode_Bool_1_argbuf_r && lizzieLet0_4MQNode_4QNode_Bool_12QNode_Bool_bufchan_buf[0]))
        lizzieLet0_4MQNode_4QNode_Bool_12QNode_Bool_bufchan_buf <= {16'd0,
                                                                    1'd0};
      else if (((! lizzieLet0_4MQNode_4QNode_Bool_12QNode_Bool_1_argbuf_r) && (! lizzieLet0_4MQNode_4QNode_Bool_12QNode_Bool_bufchan_buf[0])))
        lizzieLet0_4MQNode_4QNode_Bool_12QNode_Bool_bufchan_buf <= lizzieLet0_4MQNode_4QNode_Bool_12QNode_Bool_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (lizzieLet0_4MQNode_4QNode_Bool_12QNone_Bool,Pointer_QTree_Bool) > (lizzieLet0_4MQNode_4QNode_Bool_12QNone_Bool_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t lizzieLet0_4MQNode_4QNode_Bool_12QNone_Bool_bufchan_d;
  logic lizzieLet0_4MQNode_4QNode_Bool_12QNone_Bool_bufchan_r;
  assign lizzieLet0_4MQNode_4QNode_Bool_12QNone_Bool_r = ((! lizzieLet0_4MQNode_4QNode_Bool_12QNone_Bool_bufchan_d[0]) || lizzieLet0_4MQNode_4QNode_Bool_12QNone_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QNode_Bool_12QNone_Bool_bufchan_d <= {16'd0,
                                                                1'd0};
    else
      if (lizzieLet0_4MQNode_4QNode_Bool_12QNone_Bool_r)
        lizzieLet0_4MQNode_4QNode_Bool_12QNone_Bool_bufchan_d <= lizzieLet0_4MQNode_4QNode_Bool_12QNone_Bool_d;
  Pointer_QTree_Bool_t lizzieLet0_4MQNode_4QNode_Bool_12QNone_Bool_bufchan_buf;
  assign lizzieLet0_4MQNode_4QNode_Bool_12QNone_Bool_bufchan_r = (! lizzieLet0_4MQNode_4QNode_Bool_12QNone_Bool_bufchan_buf[0]);
  assign lizzieLet0_4MQNode_4QNode_Bool_12QNone_Bool_1_argbuf_d = (lizzieLet0_4MQNode_4QNode_Bool_12QNone_Bool_bufchan_buf[0] ? lizzieLet0_4MQNode_4QNode_Bool_12QNone_Bool_bufchan_buf :
                                                                   lizzieLet0_4MQNode_4QNode_Bool_12QNone_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QNode_Bool_12QNone_Bool_bufchan_buf <= {16'd0,
                                                                  1'd0};
    else
      if ((lizzieLet0_4MQNode_4QNode_Bool_12QNone_Bool_1_argbuf_r && lizzieLet0_4MQNode_4QNode_Bool_12QNone_Bool_bufchan_buf[0]))
        lizzieLet0_4MQNode_4QNode_Bool_12QNone_Bool_bufchan_buf <= {16'd0,
                                                                    1'd0};
      else if (((! lizzieLet0_4MQNode_4QNode_Bool_12QNone_Bool_1_argbuf_r) && (! lizzieLet0_4MQNode_4QNode_Bool_12QNone_Bool_bufchan_buf[0])))
        lizzieLet0_4MQNode_4QNode_Bool_12QNone_Bool_bufchan_buf <= lizzieLet0_4MQNode_4QNode_Bool_12QNone_Bool_bufchan_d;
  
  /* destruct (Ty QTree_Bool,
          Dcon QNode_Bool) : (lizzieLet0_4MQNode_4QNode_Bool_1QNode_Bool,QTree_Bool) > [(t1a8s_destruct,Pointer_QTree_Bool),
                                                                                        (t2a8t_destruct,Pointer_QTree_Bool),
                                                                                        (t3a8u_destruct,Pointer_QTree_Bool),
                                                                                        (t4a8v_destruct,Pointer_QTree_Bool)] */
  logic [3:0] lizzieLet0_4MQNode_4QNode_Bool_1QNode_Bool_emitted;
  logic [3:0] lizzieLet0_4MQNode_4QNode_Bool_1QNode_Bool_done;
  assign t1a8s_destruct_d = {lizzieLet0_4MQNode_4QNode_Bool_1QNode_Bool_d[18:3],
                             (lizzieLet0_4MQNode_4QNode_Bool_1QNode_Bool_d[0] && (! lizzieLet0_4MQNode_4QNode_Bool_1QNode_Bool_emitted[0]))};
  assign t2a8t_destruct_d = {lizzieLet0_4MQNode_4QNode_Bool_1QNode_Bool_d[34:19],
                             (lizzieLet0_4MQNode_4QNode_Bool_1QNode_Bool_d[0] && (! lizzieLet0_4MQNode_4QNode_Bool_1QNode_Bool_emitted[1]))};
  assign t3a8u_destruct_d = {lizzieLet0_4MQNode_4QNode_Bool_1QNode_Bool_d[50:35],
                             (lizzieLet0_4MQNode_4QNode_Bool_1QNode_Bool_d[0] && (! lizzieLet0_4MQNode_4QNode_Bool_1QNode_Bool_emitted[2]))};
  assign t4a8v_destruct_d = {lizzieLet0_4MQNode_4QNode_Bool_1QNode_Bool_d[66:51],
                             (lizzieLet0_4MQNode_4QNode_Bool_1QNode_Bool_d[0] && (! lizzieLet0_4MQNode_4QNode_Bool_1QNode_Bool_emitted[3]))};
  assign lizzieLet0_4MQNode_4QNode_Bool_1QNode_Bool_done = (lizzieLet0_4MQNode_4QNode_Bool_1QNode_Bool_emitted | ({t4a8v_destruct_d[0],
                                                                                                                   t3a8u_destruct_d[0],
                                                                                                                   t2a8t_destruct_d[0],
                                                                                                                   t1a8s_destruct_d[0]} & {t4a8v_destruct_r,
                                                                                                                                           t3a8u_destruct_r,
                                                                                                                                           t2a8t_destruct_r,
                                                                                                                                           t1a8s_destruct_r}));
  assign lizzieLet0_4MQNode_4QNode_Bool_1QNode_Bool_r = (& lizzieLet0_4MQNode_4QNode_Bool_1QNode_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QNode_Bool_1QNode_Bool_emitted <= 4'd0;
    else
      lizzieLet0_4MQNode_4QNode_Bool_1QNode_Bool_emitted <= (lizzieLet0_4MQNode_4QNode_Bool_1QNode_Bool_r ? 4'd0 :
                                                             lizzieLet0_4MQNode_4QNode_Bool_1QNode_Bool_done);
  
  /* demux (Ty QTree_Bool,
       Ty QTree_Bool) : (lizzieLet0_4MQNode_4QNode_Bool_2,QTree_Bool) (lizzieLet0_4MQNode_4QNode_Bool_1,QTree_Bool) > [(_112,QTree_Bool),
                                                                                                                       (_111,QTree_Bool),
                                                                                                                       (lizzieLet0_4MQNode_4QNode_Bool_1QNode_Bool,QTree_Bool),
                                                                                                                       (_110,QTree_Bool)] */
  logic [3:0] lizzieLet0_4MQNode_4QNode_Bool_1_onehotd;
  always_comb
    if ((lizzieLet0_4MQNode_4QNode_Bool_2_d[0] && lizzieLet0_4MQNode_4QNode_Bool_1_d[0]))
      unique case (lizzieLet0_4MQNode_4QNode_Bool_2_d[2:1])
        2'd0: lizzieLet0_4MQNode_4QNode_Bool_1_onehotd = 4'd1;
        2'd1: lizzieLet0_4MQNode_4QNode_Bool_1_onehotd = 4'd2;
        2'd2: lizzieLet0_4MQNode_4QNode_Bool_1_onehotd = 4'd4;
        2'd3: lizzieLet0_4MQNode_4QNode_Bool_1_onehotd = 4'd8;
        default: lizzieLet0_4MQNode_4QNode_Bool_1_onehotd = 4'd0;
      endcase
    else lizzieLet0_4MQNode_4QNode_Bool_1_onehotd = 4'd0;
  assign _112_d = {lizzieLet0_4MQNode_4QNode_Bool_1_d[66:1],
                   lizzieLet0_4MQNode_4QNode_Bool_1_onehotd[0]};
  assign _111_d = {lizzieLet0_4MQNode_4QNode_Bool_1_d[66:1],
                   lizzieLet0_4MQNode_4QNode_Bool_1_onehotd[1]};
  assign lizzieLet0_4MQNode_4QNode_Bool_1QNode_Bool_d = {lizzieLet0_4MQNode_4QNode_Bool_1_d[66:1],
                                                         lizzieLet0_4MQNode_4QNode_Bool_1_onehotd[2]};
  assign _110_d = {lizzieLet0_4MQNode_4QNode_Bool_1_d[66:1],
                   lizzieLet0_4MQNode_4QNode_Bool_1_onehotd[3]};
  assign lizzieLet0_4MQNode_4QNode_Bool_1_r = (| (lizzieLet0_4MQNode_4QNode_Bool_1_onehotd & {_110_r,
                                                                                              lizzieLet0_4MQNode_4QNode_Bool_1QNode_Bool_r,
                                                                                              _111_r,
                                                                                              _112_r}));
  assign lizzieLet0_4MQNode_4QNode_Bool_2_r = lizzieLet0_4MQNode_4QNode_Bool_1_r;
  
  /* demux (Ty QTree_Bool,
       Ty Go) : (lizzieLet0_4MQNode_4QNode_Bool_3,QTree_Bool) (lizzieLet0_4MQNode_3QNode_Bool,Go) > [(lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool,Go),
                                                                                                     (lizzieLet0_4MQNode_4QNode_Bool_3QVal_Bool,Go),
                                                                                                     (lizzieLet0_4MQNode_4QNode_Bool_3QNode_Bool,Go),
                                                                                                     (lizzieLet0_4MQNode_4QNode_Bool_3QError_Bool,Go)] */
  logic [3:0] lizzieLet0_4MQNode_3QNode_Bool_onehotd;
  always_comb
    if ((lizzieLet0_4MQNode_4QNode_Bool_3_d[0] && lizzieLet0_4MQNode_3QNode_Bool_d[0]))
      unique case (lizzieLet0_4MQNode_4QNode_Bool_3_d[2:1])
        2'd0: lizzieLet0_4MQNode_3QNode_Bool_onehotd = 4'd1;
        2'd1: lizzieLet0_4MQNode_3QNode_Bool_onehotd = 4'd2;
        2'd2: lizzieLet0_4MQNode_3QNode_Bool_onehotd = 4'd4;
        2'd3: lizzieLet0_4MQNode_3QNode_Bool_onehotd = 4'd8;
        default: lizzieLet0_4MQNode_3QNode_Bool_onehotd = 4'd0;
      endcase
    else lizzieLet0_4MQNode_3QNode_Bool_onehotd = 4'd0;
  assign lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_d = lizzieLet0_4MQNode_3QNode_Bool_onehotd[0];
  assign lizzieLet0_4MQNode_4QNode_Bool_3QVal_Bool_d = lizzieLet0_4MQNode_3QNode_Bool_onehotd[1];
  assign lizzieLet0_4MQNode_4QNode_Bool_3QNode_Bool_d = lizzieLet0_4MQNode_3QNode_Bool_onehotd[2];
  assign lizzieLet0_4MQNode_4QNode_Bool_3QError_Bool_d = lizzieLet0_4MQNode_3QNode_Bool_onehotd[3];
  assign lizzieLet0_4MQNode_3QNode_Bool_r = (| (lizzieLet0_4MQNode_3QNode_Bool_onehotd & {lizzieLet0_4MQNode_4QNode_Bool_3QError_Bool_r,
                                                                                          lizzieLet0_4MQNode_4QNode_Bool_3QNode_Bool_r,
                                                                                          lizzieLet0_4MQNode_4QNode_Bool_3QVal_Bool_r,
                                                                                          lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_r}));
  assign lizzieLet0_4MQNode_4QNode_Bool_3_r = lizzieLet0_4MQNode_3QNode_Bool_r;
  
  /* fork (Ty Go) : (lizzieLet0_4MQNode_4QNode_Bool_3QError_Bool,Go) > [(lizzieLet0_4MQNode_4QNode_Bool_3QError_Bool_1,Go),
                                                                   (lizzieLet0_4MQNode_4QNode_Bool_3QError_Bool_2,Go)] */
  logic [1:0] lizzieLet0_4MQNode_4QNode_Bool_3QError_Bool_emitted;
  logic [1:0] lizzieLet0_4MQNode_4QNode_Bool_3QError_Bool_done;
  assign lizzieLet0_4MQNode_4QNode_Bool_3QError_Bool_1_d = (lizzieLet0_4MQNode_4QNode_Bool_3QError_Bool_d[0] && (! lizzieLet0_4MQNode_4QNode_Bool_3QError_Bool_emitted[0]));
  assign lizzieLet0_4MQNode_4QNode_Bool_3QError_Bool_2_d = (lizzieLet0_4MQNode_4QNode_Bool_3QError_Bool_d[0] && (! lizzieLet0_4MQNode_4QNode_Bool_3QError_Bool_emitted[1]));
  assign lizzieLet0_4MQNode_4QNode_Bool_3QError_Bool_done = (lizzieLet0_4MQNode_4QNode_Bool_3QError_Bool_emitted | ({lizzieLet0_4MQNode_4QNode_Bool_3QError_Bool_2_d[0],
                                                                                                                     lizzieLet0_4MQNode_4QNode_Bool_3QError_Bool_1_d[0]} & {lizzieLet0_4MQNode_4QNode_Bool_3QError_Bool_2_r,
                                                                                                                                                                            lizzieLet0_4MQNode_4QNode_Bool_3QError_Bool_1_r}));
  assign lizzieLet0_4MQNode_4QNode_Bool_3QError_Bool_r = (& lizzieLet0_4MQNode_4QNode_Bool_3QError_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QNode_Bool_3QError_Bool_emitted <= 2'd0;
    else
      lizzieLet0_4MQNode_4QNode_Bool_3QError_Bool_emitted <= (lizzieLet0_4MQNode_4QNode_Bool_3QError_Bool_r ? 2'd0 :
                                                              lizzieLet0_4MQNode_4QNode_Bool_3QError_Bool_done);
  
  /* dcon (Ty QTree_Bool,
      Dcon QError_Bool) : [(lizzieLet0_4MQNode_4QNode_Bool_3QError_Bool_1,Go)] > (lizzieLet0_4MQNode_4QNode_Bool_3QError_Bool_1QError_Bool,QTree_Bool) */
  assign lizzieLet0_4MQNode_4QNode_Bool_3QError_Bool_1QError_Bool_d = QError_Bool_dc((& {lizzieLet0_4MQNode_4QNode_Bool_3QError_Bool_1_d[0]}), lizzieLet0_4MQNode_4QNode_Bool_3QError_Bool_1_d);
  assign {lizzieLet0_4MQNode_4QNode_Bool_3QError_Bool_1_r} = {1 {(lizzieLet0_4MQNode_4QNode_Bool_3QError_Bool_1QError_Bool_r && lizzieLet0_4MQNode_4QNode_Bool_3QError_Bool_1QError_Bool_d[0])}};
  
  /* buf (Ty QTree_Bool) : (lizzieLet0_4MQNode_4QNode_Bool_3QError_Bool_1QError_Bool,QTree_Bool) > (lizzieLet18_1_1_argbuf,QTree_Bool) */
  QTree_Bool_t lizzieLet0_4MQNode_4QNode_Bool_3QError_Bool_1QError_Bool_bufchan_d;
  logic lizzieLet0_4MQNode_4QNode_Bool_3QError_Bool_1QError_Bool_bufchan_r;
  assign lizzieLet0_4MQNode_4QNode_Bool_3QError_Bool_1QError_Bool_r = ((! lizzieLet0_4MQNode_4QNode_Bool_3QError_Bool_1QError_Bool_bufchan_d[0]) || lizzieLet0_4MQNode_4QNode_Bool_3QError_Bool_1QError_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QNode_Bool_3QError_Bool_1QError_Bool_bufchan_d <= {66'd0,
                                                                             1'd0};
    else
      if (lizzieLet0_4MQNode_4QNode_Bool_3QError_Bool_1QError_Bool_r)
        lizzieLet0_4MQNode_4QNode_Bool_3QError_Bool_1QError_Bool_bufchan_d <= lizzieLet0_4MQNode_4QNode_Bool_3QError_Bool_1QError_Bool_d;
  QTree_Bool_t lizzieLet0_4MQNode_4QNode_Bool_3QError_Bool_1QError_Bool_bufchan_buf;
  assign lizzieLet0_4MQNode_4QNode_Bool_3QError_Bool_1QError_Bool_bufchan_r = (! lizzieLet0_4MQNode_4QNode_Bool_3QError_Bool_1QError_Bool_bufchan_buf[0]);
  assign lizzieLet18_1_1_argbuf_d = (lizzieLet0_4MQNode_4QNode_Bool_3QError_Bool_1QError_Bool_bufchan_buf[0] ? lizzieLet0_4MQNode_4QNode_Bool_3QError_Bool_1QError_Bool_bufchan_buf :
                                     lizzieLet0_4MQNode_4QNode_Bool_3QError_Bool_1QError_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QNode_Bool_3QError_Bool_1QError_Bool_bufchan_buf <= {66'd0,
                                                                               1'd0};
    else
      if ((lizzieLet18_1_1_argbuf_r && lizzieLet0_4MQNode_4QNode_Bool_3QError_Bool_1QError_Bool_bufchan_buf[0]))
        lizzieLet0_4MQNode_4QNode_Bool_3QError_Bool_1QError_Bool_bufchan_buf <= {66'd0,
                                                                                 1'd0};
      else if (((! lizzieLet18_1_1_argbuf_r) && (! lizzieLet0_4MQNode_4QNode_Bool_3QError_Bool_1QError_Bool_bufchan_buf[0])))
        lizzieLet0_4MQNode_4QNode_Bool_3QError_Bool_1QError_Bool_bufchan_buf <= lizzieLet0_4MQNode_4QNode_Bool_3QError_Bool_1QError_Bool_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet0_4MQNode_4QNode_Bool_3QError_Bool_2,Go) > (lizzieLet0_4MQNode_4QNode_Bool_3QError_Bool_2_argbuf,Go) */
  Go_t lizzieLet0_4MQNode_4QNode_Bool_3QError_Bool_2_bufchan_d;
  logic lizzieLet0_4MQNode_4QNode_Bool_3QError_Bool_2_bufchan_r;
  assign lizzieLet0_4MQNode_4QNode_Bool_3QError_Bool_2_r = ((! lizzieLet0_4MQNode_4QNode_Bool_3QError_Bool_2_bufchan_d[0]) || lizzieLet0_4MQNode_4QNode_Bool_3QError_Bool_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QNode_Bool_3QError_Bool_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet0_4MQNode_4QNode_Bool_3QError_Bool_2_r)
        lizzieLet0_4MQNode_4QNode_Bool_3QError_Bool_2_bufchan_d <= lizzieLet0_4MQNode_4QNode_Bool_3QError_Bool_2_d;
  Go_t lizzieLet0_4MQNode_4QNode_Bool_3QError_Bool_2_bufchan_buf;
  assign lizzieLet0_4MQNode_4QNode_Bool_3QError_Bool_2_bufchan_r = (! lizzieLet0_4MQNode_4QNode_Bool_3QError_Bool_2_bufchan_buf[0]);
  assign lizzieLet0_4MQNode_4QNode_Bool_3QError_Bool_2_argbuf_d = (lizzieLet0_4MQNode_4QNode_Bool_3QError_Bool_2_bufchan_buf[0] ? lizzieLet0_4MQNode_4QNode_Bool_3QError_Bool_2_bufchan_buf :
                                                                   lizzieLet0_4MQNode_4QNode_Bool_3QError_Bool_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QNode_Bool_3QError_Bool_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet0_4MQNode_4QNode_Bool_3QError_Bool_2_argbuf_r && lizzieLet0_4MQNode_4QNode_Bool_3QError_Bool_2_bufchan_buf[0]))
        lizzieLet0_4MQNode_4QNode_Bool_3QError_Bool_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet0_4MQNode_4QNode_Bool_3QError_Bool_2_argbuf_r) && (! lizzieLet0_4MQNode_4QNode_Bool_3QError_Bool_2_bufchan_buf[0])))
        lizzieLet0_4MQNode_4QNode_Bool_3QError_Bool_2_bufchan_buf <= lizzieLet0_4MQNode_4QNode_Bool_3QError_Bool_2_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet0_4MQNode_4QNode_Bool_3QNode_Bool,Go) > (lizzieLet0_4MQNode_4QNode_Bool_3QNode_Bool_1_argbuf,Go) */
  Go_t lizzieLet0_4MQNode_4QNode_Bool_3QNode_Bool_bufchan_d;
  logic lizzieLet0_4MQNode_4QNode_Bool_3QNode_Bool_bufchan_r;
  assign lizzieLet0_4MQNode_4QNode_Bool_3QNode_Bool_r = ((! lizzieLet0_4MQNode_4QNode_Bool_3QNode_Bool_bufchan_d[0]) || lizzieLet0_4MQNode_4QNode_Bool_3QNode_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QNode_Bool_3QNode_Bool_bufchan_d <= 1'd0;
    else
      if (lizzieLet0_4MQNode_4QNode_Bool_3QNode_Bool_r)
        lizzieLet0_4MQNode_4QNode_Bool_3QNode_Bool_bufchan_d <= lizzieLet0_4MQNode_4QNode_Bool_3QNode_Bool_d;
  Go_t lizzieLet0_4MQNode_4QNode_Bool_3QNode_Bool_bufchan_buf;
  assign lizzieLet0_4MQNode_4QNode_Bool_3QNode_Bool_bufchan_r = (! lizzieLet0_4MQNode_4QNode_Bool_3QNode_Bool_bufchan_buf[0]);
  assign lizzieLet0_4MQNode_4QNode_Bool_3QNode_Bool_1_argbuf_d = (lizzieLet0_4MQNode_4QNode_Bool_3QNode_Bool_bufchan_buf[0] ? lizzieLet0_4MQNode_4QNode_Bool_3QNode_Bool_bufchan_buf :
                                                                  lizzieLet0_4MQNode_4QNode_Bool_3QNode_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QNode_Bool_3QNode_Bool_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet0_4MQNode_4QNode_Bool_3QNode_Bool_1_argbuf_r && lizzieLet0_4MQNode_4QNode_Bool_3QNode_Bool_bufchan_buf[0]))
        lizzieLet0_4MQNode_4QNode_Bool_3QNode_Bool_bufchan_buf <= 1'd0;
      else if (((! lizzieLet0_4MQNode_4QNode_Bool_3QNode_Bool_1_argbuf_r) && (! lizzieLet0_4MQNode_4QNode_Bool_3QNode_Bool_bufchan_buf[0])))
        lizzieLet0_4MQNode_4QNode_Bool_3QNode_Bool_bufchan_buf <= lizzieLet0_4MQNode_4QNode_Bool_3QNode_Bool_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool,Go) > [(lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_1,Go),
                                                                  (lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_2,Go),
                                                                  (lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_3,Go),
                                                                  (lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_4,Go),
                                                                  (lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_5,Go)] */
  logic [4:0] lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_emitted;
  logic [4:0] lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_done;
  assign lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_1_d = (lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_d[0] && (! lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_emitted[0]));
  assign lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_2_d = (lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_d[0] && (! lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_emitted[1]));
  assign lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_3_d = (lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_d[0] && (! lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_emitted[2]));
  assign lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_4_d = (lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_d[0] && (! lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_emitted[3]));
  assign lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_5_d = (lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_d[0] && (! lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_emitted[4]));
  assign lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_done = (lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_emitted | ({lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_5_d[0],
                                                                                                                   lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_4_d[0],
                                                                                                                   lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_3_d[0],
                                                                                                                   lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_2_d[0],
                                                                                                                   lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_1_d[0]} & {lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_5_r,
                                                                                                                                                                         lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_4_r,
                                                                                                                                                                         lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_3_r,
                                                                                                                                                                         lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_2_r,
                                                                                                                                                                         lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_1_r}));
  assign lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_r = (& lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_emitted <= 5'd0;
    else
      lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_emitted <= (lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_r ? 5'd0 :
                                                             lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_done);
  
  /* buf (Ty Go) : (lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_1,Go) > (lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_1_argbuf,Go) */
  Go_t lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_1_bufchan_d;
  logic lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_1_bufchan_r;
  assign lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_1_r = ((! lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_1_bufchan_d[0]) || lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_1_bufchan_d <= 1'd0;
    else
      if (lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_1_r)
        lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_1_bufchan_d <= lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_1_d;
  Go_t lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_1_bufchan_buf;
  assign lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_1_bufchan_r = (! lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_1_bufchan_buf[0]);
  assign lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_1_argbuf_d = (lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_1_bufchan_buf[0] ? lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_1_bufchan_buf :
                                                                  lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_1_argbuf_r && lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_1_bufchan_buf[0]))
        lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_1_argbuf_r) && (! lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_1_bufchan_buf[0])))
        lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_1_bufchan_buf <= lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_1_bufchan_d;
  
  /* dcon (Ty TupGo___Pointer_MaskQTree___Pointer_QTree_Bool,
      Dcon TupGo___Pointer_MaskQTree___Pointer_QTree_Bool) : [(lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_1_argbuf,Go),
                                                              (lizzieLet0_4MQNode_4QNode_Bool_8QNone_Bool_1_argbuf,Pointer_MaskQTree),
                                                              (lizzieLet0_4MQNode_4QNode_Bool_12QNone_Bool_1_argbuf,Pointer_QTree_Bool)] > (f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool5,TupGo___Pointer_MaskQTree___Pointer_QTree_Bool) */
  assign \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool5_d  = TupGo___Pointer_MaskQTree___Pointer_QTree_Bool_dc((& {lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_1_argbuf_d[0],
                                                                                                                                               lizzieLet0_4MQNode_4QNode_Bool_8QNone_Bool_1_argbuf_d[0],
                                                                                                                                               lizzieLet0_4MQNode_4QNode_Bool_12QNone_Bool_1_argbuf_d[0]}), lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_1_argbuf_d, lizzieLet0_4MQNode_4QNode_Bool_8QNone_Bool_1_argbuf_d, lizzieLet0_4MQNode_4QNode_Bool_12QNone_Bool_1_argbuf_d);
  assign {lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_1_argbuf_r,
          lizzieLet0_4MQNode_4QNode_Bool_8QNone_Bool_1_argbuf_r,
          lizzieLet0_4MQNode_4QNode_Bool_12QNone_Bool_1_argbuf_r} = {3 {(\f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool5_r  && \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool5_d [0])}};
  
  /* buf (Ty Go) : (lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_2,Go) > (lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_2_argbuf,Go) */
  Go_t lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_2_bufchan_d;
  logic lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_2_bufchan_r;
  assign lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_2_r = ((! lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_2_bufchan_d[0]) || lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_2_r)
        lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_2_bufchan_d <= lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_2_d;
  Go_t lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_2_bufchan_buf;
  assign lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_2_bufchan_r = (! lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_2_bufchan_buf[0]);
  assign lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_2_argbuf_d = (lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_2_bufchan_buf[0] ? lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_2_bufchan_buf :
                                                                  lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_2_argbuf_r && lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_2_bufchan_buf[0]))
        lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_2_argbuf_r) && (! lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_2_bufchan_buf[0])))
        lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_2_bufchan_buf <= lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_2_bufchan_d;
  
  /* dcon (Ty TupGo___Pointer_MaskQTree___Pointer_QTree_Bool,
      Dcon TupGo___Pointer_MaskQTree___Pointer_QTree_Bool) : [(lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_2_argbuf,Go),
                                                              (lizzieLet0_4MQNode_4QNode_Bool_7QNone_Bool_1_argbuf,Pointer_MaskQTree),
                                                              (lizzieLet0_4MQNode_4QNode_Bool_11QNone_Bool_1_argbuf,Pointer_QTree_Bool)] > (f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool6,TupGo___Pointer_MaskQTree___Pointer_QTree_Bool) */
  assign \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool6_d  = TupGo___Pointer_MaskQTree___Pointer_QTree_Bool_dc((& {lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_2_argbuf_d[0],
                                                                                                                                               lizzieLet0_4MQNode_4QNode_Bool_7QNone_Bool_1_argbuf_d[0],
                                                                                                                                               lizzieLet0_4MQNode_4QNode_Bool_11QNone_Bool_1_argbuf_d[0]}), lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_2_argbuf_d, lizzieLet0_4MQNode_4QNode_Bool_7QNone_Bool_1_argbuf_d, lizzieLet0_4MQNode_4QNode_Bool_11QNone_Bool_1_argbuf_d);
  assign {lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_2_argbuf_r,
          lizzieLet0_4MQNode_4QNode_Bool_7QNone_Bool_1_argbuf_r,
          lizzieLet0_4MQNode_4QNode_Bool_11QNone_Bool_1_argbuf_r} = {3 {(\f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool6_r  && \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool6_d [0])}};
  
  /* buf (Ty Go) : (lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_3,Go) > (lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_3_argbuf,Go) */
  Go_t lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_3_bufchan_d;
  logic lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_3_bufchan_r;
  assign lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_3_r = ((! lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_3_bufchan_d[0]) || lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_3_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_3_bufchan_d <= 1'd0;
    else
      if (lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_3_r)
        lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_3_bufchan_d <= lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_3_d;
  Go_t lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_3_bufchan_buf;
  assign lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_3_bufchan_r = (! lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_3_bufchan_buf[0]);
  assign lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_3_argbuf_d = (lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_3_bufchan_buf[0] ? lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_3_bufchan_buf :
                                                                  lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_3_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_3_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_3_argbuf_r && lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_3_bufchan_buf[0]))
        lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_3_bufchan_buf <= 1'd0;
      else if (((! lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_3_argbuf_r) && (! lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_3_bufchan_buf[0])))
        lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_3_bufchan_buf <= lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_3_bufchan_d;
  
  /* dcon (Ty TupGo___Pointer_MaskQTree___Pointer_QTree_Bool,
      Dcon TupGo___Pointer_MaskQTree___Pointer_QTree_Bool) : [(lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_3_argbuf,Go),
                                                              (lizzieLet0_4MQNode_4QNode_Bool_6QNone_Bool_1_argbuf,Pointer_MaskQTree),
                                                              (lizzieLet0_4MQNode_4QNode_Bool_10QNone_Bool_1_argbuf,Pointer_QTree_Bool)] > (f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool7,TupGo___Pointer_MaskQTree___Pointer_QTree_Bool) */
  assign \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool7_d  = TupGo___Pointer_MaskQTree___Pointer_QTree_Bool_dc((& {lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_3_argbuf_d[0],
                                                                                                                                               lizzieLet0_4MQNode_4QNode_Bool_6QNone_Bool_1_argbuf_d[0],
                                                                                                                                               lizzieLet0_4MQNode_4QNode_Bool_10QNone_Bool_1_argbuf_d[0]}), lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_3_argbuf_d, lizzieLet0_4MQNode_4QNode_Bool_6QNone_Bool_1_argbuf_d, lizzieLet0_4MQNode_4QNode_Bool_10QNone_Bool_1_argbuf_d);
  assign {lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_3_argbuf_r,
          lizzieLet0_4MQNode_4QNode_Bool_6QNone_Bool_1_argbuf_r,
          lizzieLet0_4MQNode_4QNode_Bool_10QNone_Bool_1_argbuf_r} = {3 {(\f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool7_r  && \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool7_d [0])}};
  
  /* buf (Ty Go) : (lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_4,Go) > (lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_4_argbuf,Go) */
  Go_t lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_4_bufchan_d;
  logic lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_4_bufchan_r;
  assign lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_4_r = ((! lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_4_bufchan_d[0]) || lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_4_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_4_bufchan_d <= 1'd0;
    else
      if (lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_4_r)
        lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_4_bufchan_d <= lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_4_d;
  Go_t lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_4_bufchan_buf;
  assign lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_4_bufchan_r = (! lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_4_bufchan_buf[0]);
  assign lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_4_argbuf_d = (lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_4_bufchan_buf[0] ? lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_4_bufchan_buf :
                                                                  lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_4_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_4_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_4_argbuf_r && lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_4_bufchan_buf[0]))
        lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_4_bufchan_buf <= 1'd0;
      else if (((! lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_4_argbuf_r) && (! lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_4_bufchan_buf[0])))
        lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_4_bufchan_buf <= lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_4_bufchan_d;
  
  /* dcon (Ty TupGo___Pointer_MaskQTree___Pointer_QTree_Bool,
      Dcon TupGo___Pointer_MaskQTree___Pointer_QTree_Bool) : [(lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_4_argbuf,Go),
                                                              (lizzieLet0_4MQNode_4QNode_Bool_5QNone_Bool_1_argbuf,Pointer_MaskQTree),
                                                              (lizzieLet0_4MQNode_4QNode_Bool_9QNone_Bool_1_argbuf,Pointer_QTree_Bool)] > (f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool8,TupGo___Pointer_MaskQTree___Pointer_QTree_Bool) */
  assign \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool8_d  = TupGo___Pointer_MaskQTree___Pointer_QTree_Bool_dc((& {lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_4_argbuf_d[0],
                                                                                                                                               lizzieLet0_4MQNode_4QNode_Bool_5QNone_Bool_1_argbuf_d[0],
                                                                                                                                               lizzieLet0_4MQNode_4QNode_Bool_9QNone_Bool_1_argbuf_d[0]}), lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_4_argbuf_d, lizzieLet0_4MQNode_4QNode_Bool_5QNone_Bool_1_argbuf_d, lizzieLet0_4MQNode_4QNode_Bool_9QNone_Bool_1_argbuf_d);
  assign {lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_4_argbuf_r,
          lizzieLet0_4MQNode_4QNode_Bool_5QNone_Bool_1_argbuf_r,
          lizzieLet0_4MQNode_4QNode_Bool_9QNone_Bool_1_argbuf_r} = {3 {(\f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool8_r  && \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool8_d [0])}};
  
  /* buf (Ty Go) : (lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_5,Go) > (lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_5_argbuf,Go) */
  Go_t lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_5_bufchan_d;
  logic lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_5_bufchan_r;
  assign lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_5_r = ((! lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_5_bufchan_d[0]) || lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_5_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_5_bufchan_d <= 1'd0;
    else
      if (lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_5_r)
        lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_5_bufchan_d <= lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_5_d;
  Go_t lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_5_bufchan_buf;
  assign lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_5_bufchan_r = (! lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_5_bufchan_buf[0]);
  assign lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_5_argbuf_d = (lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_5_bufchan_buf[0] ? lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_5_bufchan_buf :
                                                                  lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_5_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_5_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_5_argbuf_r && lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_5_bufchan_buf[0]))
        lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_5_bufchan_buf <= 1'd0;
      else if (((! lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_5_argbuf_r) && (! lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_5_bufchan_buf[0])))
        lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_5_bufchan_buf <= lizzieLet0_4MQNode_4QNode_Bool_3QNone_Bool_5_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet0_4MQNode_4QNode_Bool_3QVal_Bool,Go) > [(lizzieLet0_4MQNode_4QNode_Bool_3QVal_Bool_1,Go),
                                                                 (lizzieLet0_4MQNode_4QNode_Bool_3QVal_Bool_2,Go)] */
  logic [1:0] lizzieLet0_4MQNode_4QNode_Bool_3QVal_Bool_emitted;
  logic [1:0] lizzieLet0_4MQNode_4QNode_Bool_3QVal_Bool_done;
  assign lizzieLet0_4MQNode_4QNode_Bool_3QVal_Bool_1_d = (lizzieLet0_4MQNode_4QNode_Bool_3QVal_Bool_d[0] && (! lizzieLet0_4MQNode_4QNode_Bool_3QVal_Bool_emitted[0]));
  assign lizzieLet0_4MQNode_4QNode_Bool_3QVal_Bool_2_d = (lizzieLet0_4MQNode_4QNode_Bool_3QVal_Bool_d[0] && (! lizzieLet0_4MQNode_4QNode_Bool_3QVal_Bool_emitted[1]));
  assign lizzieLet0_4MQNode_4QNode_Bool_3QVal_Bool_done = (lizzieLet0_4MQNode_4QNode_Bool_3QVal_Bool_emitted | ({lizzieLet0_4MQNode_4QNode_Bool_3QVal_Bool_2_d[0],
                                                                                                                 lizzieLet0_4MQNode_4QNode_Bool_3QVal_Bool_1_d[0]} & {lizzieLet0_4MQNode_4QNode_Bool_3QVal_Bool_2_r,
                                                                                                                                                                      lizzieLet0_4MQNode_4QNode_Bool_3QVal_Bool_1_r}));
  assign lizzieLet0_4MQNode_4QNode_Bool_3QVal_Bool_r = (& lizzieLet0_4MQNode_4QNode_Bool_3QVal_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QNode_Bool_3QVal_Bool_emitted <= 2'd0;
    else
      lizzieLet0_4MQNode_4QNode_Bool_3QVal_Bool_emitted <= (lizzieLet0_4MQNode_4QNode_Bool_3QVal_Bool_r ? 2'd0 :
                                                            lizzieLet0_4MQNode_4QNode_Bool_3QVal_Bool_done);
  
  /* dcon (Ty QTree_Bool,
      Dcon QError_Bool) : [(lizzieLet0_4MQNode_4QNode_Bool_3QVal_Bool_1,Go)] > (lizzieLet0_4MQNode_4QNode_Bool_3QVal_Bool_1QError_Bool,QTree_Bool) */
  assign lizzieLet0_4MQNode_4QNode_Bool_3QVal_Bool_1QError_Bool_d = QError_Bool_dc((& {lizzieLet0_4MQNode_4QNode_Bool_3QVal_Bool_1_d[0]}), lizzieLet0_4MQNode_4QNode_Bool_3QVal_Bool_1_d);
  assign {lizzieLet0_4MQNode_4QNode_Bool_3QVal_Bool_1_r} = {1 {(lizzieLet0_4MQNode_4QNode_Bool_3QVal_Bool_1QError_Bool_r && lizzieLet0_4MQNode_4QNode_Bool_3QVal_Bool_1QError_Bool_d[0])}};
  
  /* buf (Ty QTree_Bool) : (lizzieLet0_4MQNode_4QNode_Bool_3QVal_Bool_1QError_Bool,QTree_Bool) > (lizzieLet16_1_1_argbuf,QTree_Bool) */
  QTree_Bool_t lizzieLet0_4MQNode_4QNode_Bool_3QVal_Bool_1QError_Bool_bufchan_d;
  logic lizzieLet0_4MQNode_4QNode_Bool_3QVal_Bool_1QError_Bool_bufchan_r;
  assign lizzieLet0_4MQNode_4QNode_Bool_3QVal_Bool_1QError_Bool_r = ((! lizzieLet0_4MQNode_4QNode_Bool_3QVal_Bool_1QError_Bool_bufchan_d[0]) || lizzieLet0_4MQNode_4QNode_Bool_3QVal_Bool_1QError_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QNode_Bool_3QVal_Bool_1QError_Bool_bufchan_d <= {66'd0,
                                                                           1'd0};
    else
      if (lizzieLet0_4MQNode_4QNode_Bool_3QVal_Bool_1QError_Bool_r)
        lizzieLet0_4MQNode_4QNode_Bool_3QVal_Bool_1QError_Bool_bufchan_d <= lizzieLet0_4MQNode_4QNode_Bool_3QVal_Bool_1QError_Bool_d;
  QTree_Bool_t lizzieLet0_4MQNode_4QNode_Bool_3QVal_Bool_1QError_Bool_bufchan_buf;
  assign lizzieLet0_4MQNode_4QNode_Bool_3QVal_Bool_1QError_Bool_bufchan_r = (! lizzieLet0_4MQNode_4QNode_Bool_3QVal_Bool_1QError_Bool_bufchan_buf[0]);
  assign lizzieLet16_1_1_argbuf_d = (lizzieLet0_4MQNode_4QNode_Bool_3QVal_Bool_1QError_Bool_bufchan_buf[0] ? lizzieLet0_4MQNode_4QNode_Bool_3QVal_Bool_1QError_Bool_bufchan_buf :
                                     lizzieLet0_4MQNode_4QNode_Bool_3QVal_Bool_1QError_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QNode_Bool_3QVal_Bool_1QError_Bool_bufchan_buf <= {66'd0,
                                                                             1'd0};
    else
      if ((lizzieLet16_1_1_argbuf_r && lizzieLet0_4MQNode_4QNode_Bool_3QVal_Bool_1QError_Bool_bufchan_buf[0]))
        lizzieLet0_4MQNode_4QNode_Bool_3QVal_Bool_1QError_Bool_bufchan_buf <= {66'd0,
                                                                               1'd0};
      else if (((! lizzieLet16_1_1_argbuf_r) && (! lizzieLet0_4MQNode_4QNode_Bool_3QVal_Bool_1QError_Bool_bufchan_buf[0])))
        lizzieLet0_4MQNode_4QNode_Bool_3QVal_Bool_1QError_Bool_bufchan_buf <= lizzieLet0_4MQNode_4QNode_Bool_3QVal_Bool_1QError_Bool_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet0_4MQNode_4QNode_Bool_3QVal_Bool_2,Go) > (lizzieLet0_4MQNode_4QNode_Bool_3QVal_Bool_2_argbuf,Go) */
  Go_t lizzieLet0_4MQNode_4QNode_Bool_3QVal_Bool_2_bufchan_d;
  logic lizzieLet0_4MQNode_4QNode_Bool_3QVal_Bool_2_bufchan_r;
  assign lizzieLet0_4MQNode_4QNode_Bool_3QVal_Bool_2_r = ((! lizzieLet0_4MQNode_4QNode_Bool_3QVal_Bool_2_bufchan_d[0]) || lizzieLet0_4MQNode_4QNode_Bool_3QVal_Bool_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QNode_Bool_3QVal_Bool_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet0_4MQNode_4QNode_Bool_3QVal_Bool_2_r)
        lizzieLet0_4MQNode_4QNode_Bool_3QVal_Bool_2_bufchan_d <= lizzieLet0_4MQNode_4QNode_Bool_3QVal_Bool_2_d;
  Go_t lizzieLet0_4MQNode_4QNode_Bool_3QVal_Bool_2_bufchan_buf;
  assign lizzieLet0_4MQNode_4QNode_Bool_3QVal_Bool_2_bufchan_r = (! lizzieLet0_4MQNode_4QNode_Bool_3QVal_Bool_2_bufchan_buf[0]);
  assign lizzieLet0_4MQNode_4QNode_Bool_3QVal_Bool_2_argbuf_d = (lizzieLet0_4MQNode_4QNode_Bool_3QVal_Bool_2_bufchan_buf[0] ? lizzieLet0_4MQNode_4QNode_Bool_3QVal_Bool_2_bufchan_buf :
                                                                 lizzieLet0_4MQNode_4QNode_Bool_3QVal_Bool_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QNode_Bool_3QVal_Bool_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet0_4MQNode_4QNode_Bool_3QVal_Bool_2_argbuf_r && lizzieLet0_4MQNode_4QNode_Bool_3QVal_Bool_2_bufchan_buf[0]))
        lizzieLet0_4MQNode_4QNode_Bool_3QVal_Bool_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet0_4MQNode_4QNode_Bool_3QVal_Bool_2_argbuf_r) && (! lizzieLet0_4MQNode_4QNode_Bool_3QVal_Bool_2_bufchan_buf[0])))
        lizzieLet0_4MQNode_4QNode_Bool_3QVal_Bool_2_bufchan_buf <= lizzieLet0_4MQNode_4QNode_Bool_3QVal_Bool_2_bufchan_d;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_CTf) : (lizzieLet0_4MQNode_4QNode_Bool_4,QTree_Bool) (lizzieLet0_4MQNode_5QNode_Bool,Pointer_CTf) > [(lizzieLet0_4MQNode_4QNode_Bool_4QNone_Bool,Pointer_CTf),
                                                                                                                       (lizzieLet0_4MQNode_4QNode_Bool_4QVal_Bool,Pointer_CTf),
                                                                                                                       (lizzieLet0_4MQNode_4QNode_Bool_4QNode_Bool,Pointer_CTf),
                                                                                                                       (lizzieLet0_4MQNode_4QNode_Bool_4QError_Bool,Pointer_CTf)] */
  logic [3:0] lizzieLet0_4MQNode_5QNode_Bool_onehotd;
  always_comb
    if ((lizzieLet0_4MQNode_4QNode_Bool_4_d[0] && lizzieLet0_4MQNode_5QNode_Bool_d[0]))
      unique case (lizzieLet0_4MQNode_4QNode_Bool_4_d[2:1])
        2'd0: lizzieLet0_4MQNode_5QNode_Bool_onehotd = 4'd1;
        2'd1: lizzieLet0_4MQNode_5QNode_Bool_onehotd = 4'd2;
        2'd2: lizzieLet0_4MQNode_5QNode_Bool_onehotd = 4'd4;
        2'd3: lizzieLet0_4MQNode_5QNode_Bool_onehotd = 4'd8;
        default: lizzieLet0_4MQNode_5QNode_Bool_onehotd = 4'd0;
      endcase
    else lizzieLet0_4MQNode_5QNode_Bool_onehotd = 4'd0;
  assign lizzieLet0_4MQNode_4QNode_Bool_4QNone_Bool_d = {lizzieLet0_4MQNode_5QNode_Bool_d[16:1],
                                                         lizzieLet0_4MQNode_5QNode_Bool_onehotd[0]};
  assign lizzieLet0_4MQNode_4QNode_Bool_4QVal_Bool_d = {lizzieLet0_4MQNode_5QNode_Bool_d[16:1],
                                                        lizzieLet0_4MQNode_5QNode_Bool_onehotd[1]};
  assign lizzieLet0_4MQNode_4QNode_Bool_4QNode_Bool_d = {lizzieLet0_4MQNode_5QNode_Bool_d[16:1],
                                                         lizzieLet0_4MQNode_5QNode_Bool_onehotd[2]};
  assign lizzieLet0_4MQNode_4QNode_Bool_4QError_Bool_d = {lizzieLet0_4MQNode_5QNode_Bool_d[16:1],
                                                          lizzieLet0_4MQNode_5QNode_Bool_onehotd[3]};
  assign lizzieLet0_4MQNode_5QNode_Bool_r = (| (lizzieLet0_4MQNode_5QNode_Bool_onehotd & {lizzieLet0_4MQNode_4QNode_Bool_4QError_Bool_r,
                                                                                          lizzieLet0_4MQNode_4QNode_Bool_4QNode_Bool_r,
                                                                                          lizzieLet0_4MQNode_4QNode_Bool_4QVal_Bool_r,
                                                                                          lizzieLet0_4MQNode_4QNode_Bool_4QNone_Bool_r}));
  assign lizzieLet0_4MQNode_4QNode_Bool_4_r = lizzieLet0_4MQNode_5QNode_Bool_r;
  
  /* buf (Ty Pointer_CTf) : (lizzieLet0_4MQNode_4QNode_Bool_4QError_Bool,Pointer_CTf) > (lizzieLet0_4MQNode_4QNode_Bool_4QError_Bool_1_argbuf,Pointer_CTf) */
  Pointer_CTf_t lizzieLet0_4MQNode_4QNode_Bool_4QError_Bool_bufchan_d;
  logic lizzieLet0_4MQNode_4QNode_Bool_4QError_Bool_bufchan_r;
  assign lizzieLet0_4MQNode_4QNode_Bool_4QError_Bool_r = ((! lizzieLet0_4MQNode_4QNode_Bool_4QError_Bool_bufchan_d[0]) || lizzieLet0_4MQNode_4QNode_Bool_4QError_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QNode_Bool_4QError_Bool_bufchan_d <= {16'd0,
                                                                1'd0};
    else
      if (lizzieLet0_4MQNode_4QNode_Bool_4QError_Bool_r)
        lizzieLet0_4MQNode_4QNode_Bool_4QError_Bool_bufchan_d <= lizzieLet0_4MQNode_4QNode_Bool_4QError_Bool_d;
  Pointer_CTf_t lizzieLet0_4MQNode_4QNode_Bool_4QError_Bool_bufchan_buf;
  assign lizzieLet0_4MQNode_4QNode_Bool_4QError_Bool_bufchan_r = (! lizzieLet0_4MQNode_4QNode_Bool_4QError_Bool_bufchan_buf[0]);
  assign lizzieLet0_4MQNode_4QNode_Bool_4QError_Bool_1_argbuf_d = (lizzieLet0_4MQNode_4QNode_Bool_4QError_Bool_bufchan_buf[0] ? lizzieLet0_4MQNode_4QNode_Bool_4QError_Bool_bufchan_buf :
                                                                   lizzieLet0_4MQNode_4QNode_Bool_4QError_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QNode_Bool_4QError_Bool_bufchan_buf <= {16'd0,
                                                                  1'd0};
    else
      if ((lizzieLet0_4MQNode_4QNode_Bool_4QError_Bool_1_argbuf_r && lizzieLet0_4MQNode_4QNode_Bool_4QError_Bool_bufchan_buf[0]))
        lizzieLet0_4MQNode_4QNode_Bool_4QError_Bool_bufchan_buf <= {16'd0,
                                                                    1'd0};
      else if (((! lizzieLet0_4MQNode_4QNode_Bool_4QError_Bool_1_argbuf_r) && (! lizzieLet0_4MQNode_4QNode_Bool_4QError_Bool_bufchan_buf[0])))
        lizzieLet0_4MQNode_4QNode_Bool_4QError_Bool_bufchan_buf <= lizzieLet0_4MQNode_4QNode_Bool_4QError_Bool_bufchan_d;
  
  /* dcon (Ty CTf,
      Dcon Lcall_f3) : [(lizzieLet0_4MQNode_4QNode_Bool_4QNode_Bool,Pointer_CTf),
                        (lizzieLet0_4MQNode_4QNode_Bool_5QNode_Bool,Pointer_MaskQTree),
                        (lizzieLet0_4MQNode_4QNode_Bool_9QNode_Bool,Pointer_QTree_Bool),
                        (t1a8s_destruct,Pointer_QTree_Bool),
                        (lizzieLet0_4MQNode_4QNode_Bool_6QNode_Bool,Pointer_MaskQTree),
                        (lizzieLet0_4MQNode_4QNode_Bool_10QNode_Bool,Pointer_QTree_Bool),
                        (t2a8t_destruct,Pointer_QTree_Bool),
                        (lizzieLet0_4MQNode_4QNode_Bool_7QNode_Bool,Pointer_MaskQTree),
                        (lizzieLet0_4MQNode_4QNode_Bool_11QNode_Bool,Pointer_QTree_Bool),
                        (t3a8u_destruct,Pointer_QTree_Bool)] > (lizzieLet0_4MQNode_4QNode_Bool_4QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_5QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_9QNode_Bool_1t1a8s_1lizzieLet0_4MQNode_4QNode_Bool_6QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_10QNode_Bool_1t2a8t_1lizzieLet0_4MQNode_4QNode_Bool_7QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_11QNode_Bool_1t3a8u_1Lcall_f3,CTf) */
  assign lizzieLet0_4MQNode_4QNode_Bool_4QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_5QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_9QNode_Bool_1t1a8s_1lizzieLet0_4MQNode_4QNode_Bool_6QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_10QNode_Bool_1t2a8t_1lizzieLet0_4MQNode_4QNode_Bool_7QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_11QNode_Bool_1t3a8u_1Lcall_f3_d = Lcall_f3_dc((& {lizzieLet0_4MQNode_4QNode_Bool_4QNode_Bool_d[0],
                                                                                                                                                                                                                                                                                                                                                                                 lizzieLet0_4MQNode_4QNode_Bool_5QNode_Bool_d[0],
                                                                                                                                                                                                                                                                                                                                                                                 lizzieLet0_4MQNode_4QNode_Bool_9QNode_Bool_d[0],
                                                                                                                                                                                                                                                                                                                                                                                 t1a8s_destruct_d[0],
                                                                                                                                                                                                                                                                                                                                                                                 lizzieLet0_4MQNode_4QNode_Bool_6QNode_Bool_d[0],
                                                                                                                                                                                                                                                                                                                                                                                 lizzieLet0_4MQNode_4QNode_Bool_10QNode_Bool_d[0],
                                                                                                                                                                                                                                                                                                                                                                                 t2a8t_destruct_d[0],
                                                                                                                                                                                                                                                                                                                                                                                 lizzieLet0_4MQNode_4QNode_Bool_7QNode_Bool_d[0],
                                                                                                                                                                                                                                                                                                                                                                                 lizzieLet0_4MQNode_4QNode_Bool_11QNode_Bool_d[0],
                                                                                                                                                                                                                                                                                                                                                                                 t3a8u_destruct_d[0]}), lizzieLet0_4MQNode_4QNode_Bool_4QNode_Bool_d, lizzieLet0_4MQNode_4QNode_Bool_5QNode_Bool_d, lizzieLet0_4MQNode_4QNode_Bool_9QNode_Bool_d, t1a8s_destruct_d, lizzieLet0_4MQNode_4QNode_Bool_6QNode_Bool_d, lizzieLet0_4MQNode_4QNode_Bool_10QNode_Bool_d, t2a8t_destruct_d, lizzieLet0_4MQNode_4QNode_Bool_7QNode_Bool_d, lizzieLet0_4MQNode_4QNode_Bool_11QNode_Bool_d, t3a8u_destruct_d);
  assign {lizzieLet0_4MQNode_4QNode_Bool_4QNode_Bool_r,
          lizzieLet0_4MQNode_4QNode_Bool_5QNode_Bool_r,
          lizzieLet0_4MQNode_4QNode_Bool_9QNode_Bool_r,
          t1a8s_destruct_r,
          lizzieLet0_4MQNode_4QNode_Bool_6QNode_Bool_r,
          lizzieLet0_4MQNode_4QNode_Bool_10QNode_Bool_r,
          t2a8t_destruct_r,
          lizzieLet0_4MQNode_4QNode_Bool_7QNode_Bool_r,
          lizzieLet0_4MQNode_4QNode_Bool_11QNode_Bool_r,
          t3a8u_destruct_r} = {10 {(lizzieLet0_4MQNode_4QNode_Bool_4QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_5QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_9QNode_Bool_1t1a8s_1lizzieLet0_4MQNode_4QNode_Bool_6QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_10QNode_Bool_1t2a8t_1lizzieLet0_4MQNode_4QNode_Bool_7QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_11QNode_Bool_1t3a8u_1Lcall_f3_r && lizzieLet0_4MQNode_4QNode_Bool_4QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_5QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_9QNode_Bool_1t1a8s_1lizzieLet0_4MQNode_4QNode_Bool_6QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_10QNode_Bool_1t2a8t_1lizzieLet0_4MQNode_4QNode_Bool_7QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_11QNode_Bool_1t3a8u_1Lcall_f3_d[0])}};
  
  /* buf (Ty CTf) : (lizzieLet0_4MQNode_4QNode_Bool_4QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_5QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_9QNode_Bool_1t1a8s_1lizzieLet0_4MQNode_4QNode_Bool_6QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_10QNode_Bool_1t2a8t_1lizzieLet0_4MQNode_4QNode_Bool_7QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_11QNode_Bool_1t3a8u_1Lcall_f3,CTf) > (lizzieLet17_1_1_argbuf,CTf) */
  CTf_t lizzieLet0_4MQNode_4QNode_Bool_4QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_5QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_9QNode_Bool_1t1a8s_1lizzieLet0_4MQNode_4QNode_Bool_6QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_10QNode_Bool_1t2a8t_1lizzieLet0_4MQNode_4QNode_Bool_7QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_11QNode_Bool_1t3a8u_1Lcall_f3_bufchan_d;
  logic lizzieLet0_4MQNode_4QNode_Bool_4QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_5QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_9QNode_Bool_1t1a8s_1lizzieLet0_4MQNode_4QNode_Bool_6QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_10QNode_Bool_1t2a8t_1lizzieLet0_4MQNode_4QNode_Bool_7QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_11QNode_Bool_1t3a8u_1Lcall_f3_bufchan_r;
  assign lizzieLet0_4MQNode_4QNode_Bool_4QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_5QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_9QNode_Bool_1t1a8s_1lizzieLet0_4MQNode_4QNode_Bool_6QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_10QNode_Bool_1t2a8t_1lizzieLet0_4MQNode_4QNode_Bool_7QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_11QNode_Bool_1t3a8u_1Lcall_f3_r = ((! lizzieLet0_4MQNode_4QNode_Bool_4QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_5QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_9QNode_Bool_1t1a8s_1lizzieLet0_4MQNode_4QNode_Bool_6QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_10QNode_Bool_1t2a8t_1lizzieLet0_4MQNode_4QNode_Bool_7QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_11QNode_Bool_1t3a8u_1Lcall_f3_bufchan_d[0]) || lizzieLet0_4MQNode_4QNode_Bool_4QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_5QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_9QNode_Bool_1t1a8s_1lizzieLet0_4MQNode_4QNode_Bool_6QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_10QNode_Bool_1t2a8t_1lizzieLet0_4MQNode_4QNode_Bool_7QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_11QNode_Bool_1t3a8u_1Lcall_f3_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QNode_Bool_4QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_5QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_9QNode_Bool_1t1a8s_1lizzieLet0_4MQNode_4QNode_Bool_6QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_10QNode_Bool_1t2a8t_1lizzieLet0_4MQNode_4QNode_Bool_7QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_11QNode_Bool_1t3a8u_1Lcall_f3_bufchan_d <= {163'd0,
                                                                                                                                                                                                                                                                                                                                                                        1'd0};
    else
      if (lizzieLet0_4MQNode_4QNode_Bool_4QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_5QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_9QNode_Bool_1t1a8s_1lizzieLet0_4MQNode_4QNode_Bool_6QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_10QNode_Bool_1t2a8t_1lizzieLet0_4MQNode_4QNode_Bool_7QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_11QNode_Bool_1t3a8u_1Lcall_f3_r)
        lizzieLet0_4MQNode_4QNode_Bool_4QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_5QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_9QNode_Bool_1t1a8s_1lizzieLet0_4MQNode_4QNode_Bool_6QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_10QNode_Bool_1t2a8t_1lizzieLet0_4MQNode_4QNode_Bool_7QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_11QNode_Bool_1t3a8u_1Lcall_f3_bufchan_d <= lizzieLet0_4MQNode_4QNode_Bool_4QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_5QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_9QNode_Bool_1t1a8s_1lizzieLet0_4MQNode_4QNode_Bool_6QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_10QNode_Bool_1t2a8t_1lizzieLet0_4MQNode_4QNode_Bool_7QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_11QNode_Bool_1t3a8u_1Lcall_f3_d;
  CTf_t lizzieLet0_4MQNode_4QNode_Bool_4QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_5QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_9QNode_Bool_1t1a8s_1lizzieLet0_4MQNode_4QNode_Bool_6QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_10QNode_Bool_1t2a8t_1lizzieLet0_4MQNode_4QNode_Bool_7QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_11QNode_Bool_1t3a8u_1Lcall_f3_bufchan_buf;
  assign lizzieLet0_4MQNode_4QNode_Bool_4QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_5QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_9QNode_Bool_1t1a8s_1lizzieLet0_4MQNode_4QNode_Bool_6QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_10QNode_Bool_1t2a8t_1lizzieLet0_4MQNode_4QNode_Bool_7QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_11QNode_Bool_1t3a8u_1Lcall_f3_bufchan_r = (! lizzieLet0_4MQNode_4QNode_Bool_4QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_5QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_9QNode_Bool_1t1a8s_1lizzieLet0_4MQNode_4QNode_Bool_6QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_10QNode_Bool_1t2a8t_1lizzieLet0_4MQNode_4QNode_Bool_7QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_11QNode_Bool_1t3a8u_1Lcall_f3_bufchan_buf[0]);
  assign lizzieLet17_1_1_argbuf_d = (lizzieLet0_4MQNode_4QNode_Bool_4QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_5QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_9QNode_Bool_1t1a8s_1lizzieLet0_4MQNode_4QNode_Bool_6QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_10QNode_Bool_1t2a8t_1lizzieLet0_4MQNode_4QNode_Bool_7QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_11QNode_Bool_1t3a8u_1Lcall_f3_bufchan_buf[0] ? lizzieLet0_4MQNode_4QNode_Bool_4QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_5QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_9QNode_Bool_1t1a8s_1lizzieLet0_4MQNode_4QNode_Bool_6QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_10QNode_Bool_1t2a8t_1lizzieLet0_4MQNode_4QNode_Bool_7QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_11QNode_Bool_1t3a8u_1Lcall_f3_bufchan_buf :
                                     lizzieLet0_4MQNode_4QNode_Bool_4QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_5QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_9QNode_Bool_1t1a8s_1lizzieLet0_4MQNode_4QNode_Bool_6QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_10QNode_Bool_1t2a8t_1lizzieLet0_4MQNode_4QNode_Bool_7QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_11QNode_Bool_1t3a8u_1Lcall_f3_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QNode_Bool_4QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_5QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_9QNode_Bool_1t1a8s_1lizzieLet0_4MQNode_4QNode_Bool_6QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_10QNode_Bool_1t2a8t_1lizzieLet0_4MQNode_4QNode_Bool_7QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_11QNode_Bool_1t3a8u_1Lcall_f3_bufchan_buf <= {163'd0,
                                                                                                                                                                                                                                                                                                                                                                          1'd0};
    else
      if ((lizzieLet17_1_1_argbuf_r && lizzieLet0_4MQNode_4QNode_Bool_4QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_5QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_9QNode_Bool_1t1a8s_1lizzieLet0_4MQNode_4QNode_Bool_6QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_10QNode_Bool_1t2a8t_1lizzieLet0_4MQNode_4QNode_Bool_7QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_11QNode_Bool_1t3a8u_1Lcall_f3_bufchan_buf[0]))
        lizzieLet0_4MQNode_4QNode_Bool_4QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_5QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_9QNode_Bool_1t1a8s_1lizzieLet0_4MQNode_4QNode_Bool_6QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_10QNode_Bool_1t2a8t_1lizzieLet0_4MQNode_4QNode_Bool_7QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_11QNode_Bool_1t3a8u_1Lcall_f3_bufchan_buf <= {163'd0,
                                                                                                                                                                                                                                                                                                                                                                            1'd0};
      else if (((! lizzieLet17_1_1_argbuf_r) && (! lizzieLet0_4MQNode_4QNode_Bool_4QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_5QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_9QNode_Bool_1t1a8s_1lizzieLet0_4MQNode_4QNode_Bool_6QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_10QNode_Bool_1t2a8t_1lizzieLet0_4MQNode_4QNode_Bool_7QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_11QNode_Bool_1t3a8u_1Lcall_f3_bufchan_buf[0])))
        lizzieLet0_4MQNode_4QNode_Bool_4QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_5QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_9QNode_Bool_1t1a8s_1lizzieLet0_4MQNode_4QNode_Bool_6QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_10QNode_Bool_1t2a8t_1lizzieLet0_4MQNode_4QNode_Bool_7QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_11QNode_Bool_1t3a8u_1Lcall_f3_bufchan_buf <= lizzieLet0_4MQNode_4QNode_Bool_4QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_5QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_9QNode_Bool_1t1a8s_1lizzieLet0_4MQNode_4QNode_Bool_6QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_10QNode_Bool_1t2a8t_1lizzieLet0_4MQNode_4QNode_Bool_7QNode_Bool_1lizzieLet0_4MQNode_4QNode_Bool_11QNode_Bool_1t3a8u_1Lcall_f3_bufchan_d;
  
  /* buf (Ty Pointer_CTf) : (lizzieLet0_4MQNode_4QNode_Bool_4QNone_Bool,Pointer_CTf) > (lizzieLet0_4MQNode_4QNode_Bool_4QNone_Bool_1_argbuf,Pointer_CTf) */
  Pointer_CTf_t lizzieLet0_4MQNode_4QNode_Bool_4QNone_Bool_bufchan_d;
  logic lizzieLet0_4MQNode_4QNode_Bool_4QNone_Bool_bufchan_r;
  assign lizzieLet0_4MQNode_4QNode_Bool_4QNone_Bool_r = ((! lizzieLet0_4MQNode_4QNode_Bool_4QNone_Bool_bufchan_d[0]) || lizzieLet0_4MQNode_4QNode_Bool_4QNone_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QNode_Bool_4QNone_Bool_bufchan_d <= {16'd0,
                                                               1'd0};
    else
      if (lizzieLet0_4MQNode_4QNode_Bool_4QNone_Bool_r)
        lizzieLet0_4MQNode_4QNode_Bool_4QNone_Bool_bufchan_d <= lizzieLet0_4MQNode_4QNode_Bool_4QNone_Bool_d;
  Pointer_CTf_t lizzieLet0_4MQNode_4QNode_Bool_4QNone_Bool_bufchan_buf;
  assign lizzieLet0_4MQNode_4QNode_Bool_4QNone_Bool_bufchan_r = (! lizzieLet0_4MQNode_4QNode_Bool_4QNone_Bool_bufchan_buf[0]);
  assign lizzieLet0_4MQNode_4QNode_Bool_4QNone_Bool_1_argbuf_d = (lizzieLet0_4MQNode_4QNode_Bool_4QNone_Bool_bufchan_buf[0] ? lizzieLet0_4MQNode_4QNode_Bool_4QNone_Bool_bufchan_buf :
                                                                  lizzieLet0_4MQNode_4QNode_Bool_4QNone_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QNode_Bool_4QNone_Bool_bufchan_buf <= {16'd0,
                                                                 1'd0};
    else
      if ((lizzieLet0_4MQNode_4QNode_Bool_4QNone_Bool_1_argbuf_r && lizzieLet0_4MQNode_4QNode_Bool_4QNone_Bool_bufchan_buf[0]))
        lizzieLet0_4MQNode_4QNode_Bool_4QNone_Bool_bufchan_buf <= {16'd0,
                                                                   1'd0};
      else if (((! lizzieLet0_4MQNode_4QNode_Bool_4QNone_Bool_1_argbuf_r) && (! lizzieLet0_4MQNode_4QNode_Bool_4QNone_Bool_bufchan_buf[0])))
        lizzieLet0_4MQNode_4QNode_Bool_4QNone_Bool_bufchan_buf <= lizzieLet0_4MQNode_4QNode_Bool_4QNone_Bool_bufchan_d;
  
  /* buf (Ty Pointer_CTf) : (lizzieLet0_4MQNode_4QNode_Bool_4QVal_Bool,Pointer_CTf) > (lizzieLet0_4MQNode_4QNode_Bool_4QVal_Bool_1_argbuf,Pointer_CTf) */
  Pointer_CTf_t lizzieLet0_4MQNode_4QNode_Bool_4QVal_Bool_bufchan_d;
  logic lizzieLet0_4MQNode_4QNode_Bool_4QVal_Bool_bufchan_r;
  assign lizzieLet0_4MQNode_4QNode_Bool_4QVal_Bool_r = ((! lizzieLet0_4MQNode_4QNode_Bool_4QVal_Bool_bufchan_d[0]) || lizzieLet0_4MQNode_4QNode_Bool_4QVal_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QNode_Bool_4QVal_Bool_bufchan_d <= {16'd0,
                                                              1'd0};
    else
      if (lizzieLet0_4MQNode_4QNode_Bool_4QVal_Bool_r)
        lizzieLet0_4MQNode_4QNode_Bool_4QVal_Bool_bufchan_d <= lizzieLet0_4MQNode_4QNode_Bool_4QVal_Bool_d;
  Pointer_CTf_t lizzieLet0_4MQNode_4QNode_Bool_4QVal_Bool_bufchan_buf;
  assign lizzieLet0_4MQNode_4QNode_Bool_4QVal_Bool_bufchan_r = (! lizzieLet0_4MQNode_4QNode_Bool_4QVal_Bool_bufchan_buf[0]);
  assign lizzieLet0_4MQNode_4QNode_Bool_4QVal_Bool_1_argbuf_d = (lizzieLet0_4MQNode_4QNode_Bool_4QVal_Bool_bufchan_buf[0] ? lizzieLet0_4MQNode_4QNode_Bool_4QVal_Bool_bufchan_buf :
                                                                 lizzieLet0_4MQNode_4QNode_Bool_4QVal_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QNode_Bool_4QVal_Bool_bufchan_buf <= {16'd0,
                                                                1'd0};
    else
      if ((lizzieLet0_4MQNode_4QNode_Bool_4QVal_Bool_1_argbuf_r && lizzieLet0_4MQNode_4QNode_Bool_4QVal_Bool_bufchan_buf[0]))
        lizzieLet0_4MQNode_4QNode_Bool_4QVal_Bool_bufchan_buf <= {16'd0,
                                                                  1'd0};
      else if (((! lizzieLet0_4MQNode_4QNode_Bool_4QVal_Bool_1_argbuf_r) && (! lizzieLet0_4MQNode_4QNode_Bool_4QVal_Bool_bufchan_buf[0])))
        lizzieLet0_4MQNode_4QNode_Bool_4QVal_Bool_bufchan_buf <= lizzieLet0_4MQNode_4QNode_Bool_4QVal_Bool_bufchan_d;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_MaskQTree) : (lizzieLet0_4MQNode_4QNode_Bool_5,QTree_Bool) (lizzieLet0_4MQNode_6QNode_Bool,Pointer_MaskQTree) > [(lizzieLet0_4MQNode_4QNode_Bool_5QNone_Bool,Pointer_MaskQTree),
                                                                                                                                   (_109,Pointer_MaskQTree),
                                                                                                                                   (lizzieLet0_4MQNode_4QNode_Bool_5QNode_Bool,Pointer_MaskQTree),
                                                                                                                                   (_108,Pointer_MaskQTree)] */
  logic [3:0] lizzieLet0_4MQNode_6QNode_Bool_onehotd;
  always_comb
    if ((lizzieLet0_4MQNode_4QNode_Bool_5_d[0] && lizzieLet0_4MQNode_6QNode_Bool_d[0]))
      unique case (lizzieLet0_4MQNode_4QNode_Bool_5_d[2:1])
        2'd0: lizzieLet0_4MQNode_6QNode_Bool_onehotd = 4'd1;
        2'd1: lizzieLet0_4MQNode_6QNode_Bool_onehotd = 4'd2;
        2'd2: lizzieLet0_4MQNode_6QNode_Bool_onehotd = 4'd4;
        2'd3: lizzieLet0_4MQNode_6QNode_Bool_onehotd = 4'd8;
        default: lizzieLet0_4MQNode_6QNode_Bool_onehotd = 4'd0;
      endcase
    else lizzieLet0_4MQNode_6QNode_Bool_onehotd = 4'd0;
  assign lizzieLet0_4MQNode_4QNode_Bool_5QNone_Bool_d = {lizzieLet0_4MQNode_6QNode_Bool_d[16:1],
                                                         lizzieLet0_4MQNode_6QNode_Bool_onehotd[0]};
  assign _109_d = {lizzieLet0_4MQNode_6QNode_Bool_d[16:1],
                   lizzieLet0_4MQNode_6QNode_Bool_onehotd[1]};
  assign lizzieLet0_4MQNode_4QNode_Bool_5QNode_Bool_d = {lizzieLet0_4MQNode_6QNode_Bool_d[16:1],
                                                         lizzieLet0_4MQNode_6QNode_Bool_onehotd[2]};
  assign _108_d = {lizzieLet0_4MQNode_6QNode_Bool_d[16:1],
                   lizzieLet0_4MQNode_6QNode_Bool_onehotd[3]};
  assign lizzieLet0_4MQNode_6QNode_Bool_r = (| (lizzieLet0_4MQNode_6QNode_Bool_onehotd & {_108_r,
                                                                                          lizzieLet0_4MQNode_4QNode_Bool_5QNode_Bool_r,
                                                                                          _109_r,
                                                                                          lizzieLet0_4MQNode_4QNode_Bool_5QNone_Bool_r}));
  assign lizzieLet0_4MQNode_4QNode_Bool_5_r = lizzieLet0_4MQNode_6QNode_Bool_r;
  
  /* buf (Ty Pointer_MaskQTree) : (lizzieLet0_4MQNode_4QNode_Bool_5QNone_Bool,Pointer_MaskQTree) > (lizzieLet0_4MQNode_4QNode_Bool_5QNone_Bool_1_argbuf,Pointer_MaskQTree) */
  Pointer_MaskQTree_t lizzieLet0_4MQNode_4QNode_Bool_5QNone_Bool_bufchan_d;
  logic lizzieLet0_4MQNode_4QNode_Bool_5QNone_Bool_bufchan_r;
  assign lizzieLet0_4MQNode_4QNode_Bool_5QNone_Bool_r = ((! lizzieLet0_4MQNode_4QNode_Bool_5QNone_Bool_bufchan_d[0]) || lizzieLet0_4MQNode_4QNode_Bool_5QNone_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QNode_Bool_5QNone_Bool_bufchan_d <= {16'd0,
                                                               1'd0};
    else
      if (lizzieLet0_4MQNode_4QNode_Bool_5QNone_Bool_r)
        lizzieLet0_4MQNode_4QNode_Bool_5QNone_Bool_bufchan_d <= lizzieLet0_4MQNode_4QNode_Bool_5QNone_Bool_d;
  Pointer_MaskQTree_t lizzieLet0_4MQNode_4QNode_Bool_5QNone_Bool_bufchan_buf;
  assign lizzieLet0_4MQNode_4QNode_Bool_5QNone_Bool_bufchan_r = (! lizzieLet0_4MQNode_4QNode_Bool_5QNone_Bool_bufchan_buf[0]);
  assign lizzieLet0_4MQNode_4QNode_Bool_5QNone_Bool_1_argbuf_d = (lizzieLet0_4MQNode_4QNode_Bool_5QNone_Bool_bufchan_buf[0] ? lizzieLet0_4MQNode_4QNode_Bool_5QNone_Bool_bufchan_buf :
                                                                  lizzieLet0_4MQNode_4QNode_Bool_5QNone_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QNode_Bool_5QNone_Bool_bufchan_buf <= {16'd0,
                                                                 1'd0};
    else
      if ((lizzieLet0_4MQNode_4QNode_Bool_5QNone_Bool_1_argbuf_r && lizzieLet0_4MQNode_4QNode_Bool_5QNone_Bool_bufchan_buf[0]))
        lizzieLet0_4MQNode_4QNode_Bool_5QNone_Bool_bufchan_buf <= {16'd0,
                                                                   1'd0};
      else if (((! lizzieLet0_4MQNode_4QNode_Bool_5QNone_Bool_1_argbuf_r) && (! lizzieLet0_4MQNode_4QNode_Bool_5QNone_Bool_bufchan_buf[0])))
        lizzieLet0_4MQNode_4QNode_Bool_5QNone_Bool_bufchan_buf <= lizzieLet0_4MQNode_4QNode_Bool_5QNone_Bool_bufchan_d;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_MaskQTree) : (lizzieLet0_4MQNode_4QNode_Bool_6,QTree_Bool) (lizzieLet0_4MQNode_7QNode_Bool,Pointer_MaskQTree) > [(lizzieLet0_4MQNode_4QNode_Bool_6QNone_Bool,Pointer_MaskQTree),
                                                                                                                                   (_107,Pointer_MaskQTree),
                                                                                                                                   (lizzieLet0_4MQNode_4QNode_Bool_6QNode_Bool,Pointer_MaskQTree),
                                                                                                                                   (_106,Pointer_MaskQTree)] */
  logic [3:0] lizzieLet0_4MQNode_7QNode_Bool_onehotd;
  always_comb
    if ((lizzieLet0_4MQNode_4QNode_Bool_6_d[0] && lizzieLet0_4MQNode_7QNode_Bool_d[0]))
      unique case (lizzieLet0_4MQNode_4QNode_Bool_6_d[2:1])
        2'd0: lizzieLet0_4MQNode_7QNode_Bool_onehotd = 4'd1;
        2'd1: lizzieLet0_4MQNode_7QNode_Bool_onehotd = 4'd2;
        2'd2: lizzieLet0_4MQNode_7QNode_Bool_onehotd = 4'd4;
        2'd3: lizzieLet0_4MQNode_7QNode_Bool_onehotd = 4'd8;
        default: lizzieLet0_4MQNode_7QNode_Bool_onehotd = 4'd0;
      endcase
    else lizzieLet0_4MQNode_7QNode_Bool_onehotd = 4'd0;
  assign lizzieLet0_4MQNode_4QNode_Bool_6QNone_Bool_d = {lizzieLet0_4MQNode_7QNode_Bool_d[16:1],
                                                         lizzieLet0_4MQNode_7QNode_Bool_onehotd[0]};
  assign _107_d = {lizzieLet0_4MQNode_7QNode_Bool_d[16:1],
                   lizzieLet0_4MQNode_7QNode_Bool_onehotd[1]};
  assign lizzieLet0_4MQNode_4QNode_Bool_6QNode_Bool_d = {lizzieLet0_4MQNode_7QNode_Bool_d[16:1],
                                                         lizzieLet0_4MQNode_7QNode_Bool_onehotd[2]};
  assign _106_d = {lizzieLet0_4MQNode_7QNode_Bool_d[16:1],
                   lizzieLet0_4MQNode_7QNode_Bool_onehotd[3]};
  assign lizzieLet0_4MQNode_7QNode_Bool_r = (| (lizzieLet0_4MQNode_7QNode_Bool_onehotd & {_106_r,
                                                                                          lizzieLet0_4MQNode_4QNode_Bool_6QNode_Bool_r,
                                                                                          _107_r,
                                                                                          lizzieLet0_4MQNode_4QNode_Bool_6QNone_Bool_r}));
  assign lizzieLet0_4MQNode_4QNode_Bool_6_r = lizzieLet0_4MQNode_7QNode_Bool_r;
  
  /* buf (Ty Pointer_MaskQTree) : (lizzieLet0_4MQNode_4QNode_Bool_6QNone_Bool,Pointer_MaskQTree) > (lizzieLet0_4MQNode_4QNode_Bool_6QNone_Bool_1_argbuf,Pointer_MaskQTree) */
  Pointer_MaskQTree_t lizzieLet0_4MQNode_4QNode_Bool_6QNone_Bool_bufchan_d;
  logic lizzieLet0_4MQNode_4QNode_Bool_6QNone_Bool_bufchan_r;
  assign lizzieLet0_4MQNode_4QNode_Bool_6QNone_Bool_r = ((! lizzieLet0_4MQNode_4QNode_Bool_6QNone_Bool_bufchan_d[0]) || lizzieLet0_4MQNode_4QNode_Bool_6QNone_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QNode_Bool_6QNone_Bool_bufchan_d <= {16'd0,
                                                               1'd0};
    else
      if (lizzieLet0_4MQNode_4QNode_Bool_6QNone_Bool_r)
        lizzieLet0_4MQNode_4QNode_Bool_6QNone_Bool_bufchan_d <= lizzieLet0_4MQNode_4QNode_Bool_6QNone_Bool_d;
  Pointer_MaskQTree_t lizzieLet0_4MQNode_4QNode_Bool_6QNone_Bool_bufchan_buf;
  assign lizzieLet0_4MQNode_4QNode_Bool_6QNone_Bool_bufchan_r = (! lizzieLet0_4MQNode_4QNode_Bool_6QNone_Bool_bufchan_buf[0]);
  assign lizzieLet0_4MQNode_4QNode_Bool_6QNone_Bool_1_argbuf_d = (lizzieLet0_4MQNode_4QNode_Bool_6QNone_Bool_bufchan_buf[0] ? lizzieLet0_4MQNode_4QNode_Bool_6QNone_Bool_bufchan_buf :
                                                                  lizzieLet0_4MQNode_4QNode_Bool_6QNone_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QNode_Bool_6QNone_Bool_bufchan_buf <= {16'd0,
                                                                 1'd0};
    else
      if ((lizzieLet0_4MQNode_4QNode_Bool_6QNone_Bool_1_argbuf_r && lizzieLet0_4MQNode_4QNode_Bool_6QNone_Bool_bufchan_buf[0]))
        lizzieLet0_4MQNode_4QNode_Bool_6QNone_Bool_bufchan_buf <= {16'd0,
                                                                   1'd0};
      else if (((! lizzieLet0_4MQNode_4QNode_Bool_6QNone_Bool_1_argbuf_r) && (! lizzieLet0_4MQNode_4QNode_Bool_6QNone_Bool_bufchan_buf[0])))
        lizzieLet0_4MQNode_4QNode_Bool_6QNone_Bool_bufchan_buf <= lizzieLet0_4MQNode_4QNode_Bool_6QNone_Bool_bufchan_d;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_MaskQTree) : (lizzieLet0_4MQNode_4QNode_Bool_7,QTree_Bool) (lizzieLet0_4MQNode_8QNode_Bool,Pointer_MaskQTree) > [(lizzieLet0_4MQNode_4QNode_Bool_7QNone_Bool,Pointer_MaskQTree),
                                                                                                                                   (_105,Pointer_MaskQTree),
                                                                                                                                   (lizzieLet0_4MQNode_4QNode_Bool_7QNode_Bool,Pointer_MaskQTree),
                                                                                                                                   (_104,Pointer_MaskQTree)] */
  logic [3:0] lizzieLet0_4MQNode_8QNode_Bool_onehotd;
  always_comb
    if ((lizzieLet0_4MQNode_4QNode_Bool_7_d[0] && lizzieLet0_4MQNode_8QNode_Bool_d[0]))
      unique case (lizzieLet0_4MQNode_4QNode_Bool_7_d[2:1])
        2'd0: lizzieLet0_4MQNode_8QNode_Bool_onehotd = 4'd1;
        2'd1: lizzieLet0_4MQNode_8QNode_Bool_onehotd = 4'd2;
        2'd2: lizzieLet0_4MQNode_8QNode_Bool_onehotd = 4'd4;
        2'd3: lizzieLet0_4MQNode_8QNode_Bool_onehotd = 4'd8;
        default: lizzieLet0_4MQNode_8QNode_Bool_onehotd = 4'd0;
      endcase
    else lizzieLet0_4MQNode_8QNode_Bool_onehotd = 4'd0;
  assign lizzieLet0_4MQNode_4QNode_Bool_7QNone_Bool_d = {lizzieLet0_4MQNode_8QNode_Bool_d[16:1],
                                                         lizzieLet0_4MQNode_8QNode_Bool_onehotd[0]};
  assign _105_d = {lizzieLet0_4MQNode_8QNode_Bool_d[16:1],
                   lizzieLet0_4MQNode_8QNode_Bool_onehotd[1]};
  assign lizzieLet0_4MQNode_4QNode_Bool_7QNode_Bool_d = {lizzieLet0_4MQNode_8QNode_Bool_d[16:1],
                                                         lizzieLet0_4MQNode_8QNode_Bool_onehotd[2]};
  assign _104_d = {lizzieLet0_4MQNode_8QNode_Bool_d[16:1],
                   lizzieLet0_4MQNode_8QNode_Bool_onehotd[3]};
  assign lizzieLet0_4MQNode_8QNode_Bool_r = (| (lizzieLet0_4MQNode_8QNode_Bool_onehotd & {_104_r,
                                                                                          lizzieLet0_4MQNode_4QNode_Bool_7QNode_Bool_r,
                                                                                          _105_r,
                                                                                          lizzieLet0_4MQNode_4QNode_Bool_7QNone_Bool_r}));
  assign lizzieLet0_4MQNode_4QNode_Bool_7_r = lizzieLet0_4MQNode_8QNode_Bool_r;
  
  /* buf (Ty Pointer_MaskQTree) : (lizzieLet0_4MQNode_4QNode_Bool_7QNone_Bool,Pointer_MaskQTree) > (lizzieLet0_4MQNode_4QNode_Bool_7QNone_Bool_1_argbuf,Pointer_MaskQTree) */
  Pointer_MaskQTree_t lizzieLet0_4MQNode_4QNode_Bool_7QNone_Bool_bufchan_d;
  logic lizzieLet0_4MQNode_4QNode_Bool_7QNone_Bool_bufchan_r;
  assign lizzieLet0_4MQNode_4QNode_Bool_7QNone_Bool_r = ((! lizzieLet0_4MQNode_4QNode_Bool_7QNone_Bool_bufchan_d[0]) || lizzieLet0_4MQNode_4QNode_Bool_7QNone_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QNode_Bool_7QNone_Bool_bufchan_d <= {16'd0,
                                                               1'd0};
    else
      if (lizzieLet0_4MQNode_4QNode_Bool_7QNone_Bool_r)
        lizzieLet0_4MQNode_4QNode_Bool_7QNone_Bool_bufchan_d <= lizzieLet0_4MQNode_4QNode_Bool_7QNone_Bool_d;
  Pointer_MaskQTree_t lizzieLet0_4MQNode_4QNode_Bool_7QNone_Bool_bufchan_buf;
  assign lizzieLet0_4MQNode_4QNode_Bool_7QNone_Bool_bufchan_r = (! lizzieLet0_4MQNode_4QNode_Bool_7QNone_Bool_bufchan_buf[0]);
  assign lizzieLet0_4MQNode_4QNode_Bool_7QNone_Bool_1_argbuf_d = (lizzieLet0_4MQNode_4QNode_Bool_7QNone_Bool_bufchan_buf[0] ? lizzieLet0_4MQNode_4QNode_Bool_7QNone_Bool_bufchan_buf :
                                                                  lizzieLet0_4MQNode_4QNode_Bool_7QNone_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QNode_Bool_7QNone_Bool_bufchan_buf <= {16'd0,
                                                                 1'd0};
    else
      if ((lizzieLet0_4MQNode_4QNode_Bool_7QNone_Bool_1_argbuf_r && lizzieLet0_4MQNode_4QNode_Bool_7QNone_Bool_bufchan_buf[0]))
        lizzieLet0_4MQNode_4QNode_Bool_7QNone_Bool_bufchan_buf <= {16'd0,
                                                                   1'd0};
      else if (((! lizzieLet0_4MQNode_4QNode_Bool_7QNone_Bool_1_argbuf_r) && (! lizzieLet0_4MQNode_4QNode_Bool_7QNone_Bool_bufchan_buf[0])))
        lizzieLet0_4MQNode_4QNode_Bool_7QNone_Bool_bufchan_buf <= lizzieLet0_4MQNode_4QNode_Bool_7QNone_Bool_bufchan_d;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_MaskQTree) : (lizzieLet0_4MQNode_4QNode_Bool_8,QTree_Bool) (lizzieLet0_4MQNode_9QNode_Bool,Pointer_MaskQTree) > [(lizzieLet0_4MQNode_4QNode_Bool_8QNone_Bool,Pointer_MaskQTree),
                                                                                                                                   (_103,Pointer_MaskQTree),
                                                                                                                                   (lizzieLet0_4MQNode_4QNode_Bool_8QNode_Bool,Pointer_MaskQTree),
                                                                                                                                   (_102,Pointer_MaskQTree)] */
  logic [3:0] lizzieLet0_4MQNode_9QNode_Bool_onehotd;
  always_comb
    if ((lizzieLet0_4MQNode_4QNode_Bool_8_d[0] && lizzieLet0_4MQNode_9QNode_Bool_d[0]))
      unique case (lizzieLet0_4MQNode_4QNode_Bool_8_d[2:1])
        2'd0: lizzieLet0_4MQNode_9QNode_Bool_onehotd = 4'd1;
        2'd1: lizzieLet0_4MQNode_9QNode_Bool_onehotd = 4'd2;
        2'd2: lizzieLet0_4MQNode_9QNode_Bool_onehotd = 4'd4;
        2'd3: lizzieLet0_4MQNode_9QNode_Bool_onehotd = 4'd8;
        default: lizzieLet0_4MQNode_9QNode_Bool_onehotd = 4'd0;
      endcase
    else lizzieLet0_4MQNode_9QNode_Bool_onehotd = 4'd0;
  assign lizzieLet0_4MQNode_4QNode_Bool_8QNone_Bool_d = {lizzieLet0_4MQNode_9QNode_Bool_d[16:1],
                                                         lizzieLet0_4MQNode_9QNode_Bool_onehotd[0]};
  assign _103_d = {lizzieLet0_4MQNode_9QNode_Bool_d[16:1],
                   lizzieLet0_4MQNode_9QNode_Bool_onehotd[1]};
  assign lizzieLet0_4MQNode_4QNode_Bool_8QNode_Bool_d = {lizzieLet0_4MQNode_9QNode_Bool_d[16:1],
                                                         lizzieLet0_4MQNode_9QNode_Bool_onehotd[2]};
  assign _102_d = {lizzieLet0_4MQNode_9QNode_Bool_d[16:1],
                   lizzieLet0_4MQNode_9QNode_Bool_onehotd[3]};
  assign lizzieLet0_4MQNode_9QNode_Bool_r = (| (lizzieLet0_4MQNode_9QNode_Bool_onehotd & {_102_r,
                                                                                          lizzieLet0_4MQNode_4QNode_Bool_8QNode_Bool_r,
                                                                                          _103_r,
                                                                                          lizzieLet0_4MQNode_4QNode_Bool_8QNone_Bool_r}));
  assign lizzieLet0_4MQNode_4QNode_Bool_8_r = lizzieLet0_4MQNode_9QNode_Bool_r;
  
  /* buf (Ty Pointer_MaskQTree) : (lizzieLet0_4MQNode_4QNode_Bool_8QNode_Bool,Pointer_MaskQTree) > (lizzieLet0_4MQNode_4QNode_Bool_8QNode_Bool_1_argbuf,Pointer_MaskQTree) */
  Pointer_MaskQTree_t lizzieLet0_4MQNode_4QNode_Bool_8QNode_Bool_bufchan_d;
  logic lizzieLet0_4MQNode_4QNode_Bool_8QNode_Bool_bufchan_r;
  assign lizzieLet0_4MQNode_4QNode_Bool_8QNode_Bool_r = ((! lizzieLet0_4MQNode_4QNode_Bool_8QNode_Bool_bufchan_d[0]) || lizzieLet0_4MQNode_4QNode_Bool_8QNode_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QNode_Bool_8QNode_Bool_bufchan_d <= {16'd0,
                                                               1'd0};
    else
      if (lizzieLet0_4MQNode_4QNode_Bool_8QNode_Bool_r)
        lizzieLet0_4MQNode_4QNode_Bool_8QNode_Bool_bufchan_d <= lizzieLet0_4MQNode_4QNode_Bool_8QNode_Bool_d;
  Pointer_MaskQTree_t lizzieLet0_4MQNode_4QNode_Bool_8QNode_Bool_bufchan_buf;
  assign lizzieLet0_4MQNode_4QNode_Bool_8QNode_Bool_bufchan_r = (! lizzieLet0_4MQNode_4QNode_Bool_8QNode_Bool_bufchan_buf[0]);
  assign lizzieLet0_4MQNode_4QNode_Bool_8QNode_Bool_1_argbuf_d = (lizzieLet0_4MQNode_4QNode_Bool_8QNode_Bool_bufchan_buf[0] ? lizzieLet0_4MQNode_4QNode_Bool_8QNode_Bool_bufchan_buf :
                                                                  lizzieLet0_4MQNode_4QNode_Bool_8QNode_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QNode_Bool_8QNode_Bool_bufchan_buf <= {16'd0,
                                                                 1'd0};
    else
      if ((lizzieLet0_4MQNode_4QNode_Bool_8QNode_Bool_1_argbuf_r && lizzieLet0_4MQNode_4QNode_Bool_8QNode_Bool_bufchan_buf[0]))
        lizzieLet0_4MQNode_4QNode_Bool_8QNode_Bool_bufchan_buf <= {16'd0,
                                                                   1'd0};
      else if (((! lizzieLet0_4MQNode_4QNode_Bool_8QNode_Bool_1_argbuf_r) && (! lizzieLet0_4MQNode_4QNode_Bool_8QNode_Bool_bufchan_buf[0])))
        lizzieLet0_4MQNode_4QNode_Bool_8QNode_Bool_bufchan_buf <= lizzieLet0_4MQNode_4QNode_Bool_8QNode_Bool_bufchan_d;
  
  /* buf (Ty Pointer_MaskQTree) : (lizzieLet0_4MQNode_4QNode_Bool_8QNone_Bool,Pointer_MaskQTree) > (lizzieLet0_4MQNode_4QNode_Bool_8QNone_Bool_1_argbuf,Pointer_MaskQTree) */
  Pointer_MaskQTree_t lizzieLet0_4MQNode_4QNode_Bool_8QNone_Bool_bufchan_d;
  logic lizzieLet0_4MQNode_4QNode_Bool_8QNone_Bool_bufchan_r;
  assign lizzieLet0_4MQNode_4QNode_Bool_8QNone_Bool_r = ((! lizzieLet0_4MQNode_4QNode_Bool_8QNone_Bool_bufchan_d[0]) || lizzieLet0_4MQNode_4QNode_Bool_8QNone_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QNode_Bool_8QNone_Bool_bufchan_d <= {16'd0,
                                                               1'd0};
    else
      if (lizzieLet0_4MQNode_4QNode_Bool_8QNone_Bool_r)
        lizzieLet0_4MQNode_4QNode_Bool_8QNone_Bool_bufchan_d <= lizzieLet0_4MQNode_4QNode_Bool_8QNone_Bool_d;
  Pointer_MaskQTree_t lizzieLet0_4MQNode_4QNode_Bool_8QNone_Bool_bufchan_buf;
  assign lizzieLet0_4MQNode_4QNode_Bool_8QNone_Bool_bufchan_r = (! lizzieLet0_4MQNode_4QNode_Bool_8QNone_Bool_bufchan_buf[0]);
  assign lizzieLet0_4MQNode_4QNode_Bool_8QNone_Bool_1_argbuf_d = (lizzieLet0_4MQNode_4QNode_Bool_8QNone_Bool_bufchan_buf[0] ? lizzieLet0_4MQNode_4QNode_Bool_8QNone_Bool_bufchan_buf :
                                                                  lizzieLet0_4MQNode_4QNode_Bool_8QNone_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QNode_Bool_8QNone_Bool_bufchan_buf <= {16'd0,
                                                                 1'd0};
    else
      if ((lizzieLet0_4MQNode_4QNode_Bool_8QNone_Bool_1_argbuf_r && lizzieLet0_4MQNode_4QNode_Bool_8QNone_Bool_bufchan_buf[0]))
        lizzieLet0_4MQNode_4QNode_Bool_8QNone_Bool_bufchan_buf <= {16'd0,
                                                                   1'd0};
      else if (((! lizzieLet0_4MQNode_4QNode_Bool_8QNone_Bool_1_argbuf_r) && (! lizzieLet0_4MQNode_4QNode_Bool_8QNone_Bool_bufchan_buf[0])))
        lizzieLet0_4MQNode_4QNode_Bool_8QNone_Bool_bufchan_buf <= lizzieLet0_4MQNode_4QNode_Bool_8QNone_Bool_bufchan_d;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_QTree_Bool) : (lizzieLet0_4MQNode_4QNode_Bool_9,QTree_Bool) (q1'a8n_destruct,Pointer_QTree_Bool) > [(lizzieLet0_4MQNode_4QNode_Bool_9QNone_Bool,Pointer_QTree_Bool),
                                                                                                                      (_101,Pointer_QTree_Bool),
                                                                                                                      (lizzieLet0_4MQNode_4QNode_Bool_9QNode_Bool,Pointer_QTree_Bool),
                                                                                                                      (_100,Pointer_QTree_Bool)] */
  logic [3:0] \q1'a8n_destruct_onehotd ;
  always_comb
    if ((lizzieLet0_4MQNode_4QNode_Bool_9_d[0] && \q1'a8n_destruct_d [0]))
      unique case (lizzieLet0_4MQNode_4QNode_Bool_9_d[2:1])
        2'd0: \q1'a8n_destruct_onehotd  = 4'd1;
        2'd1: \q1'a8n_destruct_onehotd  = 4'd2;
        2'd2: \q1'a8n_destruct_onehotd  = 4'd4;
        2'd3: \q1'a8n_destruct_onehotd  = 4'd8;
        default: \q1'a8n_destruct_onehotd  = 4'd0;
      endcase
    else \q1'a8n_destruct_onehotd  = 4'd0;
  assign lizzieLet0_4MQNode_4QNode_Bool_9QNone_Bool_d = {\q1'a8n_destruct_d [16:1],
                                                         \q1'a8n_destruct_onehotd [0]};
  assign _101_d = {\q1'a8n_destruct_d [16:1],
                   \q1'a8n_destruct_onehotd [1]};
  assign lizzieLet0_4MQNode_4QNode_Bool_9QNode_Bool_d = {\q1'a8n_destruct_d [16:1],
                                                         \q1'a8n_destruct_onehotd [2]};
  assign _100_d = {\q1'a8n_destruct_d [16:1],
                   \q1'a8n_destruct_onehotd [3]};
  assign \q1'a8n_destruct_r  = (| (\q1'a8n_destruct_onehotd  & {_100_r,
                                                                lizzieLet0_4MQNode_4QNode_Bool_9QNode_Bool_r,
                                                                _101_r,
                                                                lizzieLet0_4MQNode_4QNode_Bool_9QNone_Bool_r}));
  assign lizzieLet0_4MQNode_4QNode_Bool_9_r = \q1'a8n_destruct_r ;
  
  /* buf (Ty Pointer_QTree_Bool) : (lizzieLet0_4MQNode_4QNode_Bool_9QNone_Bool,Pointer_QTree_Bool) > (lizzieLet0_4MQNode_4QNode_Bool_9QNone_Bool_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t lizzieLet0_4MQNode_4QNode_Bool_9QNone_Bool_bufchan_d;
  logic lizzieLet0_4MQNode_4QNode_Bool_9QNone_Bool_bufchan_r;
  assign lizzieLet0_4MQNode_4QNode_Bool_9QNone_Bool_r = ((! lizzieLet0_4MQNode_4QNode_Bool_9QNone_Bool_bufchan_d[0]) || lizzieLet0_4MQNode_4QNode_Bool_9QNone_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QNode_Bool_9QNone_Bool_bufchan_d <= {16'd0,
                                                               1'd0};
    else
      if (lizzieLet0_4MQNode_4QNode_Bool_9QNone_Bool_r)
        lizzieLet0_4MQNode_4QNode_Bool_9QNone_Bool_bufchan_d <= lizzieLet0_4MQNode_4QNode_Bool_9QNone_Bool_d;
  Pointer_QTree_Bool_t lizzieLet0_4MQNode_4QNode_Bool_9QNone_Bool_bufchan_buf;
  assign lizzieLet0_4MQNode_4QNode_Bool_9QNone_Bool_bufchan_r = (! lizzieLet0_4MQNode_4QNode_Bool_9QNone_Bool_bufchan_buf[0]);
  assign lizzieLet0_4MQNode_4QNode_Bool_9QNone_Bool_1_argbuf_d = (lizzieLet0_4MQNode_4QNode_Bool_9QNone_Bool_bufchan_buf[0] ? lizzieLet0_4MQNode_4QNode_Bool_9QNone_Bool_bufchan_buf :
                                                                  lizzieLet0_4MQNode_4QNode_Bool_9QNone_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QNode_Bool_9QNone_Bool_bufchan_buf <= {16'd0,
                                                                 1'd0};
    else
      if ((lizzieLet0_4MQNode_4QNode_Bool_9QNone_Bool_1_argbuf_r && lizzieLet0_4MQNode_4QNode_Bool_9QNone_Bool_bufchan_buf[0]))
        lizzieLet0_4MQNode_4QNode_Bool_9QNone_Bool_bufchan_buf <= {16'd0,
                                                                   1'd0};
      else if (((! lizzieLet0_4MQNode_4QNode_Bool_9QNone_Bool_1_argbuf_r) && (! lizzieLet0_4MQNode_4QNode_Bool_9QNone_Bool_bufchan_buf[0])))
        lizzieLet0_4MQNode_4QNode_Bool_9QNone_Bool_bufchan_buf <= lizzieLet0_4MQNode_4QNode_Bool_9QNone_Bool_bufchan_d;
  
  /* fork (Ty QTree_Bool) : (lizzieLet0_4MQNode_4QNone_Bool,QTree_Bool) > [(lizzieLet0_4MQNode_4QNone_Bool_1,QTree_Bool),
                                                                      (lizzieLet0_4MQNode_4QNone_Bool_2,QTree_Bool),
                                                                      (lizzieLet0_4MQNode_4QNone_Bool_3,QTree_Bool),
                                                                      (lizzieLet0_4MQNode_4QNone_Bool_4,QTree_Bool),
                                                                      (lizzieLet0_4MQNode_4QNone_Bool_5,QTree_Bool),
                                                                      (lizzieLet0_4MQNode_4QNone_Bool_6,QTree_Bool),
                                                                      (lizzieLet0_4MQNode_4QNone_Bool_7,QTree_Bool),
                                                                      (lizzieLet0_4MQNode_4QNone_Bool_8,QTree_Bool)] */
  logic [7:0] lizzieLet0_4MQNode_4QNone_Bool_emitted;
  logic [7:0] lizzieLet0_4MQNode_4QNone_Bool_done;
  assign lizzieLet0_4MQNode_4QNone_Bool_1_d = {lizzieLet0_4MQNode_4QNone_Bool_d[66:1],
                                               (lizzieLet0_4MQNode_4QNone_Bool_d[0] && (! lizzieLet0_4MQNode_4QNone_Bool_emitted[0]))};
  assign lizzieLet0_4MQNode_4QNone_Bool_2_d = {lizzieLet0_4MQNode_4QNone_Bool_d[66:1],
                                               (lizzieLet0_4MQNode_4QNone_Bool_d[0] && (! lizzieLet0_4MQNode_4QNone_Bool_emitted[1]))};
  assign lizzieLet0_4MQNode_4QNone_Bool_3_d = {lizzieLet0_4MQNode_4QNone_Bool_d[66:1],
                                               (lizzieLet0_4MQNode_4QNone_Bool_d[0] && (! lizzieLet0_4MQNode_4QNone_Bool_emitted[2]))};
  assign lizzieLet0_4MQNode_4QNone_Bool_4_d = {lizzieLet0_4MQNode_4QNone_Bool_d[66:1],
                                               (lizzieLet0_4MQNode_4QNone_Bool_d[0] && (! lizzieLet0_4MQNode_4QNone_Bool_emitted[3]))};
  assign lizzieLet0_4MQNode_4QNone_Bool_5_d = {lizzieLet0_4MQNode_4QNone_Bool_d[66:1],
                                               (lizzieLet0_4MQNode_4QNone_Bool_d[0] && (! lizzieLet0_4MQNode_4QNone_Bool_emitted[4]))};
  assign lizzieLet0_4MQNode_4QNone_Bool_6_d = {lizzieLet0_4MQNode_4QNone_Bool_d[66:1],
                                               (lizzieLet0_4MQNode_4QNone_Bool_d[0] && (! lizzieLet0_4MQNode_4QNone_Bool_emitted[5]))};
  assign lizzieLet0_4MQNode_4QNone_Bool_7_d = {lizzieLet0_4MQNode_4QNone_Bool_d[66:1],
                                               (lizzieLet0_4MQNode_4QNone_Bool_d[0] && (! lizzieLet0_4MQNode_4QNone_Bool_emitted[6]))};
  assign lizzieLet0_4MQNode_4QNone_Bool_8_d = {lizzieLet0_4MQNode_4QNone_Bool_d[66:1],
                                               (lizzieLet0_4MQNode_4QNone_Bool_d[0] && (! lizzieLet0_4MQNode_4QNone_Bool_emitted[7]))};
  assign lizzieLet0_4MQNode_4QNone_Bool_done = (lizzieLet0_4MQNode_4QNone_Bool_emitted | ({lizzieLet0_4MQNode_4QNone_Bool_8_d[0],
                                                                                           lizzieLet0_4MQNode_4QNone_Bool_7_d[0],
                                                                                           lizzieLet0_4MQNode_4QNone_Bool_6_d[0],
                                                                                           lizzieLet0_4MQNode_4QNone_Bool_5_d[0],
                                                                                           lizzieLet0_4MQNode_4QNone_Bool_4_d[0],
                                                                                           lizzieLet0_4MQNode_4QNone_Bool_3_d[0],
                                                                                           lizzieLet0_4MQNode_4QNone_Bool_2_d[0],
                                                                                           lizzieLet0_4MQNode_4QNone_Bool_1_d[0]} & {lizzieLet0_4MQNode_4QNone_Bool_8_r,
                                                                                                                                     lizzieLet0_4MQNode_4QNone_Bool_7_r,
                                                                                                                                     lizzieLet0_4MQNode_4QNone_Bool_6_r,
                                                                                                                                     lizzieLet0_4MQNode_4QNone_Bool_5_r,
                                                                                                                                     lizzieLet0_4MQNode_4QNone_Bool_4_r,
                                                                                                                                     lizzieLet0_4MQNode_4QNone_Bool_3_r,
                                                                                                                                     lizzieLet0_4MQNode_4QNone_Bool_2_r,
                                                                                                                                     lizzieLet0_4MQNode_4QNone_Bool_1_r}));
  assign lizzieLet0_4MQNode_4QNone_Bool_r = (& lizzieLet0_4MQNode_4QNone_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QNone_Bool_emitted <= 8'd0;
    else
      lizzieLet0_4MQNode_4QNone_Bool_emitted <= (lizzieLet0_4MQNode_4QNone_Bool_r ? 8'd0 :
                                                 lizzieLet0_4MQNode_4QNone_Bool_done);
  
  /* destruct (Ty QTree_Bool,
          Dcon QNode_Bool) : (lizzieLet0_4MQNode_4QNone_Bool_1QNode_Bool,QTree_Bool) > [(t1a8d_destruct,Pointer_QTree_Bool),
                                                                                        (t2a8e_destruct,Pointer_QTree_Bool),
                                                                                        (t3a8f_destruct,Pointer_QTree_Bool),
                                                                                        (t4a8g_destruct,Pointer_QTree_Bool)] */
  logic [3:0] lizzieLet0_4MQNode_4QNone_Bool_1QNode_Bool_emitted;
  logic [3:0] lizzieLet0_4MQNode_4QNone_Bool_1QNode_Bool_done;
  assign t1a8d_destruct_d = {lizzieLet0_4MQNode_4QNone_Bool_1QNode_Bool_d[18:3],
                             (lizzieLet0_4MQNode_4QNone_Bool_1QNode_Bool_d[0] && (! lizzieLet0_4MQNode_4QNone_Bool_1QNode_Bool_emitted[0]))};
  assign t2a8e_destruct_d = {lizzieLet0_4MQNode_4QNone_Bool_1QNode_Bool_d[34:19],
                             (lizzieLet0_4MQNode_4QNone_Bool_1QNode_Bool_d[0] && (! lizzieLet0_4MQNode_4QNone_Bool_1QNode_Bool_emitted[1]))};
  assign t3a8f_destruct_d = {lizzieLet0_4MQNode_4QNone_Bool_1QNode_Bool_d[50:35],
                             (lizzieLet0_4MQNode_4QNone_Bool_1QNode_Bool_d[0] && (! lizzieLet0_4MQNode_4QNone_Bool_1QNode_Bool_emitted[2]))};
  assign t4a8g_destruct_d = {lizzieLet0_4MQNode_4QNone_Bool_1QNode_Bool_d[66:51],
                             (lizzieLet0_4MQNode_4QNone_Bool_1QNode_Bool_d[0] && (! lizzieLet0_4MQNode_4QNone_Bool_1QNode_Bool_emitted[3]))};
  assign lizzieLet0_4MQNode_4QNone_Bool_1QNode_Bool_done = (lizzieLet0_4MQNode_4QNone_Bool_1QNode_Bool_emitted | ({t4a8g_destruct_d[0],
                                                                                                                   t3a8f_destruct_d[0],
                                                                                                                   t2a8e_destruct_d[0],
                                                                                                                   t1a8d_destruct_d[0]} & {t4a8g_destruct_r,
                                                                                                                                           t3a8f_destruct_r,
                                                                                                                                           t2a8e_destruct_r,
                                                                                                                                           t1a8d_destruct_r}));
  assign lizzieLet0_4MQNode_4QNone_Bool_1QNode_Bool_r = (& lizzieLet0_4MQNode_4QNone_Bool_1QNode_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QNone_Bool_1QNode_Bool_emitted <= 4'd0;
    else
      lizzieLet0_4MQNode_4QNone_Bool_1QNode_Bool_emitted <= (lizzieLet0_4MQNode_4QNone_Bool_1QNode_Bool_r ? 4'd0 :
                                                             lizzieLet0_4MQNode_4QNone_Bool_1QNode_Bool_done);
  
  /* demux (Ty QTree_Bool,
       Ty QTree_Bool) : (lizzieLet0_4MQNode_4QNone_Bool_2,QTree_Bool) (lizzieLet0_4MQNode_4QNone_Bool_1,QTree_Bool) > [(_99,QTree_Bool),
                                                                                                                       (_98,QTree_Bool),
                                                                                                                       (lizzieLet0_4MQNode_4QNone_Bool_1QNode_Bool,QTree_Bool),
                                                                                                                       (_97,QTree_Bool)] */
  logic [3:0] lizzieLet0_4MQNode_4QNone_Bool_1_onehotd;
  always_comb
    if ((lizzieLet0_4MQNode_4QNone_Bool_2_d[0] && lizzieLet0_4MQNode_4QNone_Bool_1_d[0]))
      unique case (lizzieLet0_4MQNode_4QNone_Bool_2_d[2:1])
        2'd0: lizzieLet0_4MQNode_4QNone_Bool_1_onehotd = 4'd1;
        2'd1: lizzieLet0_4MQNode_4QNone_Bool_1_onehotd = 4'd2;
        2'd2: lizzieLet0_4MQNode_4QNone_Bool_1_onehotd = 4'd4;
        2'd3: lizzieLet0_4MQNode_4QNone_Bool_1_onehotd = 4'd8;
        default: lizzieLet0_4MQNode_4QNone_Bool_1_onehotd = 4'd0;
      endcase
    else lizzieLet0_4MQNode_4QNone_Bool_1_onehotd = 4'd0;
  assign _99_d = {lizzieLet0_4MQNode_4QNone_Bool_1_d[66:1],
                  lizzieLet0_4MQNode_4QNone_Bool_1_onehotd[0]};
  assign _98_d = {lizzieLet0_4MQNode_4QNone_Bool_1_d[66:1],
                  lizzieLet0_4MQNode_4QNone_Bool_1_onehotd[1]};
  assign lizzieLet0_4MQNode_4QNone_Bool_1QNode_Bool_d = {lizzieLet0_4MQNode_4QNone_Bool_1_d[66:1],
                                                         lizzieLet0_4MQNode_4QNone_Bool_1_onehotd[2]};
  assign _97_d = {lizzieLet0_4MQNode_4QNone_Bool_1_d[66:1],
                  lizzieLet0_4MQNode_4QNone_Bool_1_onehotd[3]};
  assign lizzieLet0_4MQNode_4QNone_Bool_1_r = (| (lizzieLet0_4MQNode_4QNone_Bool_1_onehotd & {_97_r,
                                                                                              lizzieLet0_4MQNode_4QNone_Bool_1QNode_Bool_r,
                                                                                              _98_r,
                                                                                              _99_r}));
  assign lizzieLet0_4MQNode_4QNone_Bool_2_r = lizzieLet0_4MQNode_4QNone_Bool_1_r;
  
  /* demux (Ty QTree_Bool,
       Ty Go) : (lizzieLet0_4MQNode_4QNone_Bool_3,QTree_Bool) (lizzieLet0_4MQNode_3QNone_Bool,Go) > [(lizzieLet0_4MQNode_4QNone_Bool_3QNone_Bool,Go),
                                                                                                     (lizzieLet0_4MQNode_4QNone_Bool_3QVal_Bool,Go),
                                                                                                     (lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool,Go),
                                                                                                     (lizzieLet0_4MQNode_4QNone_Bool_3QError_Bool,Go)] */
  logic [3:0] lizzieLet0_4MQNode_3QNone_Bool_onehotd;
  always_comb
    if ((lizzieLet0_4MQNode_4QNone_Bool_3_d[0] && lizzieLet0_4MQNode_3QNone_Bool_d[0]))
      unique case (lizzieLet0_4MQNode_4QNone_Bool_3_d[2:1])
        2'd0: lizzieLet0_4MQNode_3QNone_Bool_onehotd = 4'd1;
        2'd1: lizzieLet0_4MQNode_3QNone_Bool_onehotd = 4'd2;
        2'd2: lizzieLet0_4MQNode_3QNone_Bool_onehotd = 4'd4;
        2'd3: lizzieLet0_4MQNode_3QNone_Bool_onehotd = 4'd8;
        default: lizzieLet0_4MQNode_3QNone_Bool_onehotd = 4'd0;
      endcase
    else lizzieLet0_4MQNode_3QNone_Bool_onehotd = 4'd0;
  assign lizzieLet0_4MQNode_4QNone_Bool_3QNone_Bool_d = lizzieLet0_4MQNode_3QNone_Bool_onehotd[0];
  assign lizzieLet0_4MQNode_4QNone_Bool_3QVal_Bool_d = lizzieLet0_4MQNode_3QNone_Bool_onehotd[1];
  assign lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_d = lizzieLet0_4MQNode_3QNone_Bool_onehotd[2];
  assign lizzieLet0_4MQNode_4QNone_Bool_3QError_Bool_d = lizzieLet0_4MQNode_3QNone_Bool_onehotd[3];
  assign lizzieLet0_4MQNode_3QNone_Bool_r = (| (lizzieLet0_4MQNode_3QNone_Bool_onehotd & {lizzieLet0_4MQNode_4QNone_Bool_3QError_Bool_r,
                                                                                          lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_r,
                                                                                          lizzieLet0_4MQNode_4QNone_Bool_3QVal_Bool_r,
                                                                                          lizzieLet0_4MQNode_4QNone_Bool_3QNone_Bool_r}));
  assign lizzieLet0_4MQNode_4QNone_Bool_3_r = lizzieLet0_4MQNode_3QNone_Bool_r;
  
  /* fork (Ty Go) : (lizzieLet0_4MQNode_4QNone_Bool_3QError_Bool,Go) > [(lizzieLet0_4MQNode_4QNone_Bool_3QError_Bool_1,Go),
                                                                   (lizzieLet0_4MQNode_4QNone_Bool_3QError_Bool_2,Go)] */
  logic [1:0] lizzieLet0_4MQNode_4QNone_Bool_3QError_Bool_emitted;
  logic [1:0] lizzieLet0_4MQNode_4QNone_Bool_3QError_Bool_done;
  assign lizzieLet0_4MQNode_4QNone_Bool_3QError_Bool_1_d = (lizzieLet0_4MQNode_4QNone_Bool_3QError_Bool_d[0] && (! lizzieLet0_4MQNode_4QNone_Bool_3QError_Bool_emitted[0]));
  assign lizzieLet0_4MQNode_4QNone_Bool_3QError_Bool_2_d = (lizzieLet0_4MQNode_4QNone_Bool_3QError_Bool_d[0] && (! lizzieLet0_4MQNode_4QNone_Bool_3QError_Bool_emitted[1]));
  assign lizzieLet0_4MQNode_4QNone_Bool_3QError_Bool_done = (lizzieLet0_4MQNode_4QNone_Bool_3QError_Bool_emitted | ({lizzieLet0_4MQNode_4QNone_Bool_3QError_Bool_2_d[0],
                                                                                                                     lizzieLet0_4MQNode_4QNone_Bool_3QError_Bool_1_d[0]} & {lizzieLet0_4MQNode_4QNone_Bool_3QError_Bool_2_r,
                                                                                                                                                                            lizzieLet0_4MQNode_4QNone_Bool_3QError_Bool_1_r}));
  assign lizzieLet0_4MQNode_4QNone_Bool_3QError_Bool_r = (& lizzieLet0_4MQNode_4QNone_Bool_3QError_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QNone_Bool_3QError_Bool_emitted <= 2'd0;
    else
      lizzieLet0_4MQNode_4QNone_Bool_3QError_Bool_emitted <= (lizzieLet0_4MQNode_4QNone_Bool_3QError_Bool_r ? 2'd0 :
                                                              lizzieLet0_4MQNode_4QNone_Bool_3QError_Bool_done);
  
  /* dcon (Ty QTree_Bool,
      Dcon QError_Bool) : [(lizzieLet0_4MQNode_4QNone_Bool_3QError_Bool_1,Go)] > (lizzieLet0_4MQNode_4QNone_Bool_3QError_Bool_1QError_Bool,QTree_Bool) */
  assign lizzieLet0_4MQNode_4QNone_Bool_3QError_Bool_1QError_Bool_d = QError_Bool_dc((& {lizzieLet0_4MQNode_4QNone_Bool_3QError_Bool_1_d[0]}), lizzieLet0_4MQNode_4QNone_Bool_3QError_Bool_1_d);
  assign {lizzieLet0_4MQNode_4QNone_Bool_3QError_Bool_1_r} = {1 {(lizzieLet0_4MQNode_4QNone_Bool_3QError_Bool_1QError_Bool_r && lizzieLet0_4MQNode_4QNone_Bool_3QError_Bool_1QError_Bool_d[0])}};
  
  /* buf (Ty QTree_Bool) : (lizzieLet0_4MQNode_4QNone_Bool_3QError_Bool_1QError_Bool,QTree_Bool) > (lizzieLet7_1_argbuf,QTree_Bool) */
  QTree_Bool_t lizzieLet0_4MQNode_4QNone_Bool_3QError_Bool_1QError_Bool_bufchan_d;
  logic lizzieLet0_4MQNode_4QNone_Bool_3QError_Bool_1QError_Bool_bufchan_r;
  assign lizzieLet0_4MQNode_4QNone_Bool_3QError_Bool_1QError_Bool_r = ((! lizzieLet0_4MQNode_4QNone_Bool_3QError_Bool_1QError_Bool_bufchan_d[0]) || lizzieLet0_4MQNode_4QNone_Bool_3QError_Bool_1QError_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QNone_Bool_3QError_Bool_1QError_Bool_bufchan_d <= {66'd0,
                                                                             1'd0};
    else
      if (lizzieLet0_4MQNode_4QNone_Bool_3QError_Bool_1QError_Bool_r)
        lizzieLet0_4MQNode_4QNone_Bool_3QError_Bool_1QError_Bool_bufchan_d <= lizzieLet0_4MQNode_4QNone_Bool_3QError_Bool_1QError_Bool_d;
  QTree_Bool_t lizzieLet0_4MQNode_4QNone_Bool_3QError_Bool_1QError_Bool_bufchan_buf;
  assign lizzieLet0_4MQNode_4QNone_Bool_3QError_Bool_1QError_Bool_bufchan_r = (! lizzieLet0_4MQNode_4QNone_Bool_3QError_Bool_1QError_Bool_bufchan_buf[0]);
  assign lizzieLet7_1_argbuf_d = (lizzieLet0_4MQNode_4QNone_Bool_3QError_Bool_1QError_Bool_bufchan_buf[0] ? lizzieLet0_4MQNode_4QNone_Bool_3QError_Bool_1QError_Bool_bufchan_buf :
                                  lizzieLet0_4MQNode_4QNone_Bool_3QError_Bool_1QError_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QNone_Bool_3QError_Bool_1QError_Bool_bufchan_buf <= {66'd0,
                                                                               1'd0};
    else
      if ((lizzieLet7_1_argbuf_r && lizzieLet0_4MQNode_4QNone_Bool_3QError_Bool_1QError_Bool_bufchan_buf[0]))
        lizzieLet0_4MQNode_4QNone_Bool_3QError_Bool_1QError_Bool_bufchan_buf <= {66'd0,
                                                                                 1'd0};
      else if (((! lizzieLet7_1_argbuf_r) && (! lizzieLet0_4MQNode_4QNone_Bool_3QError_Bool_1QError_Bool_bufchan_buf[0])))
        lizzieLet0_4MQNode_4QNone_Bool_3QError_Bool_1QError_Bool_bufchan_buf <= lizzieLet0_4MQNode_4QNone_Bool_3QError_Bool_1QError_Bool_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet0_4MQNode_4QNone_Bool_3QError_Bool_2,Go) > (lizzieLet0_4MQNode_4QNone_Bool_3QError_Bool_2_argbuf,Go) */
  Go_t lizzieLet0_4MQNode_4QNone_Bool_3QError_Bool_2_bufchan_d;
  logic lizzieLet0_4MQNode_4QNone_Bool_3QError_Bool_2_bufchan_r;
  assign lizzieLet0_4MQNode_4QNone_Bool_3QError_Bool_2_r = ((! lizzieLet0_4MQNode_4QNone_Bool_3QError_Bool_2_bufchan_d[0]) || lizzieLet0_4MQNode_4QNone_Bool_3QError_Bool_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QNone_Bool_3QError_Bool_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet0_4MQNode_4QNone_Bool_3QError_Bool_2_r)
        lizzieLet0_4MQNode_4QNone_Bool_3QError_Bool_2_bufchan_d <= lizzieLet0_4MQNode_4QNone_Bool_3QError_Bool_2_d;
  Go_t lizzieLet0_4MQNode_4QNone_Bool_3QError_Bool_2_bufchan_buf;
  assign lizzieLet0_4MQNode_4QNone_Bool_3QError_Bool_2_bufchan_r = (! lizzieLet0_4MQNode_4QNone_Bool_3QError_Bool_2_bufchan_buf[0]);
  assign lizzieLet0_4MQNode_4QNone_Bool_3QError_Bool_2_argbuf_d = (lizzieLet0_4MQNode_4QNone_Bool_3QError_Bool_2_bufchan_buf[0] ? lizzieLet0_4MQNode_4QNone_Bool_3QError_Bool_2_bufchan_buf :
                                                                   lizzieLet0_4MQNode_4QNone_Bool_3QError_Bool_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QNone_Bool_3QError_Bool_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet0_4MQNode_4QNone_Bool_3QError_Bool_2_argbuf_r && lizzieLet0_4MQNode_4QNone_Bool_3QError_Bool_2_bufchan_buf[0]))
        lizzieLet0_4MQNode_4QNone_Bool_3QError_Bool_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet0_4MQNode_4QNone_Bool_3QError_Bool_2_argbuf_r) && (! lizzieLet0_4MQNode_4QNone_Bool_3QError_Bool_2_bufchan_buf[0])))
        lizzieLet0_4MQNode_4QNone_Bool_3QError_Bool_2_bufchan_buf <= lizzieLet0_4MQNode_4QNone_Bool_3QError_Bool_2_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool,Go) > [(lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_1,Go),
                                                                  (lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_2,Go),
                                                                  (lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_3,Go),
                                                                  (lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_4,Go),
                                                                  (lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_5,Go)] */
  logic [4:0] lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_emitted;
  logic [4:0] lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_done;
  assign lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_1_d = (lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_d[0] && (! lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_emitted[0]));
  assign lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_2_d = (lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_d[0] && (! lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_emitted[1]));
  assign lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_3_d = (lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_d[0] && (! lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_emitted[2]));
  assign lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_4_d = (lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_d[0] && (! lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_emitted[3]));
  assign lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_5_d = (lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_d[0] && (! lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_emitted[4]));
  assign lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_done = (lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_emitted | ({lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_5_d[0],
                                                                                                                   lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_4_d[0],
                                                                                                                   lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_3_d[0],
                                                                                                                   lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_2_d[0],
                                                                                                                   lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_1_d[0]} & {lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_5_r,
                                                                                                                                                                         lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_4_r,
                                                                                                                                                                         lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_3_r,
                                                                                                                                                                         lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_2_r,
                                                                                                                                                                         lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_1_r}));
  assign lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_r = (& lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_emitted <= 5'd0;
    else
      lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_emitted <= (lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_r ? 5'd0 :
                                                             lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_done);
  
  /* buf (Ty Go) : (lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_1,Go) > (lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_1_argbuf,Go) */
  Go_t lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_1_bufchan_d;
  logic lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_1_bufchan_r;
  assign lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_1_r = ((! lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_1_bufchan_d[0]) || lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_1_bufchan_d <= 1'd0;
    else
      if (lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_1_r)
        lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_1_bufchan_d <= lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_1_d;
  Go_t lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_1_bufchan_buf;
  assign lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_1_bufchan_r = (! lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_1_bufchan_buf[0]);
  assign lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_1_argbuf_d = (lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_1_bufchan_buf[0] ? lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_1_bufchan_buf :
                                                                  lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_1_argbuf_r && lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_1_bufchan_buf[0]))
        lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_1_argbuf_r) && (! lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_1_bufchan_buf[0])))
        lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_1_bufchan_buf <= lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_1_bufchan_d;
  
  /* dcon (Ty TupGo___Pointer_MaskQTree___Pointer_QTree_Bool,
      Dcon TupGo___Pointer_MaskQTree___Pointer_QTree_Bool) : [(lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_1_argbuf,Go),
                                                              (lizzieLet0_4MQNode_4QNone_Bool_8QNode_Bool_1_argbuf,Pointer_MaskQTree),
                                                              (t4a8g_1_argbuf,Pointer_QTree_Bool)] > (f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool_1,TupGo___Pointer_MaskQTree___Pointer_QTree_Bool) */
  assign \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool_1_d  = TupGo___Pointer_MaskQTree___Pointer_QTree_Bool_dc((& {lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_1_argbuf_d[0],
                                                                                                                                                lizzieLet0_4MQNode_4QNone_Bool_8QNode_Bool_1_argbuf_d[0],
                                                                                                                                                t4a8g_1_argbuf_d[0]}), lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_1_argbuf_d, lizzieLet0_4MQNode_4QNone_Bool_8QNode_Bool_1_argbuf_d, t4a8g_1_argbuf_d);
  assign {lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_1_argbuf_r,
          lizzieLet0_4MQNode_4QNone_Bool_8QNode_Bool_1_argbuf_r,
          t4a8g_1_argbuf_r} = {3 {(\f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool_1_r  && \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool_1_d [0])}};
  
  /* buf (Ty Go) : (lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_2,Go) > (lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_2_argbuf,Go) */
  Go_t lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_2_bufchan_d;
  logic lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_2_bufchan_r;
  assign lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_2_r = ((! lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_2_bufchan_d[0]) || lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_2_r)
        lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_2_bufchan_d <= lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_2_d;
  Go_t lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_2_bufchan_buf;
  assign lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_2_bufchan_r = (! lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_2_bufchan_buf[0]);
  assign lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_2_argbuf_d = (lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_2_bufchan_buf[0] ? lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_2_bufchan_buf :
                                                                  lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_2_argbuf_r && lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_2_bufchan_buf[0]))
        lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_2_argbuf_r) && (! lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_2_bufchan_buf[0])))
        lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_2_bufchan_buf <= lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_2_bufchan_d;
  
  /* dcon (Ty TupGo___Pointer_MaskQTree___Pointer_QTree_Bool,
      Dcon TupGo___Pointer_MaskQTree___Pointer_QTree_Bool) : [(lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_2_argbuf,Go),
                                                              (lizzieLet0_4MQNode_4QNone_Bool_7QNode_Bool_1_argbuf,Pointer_MaskQTree),
                                                              (t3a8f_1_argbuf,Pointer_QTree_Bool)] > (f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool2,TupGo___Pointer_MaskQTree___Pointer_QTree_Bool) */
  assign \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool2_d  = TupGo___Pointer_MaskQTree___Pointer_QTree_Bool_dc((& {lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_2_argbuf_d[0],
                                                                                                                                               lizzieLet0_4MQNode_4QNone_Bool_7QNode_Bool_1_argbuf_d[0],
                                                                                                                                               t3a8f_1_argbuf_d[0]}), lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_2_argbuf_d, lizzieLet0_4MQNode_4QNone_Bool_7QNode_Bool_1_argbuf_d, t3a8f_1_argbuf_d);
  assign {lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_2_argbuf_r,
          lizzieLet0_4MQNode_4QNone_Bool_7QNode_Bool_1_argbuf_r,
          t3a8f_1_argbuf_r} = {3 {(\f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool2_r  && \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool2_d [0])}};
  
  /* buf (Ty Go) : (lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_3,Go) > (lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_3_argbuf,Go) */
  Go_t lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_3_bufchan_d;
  logic lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_3_bufchan_r;
  assign lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_3_r = ((! lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_3_bufchan_d[0]) || lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_3_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_3_bufchan_d <= 1'd0;
    else
      if (lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_3_r)
        lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_3_bufchan_d <= lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_3_d;
  Go_t lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_3_bufchan_buf;
  assign lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_3_bufchan_r = (! lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_3_bufchan_buf[0]);
  assign lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_3_argbuf_d = (lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_3_bufchan_buf[0] ? lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_3_bufchan_buf :
                                                                  lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_3_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_3_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_3_argbuf_r && lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_3_bufchan_buf[0]))
        lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_3_bufchan_buf <= 1'd0;
      else if (((! lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_3_argbuf_r) && (! lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_3_bufchan_buf[0])))
        lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_3_bufchan_buf <= lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_3_bufchan_d;
  
  /* dcon (Ty TupGo___Pointer_MaskQTree___Pointer_QTree_Bool,
      Dcon TupGo___Pointer_MaskQTree___Pointer_QTree_Bool) : [(lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_3_argbuf,Go),
                                                              (lizzieLet0_4MQNode_4QNone_Bool_6QNode_Bool_1_argbuf,Pointer_MaskQTree),
                                                              (t2a8e_1_argbuf,Pointer_QTree_Bool)] > (f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool3,TupGo___Pointer_MaskQTree___Pointer_QTree_Bool) */
  assign \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool3_d  = TupGo___Pointer_MaskQTree___Pointer_QTree_Bool_dc((& {lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_3_argbuf_d[0],
                                                                                                                                               lizzieLet0_4MQNode_4QNone_Bool_6QNode_Bool_1_argbuf_d[0],
                                                                                                                                               t2a8e_1_argbuf_d[0]}), lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_3_argbuf_d, lizzieLet0_4MQNode_4QNone_Bool_6QNode_Bool_1_argbuf_d, t2a8e_1_argbuf_d);
  assign {lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_3_argbuf_r,
          lizzieLet0_4MQNode_4QNone_Bool_6QNode_Bool_1_argbuf_r,
          t2a8e_1_argbuf_r} = {3 {(\f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool3_r  && \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool3_d [0])}};
  
  /* buf (Ty Go) : (lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_4,Go) > (lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_4_argbuf,Go) */
  Go_t lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_4_bufchan_d;
  logic lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_4_bufchan_r;
  assign lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_4_r = ((! lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_4_bufchan_d[0]) || lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_4_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_4_bufchan_d <= 1'd0;
    else
      if (lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_4_r)
        lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_4_bufchan_d <= lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_4_d;
  Go_t lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_4_bufchan_buf;
  assign lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_4_bufchan_r = (! lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_4_bufchan_buf[0]);
  assign lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_4_argbuf_d = (lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_4_bufchan_buf[0] ? lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_4_bufchan_buf :
                                                                  lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_4_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_4_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_4_argbuf_r && lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_4_bufchan_buf[0]))
        lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_4_bufchan_buf <= 1'd0;
      else if (((! lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_4_argbuf_r) && (! lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_4_bufchan_buf[0])))
        lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_4_bufchan_buf <= lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_4_bufchan_d;
  
  /* dcon (Ty TupGo___Pointer_MaskQTree___Pointer_QTree_Bool,
      Dcon TupGo___Pointer_MaskQTree___Pointer_QTree_Bool) : [(lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_4_argbuf,Go),
                                                              (lizzieLet0_4MQNode_4QNone_Bool_5QNode_Bool_1_argbuf,Pointer_MaskQTree),
                                                              (t1a8d_1_argbuf,Pointer_QTree_Bool)] > (f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool4,TupGo___Pointer_MaskQTree___Pointer_QTree_Bool) */
  assign \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool4_d  = TupGo___Pointer_MaskQTree___Pointer_QTree_Bool_dc((& {lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_4_argbuf_d[0],
                                                                                                                                               lizzieLet0_4MQNode_4QNone_Bool_5QNode_Bool_1_argbuf_d[0],
                                                                                                                                               t1a8d_1_argbuf_d[0]}), lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_4_argbuf_d, lizzieLet0_4MQNode_4QNone_Bool_5QNode_Bool_1_argbuf_d, t1a8d_1_argbuf_d);
  assign {lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_4_argbuf_r,
          lizzieLet0_4MQNode_4QNone_Bool_5QNode_Bool_1_argbuf_r,
          t1a8d_1_argbuf_r} = {3 {(\f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool4_r  && \f'''''''''_f'''''''''_BoolTupGo___Pointer_MaskQTree___Pointer_QTree_Bool4_d [0])}};
  
  /* buf (Ty Go) : (lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_5,Go) > (lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_5_argbuf,Go) */
  Go_t lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_5_bufchan_d;
  logic lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_5_bufchan_r;
  assign lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_5_r = ((! lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_5_bufchan_d[0]) || lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_5_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_5_bufchan_d <= 1'd0;
    else
      if (lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_5_r)
        lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_5_bufchan_d <= lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_5_d;
  Go_t lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_5_bufchan_buf;
  assign lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_5_bufchan_r = (! lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_5_bufchan_buf[0]);
  assign lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_5_argbuf_d = (lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_5_bufchan_buf[0] ? lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_5_bufchan_buf :
                                                                  lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_5_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_5_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_5_argbuf_r && lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_5_bufchan_buf[0]))
        lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_5_bufchan_buf <= 1'd0;
      else if (((! lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_5_argbuf_r) && (! lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_5_bufchan_buf[0])))
        lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_5_bufchan_buf <= lizzieLet0_4MQNode_4QNone_Bool_3QNode_Bool_5_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet0_4MQNode_4QNone_Bool_3QNone_Bool,Go) > [(lizzieLet0_4MQNode_4QNone_Bool_3QNone_Bool_1,Go),
                                                                  (lizzieLet0_4MQNode_4QNone_Bool_3QNone_Bool_2,Go)] */
  logic [1:0] lizzieLet0_4MQNode_4QNone_Bool_3QNone_Bool_emitted;
  logic [1:0] lizzieLet0_4MQNode_4QNone_Bool_3QNone_Bool_done;
  assign lizzieLet0_4MQNode_4QNone_Bool_3QNone_Bool_1_d = (lizzieLet0_4MQNode_4QNone_Bool_3QNone_Bool_d[0] && (! lizzieLet0_4MQNode_4QNone_Bool_3QNone_Bool_emitted[0]));
  assign lizzieLet0_4MQNode_4QNone_Bool_3QNone_Bool_2_d = (lizzieLet0_4MQNode_4QNone_Bool_3QNone_Bool_d[0] && (! lizzieLet0_4MQNode_4QNone_Bool_3QNone_Bool_emitted[1]));
  assign lizzieLet0_4MQNode_4QNone_Bool_3QNone_Bool_done = (lizzieLet0_4MQNode_4QNone_Bool_3QNone_Bool_emitted | ({lizzieLet0_4MQNode_4QNone_Bool_3QNone_Bool_2_d[0],
                                                                                                                   lizzieLet0_4MQNode_4QNone_Bool_3QNone_Bool_1_d[0]} & {lizzieLet0_4MQNode_4QNone_Bool_3QNone_Bool_2_r,
                                                                                                                                                                         lizzieLet0_4MQNode_4QNone_Bool_3QNone_Bool_1_r}));
  assign lizzieLet0_4MQNode_4QNone_Bool_3QNone_Bool_r = (& lizzieLet0_4MQNode_4QNone_Bool_3QNone_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QNone_Bool_3QNone_Bool_emitted <= 2'd0;
    else
      lizzieLet0_4MQNode_4QNone_Bool_3QNone_Bool_emitted <= (lizzieLet0_4MQNode_4QNone_Bool_3QNone_Bool_r ? 2'd0 :
                                                             lizzieLet0_4MQNode_4QNone_Bool_3QNone_Bool_done);
  
  /* dcon (Ty QTree_Bool,
      Dcon QNone_Bool) : [(lizzieLet0_4MQNode_4QNone_Bool_3QNone_Bool_1,Go)] > (lizzieLet0_4MQNode_4QNone_Bool_3QNone_Bool_1QNone_Bool,QTree_Bool) */
  assign lizzieLet0_4MQNode_4QNone_Bool_3QNone_Bool_1QNone_Bool_d = QNone_Bool_dc((& {lizzieLet0_4MQNode_4QNone_Bool_3QNone_Bool_1_d[0]}), lizzieLet0_4MQNode_4QNone_Bool_3QNone_Bool_1_d);
  assign {lizzieLet0_4MQNode_4QNone_Bool_3QNone_Bool_1_r} = {1 {(lizzieLet0_4MQNode_4QNone_Bool_3QNone_Bool_1QNone_Bool_r && lizzieLet0_4MQNode_4QNone_Bool_3QNone_Bool_1QNone_Bool_d[0])}};
  
  /* buf (Ty QTree_Bool) : (lizzieLet0_4MQNode_4QNone_Bool_3QNone_Bool_1QNone_Bool,QTree_Bool) > (lizzieLet4_1_argbuf,QTree_Bool) */
  QTree_Bool_t lizzieLet0_4MQNode_4QNone_Bool_3QNone_Bool_1QNone_Bool_bufchan_d;
  logic lizzieLet0_4MQNode_4QNone_Bool_3QNone_Bool_1QNone_Bool_bufchan_r;
  assign lizzieLet0_4MQNode_4QNone_Bool_3QNone_Bool_1QNone_Bool_r = ((! lizzieLet0_4MQNode_4QNone_Bool_3QNone_Bool_1QNone_Bool_bufchan_d[0]) || lizzieLet0_4MQNode_4QNone_Bool_3QNone_Bool_1QNone_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QNone_Bool_3QNone_Bool_1QNone_Bool_bufchan_d <= {66'd0,
                                                                           1'd0};
    else
      if (lizzieLet0_4MQNode_4QNone_Bool_3QNone_Bool_1QNone_Bool_r)
        lizzieLet0_4MQNode_4QNone_Bool_3QNone_Bool_1QNone_Bool_bufchan_d <= lizzieLet0_4MQNode_4QNone_Bool_3QNone_Bool_1QNone_Bool_d;
  QTree_Bool_t lizzieLet0_4MQNode_4QNone_Bool_3QNone_Bool_1QNone_Bool_bufchan_buf;
  assign lizzieLet0_4MQNode_4QNone_Bool_3QNone_Bool_1QNone_Bool_bufchan_r = (! lizzieLet0_4MQNode_4QNone_Bool_3QNone_Bool_1QNone_Bool_bufchan_buf[0]);
  assign lizzieLet4_1_argbuf_d = (lizzieLet0_4MQNode_4QNone_Bool_3QNone_Bool_1QNone_Bool_bufchan_buf[0] ? lizzieLet0_4MQNode_4QNone_Bool_3QNone_Bool_1QNone_Bool_bufchan_buf :
                                  lizzieLet0_4MQNode_4QNone_Bool_3QNone_Bool_1QNone_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QNone_Bool_3QNone_Bool_1QNone_Bool_bufchan_buf <= {66'd0,
                                                                             1'd0};
    else
      if ((lizzieLet4_1_argbuf_r && lizzieLet0_4MQNode_4QNone_Bool_3QNone_Bool_1QNone_Bool_bufchan_buf[0]))
        lizzieLet0_4MQNode_4QNone_Bool_3QNone_Bool_1QNone_Bool_bufchan_buf <= {66'd0,
                                                                               1'd0};
      else if (((! lizzieLet4_1_argbuf_r) && (! lizzieLet0_4MQNode_4QNone_Bool_3QNone_Bool_1QNone_Bool_bufchan_buf[0])))
        lizzieLet0_4MQNode_4QNone_Bool_3QNone_Bool_1QNone_Bool_bufchan_buf <= lizzieLet0_4MQNode_4QNone_Bool_3QNone_Bool_1QNone_Bool_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet0_4MQNode_4QNone_Bool_3QNone_Bool_2,Go) > (lizzieLet0_4MQNode_4QNone_Bool_3QNone_Bool_2_argbuf,Go) */
  Go_t lizzieLet0_4MQNode_4QNone_Bool_3QNone_Bool_2_bufchan_d;
  logic lizzieLet0_4MQNode_4QNone_Bool_3QNone_Bool_2_bufchan_r;
  assign lizzieLet0_4MQNode_4QNone_Bool_3QNone_Bool_2_r = ((! lizzieLet0_4MQNode_4QNone_Bool_3QNone_Bool_2_bufchan_d[0]) || lizzieLet0_4MQNode_4QNone_Bool_3QNone_Bool_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QNone_Bool_3QNone_Bool_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet0_4MQNode_4QNone_Bool_3QNone_Bool_2_r)
        lizzieLet0_4MQNode_4QNone_Bool_3QNone_Bool_2_bufchan_d <= lizzieLet0_4MQNode_4QNone_Bool_3QNone_Bool_2_d;
  Go_t lizzieLet0_4MQNode_4QNone_Bool_3QNone_Bool_2_bufchan_buf;
  assign lizzieLet0_4MQNode_4QNone_Bool_3QNone_Bool_2_bufchan_r = (! lizzieLet0_4MQNode_4QNone_Bool_3QNone_Bool_2_bufchan_buf[0]);
  assign lizzieLet0_4MQNode_4QNone_Bool_3QNone_Bool_2_argbuf_d = (lizzieLet0_4MQNode_4QNone_Bool_3QNone_Bool_2_bufchan_buf[0] ? lizzieLet0_4MQNode_4QNone_Bool_3QNone_Bool_2_bufchan_buf :
                                                                  lizzieLet0_4MQNode_4QNone_Bool_3QNone_Bool_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QNone_Bool_3QNone_Bool_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet0_4MQNode_4QNone_Bool_3QNone_Bool_2_argbuf_r && lizzieLet0_4MQNode_4QNone_Bool_3QNone_Bool_2_bufchan_buf[0]))
        lizzieLet0_4MQNode_4QNone_Bool_3QNone_Bool_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet0_4MQNode_4QNone_Bool_3QNone_Bool_2_argbuf_r) && (! lizzieLet0_4MQNode_4QNone_Bool_3QNone_Bool_2_bufchan_buf[0])))
        lizzieLet0_4MQNode_4QNone_Bool_3QNone_Bool_2_bufchan_buf <= lizzieLet0_4MQNode_4QNone_Bool_3QNone_Bool_2_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet0_4MQNode_4QNone_Bool_3QVal_Bool,Go) > [(lizzieLet0_4MQNode_4QNone_Bool_3QVal_Bool_1,Go),
                                                                 (lizzieLet0_4MQNode_4QNone_Bool_3QVal_Bool_2,Go)] */
  logic [1:0] lizzieLet0_4MQNode_4QNone_Bool_3QVal_Bool_emitted;
  logic [1:0] lizzieLet0_4MQNode_4QNone_Bool_3QVal_Bool_done;
  assign lizzieLet0_4MQNode_4QNone_Bool_3QVal_Bool_1_d = (lizzieLet0_4MQNode_4QNone_Bool_3QVal_Bool_d[0] && (! lizzieLet0_4MQNode_4QNone_Bool_3QVal_Bool_emitted[0]));
  assign lizzieLet0_4MQNode_4QNone_Bool_3QVal_Bool_2_d = (lizzieLet0_4MQNode_4QNone_Bool_3QVal_Bool_d[0] && (! lizzieLet0_4MQNode_4QNone_Bool_3QVal_Bool_emitted[1]));
  assign lizzieLet0_4MQNode_4QNone_Bool_3QVal_Bool_done = (lizzieLet0_4MQNode_4QNone_Bool_3QVal_Bool_emitted | ({lizzieLet0_4MQNode_4QNone_Bool_3QVal_Bool_2_d[0],
                                                                                                                 lizzieLet0_4MQNode_4QNone_Bool_3QVal_Bool_1_d[0]} & {lizzieLet0_4MQNode_4QNone_Bool_3QVal_Bool_2_r,
                                                                                                                                                                      lizzieLet0_4MQNode_4QNone_Bool_3QVal_Bool_1_r}));
  assign lizzieLet0_4MQNode_4QNone_Bool_3QVal_Bool_r = (& lizzieLet0_4MQNode_4QNone_Bool_3QVal_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QNone_Bool_3QVal_Bool_emitted <= 2'd0;
    else
      lizzieLet0_4MQNode_4QNone_Bool_3QVal_Bool_emitted <= (lizzieLet0_4MQNode_4QNone_Bool_3QVal_Bool_r ? 2'd0 :
                                                            lizzieLet0_4MQNode_4QNone_Bool_3QVal_Bool_done);
  
  /* dcon (Ty QTree_Bool,
      Dcon QError_Bool) : [(lizzieLet0_4MQNode_4QNone_Bool_3QVal_Bool_1,Go)] > (lizzieLet0_4MQNode_4QNone_Bool_3QVal_Bool_1QError_Bool,QTree_Bool) */
  assign lizzieLet0_4MQNode_4QNone_Bool_3QVal_Bool_1QError_Bool_d = QError_Bool_dc((& {lizzieLet0_4MQNode_4QNone_Bool_3QVal_Bool_1_d[0]}), lizzieLet0_4MQNode_4QNone_Bool_3QVal_Bool_1_d);
  assign {lizzieLet0_4MQNode_4QNone_Bool_3QVal_Bool_1_r} = {1 {(lizzieLet0_4MQNode_4QNone_Bool_3QVal_Bool_1QError_Bool_r && lizzieLet0_4MQNode_4QNone_Bool_3QVal_Bool_1QError_Bool_d[0])}};
  
  /* buf (Ty QTree_Bool) : (lizzieLet0_4MQNode_4QNone_Bool_3QVal_Bool_1QError_Bool,QTree_Bool) > (lizzieLet5_1_argbuf,QTree_Bool) */
  QTree_Bool_t lizzieLet0_4MQNode_4QNone_Bool_3QVal_Bool_1QError_Bool_bufchan_d;
  logic lizzieLet0_4MQNode_4QNone_Bool_3QVal_Bool_1QError_Bool_bufchan_r;
  assign lizzieLet0_4MQNode_4QNone_Bool_3QVal_Bool_1QError_Bool_r = ((! lizzieLet0_4MQNode_4QNone_Bool_3QVal_Bool_1QError_Bool_bufchan_d[0]) || lizzieLet0_4MQNode_4QNone_Bool_3QVal_Bool_1QError_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QNone_Bool_3QVal_Bool_1QError_Bool_bufchan_d <= {66'd0,
                                                                           1'd0};
    else
      if (lizzieLet0_4MQNode_4QNone_Bool_3QVal_Bool_1QError_Bool_r)
        lizzieLet0_4MQNode_4QNone_Bool_3QVal_Bool_1QError_Bool_bufchan_d <= lizzieLet0_4MQNode_4QNone_Bool_3QVal_Bool_1QError_Bool_d;
  QTree_Bool_t lizzieLet0_4MQNode_4QNone_Bool_3QVal_Bool_1QError_Bool_bufchan_buf;
  assign lizzieLet0_4MQNode_4QNone_Bool_3QVal_Bool_1QError_Bool_bufchan_r = (! lizzieLet0_4MQNode_4QNone_Bool_3QVal_Bool_1QError_Bool_bufchan_buf[0]);
  assign lizzieLet5_1_argbuf_d = (lizzieLet0_4MQNode_4QNone_Bool_3QVal_Bool_1QError_Bool_bufchan_buf[0] ? lizzieLet0_4MQNode_4QNone_Bool_3QVal_Bool_1QError_Bool_bufchan_buf :
                                  lizzieLet0_4MQNode_4QNone_Bool_3QVal_Bool_1QError_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QNone_Bool_3QVal_Bool_1QError_Bool_bufchan_buf <= {66'd0,
                                                                             1'd0};
    else
      if ((lizzieLet5_1_argbuf_r && lizzieLet0_4MQNode_4QNone_Bool_3QVal_Bool_1QError_Bool_bufchan_buf[0]))
        lizzieLet0_4MQNode_4QNone_Bool_3QVal_Bool_1QError_Bool_bufchan_buf <= {66'd0,
                                                                               1'd0};
      else if (((! lizzieLet5_1_argbuf_r) && (! lizzieLet0_4MQNode_4QNone_Bool_3QVal_Bool_1QError_Bool_bufchan_buf[0])))
        lizzieLet0_4MQNode_4QNone_Bool_3QVal_Bool_1QError_Bool_bufchan_buf <= lizzieLet0_4MQNode_4QNone_Bool_3QVal_Bool_1QError_Bool_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet0_4MQNode_4QNone_Bool_3QVal_Bool_2,Go) > (lizzieLet0_4MQNode_4QNone_Bool_3QVal_Bool_2_argbuf,Go) */
  Go_t lizzieLet0_4MQNode_4QNone_Bool_3QVal_Bool_2_bufchan_d;
  logic lizzieLet0_4MQNode_4QNone_Bool_3QVal_Bool_2_bufchan_r;
  assign lizzieLet0_4MQNode_4QNone_Bool_3QVal_Bool_2_r = ((! lizzieLet0_4MQNode_4QNone_Bool_3QVal_Bool_2_bufchan_d[0]) || lizzieLet0_4MQNode_4QNone_Bool_3QVal_Bool_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QNone_Bool_3QVal_Bool_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet0_4MQNode_4QNone_Bool_3QVal_Bool_2_r)
        lizzieLet0_4MQNode_4QNone_Bool_3QVal_Bool_2_bufchan_d <= lizzieLet0_4MQNode_4QNone_Bool_3QVal_Bool_2_d;
  Go_t lizzieLet0_4MQNode_4QNone_Bool_3QVal_Bool_2_bufchan_buf;
  assign lizzieLet0_4MQNode_4QNone_Bool_3QVal_Bool_2_bufchan_r = (! lizzieLet0_4MQNode_4QNone_Bool_3QVal_Bool_2_bufchan_buf[0]);
  assign lizzieLet0_4MQNode_4QNone_Bool_3QVal_Bool_2_argbuf_d = (lizzieLet0_4MQNode_4QNone_Bool_3QVal_Bool_2_bufchan_buf[0] ? lizzieLet0_4MQNode_4QNone_Bool_3QVal_Bool_2_bufchan_buf :
                                                                 lizzieLet0_4MQNode_4QNone_Bool_3QVal_Bool_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QNone_Bool_3QVal_Bool_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet0_4MQNode_4QNone_Bool_3QVal_Bool_2_argbuf_r && lizzieLet0_4MQNode_4QNone_Bool_3QVal_Bool_2_bufchan_buf[0]))
        lizzieLet0_4MQNode_4QNone_Bool_3QVal_Bool_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet0_4MQNode_4QNone_Bool_3QVal_Bool_2_argbuf_r) && (! lizzieLet0_4MQNode_4QNone_Bool_3QVal_Bool_2_bufchan_buf[0])))
        lizzieLet0_4MQNode_4QNone_Bool_3QVal_Bool_2_bufchan_buf <= lizzieLet0_4MQNode_4QNone_Bool_3QVal_Bool_2_bufchan_d;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_CTf) : (lizzieLet0_4MQNode_4QNone_Bool_4,QTree_Bool) (lizzieLet0_4MQNode_5QNone_Bool,Pointer_CTf) > [(lizzieLet0_4MQNode_4QNone_Bool_4QNone_Bool,Pointer_CTf),
                                                                                                                       (lizzieLet0_4MQNode_4QNone_Bool_4QVal_Bool,Pointer_CTf),
                                                                                                                       (lizzieLet0_4MQNode_4QNone_Bool_4QNode_Bool,Pointer_CTf),
                                                                                                                       (lizzieLet0_4MQNode_4QNone_Bool_4QError_Bool,Pointer_CTf)] */
  logic [3:0] lizzieLet0_4MQNode_5QNone_Bool_onehotd;
  always_comb
    if ((lizzieLet0_4MQNode_4QNone_Bool_4_d[0] && lizzieLet0_4MQNode_5QNone_Bool_d[0]))
      unique case (lizzieLet0_4MQNode_4QNone_Bool_4_d[2:1])
        2'd0: lizzieLet0_4MQNode_5QNone_Bool_onehotd = 4'd1;
        2'd1: lizzieLet0_4MQNode_5QNone_Bool_onehotd = 4'd2;
        2'd2: lizzieLet0_4MQNode_5QNone_Bool_onehotd = 4'd4;
        2'd3: lizzieLet0_4MQNode_5QNone_Bool_onehotd = 4'd8;
        default: lizzieLet0_4MQNode_5QNone_Bool_onehotd = 4'd0;
      endcase
    else lizzieLet0_4MQNode_5QNone_Bool_onehotd = 4'd0;
  assign lizzieLet0_4MQNode_4QNone_Bool_4QNone_Bool_d = {lizzieLet0_4MQNode_5QNone_Bool_d[16:1],
                                                         lizzieLet0_4MQNode_5QNone_Bool_onehotd[0]};
  assign lizzieLet0_4MQNode_4QNone_Bool_4QVal_Bool_d = {lizzieLet0_4MQNode_5QNone_Bool_d[16:1],
                                                        lizzieLet0_4MQNode_5QNone_Bool_onehotd[1]};
  assign lizzieLet0_4MQNode_4QNone_Bool_4QNode_Bool_d = {lizzieLet0_4MQNode_5QNone_Bool_d[16:1],
                                                         lizzieLet0_4MQNode_5QNone_Bool_onehotd[2]};
  assign lizzieLet0_4MQNode_4QNone_Bool_4QError_Bool_d = {lizzieLet0_4MQNode_5QNone_Bool_d[16:1],
                                                          lizzieLet0_4MQNode_5QNone_Bool_onehotd[3]};
  assign lizzieLet0_4MQNode_5QNone_Bool_r = (| (lizzieLet0_4MQNode_5QNone_Bool_onehotd & {lizzieLet0_4MQNode_4QNone_Bool_4QError_Bool_r,
                                                                                          lizzieLet0_4MQNode_4QNone_Bool_4QNode_Bool_r,
                                                                                          lizzieLet0_4MQNode_4QNone_Bool_4QVal_Bool_r,
                                                                                          lizzieLet0_4MQNode_4QNone_Bool_4QNone_Bool_r}));
  assign lizzieLet0_4MQNode_4QNone_Bool_4_r = lizzieLet0_4MQNode_5QNone_Bool_r;
  
  /* buf (Ty Pointer_CTf) : (lizzieLet0_4MQNode_4QNone_Bool_4QError_Bool,Pointer_CTf) > (lizzieLet0_4MQNode_4QNone_Bool_4QError_Bool_1_argbuf,Pointer_CTf) */
  Pointer_CTf_t lizzieLet0_4MQNode_4QNone_Bool_4QError_Bool_bufchan_d;
  logic lizzieLet0_4MQNode_4QNone_Bool_4QError_Bool_bufchan_r;
  assign lizzieLet0_4MQNode_4QNone_Bool_4QError_Bool_r = ((! lizzieLet0_4MQNode_4QNone_Bool_4QError_Bool_bufchan_d[0]) || lizzieLet0_4MQNode_4QNone_Bool_4QError_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QNone_Bool_4QError_Bool_bufchan_d <= {16'd0,
                                                                1'd0};
    else
      if (lizzieLet0_4MQNode_4QNone_Bool_4QError_Bool_r)
        lizzieLet0_4MQNode_4QNone_Bool_4QError_Bool_bufchan_d <= lizzieLet0_4MQNode_4QNone_Bool_4QError_Bool_d;
  Pointer_CTf_t lizzieLet0_4MQNode_4QNone_Bool_4QError_Bool_bufchan_buf;
  assign lizzieLet0_4MQNode_4QNone_Bool_4QError_Bool_bufchan_r = (! lizzieLet0_4MQNode_4QNone_Bool_4QError_Bool_bufchan_buf[0]);
  assign lizzieLet0_4MQNode_4QNone_Bool_4QError_Bool_1_argbuf_d = (lizzieLet0_4MQNode_4QNone_Bool_4QError_Bool_bufchan_buf[0] ? lizzieLet0_4MQNode_4QNone_Bool_4QError_Bool_bufchan_buf :
                                                                   lizzieLet0_4MQNode_4QNone_Bool_4QError_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QNone_Bool_4QError_Bool_bufchan_buf <= {16'd0,
                                                                  1'd0};
    else
      if ((lizzieLet0_4MQNode_4QNone_Bool_4QError_Bool_1_argbuf_r && lizzieLet0_4MQNode_4QNone_Bool_4QError_Bool_bufchan_buf[0]))
        lizzieLet0_4MQNode_4QNone_Bool_4QError_Bool_bufchan_buf <= {16'd0,
                                                                    1'd0};
      else if (((! lizzieLet0_4MQNode_4QNone_Bool_4QError_Bool_1_argbuf_r) && (! lizzieLet0_4MQNode_4QNone_Bool_4QError_Bool_bufchan_buf[0])))
        lizzieLet0_4MQNode_4QNone_Bool_4QError_Bool_bufchan_buf <= lizzieLet0_4MQNode_4QNone_Bool_4QError_Bool_bufchan_d;
  
  /* buf (Ty Pointer_CTf) : (lizzieLet0_4MQNode_4QNone_Bool_4QNode_Bool,Pointer_CTf) > (lizzieLet0_4MQNode_4QNone_Bool_4QNode_Bool_1_argbuf,Pointer_CTf) */
  Pointer_CTf_t lizzieLet0_4MQNode_4QNone_Bool_4QNode_Bool_bufchan_d;
  logic lizzieLet0_4MQNode_4QNone_Bool_4QNode_Bool_bufchan_r;
  assign lizzieLet0_4MQNode_4QNone_Bool_4QNode_Bool_r = ((! lizzieLet0_4MQNode_4QNone_Bool_4QNode_Bool_bufchan_d[0]) || lizzieLet0_4MQNode_4QNone_Bool_4QNode_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QNone_Bool_4QNode_Bool_bufchan_d <= {16'd0,
                                                               1'd0};
    else
      if (lizzieLet0_4MQNode_4QNone_Bool_4QNode_Bool_r)
        lizzieLet0_4MQNode_4QNone_Bool_4QNode_Bool_bufchan_d <= lizzieLet0_4MQNode_4QNone_Bool_4QNode_Bool_d;
  Pointer_CTf_t lizzieLet0_4MQNode_4QNone_Bool_4QNode_Bool_bufchan_buf;
  assign lizzieLet0_4MQNode_4QNone_Bool_4QNode_Bool_bufchan_r = (! lizzieLet0_4MQNode_4QNone_Bool_4QNode_Bool_bufchan_buf[0]);
  assign lizzieLet0_4MQNode_4QNone_Bool_4QNode_Bool_1_argbuf_d = (lizzieLet0_4MQNode_4QNone_Bool_4QNode_Bool_bufchan_buf[0] ? lizzieLet0_4MQNode_4QNone_Bool_4QNode_Bool_bufchan_buf :
                                                                  lizzieLet0_4MQNode_4QNone_Bool_4QNode_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QNone_Bool_4QNode_Bool_bufchan_buf <= {16'd0,
                                                                 1'd0};
    else
      if ((lizzieLet0_4MQNode_4QNone_Bool_4QNode_Bool_1_argbuf_r && lizzieLet0_4MQNode_4QNone_Bool_4QNode_Bool_bufchan_buf[0]))
        lizzieLet0_4MQNode_4QNone_Bool_4QNode_Bool_bufchan_buf <= {16'd0,
                                                                   1'd0};
      else if (((! lizzieLet0_4MQNode_4QNone_Bool_4QNode_Bool_1_argbuf_r) && (! lizzieLet0_4MQNode_4QNone_Bool_4QNode_Bool_bufchan_buf[0])))
        lizzieLet0_4MQNode_4QNone_Bool_4QNode_Bool_bufchan_buf <= lizzieLet0_4MQNode_4QNone_Bool_4QNode_Bool_bufchan_d;
  
  /* buf (Ty Pointer_CTf) : (lizzieLet0_4MQNode_4QNone_Bool_4QNone_Bool,Pointer_CTf) > (lizzieLet0_4MQNode_4QNone_Bool_4QNone_Bool_1_argbuf,Pointer_CTf) */
  Pointer_CTf_t lizzieLet0_4MQNode_4QNone_Bool_4QNone_Bool_bufchan_d;
  logic lizzieLet0_4MQNode_4QNone_Bool_4QNone_Bool_bufchan_r;
  assign lizzieLet0_4MQNode_4QNone_Bool_4QNone_Bool_r = ((! lizzieLet0_4MQNode_4QNone_Bool_4QNone_Bool_bufchan_d[0]) || lizzieLet0_4MQNode_4QNone_Bool_4QNone_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QNone_Bool_4QNone_Bool_bufchan_d <= {16'd0,
                                                               1'd0};
    else
      if (lizzieLet0_4MQNode_4QNone_Bool_4QNone_Bool_r)
        lizzieLet0_4MQNode_4QNone_Bool_4QNone_Bool_bufchan_d <= lizzieLet0_4MQNode_4QNone_Bool_4QNone_Bool_d;
  Pointer_CTf_t lizzieLet0_4MQNode_4QNone_Bool_4QNone_Bool_bufchan_buf;
  assign lizzieLet0_4MQNode_4QNone_Bool_4QNone_Bool_bufchan_r = (! lizzieLet0_4MQNode_4QNone_Bool_4QNone_Bool_bufchan_buf[0]);
  assign lizzieLet0_4MQNode_4QNone_Bool_4QNone_Bool_1_argbuf_d = (lizzieLet0_4MQNode_4QNone_Bool_4QNone_Bool_bufchan_buf[0] ? lizzieLet0_4MQNode_4QNone_Bool_4QNone_Bool_bufchan_buf :
                                                                  lizzieLet0_4MQNode_4QNone_Bool_4QNone_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QNone_Bool_4QNone_Bool_bufchan_buf <= {16'd0,
                                                                 1'd0};
    else
      if ((lizzieLet0_4MQNode_4QNone_Bool_4QNone_Bool_1_argbuf_r && lizzieLet0_4MQNode_4QNone_Bool_4QNone_Bool_bufchan_buf[0]))
        lizzieLet0_4MQNode_4QNone_Bool_4QNone_Bool_bufchan_buf <= {16'd0,
                                                                   1'd0};
      else if (((! lizzieLet0_4MQNode_4QNone_Bool_4QNone_Bool_1_argbuf_r) && (! lizzieLet0_4MQNode_4QNone_Bool_4QNone_Bool_bufchan_buf[0])))
        lizzieLet0_4MQNode_4QNone_Bool_4QNone_Bool_bufchan_buf <= lizzieLet0_4MQNode_4QNone_Bool_4QNone_Bool_bufchan_d;
  
  /* buf (Ty Pointer_CTf) : (lizzieLet0_4MQNode_4QNone_Bool_4QVal_Bool,Pointer_CTf) > (lizzieLet0_4MQNode_4QNone_Bool_4QVal_Bool_1_argbuf,Pointer_CTf) */
  Pointer_CTf_t lizzieLet0_4MQNode_4QNone_Bool_4QVal_Bool_bufchan_d;
  logic lizzieLet0_4MQNode_4QNone_Bool_4QVal_Bool_bufchan_r;
  assign lizzieLet0_4MQNode_4QNone_Bool_4QVal_Bool_r = ((! lizzieLet0_4MQNode_4QNone_Bool_4QVal_Bool_bufchan_d[0]) || lizzieLet0_4MQNode_4QNone_Bool_4QVal_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QNone_Bool_4QVal_Bool_bufchan_d <= {16'd0,
                                                              1'd0};
    else
      if (lizzieLet0_4MQNode_4QNone_Bool_4QVal_Bool_r)
        lizzieLet0_4MQNode_4QNone_Bool_4QVal_Bool_bufchan_d <= lizzieLet0_4MQNode_4QNone_Bool_4QVal_Bool_d;
  Pointer_CTf_t lizzieLet0_4MQNode_4QNone_Bool_4QVal_Bool_bufchan_buf;
  assign lizzieLet0_4MQNode_4QNone_Bool_4QVal_Bool_bufchan_r = (! lizzieLet0_4MQNode_4QNone_Bool_4QVal_Bool_bufchan_buf[0]);
  assign lizzieLet0_4MQNode_4QNone_Bool_4QVal_Bool_1_argbuf_d = (lizzieLet0_4MQNode_4QNone_Bool_4QVal_Bool_bufchan_buf[0] ? lizzieLet0_4MQNode_4QNone_Bool_4QVal_Bool_bufchan_buf :
                                                                 lizzieLet0_4MQNode_4QNone_Bool_4QVal_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QNone_Bool_4QVal_Bool_bufchan_buf <= {16'd0,
                                                                1'd0};
    else
      if ((lizzieLet0_4MQNode_4QNone_Bool_4QVal_Bool_1_argbuf_r && lizzieLet0_4MQNode_4QNone_Bool_4QVal_Bool_bufchan_buf[0]))
        lizzieLet0_4MQNode_4QNone_Bool_4QVal_Bool_bufchan_buf <= {16'd0,
                                                                  1'd0};
      else if (((! lizzieLet0_4MQNode_4QNone_Bool_4QVal_Bool_1_argbuf_r) && (! lizzieLet0_4MQNode_4QNone_Bool_4QVal_Bool_bufchan_buf[0])))
        lizzieLet0_4MQNode_4QNone_Bool_4QVal_Bool_bufchan_buf <= lizzieLet0_4MQNode_4QNone_Bool_4QVal_Bool_bufchan_d;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_MaskQTree) : (lizzieLet0_4MQNode_4QNone_Bool_5,QTree_Bool) (lizzieLet0_4MQNode_6QNone_Bool,Pointer_MaskQTree) > [(_96,Pointer_MaskQTree),
                                                                                                                                   (_95,Pointer_MaskQTree),
                                                                                                                                   (lizzieLet0_4MQNode_4QNone_Bool_5QNode_Bool,Pointer_MaskQTree),
                                                                                                                                   (_94,Pointer_MaskQTree)] */
  logic [3:0] lizzieLet0_4MQNode_6QNone_Bool_onehotd;
  always_comb
    if ((lizzieLet0_4MQNode_4QNone_Bool_5_d[0] && lizzieLet0_4MQNode_6QNone_Bool_d[0]))
      unique case (lizzieLet0_4MQNode_4QNone_Bool_5_d[2:1])
        2'd0: lizzieLet0_4MQNode_6QNone_Bool_onehotd = 4'd1;
        2'd1: lizzieLet0_4MQNode_6QNone_Bool_onehotd = 4'd2;
        2'd2: lizzieLet0_4MQNode_6QNone_Bool_onehotd = 4'd4;
        2'd3: lizzieLet0_4MQNode_6QNone_Bool_onehotd = 4'd8;
        default: lizzieLet0_4MQNode_6QNone_Bool_onehotd = 4'd0;
      endcase
    else lizzieLet0_4MQNode_6QNone_Bool_onehotd = 4'd0;
  assign _96_d = {lizzieLet0_4MQNode_6QNone_Bool_d[16:1],
                  lizzieLet0_4MQNode_6QNone_Bool_onehotd[0]};
  assign _95_d = {lizzieLet0_4MQNode_6QNone_Bool_d[16:1],
                  lizzieLet0_4MQNode_6QNone_Bool_onehotd[1]};
  assign lizzieLet0_4MQNode_4QNone_Bool_5QNode_Bool_d = {lizzieLet0_4MQNode_6QNone_Bool_d[16:1],
                                                         lizzieLet0_4MQNode_6QNone_Bool_onehotd[2]};
  assign _94_d = {lizzieLet0_4MQNode_6QNone_Bool_d[16:1],
                  lizzieLet0_4MQNode_6QNone_Bool_onehotd[3]};
  assign lizzieLet0_4MQNode_6QNone_Bool_r = (| (lizzieLet0_4MQNode_6QNone_Bool_onehotd & {_94_r,
                                                                                          lizzieLet0_4MQNode_4QNone_Bool_5QNode_Bool_r,
                                                                                          _95_r,
                                                                                          _96_r}));
  assign lizzieLet0_4MQNode_4QNone_Bool_5_r = lizzieLet0_4MQNode_6QNone_Bool_r;
  
  /* buf (Ty Pointer_MaskQTree) : (lizzieLet0_4MQNode_4QNone_Bool_5QNode_Bool,Pointer_MaskQTree) > (lizzieLet0_4MQNode_4QNone_Bool_5QNode_Bool_1_argbuf,Pointer_MaskQTree) */
  Pointer_MaskQTree_t lizzieLet0_4MQNode_4QNone_Bool_5QNode_Bool_bufchan_d;
  logic lizzieLet0_4MQNode_4QNone_Bool_5QNode_Bool_bufchan_r;
  assign lizzieLet0_4MQNode_4QNone_Bool_5QNode_Bool_r = ((! lizzieLet0_4MQNode_4QNone_Bool_5QNode_Bool_bufchan_d[0]) || lizzieLet0_4MQNode_4QNone_Bool_5QNode_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QNone_Bool_5QNode_Bool_bufchan_d <= {16'd0,
                                                               1'd0};
    else
      if (lizzieLet0_4MQNode_4QNone_Bool_5QNode_Bool_r)
        lizzieLet0_4MQNode_4QNone_Bool_5QNode_Bool_bufchan_d <= lizzieLet0_4MQNode_4QNone_Bool_5QNode_Bool_d;
  Pointer_MaskQTree_t lizzieLet0_4MQNode_4QNone_Bool_5QNode_Bool_bufchan_buf;
  assign lizzieLet0_4MQNode_4QNone_Bool_5QNode_Bool_bufchan_r = (! lizzieLet0_4MQNode_4QNone_Bool_5QNode_Bool_bufchan_buf[0]);
  assign lizzieLet0_4MQNode_4QNone_Bool_5QNode_Bool_1_argbuf_d = (lizzieLet0_4MQNode_4QNone_Bool_5QNode_Bool_bufchan_buf[0] ? lizzieLet0_4MQNode_4QNone_Bool_5QNode_Bool_bufchan_buf :
                                                                  lizzieLet0_4MQNode_4QNone_Bool_5QNode_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QNone_Bool_5QNode_Bool_bufchan_buf <= {16'd0,
                                                                 1'd0};
    else
      if ((lizzieLet0_4MQNode_4QNone_Bool_5QNode_Bool_1_argbuf_r && lizzieLet0_4MQNode_4QNone_Bool_5QNode_Bool_bufchan_buf[0]))
        lizzieLet0_4MQNode_4QNone_Bool_5QNode_Bool_bufchan_buf <= {16'd0,
                                                                   1'd0};
      else if (((! lizzieLet0_4MQNode_4QNone_Bool_5QNode_Bool_1_argbuf_r) && (! lizzieLet0_4MQNode_4QNone_Bool_5QNode_Bool_bufchan_buf[0])))
        lizzieLet0_4MQNode_4QNone_Bool_5QNode_Bool_bufchan_buf <= lizzieLet0_4MQNode_4QNone_Bool_5QNode_Bool_bufchan_d;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_MaskQTree) : (lizzieLet0_4MQNode_4QNone_Bool_6,QTree_Bool) (lizzieLet0_4MQNode_7QNone_Bool,Pointer_MaskQTree) > [(_93,Pointer_MaskQTree),
                                                                                                                                   (_92,Pointer_MaskQTree),
                                                                                                                                   (lizzieLet0_4MQNode_4QNone_Bool_6QNode_Bool,Pointer_MaskQTree),
                                                                                                                                   (_91,Pointer_MaskQTree)] */
  logic [3:0] lizzieLet0_4MQNode_7QNone_Bool_onehotd;
  always_comb
    if ((lizzieLet0_4MQNode_4QNone_Bool_6_d[0] && lizzieLet0_4MQNode_7QNone_Bool_d[0]))
      unique case (lizzieLet0_4MQNode_4QNone_Bool_6_d[2:1])
        2'd0: lizzieLet0_4MQNode_7QNone_Bool_onehotd = 4'd1;
        2'd1: lizzieLet0_4MQNode_7QNone_Bool_onehotd = 4'd2;
        2'd2: lizzieLet0_4MQNode_7QNone_Bool_onehotd = 4'd4;
        2'd3: lizzieLet0_4MQNode_7QNone_Bool_onehotd = 4'd8;
        default: lizzieLet0_4MQNode_7QNone_Bool_onehotd = 4'd0;
      endcase
    else lizzieLet0_4MQNode_7QNone_Bool_onehotd = 4'd0;
  assign _93_d = {lizzieLet0_4MQNode_7QNone_Bool_d[16:1],
                  lizzieLet0_4MQNode_7QNone_Bool_onehotd[0]};
  assign _92_d = {lizzieLet0_4MQNode_7QNone_Bool_d[16:1],
                  lizzieLet0_4MQNode_7QNone_Bool_onehotd[1]};
  assign lizzieLet0_4MQNode_4QNone_Bool_6QNode_Bool_d = {lizzieLet0_4MQNode_7QNone_Bool_d[16:1],
                                                         lizzieLet0_4MQNode_7QNone_Bool_onehotd[2]};
  assign _91_d = {lizzieLet0_4MQNode_7QNone_Bool_d[16:1],
                  lizzieLet0_4MQNode_7QNone_Bool_onehotd[3]};
  assign lizzieLet0_4MQNode_7QNone_Bool_r = (| (lizzieLet0_4MQNode_7QNone_Bool_onehotd & {_91_r,
                                                                                          lizzieLet0_4MQNode_4QNone_Bool_6QNode_Bool_r,
                                                                                          _92_r,
                                                                                          _93_r}));
  assign lizzieLet0_4MQNode_4QNone_Bool_6_r = lizzieLet0_4MQNode_7QNone_Bool_r;
  
  /* buf (Ty Pointer_MaskQTree) : (lizzieLet0_4MQNode_4QNone_Bool_6QNode_Bool,Pointer_MaskQTree) > (lizzieLet0_4MQNode_4QNone_Bool_6QNode_Bool_1_argbuf,Pointer_MaskQTree) */
  Pointer_MaskQTree_t lizzieLet0_4MQNode_4QNone_Bool_6QNode_Bool_bufchan_d;
  logic lizzieLet0_4MQNode_4QNone_Bool_6QNode_Bool_bufchan_r;
  assign lizzieLet0_4MQNode_4QNone_Bool_6QNode_Bool_r = ((! lizzieLet0_4MQNode_4QNone_Bool_6QNode_Bool_bufchan_d[0]) || lizzieLet0_4MQNode_4QNone_Bool_6QNode_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QNone_Bool_6QNode_Bool_bufchan_d <= {16'd0,
                                                               1'd0};
    else
      if (lizzieLet0_4MQNode_4QNone_Bool_6QNode_Bool_r)
        lizzieLet0_4MQNode_4QNone_Bool_6QNode_Bool_bufchan_d <= lizzieLet0_4MQNode_4QNone_Bool_6QNode_Bool_d;
  Pointer_MaskQTree_t lizzieLet0_4MQNode_4QNone_Bool_6QNode_Bool_bufchan_buf;
  assign lizzieLet0_4MQNode_4QNone_Bool_6QNode_Bool_bufchan_r = (! lizzieLet0_4MQNode_4QNone_Bool_6QNode_Bool_bufchan_buf[0]);
  assign lizzieLet0_4MQNode_4QNone_Bool_6QNode_Bool_1_argbuf_d = (lizzieLet0_4MQNode_4QNone_Bool_6QNode_Bool_bufchan_buf[0] ? lizzieLet0_4MQNode_4QNone_Bool_6QNode_Bool_bufchan_buf :
                                                                  lizzieLet0_4MQNode_4QNone_Bool_6QNode_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QNone_Bool_6QNode_Bool_bufchan_buf <= {16'd0,
                                                                 1'd0};
    else
      if ((lizzieLet0_4MQNode_4QNone_Bool_6QNode_Bool_1_argbuf_r && lizzieLet0_4MQNode_4QNone_Bool_6QNode_Bool_bufchan_buf[0]))
        lizzieLet0_4MQNode_4QNone_Bool_6QNode_Bool_bufchan_buf <= {16'd0,
                                                                   1'd0};
      else if (((! lizzieLet0_4MQNode_4QNone_Bool_6QNode_Bool_1_argbuf_r) && (! lizzieLet0_4MQNode_4QNone_Bool_6QNode_Bool_bufchan_buf[0])))
        lizzieLet0_4MQNode_4QNone_Bool_6QNode_Bool_bufchan_buf <= lizzieLet0_4MQNode_4QNone_Bool_6QNode_Bool_bufchan_d;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_MaskQTree) : (lizzieLet0_4MQNode_4QNone_Bool_7,QTree_Bool) (lizzieLet0_4MQNode_8QNone_Bool,Pointer_MaskQTree) > [(_90,Pointer_MaskQTree),
                                                                                                                                   (_89,Pointer_MaskQTree),
                                                                                                                                   (lizzieLet0_4MQNode_4QNone_Bool_7QNode_Bool,Pointer_MaskQTree),
                                                                                                                                   (_88,Pointer_MaskQTree)] */
  logic [3:0] lizzieLet0_4MQNode_8QNone_Bool_onehotd;
  always_comb
    if ((lizzieLet0_4MQNode_4QNone_Bool_7_d[0] && lizzieLet0_4MQNode_8QNone_Bool_d[0]))
      unique case (lizzieLet0_4MQNode_4QNone_Bool_7_d[2:1])
        2'd0: lizzieLet0_4MQNode_8QNone_Bool_onehotd = 4'd1;
        2'd1: lizzieLet0_4MQNode_8QNone_Bool_onehotd = 4'd2;
        2'd2: lizzieLet0_4MQNode_8QNone_Bool_onehotd = 4'd4;
        2'd3: lizzieLet0_4MQNode_8QNone_Bool_onehotd = 4'd8;
        default: lizzieLet0_4MQNode_8QNone_Bool_onehotd = 4'd0;
      endcase
    else lizzieLet0_4MQNode_8QNone_Bool_onehotd = 4'd0;
  assign _90_d = {lizzieLet0_4MQNode_8QNone_Bool_d[16:1],
                  lizzieLet0_4MQNode_8QNone_Bool_onehotd[0]};
  assign _89_d = {lizzieLet0_4MQNode_8QNone_Bool_d[16:1],
                  lizzieLet0_4MQNode_8QNone_Bool_onehotd[1]};
  assign lizzieLet0_4MQNode_4QNone_Bool_7QNode_Bool_d = {lizzieLet0_4MQNode_8QNone_Bool_d[16:1],
                                                         lizzieLet0_4MQNode_8QNone_Bool_onehotd[2]};
  assign _88_d = {lizzieLet0_4MQNode_8QNone_Bool_d[16:1],
                  lizzieLet0_4MQNode_8QNone_Bool_onehotd[3]};
  assign lizzieLet0_4MQNode_8QNone_Bool_r = (| (lizzieLet0_4MQNode_8QNone_Bool_onehotd & {_88_r,
                                                                                          lizzieLet0_4MQNode_4QNone_Bool_7QNode_Bool_r,
                                                                                          _89_r,
                                                                                          _90_r}));
  assign lizzieLet0_4MQNode_4QNone_Bool_7_r = lizzieLet0_4MQNode_8QNone_Bool_r;
  
  /* buf (Ty Pointer_MaskQTree) : (lizzieLet0_4MQNode_4QNone_Bool_7QNode_Bool,Pointer_MaskQTree) > (lizzieLet0_4MQNode_4QNone_Bool_7QNode_Bool_1_argbuf,Pointer_MaskQTree) */
  Pointer_MaskQTree_t lizzieLet0_4MQNode_4QNone_Bool_7QNode_Bool_bufchan_d;
  logic lizzieLet0_4MQNode_4QNone_Bool_7QNode_Bool_bufchan_r;
  assign lizzieLet0_4MQNode_4QNone_Bool_7QNode_Bool_r = ((! lizzieLet0_4MQNode_4QNone_Bool_7QNode_Bool_bufchan_d[0]) || lizzieLet0_4MQNode_4QNone_Bool_7QNode_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QNone_Bool_7QNode_Bool_bufchan_d <= {16'd0,
                                                               1'd0};
    else
      if (lizzieLet0_4MQNode_4QNone_Bool_7QNode_Bool_r)
        lizzieLet0_4MQNode_4QNone_Bool_7QNode_Bool_bufchan_d <= lizzieLet0_4MQNode_4QNone_Bool_7QNode_Bool_d;
  Pointer_MaskQTree_t lizzieLet0_4MQNode_4QNone_Bool_7QNode_Bool_bufchan_buf;
  assign lizzieLet0_4MQNode_4QNone_Bool_7QNode_Bool_bufchan_r = (! lizzieLet0_4MQNode_4QNone_Bool_7QNode_Bool_bufchan_buf[0]);
  assign lizzieLet0_4MQNode_4QNone_Bool_7QNode_Bool_1_argbuf_d = (lizzieLet0_4MQNode_4QNone_Bool_7QNode_Bool_bufchan_buf[0] ? lizzieLet0_4MQNode_4QNone_Bool_7QNode_Bool_bufchan_buf :
                                                                  lizzieLet0_4MQNode_4QNone_Bool_7QNode_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QNone_Bool_7QNode_Bool_bufchan_buf <= {16'd0,
                                                                 1'd0};
    else
      if ((lizzieLet0_4MQNode_4QNone_Bool_7QNode_Bool_1_argbuf_r && lizzieLet0_4MQNode_4QNone_Bool_7QNode_Bool_bufchan_buf[0]))
        lizzieLet0_4MQNode_4QNone_Bool_7QNode_Bool_bufchan_buf <= {16'd0,
                                                                   1'd0};
      else if (((! lizzieLet0_4MQNode_4QNone_Bool_7QNode_Bool_1_argbuf_r) && (! lizzieLet0_4MQNode_4QNone_Bool_7QNode_Bool_bufchan_buf[0])))
        lizzieLet0_4MQNode_4QNone_Bool_7QNode_Bool_bufchan_buf <= lizzieLet0_4MQNode_4QNone_Bool_7QNode_Bool_bufchan_d;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_MaskQTree) : (lizzieLet0_4MQNode_4QNone_Bool_8,QTree_Bool) (lizzieLet0_4MQNode_9QNone_Bool,Pointer_MaskQTree) > [(_87,Pointer_MaskQTree),
                                                                                                                                   (_86,Pointer_MaskQTree),
                                                                                                                                   (lizzieLet0_4MQNode_4QNone_Bool_8QNode_Bool,Pointer_MaskQTree),
                                                                                                                                   (_85,Pointer_MaskQTree)] */
  logic [3:0] lizzieLet0_4MQNode_9QNone_Bool_onehotd;
  always_comb
    if ((lizzieLet0_4MQNode_4QNone_Bool_8_d[0] && lizzieLet0_4MQNode_9QNone_Bool_d[0]))
      unique case (lizzieLet0_4MQNode_4QNone_Bool_8_d[2:1])
        2'd0: lizzieLet0_4MQNode_9QNone_Bool_onehotd = 4'd1;
        2'd1: lizzieLet0_4MQNode_9QNone_Bool_onehotd = 4'd2;
        2'd2: lizzieLet0_4MQNode_9QNone_Bool_onehotd = 4'd4;
        2'd3: lizzieLet0_4MQNode_9QNone_Bool_onehotd = 4'd8;
        default: lizzieLet0_4MQNode_9QNone_Bool_onehotd = 4'd0;
      endcase
    else lizzieLet0_4MQNode_9QNone_Bool_onehotd = 4'd0;
  assign _87_d = {lizzieLet0_4MQNode_9QNone_Bool_d[16:1],
                  lizzieLet0_4MQNode_9QNone_Bool_onehotd[0]};
  assign _86_d = {lizzieLet0_4MQNode_9QNone_Bool_d[16:1],
                  lizzieLet0_4MQNode_9QNone_Bool_onehotd[1]};
  assign lizzieLet0_4MQNode_4QNone_Bool_8QNode_Bool_d = {lizzieLet0_4MQNode_9QNone_Bool_d[16:1],
                                                         lizzieLet0_4MQNode_9QNone_Bool_onehotd[2]};
  assign _85_d = {lizzieLet0_4MQNode_9QNone_Bool_d[16:1],
                  lizzieLet0_4MQNode_9QNone_Bool_onehotd[3]};
  assign lizzieLet0_4MQNode_9QNone_Bool_r = (| (lizzieLet0_4MQNode_9QNone_Bool_onehotd & {_85_r,
                                                                                          lizzieLet0_4MQNode_4QNone_Bool_8QNode_Bool_r,
                                                                                          _86_r,
                                                                                          _87_r}));
  assign lizzieLet0_4MQNode_4QNone_Bool_8_r = lizzieLet0_4MQNode_9QNone_Bool_r;
  
  /* buf (Ty Pointer_MaskQTree) : (lizzieLet0_4MQNode_4QNone_Bool_8QNode_Bool,Pointer_MaskQTree) > (lizzieLet0_4MQNode_4QNone_Bool_8QNode_Bool_1_argbuf,Pointer_MaskQTree) */
  Pointer_MaskQTree_t lizzieLet0_4MQNode_4QNone_Bool_8QNode_Bool_bufchan_d;
  logic lizzieLet0_4MQNode_4QNone_Bool_8QNode_Bool_bufchan_r;
  assign lizzieLet0_4MQNode_4QNone_Bool_8QNode_Bool_r = ((! lizzieLet0_4MQNode_4QNone_Bool_8QNode_Bool_bufchan_d[0]) || lizzieLet0_4MQNode_4QNone_Bool_8QNode_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QNone_Bool_8QNode_Bool_bufchan_d <= {16'd0,
                                                               1'd0};
    else
      if (lizzieLet0_4MQNode_4QNone_Bool_8QNode_Bool_r)
        lizzieLet0_4MQNode_4QNone_Bool_8QNode_Bool_bufchan_d <= lizzieLet0_4MQNode_4QNone_Bool_8QNode_Bool_d;
  Pointer_MaskQTree_t lizzieLet0_4MQNode_4QNone_Bool_8QNode_Bool_bufchan_buf;
  assign lizzieLet0_4MQNode_4QNone_Bool_8QNode_Bool_bufchan_r = (! lizzieLet0_4MQNode_4QNone_Bool_8QNode_Bool_bufchan_buf[0]);
  assign lizzieLet0_4MQNode_4QNone_Bool_8QNode_Bool_1_argbuf_d = (lizzieLet0_4MQNode_4QNone_Bool_8QNode_Bool_bufchan_buf[0] ? lizzieLet0_4MQNode_4QNone_Bool_8QNode_Bool_bufchan_buf :
                                                                  lizzieLet0_4MQNode_4QNone_Bool_8QNode_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QNone_Bool_8QNode_Bool_bufchan_buf <= {16'd0,
                                                                 1'd0};
    else
      if ((lizzieLet0_4MQNode_4QNone_Bool_8QNode_Bool_1_argbuf_r && lizzieLet0_4MQNode_4QNone_Bool_8QNode_Bool_bufchan_buf[0]))
        lizzieLet0_4MQNode_4QNone_Bool_8QNode_Bool_bufchan_buf <= {16'd0,
                                                                   1'd0};
      else if (((! lizzieLet0_4MQNode_4QNone_Bool_8QNode_Bool_1_argbuf_r) && (! lizzieLet0_4MQNode_4QNone_Bool_8QNode_Bool_bufchan_buf[0])))
        lizzieLet0_4MQNode_4QNone_Bool_8QNode_Bool_bufchan_buf <= lizzieLet0_4MQNode_4QNone_Bool_8QNode_Bool_bufchan_d;
  
  /* fork (Ty QTree_Bool) : (lizzieLet0_4MQNode_4QVal_Bool,QTree_Bool) > [(lizzieLet0_4MQNode_4QVal_Bool_1,QTree_Bool),
                                                                     (lizzieLet0_4MQNode_4QVal_Bool_2,QTree_Bool),
                                                                     (lizzieLet0_4MQNode_4QVal_Bool_3,QTree_Bool),
                                                                     (lizzieLet0_4MQNode_4QVal_Bool_4,QTree_Bool),
                                                                     (lizzieLet0_4MQNode_4QVal_Bool_5,QTree_Bool)] */
  logic [4:0] lizzieLet0_4MQNode_4QVal_Bool_emitted;
  logic [4:0] lizzieLet0_4MQNode_4QVal_Bool_done;
  assign lizzieLet0_4MQNode_4QVal_Bool_1_d = {lizzieLet0_4MQNode_4QVal_Bool_d[66:1],
                                              (lizzieLet0_4MQNode_4QVal_Bool_d[0] && (! lizzieLet0_4MQNode_4QVal_Bool_emitted[0]))};
  assign lizzieLet0_4MQNode_4QVal_Bool_2_d = {lizzieLet0_4MQNode_4QVal_Bool_d[66:1],
                                              (lizzieLet0_4MQNode_4QVal_Bool_d[0] && (! lizzieLet0_4MQNode_4QVal_Bool_emitted[1]))};
  assign lizzieLet0_4MQNode_4QVal_Bool_3_d = {lizzieLet0_4MQNode_4QVal_Bool_d[66:1],
                                              (lizzieLet0_4MQNode_4QVal_Bool_d[0] && (! lizzieLet0_4MQNode_4QVal_Bool_emitted[2]))};
  assign lizzieLet0_4MQNode_4QVal_Bool_4_d = {lizzieLet0_4MQNode_4QVal_Bool_d[66:1],
                                              (lizzieLet0_4MQNode_4QVal_Bool_d[0] && (! lizzieLet0_4MQNode_4QVal_Bool_emitted[3]))};
  assign lizzieLet0_4MQNode_4QVal_Bool_5_d = {lizzieLet0_4MQNode_4QVal_Bool_d[66:1],
                                              (lizzieLet0_4MQNode_4QVal_Bool_d[0] && (! lizzieLet0_4MQNode_4QVal_Bool_emitted[4]))};
  assign lizzieLet0_4MQNode_4QVal_Bool_done = (lizzieLet0_4MQNode_4QVal_Bool_emitted | ({lizzieLet0_4MQNode_4QVal_Bool_5_d[0],
                                                                                         lizzieLet0_4MQNode_4QVal_Bool_4_d[0],
                                                                                         lizzieLet0_4MQNode_4QVal_Bool_3_d[0],
                                                                                         lizzieLet0_4MQNode_4QVal_Bool_2_d[0],
                                                                                         lizzieLet0_4MQNode_4QVal_Bool_1_d[0]} & {lizzieLet0_4MQNode_4QVal_Bool_5_r,
                                                                                                                                  lizzieLet0_4MQNode_4QVal_Bool_4_r,
                                                                                                                                  lizzieLet0_4MQNode_4QVal_Bool_3_r,
                                                                                                                                  lizzieLet0_4MQNode_4QVal_Bool_2_r,
                                                                                                                                  lizzieLet0_4MQNode_4QVal_Bool_1_r}));
  assign lizzieLet0_4MQNode_4QVal_Bool_r = (& lizzieLet0_4MQNode_4QVal_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet0_4MQNode_4QVal_Bool_emitted <= 5'd0;
    else
      lizzieLet0_4MQNode_4QVal_Bool_emitted <= (lizzieLet0_4MQNode_4QVal_Bool_r ? 5'd0 :
                                                lizzieLet0_4MQNode_4QVal_Bool_done);
  
  /* destruct (Ty QTree_Bool,
          Dcon QVal_Bool) : (lizzieLet0_4MQNode_4QVal_Bool_1QVal_Bool,QTree_Bool) > [(va8i_destruct,MyBool)] */
  assign va8i_destruct_d = {lizzieLet0_4MQNode_4QVal_Bool_1QVal_Bool_d[3:3],
                            lizzieLet0_4MQNode_4QVal_Bool_1QVal_Bool_d[0]};
  assign lizzieLet0_4MQNode_4QVal_Bool_1QVal_Bool_r = va8i_destruct_r;
  
  /* demux (Ty QTree_Bool,
       Ty QTree_Bool) : (lizzieLet0_4MQNode_4QVal_Bool_2,QTree_Bool) (lizzieLet0_4MQNode_4QVal_Bool_1,QTree_Bool) > [(_84,QTree_Bool),
                                                                                                                     (lizzieLet0_4MQNode_4QVal_Bool_1QVal_Bool,QTree_Bool),
                                                                                                                     (_83,QTree_Bool),
                                                                                                                     (_82,QTree_Bool)] */
  logic [3:0] lizzieLet0_4MQNode_4QVal_Bool_1_onehotd;
  always_comb
    if ((lizzieLet0_4MQNode_4QVal_Bool_2_d[0] && lizzieLet0_4MQNode_4QVal_Bool_1_d[0]))
      unique case (lizzieLet0_4MQNode_4QVal_Bool_2_d[2:1])
        2'd0: lizzieLet0_4MQNode_4QVal_Bool_1_onehotd = 4'd1;
        2'd1: lizzieLet0_4MQNode_4QVal_Bool_1_onehotd = 4'd2;
        2'd2: lizzieLet0_4MQNode_4QVal_Bool_1_onehotd = 4'd4;
        2'd3: lizzieLet0_4MQNode_4QVal_Bool_1_onehotd = 4'd8;
        default: lizzieLet0_4MQNode_4QVal_Bool_1_onehotd = 4'd0;
      endcase
    else lizzieLet0_4MQNode_4QVal_Bool_1_onehotd = 4'd0;
  assign _84_d = {lizzieLet0_4MQNode_4QVal_Bool_1_d[66:1],
                  lizzieLet0_4MQNode_4QVal_Bool_1_onehotd[0]};
  assign lizzieLet0_4MQNode_4QVal_Bool_1QVal_Bool_d = {lizzieLet0_4MQNode_4QVal_Bool_1_d[66:1],
                                                       lizzieLet0_4MQNode_4QVal_Bool_1_onehotd[1]};
  assign _83_d = {lizzieLet0_4MQNode_4QVal_Bool_1_d[66:1],
                  lizzieLet0_4MQNode_4QVal_Bool_1_onehotd[2]};
  assign _82_d = {lizzieLet0_4MQNode_4QVal_Bool_1_d[66:1],
                  lizzieLet0_4MQNode_4QVal_Bool_1_onehotd[3]};
  assign lizzieLet0_4MQNode_4QVal_Bool_1_r = (| (lizzieLet0_4MQNode_4QVal_Bool_1_onehotd & {_82_r,
                                                                                            _83_r,
                                                                                            lizzieLet0_4MQNode_4QVal_Bool_1QVal_Bool_r,
                                                                                            _84_r}));
  assign lizzieLet0_4MQNode_4QVal_Bool_2_r = lizzieLet0_4MQNode_4QVal_Bool_1_r;
  
  /* demux (Ty QTree_Bool,
       Ty Go) : (lizzieLet0_4MQNode_4QVal_Bool_3,QTree_Bool) (lizzieLet0_4MQNode_3QVal_Bool,Go) > [(lizzieLet0_4MQNode_4QVal_Bool_3QNone_Bool,Go),
                                                                                                   (lizzieLet0_4MQNode_4QVal_Bool_3QVal_Bool,Go),
                                                                                                   (lizzieLet0_4MQNode_4QVal_Bool_3QNode_Bool,Go),
                                                                                                   (lizzieLet0_4MQNode_4QVal_Bool_3QError_Bool,Go)] */
  logic [3:0] lizzieLet0_4MQNode_3QVal_Bool_onehotd;
  always_comb
    if ((lizzieLet0_4MQNode_4QVal_Bool_3_d[0] && lizzieLet0_4MQNode_3QVal_Bool_d[0]))
      unique case (lizzieLet0_4MQNode_4QVal_Bool_3_d[2:1])
        2'd0: lizzieLet0_4MQNode_3QVal_Bool_onehotd = 4'd1;
        2'd1: lizzieLet0_4MQNode_3QVal_Bool_onehotd = 4'd2;
        2'd2: lizzieLet0_4MQNode_3QVal_Bool_onehotd = 4'd4;
        2'd3: lizzieLet0_4MQNode_3QVal_Bool_onehotd = 4'd8;
        default: lizzieLet0_4MQNode_3QVal_Bool_onehotd = 4'd0;
      endcase
    else lizzieLet0_4MQNode_3QVal_Bool_onehotd = 4'd0;
  assign lizzieLet0_4MQNode_4QVal_Bool_3QNone_Bool_d = lizzieLet0_4MQNode_3QVal_Bool_onehotd[0];
  assign lizzieLet0_4MQNode_4QVal_Bool_3QVal_Bool_d = lizzieLet0_4MQNode_3QVal_Bool_onehotd[1];
  assign lizzieLet0_4MQNode_4QVal_Bool_3QNode_Bool_d = lizzieLet0_4MQNode_3QVal_Bool_onehotd[2];
  assign lizzieLet0_4MQNode_4QVal_Bool_3QError_Bool_d = lizzieLet0_4MQNode_3QVal_Bool_onehotd[3];
  assign lizzieLet0_4MQNode_3QVal_Bool_r = (| (lizzieLet0_4MQNode_3QVal_Bool_onehotd & {lizzieLet0_4MQNode_4QVal_Bool_3QError_Bool_r,
                                                                                        lizzieLet0_4MQNode_4QVal_Bool_3QNode_Bool_r,
                                                                                        lizzieLet0_4MQNode_4QVal_Bool_3QVal_Bool_r,
                                                                                        lizzieLet0_4MQNode_4QVal_Bool_3QNone_Bool_r}));
  assign lizzieLet0_4MQNode_4QVal_Bool_3_r = lizzieLet0_4MQNode_3QVal_Bool_r;
  
  /* fork (Ty Go) : (lizzieLet0_4MQNode_4QVal_Bool_3QError_Bool,Go) > [(lizzieLet0_4MQNode_4QVal_Bool_3QError_Bool_1,Go),
                                                                  (lizzieLet0_4MQNode_4QVal_Bool_3QError_Bool_2,Go)] */
  logic [1:0] lizzieLet0_4MQNode_4QVal_Bool_3QError_Bool_emitted;
  logic [1:0] lizzieLet0_4MQNode_4QVal_Bool_3QError_Bool_done;
  assign lizzieLet0_4MQNode_4QVal_Bool_3QError_Bool_1_d = (lizzieLet0_4MQNode_4QVal_Bool_3QError_Bool_d[0] && (! lizzieLet0_4MQNode_4QVal_Bool_3QError_Bool_emitted[0]));
  assign lizzieLet0_4MQNode_4QVal_Bool_3QError_Bool_2_d = (lizzieLet0_4MQNode_4QVal_Bool_3QError_Bool_d[0] && (! lizzieLet0_4MQNode_4QVal_Bool_3QError_Bool_emitted[1]));
  assign lizzieLet0_4MQNode_4QVal_Bool_3QError_Bool_done = (lizzieLet0_4MQNode_4QVal_Bool_3QError_Bool_emitted | ({lizzieLet0_4MQNode_4QVal_Bool_3QError_Bool_2_d[0],
                                                                                                                   lizzieLet0_4MQNode_4QVal_Bool_3QError_Bool_1_d[0]} & {lizzieLet0_4MQNode_4QVal_Bool_3QError_Bool_2_r,
                                                                                                                                                                         lizzieLet0_4MQNode_4QVal_Bool_3QError_Bool_1_r}));
  assign lizzieLet0_4MQNode_4QVal_Bool_3QError_Bool_r = (& lizzieLet0_4MQNode_4QVal_Bool_3QError_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QVal_Bool_3QError_Bool_emitted <= 2'd0;
    else
      lizzieLet0_4MQNode_4QVal_Bool_3QError_Bool_emitted <= (lizzieLet0_4MQNode_4QVal_Bool_3QError_Bool_r ? 2'd0 :
                                                             lizzieLet0_4MQNode_4QVal_Bool_3QError_Bool_done);
  
  /* dcon (Ty QTree_Bool,
      Dcon QError_Bool) : [(lizzieLet0_4MQNode_4QVal_Bool_3QError_Bool_1,Go)] > (lizzieLet0_4MQNode_4QVal_Bool_3QError_Bool_1QError_Bool,QTree_Bool) */
  assign lizzieLet0_4MQNode_4QVal_Bool_3QError_Bool_1QError_Bool_d = QError_Bool_dc((& {lizzieLet0_4MQNode_4QVal_Bool_3QError_Bool_1_d[0]}), lizzieLet0_4MQNode_4QVal_Bool_3QError_Bool_1_d);
  assign {lizzieLet0_4MQNode_4QVal_Bool_3QError_Bool_1_r} = {1 {(lizzieLet0_4MQNode_4QVal_Bool_3QError_Bool_1QError_Bool_r && lizzieLet0_4MQNode_4QVal_Bool_3QError_Bool_1QError_Bool_d[0])}};
  
  /* buf (Ty QTree_Bool) : (lizzieLet0_4MQNode_4QVal_Bool_3QError_Bool_1QError_Bool,QTree_Bool) > (lizzieLet9_1_1_argbuf,QTree_Bool) */
  QTree_Bool_t lizzieLet0_4MQNode_4QVal_Bool_3QError_Bool_1QError_Bool_bufchan_d;
  logic lizzieLet0_4MQNode_4QVal_Bool_3QError_Bool_1QError_Bool_bufchan_r;
  assign lizzieLet0_4MQNode_4QVal_Bool_3QError_Bool_1QError_Bool_r = ((! lizzieLet0_4MQNode_4QVal_Bool_3QError_Bool_1QError_Bool_bufchan_d[0]) || lizzieLet0_4MQNode_4QVal_Bool_3QError_Bool_1QError_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QVal_Bool_3QError_Bool_1QError_Bool_bufchan_d <= {66'd0,
                                                                            1'd0};
    else
      if (lizzieLet0_4MQNode_4QVal_Bool_3QError_Bool_1QError_Bool_r)
        lizzieLet0_4MQNode_4QVal_Bool_3QError_Bool_1QError_Bool_bufchan_d <= lizzieLet0_4MQNode_4QVal_Bool_3QError_Bool_1QError_Bool_d;
  QTree_Bool_t lizzieLet0_4MQNode_4QVal_Bool_3QError_Bool_1QError_Bool_bufchan_buf;
  assign lizzieLet0_4MQNode_4QVal_Bool_3QError_Bool_1QError_Bool_bufchan_r = (! lizzieLet0_4MQNode_4QVal_Bool_3QError_Bool_1QError_Bool_bufchan_buf[0]);
  assign lizzieLet9_1_1_argbuf_d = (lizzieLet0_4MQNode_4QVal_Bool_3QError_Bool_1QError_Bool_bufchan_buf[0] ? lizzieLet0_4MQNode_4QVal_Bool_3QError_Bool_1QError_Bool_bufchan_buf :
                                    lizzieLet0_4MQNode_4QVal_Bool_3QError_Bool_1QError_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QVal_Bool_3QError_Bool_1QError_Bool_bufchan_buf <= {66'd0,
                                                                              1'd0};
    else
      if ((lizzieLet9_1_1_argbuf_r && lizzieLet0_4MQNode_4QVal_Bool_3QError_Bool_1QError_Bool_bufchan_buf[0]))
        lizzieLet0_4MQNode_4QVal_Bool_3QError_Bool_1QError_Bool_bufchan_buf <= {66'd0,
                                                                                1'd0};
      else if (((! lizzieLet9_1_1_argbuf_r) && (! lizzieLet0_4MQNode_4QVal_Bool_3QError_Bool_1QError_Bool_bufchan_buf[0])))
        lizzieLet0_4MQNode_4QVal_Bool_3QError_Bool_1QError_Bool_bufchan_buf <= lizzieLet0_4MQNode_4QVal_Bool_3QError_Bool_1QError_Bool_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet0_4MQNode_4QVal_Bool_3QError_Bool_2,Go) > (lizzieLet0_4MQNode_4QVal_Bool_3QError_Bool_2_argbuf,Go) */
  Go_t lizzieLet0_4MQNode_4QVal_Bool_3QError_Bool_2_bufchan_d;
  logic lizzieLet0_4MQNode_4QVal_Bool_3QError_Bool_2_bufchan_r;
  assign lizzieLet0_4MQNode_4QVal_Bool_3QError_Bool_2_r = ((! lizzieLet0_4MQNode_4QVal_Bool_3QError_Bool_2_bufchan_d[0]) || lizzieLet0_4MQNode_4QVal_Bool_3QError_Bool_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QVal_Bool_3QError_Bool_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet0_4MQNode_4QVal_Bool_3QError_Bool_2_r)
        lizzieLet0_4MQNode_4QVal_Bool_3QError_Bool_2_bufchan_d <= lizzieLet0_4MQNode_4QVal_Bool_3QError_Bool_2_d;
  Go_t lizzieLet0_4MQNode_4QVal_Bool_3QError_Bool_2_bufchan_buf;
  assign lizzieLet0_4MQNode_4QVal_Bool_3QError_Bool_2_bufchan_r = (! lizzieLet0_4MQNode_4QVal_Bool_3QError_Bool_2_bufchan_buf[0]);
  assign lizzieLet0_4MQNode_4QVal_Bool_3QError_Bool_2_argbuf_d = (lizzieLet0_4MQNode_4QVal_Bool_3QError_Bool_2_bufchan_buf[0] ? lizzieLet0_4MQNode_4QVal_Bool_3QError_Bool_2_bufchan_buf :
                                                                  lizzieLet0_4MQNode_4QVal_Bool_3QError_Bool_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QVal_Bool_3QError_Bool_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet0_4MQNode_4QVal_Bool_3QError_Bool_2_argbuf_r && lizzieLet0_4MQNode_4QVal_Bool_3QError_Bool_2_bufchan_buf[0]))
        lizzieLet0_4MQNode_4QVal_Bool_3QError_Bool_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet0_4MQNode_4QVal_Bool_3QError_Bool_2_argbuf_r) && (! lizzieLet0_4MQNode_4QVal_Bool_3QError_Bool_2_bufchan_buf[0])))
        lizzieLet0_4MQNode_4QVal_Bool_3QError_Bool_2_bufchan_buf <= lizzieLet0_4MQNode_4QVal_Bool_3QError_Bool_2_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet0_4MQNode_4QVal_Bool_3QNode_Bool,Go) > [(lizzieLet0_4MQNode_4QVal_Bool_3QNode_Bool_1,Go),
                                                                 (lizzieLet0_4MQNode_4QVal_Bool_3QNode_Bool_2,Go)] */
  logic [1:0] lizzieLet0_4MQNode_4QVal_Bool_3QNode_Bool_emitted;
  logic [1:0] lizzieLet0_4MQNode_4QVal_Bool_3QNode_Bool_done;
  assign lizzieLet0_4MQNode_4QVal_Bool_3QNode_Bool_1_d = (lizzieLet0_4MQNode_4QVal_Bool_3QNode_Bool_d[0] && (! lizzieLet0_4MQNode_4QVal_Bool_3QNode_Bool_emitted[0]));
  assign lizzieLet0_4MQNode_4QVal_Bool_3QNode_Bool_2_d = (lizzieLet0_4MQNode_4QVal_Bool_3QNode_Bool_d[0] && (! lizzieLet0_4MQNode_4QVal_Bool_3QNode_Bool_emitted[1]));
  assign lizzieLet0_4MQNode_4QVal_Bool_3QNode_Bool_done = (lizzieLet0_4MQNode_4QVal_Bool_3QNode_Bool_emitted | ({lizzieLet0_4MQNode_4QVal_Bool_3QNode_Bool_2_d[0],
                                                                                                                 lizzieLet0_4MQNode_4QVal_Bool_3QNode_Bool_1_d[0]} & {lizzieLet0_4MQNode_4QVal_Bool_3QNode_Bool_2_r,
                                                                                                                                                                      lizzieLet0_4MQNode_4QVal_Bool_3QNode_Bool_1_r}));
  assign lizzieLet0_4MQNode_4QVal_Bool_3QNode_Bool_r = (& lizzieLet0_4MQNode_4QVal_Bool_3QNode_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QVal_Bool_3QNode_Bool_emitted <= 2'd0;
    else
      lizzieLet0_4MQNode_4QVal_Bool_3QNode_Bool_emitted <= (lizzieLet0_4MQNode_4QVal_Bool_3QNode_Bool_r ? 2'd0 :
                                                            lizzieLet0_4MQNode_4QVal_Bool_3QNode_Bool_done);
  
  /* dcon (Ty QTree_Bool,
      Dcon QError_Bool) : [(lizzieLet0_4MQNode_4QVal_Bool_3QNode_Bool_1,Go)] > (lizzieLet0_4MQNode_4QVal_Bool_3QNode_Bool_1QError_Bool,QTree_Bool) */
  assign lizzieLet0_4MQNode_4QVal_Bool_3QNode_Bool_1QError_Bool_d = QError_Bool_dc((& {lizzieLet0_4MQNode_4QVal_Bool_3QNode_Bool_1_d[0]}), lizzieLet0_4MQNode_4QVal_Bool_3QNode_Bool_1_d);
  assign {lizzieLet0_4MQNode_4QVal_Bool_3QNode_Bool_1_r} = {1 {(lizzieLet0_4MQNode_4QVal_Bool_3QNode_Bool_1QError_Bool_r && lizzieLet0_4MQNode_4QVal_Bool_3QNode_Bool_1QError_Bool_d[0])}};
  
  /* buf (Ty QTree_Bool) : (lizzieLet0_4MQNode_4QVal_Bool_3QNode_Bool_1QError_Bool,QTree_Bool) > (lizzieLet13_1_1_argbuf,QTree_Bool) */
  QTree_Bool_t lizzieLet0_4MQNode_4QVal_Bool_3QNode_Bool_1QError_Bool_bufchan_d;
  logic lizzieLet0_4MQNode_4QVal_Bool_3QNode_Bool_1QError_Bool_bufchan_r;
  assign lizzieLet0_4MQNode_4QVal_Bool_3QNode_Bool_1QError_Bool_r = ((! lizzieLet0_4MQNode_4QVal_Bool_3QNode_Bool_1QError_Bool_bufchan_d[0]) || lizzieLet0_4MQNode_4QVal_Bool_3QNode_Bool_1QError_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QVal_Bool_3QNode_Bool_1QError_Bool_bufchan_d <= {66'd0,
                                                                           1'd0};
    else
      if (lizzieLet0_4MQNode_4QVal_Bool_3QNode_Bool_1QError_Bool_r)
        lizzieLet0_4MQNode_4QVal_Bool_3QNode_Bool_1QError_Bool_bufchan_d <= lizzieLet0_4MQNode_4QVal_Bool_3QNode_Bool_1QError_Bool_d;
  QTree_Bool_t lizzieLet0_4MQNode_4QVal_Bool_3QNode_Bool_1QError_Bool_bufchan_buf;
  assign lizzieLet0_4MQNode_4QVal_Bool_3QNode_Bool_1QError_Bool_bufchan_r = (! lizzieLet0_4MQNode_4QVal_Bool_3QNode_Bool_1QError_Bool_bufchan_buf[0]);
  assign lizzieLet13_1_1_argbuf_d = (lizzieLet0_4MQNode_4QVal_Bool_3QNode_Bool_1QError_Bool_bufchan_buf[0] ? lizzieLet0_4MQNode_4QVal_Bool_3QNode_Bool_1QError_Bool_bufchan_buf :
                                     lizzieLet0_4MQNode_4QVal_Bool_3QNode_Bool_1QError_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QVal_Bool_3QNode_Bool_1QError_Bool_bufchan_buf <= {66'd0,
                                                                             1'd0};
    else
      if ((lizzieLet13_1_1_argbuf_r && lizzieLet0_4MQNode_4QVal_Bool_3QNode_Bool_1QError_Bool_bufchan_buf[0]))
        lizzieLet0_4MQNode_4QVal_Bool_3QNode_Bool_1QError_Bool_bufchan_buf <= {66'd0,
                                                                               1'd0};
      else if (((! lizzieLet13_1_1_argbuf_r) && (! lizzieLet0_4MQNode_4QVal_Bool_3QNode_Bool_1QError_Bool_bufchan_buf[0])))
        lizzieLet0_4MQNode_4QVal_Bool_3QNode_Bool_1QError_Bool_bufchan_buf <= lizzieLet0_4MQNode_4QVal_Bool_3QNode_Bool_1QError_Bool_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet0_4MQNode_4QVal_Bool_3QNode_Bool_2,Go) > (lizzieLet0_4MQNode_4QVal_Bool_3QNode_Bool_2_argbuf,Go) */
  Go_t lizzieLet0_4MQNode_4QVal_Bool_3QNode_Bool_2_bufchan_d;
  logic lizzieLet0_4MQNode_4QVal_Bool_3QNode_Bool_2_bufchan_r;
  assign lizzieLet0_4MQNode_4QVal_Bool_3QNode_Bool_2_r = ((! lizzieLet0_4MQNode_4QVal_Bool_3QNode_Bool_2_bufchan_d[0]) || lizzieLet0_4MQNode_4QVal_Bool_3QNode_Bool_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QVal_Bool_3QNode_Bool_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet0_4MQNode_4QVal_Bool_3QNode_Bool_2_r)
        lizzieLet0_4MQNode_4QVal_Bool_3QNode_Bool_2_bufchan_d <= lizzieLet0_4MQNode_4QVal_Bool_3QNode_Bool_2_d;
  Go_t lizzieLet0_4MQNode_4QVal_Bool_3QNode_Bool_2_bufchan_buf;
  assign lizzieLet0_4MQNode_4QVal_Bool_3QNode_Bool_2_bufchan_r = (! lizzieLet0_4MQNode_4QVal_Bool_3QNode_Bool_2_bufchan_buf[0]);
  assign lizzieLet0_4MQNode_4QVal_Bool_3QNode_Bool_2_argbuf_d = (lizzieLet0_4MQNode_4QVal_Bool_3QNode_Bool_2_bufchan_buf[0] ? lizzieLet0_4MQNode_4QVal_Bool_3QNode_Bool_2_bufchan_buf :
                                                                 lizzieLet0_4MQNode_4QVal_Bool_3QNode_Bool_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QVal_Bool_3QNode_Bool_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet0_4MQNode_4QVal_Bool_3QNode_Bool_2_argbuf_r && lizzieLet0_4MQNode_4QVal_Bool_3QNode_Bool_2_bufchan_buf[0]))
        lizzieLet0_4MQNode_4QVal_Bool_3QNode_Bool_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet0_4MQNode_4QVal_Bool_3QNode_Bool_2_argbuf_r) && (! lizzieLet0_4MQNode_4QVal_Bool_3QNode_Bool_2_bufchan_buf[0])))
        lizzieLet0_4MQNode_4QVal_Bool_3QNode_Bool_2_bufchan_buf <= lizzieLet0_4MQNode_4QVal_Bool_3QNode_Bool_2_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet0_4MQNode_4QVal_Bool_3QNone_Bool,Go) > [(lizzieLet0_4MQNode_4QVal_Bool_3QNone_Bool_1,Go),
                                                                 (lizzieLet0_4MQNode_4QVal_Bool_3QNone_Bool_2,Go)] */
  logic [1:0] lizzieLet0_4MQNode_4QVal_Bool_3QNone_Bool_emitted;
  logic [1:0] lizzieLet0_4MQNode_4QVal_Bool_3QNone_Bool_done;
  assign lizzieLet0_4MQNode_4QVal_Bool_3QNone_Bool_1_d = (lizzieLet0_4MQNode_4QVal_Bool_3QNone_Bool_d[0] && (! lizzieLet0_4MQNode_4QVal_Bool_3QNone_Bool_emitted[0]));
  assign lizzieLet0_4MQNode_4QVal_Bool_3QNone_Bool_2_d = (lizzieLet0_4MQNode_4QVal_Bool_3QNone_Bool_d[0] && (! lizzieLet0_4MQNode_4QVal_Bool_3QNone_Bool_emitted[1]));
  assign lizzieLet0_4MQNode_4QVal_Bool_3QNone_Bool_done = (lizzieLet0_4MQNode_4QVal_Bool_3QNone_Bool_emitted | ({lizzieLet0_4MQNode_4QVal_Bool_3QNone_Bool_2_d[0],
                                                                                                                 lizzieLet0_4MQNode_4QVal_Bool_3QNone_Bool_1_d[0]} & {lizzieLet0_4MQNode_4QVal_Bool_3QNone_Bool_2_r,
                                                                                                                                                                      lizzieLet0_4MQNode_4QVal_Bool_3QNone_Bool_1_r}));
  assign lizzieLet0_4MQNode_4QVal_Bool_3QNone_Bool_r = (& lizzieLet0_4MQNode_4QVal_Bool_3QNone_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QVal_Bool_3QNone_Bool_emitted <= 2'd0;
    else
      lizzieLet0_4MQNode_4QVal_Bool_3QNone_Bool_emitted <= (lizzieLet0_4MQNode_4QVal_Bool_3QNone_Bool_r ? 2'd0 :
                                                            lizzieLet0_4MQNode_4QVal_Bool_3QNone_Bool_done);
  
  /* dcon (Ty QTree_Bool,
      Dcon QError_Bool) : [(lizzieLet0_4MQNode_4QVal_Bool_3QNone_Bool_1,Go)] > (lizzieLet0_4MQNode_4QVal_Bool_3QNone_Bool_1QError_Bool,QTree_Bool) */
  assign lizzieLet0_4MQNode_4QVal_Bool_3QNone_Bool_1QError_Bool_d = QError_Bool_dc((& {lizzieLet0_4MQNode_4QVal_Bool_3QNone_Bool_1_d[0]}), lizzieLet0_4MQNode_4QVal_Bool_3QNone_Bool_1_d);
  assign {lizzieLet0_4MQNode_4QVal_Bool_3QNone_Bool_1_r} = {1 {(lizzieLet0_4MQNode_4QVal_Bool_3QNone_Bool_1QError_Bool_r && lizzieLet0_4MQNode_4QVal_Bool_3QNone_Bool_1QError_Bool_d[0])}};
  
  /* buf (Ty QTree_Bool) : (lizzieLet0_4MQNode_4QVal_Bool_3QNone_Bool_1QError_Bool,QTree_Bool) > (lizzieLet9_1_argbuf,QTree_Bool) */
  QTree_Bool_t lizzieLet0_4MQNode_4QVal_Bool_3QNone_Bool_1QError_Bool_bufchan_d;
  logic lizzieLet0_4MQNode_4QVal_Bool_3QNone_Bool_1QError_Bool_bufchan_r;
  assign lizzieLet0_4MQNode_4QVal_Bool_3QNone_Bool_1QError_Bool_r = ((! lizzieLet0_4MQNode_4QVal_Bool_3QNone_Bool_1QError_Bool_bufchan_d[0]) || lizzieLet0_4MQNode_4QVal_Bool_3QNone_Bool_1QError_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QVal_Bool_3QNone_Bool_1QError_Bool_bufchan_d <= {66'd0,
                                                                           1'd0};
    else
      if (lizzieLet0_4MQNode_4QVal_Bool_3QNone_Bool_1QError_Bool_r)
        lizzieLet0_4MQNode_4QVal_Bool_3QNone_Bool_1QError_Bool_bufchan_d <= lizzieLet0_4MQNode_4QVal_Bool_3QNone_Bool_1QError_Bool_d;
  QTree_Bool_t lizzieLet0_4MQNode_4QVal_Bool_3QNone_Bool_1QError_Bool_bufchan_buf;
  assign lizzieLet0_4MQNode_4QVal_Bool_3QNone_Bool_1QError_Bool_bufchan_r = (! lizzieLet0_4MQNode_4QVal_Bool_3QNone_Bool_1QError_Bool_bufchan_buf[0]);
  assign lizzieLet9_1_argbuf_d = (lizzieLet0_4MQNode_4QVal_Bool_3QNone_Bool_1QError_Bool_bufchan_buf[0] ? lizzieLet0_4MQNode_4QVal_Bool_3QNone_Bool_1QError_Bool_bufchan_buf :
                                  lizzieLet0_4MQNode_4QVal_Bool_3QNone_Bool_1QError_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QVal_Bool_3QNone_Bool_1QError_Bool_bufchan_buf <= {66'd0,
                                                                             1'd0};
    else
      if ((lizzieLet9_1_argbuf_r && lizzieLet0_4MQNode_4QVal_Bool_3QNone_Bool_1QError_Bool_bufchan_buf[0]))
        lizzieLet0_4MQNode_4QVal_Bool_3QNone_Bool_1QError_Bool_bufchan_buf <= {66'd0,
                                                                               1'd0};
      else if (((! lizzieLet9_1_argbuf_r) && (! lizzieLet0_4MQNode_4QVal_Bool_3QNone_Bool_1QError_Bool_bufchan_buf[0])))
        lizzieLet0_4MQNode_4QVal_Bool_3QNone_Bool_1QError_Bool_bufchan_buf <= lizzieLet0_4MQNode_4QVal_Bool_3QNone_Bool_1QError_Bool_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet0_4MQNode_4QVal_Bool_3QNone_Bool_2,Go) > (lizzieLet0_4MQNode_4QVal_Bool_3QNone_Bool_2_argbuf,Go) */
  Go_t lizzieLet0_4MQNode_4QVal_Bool_3QNone_Bool_2_bufchan_d;
  logic lizzieLet0_4MQNode_4QVal_Bool_3QNone_Bool_2_bufchan_r;
  assign lizzieLet0_4MQNode_4QVal_Bool_3QNone_Bool_2_r = ((! lizzieLet0_4MQNode_4QVal_Bool_3QNone_Bool_2_bufchan_d[0]) || lizzieLet0_4MQNode_4QVal_Bool_3QNone_Bool_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QVal_Bool_3QNone_Bool_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet0_4MQNode_4QVal_Bool_3QNone_Bool_2_r)
        lizzieLet0_4MQNode_4QVal_Bool_3QNone_Bool_2_bufchan_d <= lizzieLet0_4MQNode_4QVal_Bool_3QNone_Bool_2_d;
  Go_t lizzieLet0_4MQNode_4QVal_Bool_3QNone_Bool_2_bufchan_buf;
  assign lizzieLet0_4MQNode_4QVal_Bool_3QNone_Bool_2_bufchan_r = (! lizzieLet0_4MQNode_4QVal_Bool_3QNone_Bool_2_bufchan_buf[0]);
  assign lizzieLet0_4MQNode_4QVal_Bool_3QNone_Bool_2_argbuf_d = (lizzieLet0_4MQNode_4QVal_Bool_3QNone_Bool_2_bufchan_buf[0] ? lizzieLet0_4MQNode_4QVal_Bool_3QNone_Bool_2_bufchan_buf :
                                                                 lizzieLet0_4MQNode_4QVal_Bool_3QNone_Bool_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QVal_Bool_3QNone_Bool_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet0_4MQNode_4QVal_Bool_3QNone_Bool_2_argbuf_r && lizzieLet0_4MQNode_4QVal_Bool_3QNone_Bool_2_bufchan_buf[0]))
        lizzieLet0_4MQNode_4QVal_Bool_3QNone_Bool_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet0_4MQNode_4QVal_Bool_3QNone_Bool_2_argbuf_r) && (! lizzieLet0_4MQNode_4QVal_Bool_3QNone_Bool_2_bufchan_buf[0])))
        lizzieLet0_4MQNode_4QVal_Bool_3QNone_Bool_2_bufchan_buf <= lizzieLet0_4MQNode_4QVal_Bool_3QNone_Bool_2_bufchan_d;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_CTf) : (lizzieLet0_4MQNode_4QVal_Bool_4,QTree_Bool) (lizzieLet0_4MQNode_5QVal_Bool,Pointer_CTf) > [(lizzieLet0_4MQNode_4QVal_Bool_4QNone_Bool,Pointer_CTf),
                                                                                                                     (lizzieLet0_4MQNode_4QVal_Bool_4QVal_Bool,Pointer_CTf),
                                                                                                                     (lizzieLet0_4MQNode_4QVal_Bool_4QNode_Bool,Pointer_CTf),
                                                                                                                     (lizzieLet0_4MQNode_4QVal_Bool_4QError_Bool,Pointer_CTf)] */
  logic [3:0] lizzieLet0_4MQNode_5QVal_Bool_onehotd;
  always_comb
    if ((lizzieLet0_4MQNode_4QVal_Bool_4_d[0] && lizzieLet0_4MQNode_5QVal_Bool_d[0]))
      unique case (lizzieLet0_4MQNode_4QVal_Bool_4_d[2:1])
        2'd0: lizzieLet0_4MQNode_5QVal_Bool_onehotd = 4'd1;
        2'd1: lizzieLet0_4MQNode_5QVal_Bool_onehotd = 4'd2;
        2'd2: lizzieLet0_4MQNode_5QVal_Bool_onehotd = 4'd4;
        2'd3: lizzieLet0_4MQNode_5QVal_Bool_onehotd = 4'd8;
        default: lizzieLet0_4MQNode_5QVal_Bool_onehotd = 4'd0;
      endcase
    else lizzieLet0_4MQNode_5QVal_Bool_onehotd = 4'd0;
  assign lizzieLet0_4MQNode_4QVal_Bool_4QNone_Bool_d = {lizzieLet0_4MQNode_5QVal_Bool_d[16:1],
                                                        lizzieLet0_4MQNode_5QVal_Bool_onehotd[0]};
  assign lizzieLet0_4MQNode_4QVal_Bool_4QVal_Bool_d = {lizzieLet0_4MQNode_5QVal_Bool_d[16:1],
                                                       lizzieLet0_4MQNode_5QVal_Bool_onehotd[1]};
  assign lizzieLet0_4MQNode_4QVal_Bool_4QNode_Bool_d = {lizzieLet0_4MQNode_5QVal_Bool_d[16:1],
                                                        lizzieLet0_4MQNode_5QVal_Bool_onehotd[2]};
  assign lizzieLet0_4MQNode_4QVal_Bool_4QError_Bool_d = {lizzieLet0_4MQNode_5QVal_Bool_d[16:1],
                                                         lizzieLet0_4MQNode_5QVal_Bool_onehotd[3]};
  assign lizzieLet0_4MQNode_5QVal_Bool_r = (| (lizzieLet0_4MQNode_5QVal_Bool_onehotd & {lizzieLet0_4MQNode_4QVal_Bool_4QError_Bool_r,
                                                                                        lizzieLet0_4MQNode_4QVal_Bool_4QNode_Bool_r,
                                                                                        lizzieLet0_4MQNode_4QVal_Bool_4QVal_Bool_r,
                                                                                        lizzieLet0_4MQNode_4QVal_Bool_4QNone_Bool_r}));
  assign lizzieLet0_4MQNode_4QVal_Bool_4_r = lizzieLet0_4MQNode_5QVal_Bool_r;
  
  /* buf (Ty Pointer_CTf) : (lizzieLet0_4MQNode_4QVal_Bool_4QError_Bool,Pointer_CTf) > (lizzieLet0_4MQNode_4QVal_Bool_4QError_Bool_1_argbuf,Pointer_CTf) */
  Pointer_CTf_t lizzieLet0_4MQNode_4QVal_Bool_4QError_Bool_bufchan_d;
  logic lizzieLet0_4MQNode_4QVal_Bool_4QError_Bool_bufchan_r;
  assign lizzieLet0_4MQNode_4QVal_Bool_4QError_Bool_r = ((! lizzieLet0_4MQNode_4QVal_Bool_4QError_Bool_bufchan_d[0]) || lizzieLet0_4MQNode_4QVal_Bool_4QError_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QVal_Bool_4QError_Bool_bufchan_d <= {16'd0,
                                                               1'd0};
    else
      if (lizzieLet0_4MQNode_4QVal_Bool_4QError_Bool_r)
        lizzieLet0_4MQNode_4QVal_Bool_4QError_Bool_bufchan_d <= lizzieLet0_4MQNode_4QVal_Bool_4QError_Bool_d;
  Pointer_CTf_t lizzieLet0_4MQNode_4QVal_Bool_4QError_Bool_bufchan_buf;
  assign lizzieLet0_4MQNode_4QVal_Bool_4QError_Bool_bufchan_r = (! lizzieLet0_4MQNode_4QVal_Bool_4QError_Bool_bufchan_buf[0]);
  assign lizzieLet0_4MQNode_4QVal_Bool_4QError_Bool_1_argbuf_d = (lizzieLet0_4MQNode_4QVal_Bool_4QError_Bool_bufchan_buf[0] ? lizzieLet0_4MQNode_4QVal_Bool_4QError_Bool_bufchan_buf :
                                                                  lizzieLet0_4MQNode_4QVal_Bool_4QError_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QVal_Bool_4QError_Bool_bufchan_buf <= {16'd0,
                                                                 1'd0};
    else
      if ((lizzieLet0_4MQNode_4QVal_Bool_4QError_Bool_1_argbuf_r && lizzieLet0_4MQNode_4QVal_Bool_4QError_Bool_bufchan_buf[0]))
        lizzieLet0_4MQNode_4QVal_Bool_4QError_Bool_bufchan_buf <= {16'd0,
                                                                   1'd0};
      else if (((! lizzieLet0_4MQNode_4QVal_Bool_4QError_Bool_1_argbuf_r) && (! lizzieLet0_4MQNode_4QVal_Bool_4QError_Bool_bufchan_buf[0])))
        lizzieLet0_4MQNode_4QVal_Bool_4QError_Bool_bufchan_buf <= lizzieLet0_4MQNode_4QVal_Bool_4QError_Bool_bufchan_d;
  
  /* buf (Ty Pointer_CTf) : (lizzieLet0_4MQNode_4QVal_Bool_4QNode_Bool,Pointer_CTf) > (lizzieLet0_4MQNode_4QVal_Bool_4QNode_Bool_1_argbuf,Pointer_CTf) */
  Pointer_CTf_t lizzieLet0_4MQNode_4QVal_Bool_4QNode_Bool_bufchan_d;
  logic lizzieLet0_4MQNode_4QVal_Bool_4QNode_Bool_bufchan_r;
  assign lizzieLet0_4MQNode_4QVal_Bool_4QNode_Bool_r = ((! lizzieLet0_4MQNode_4QVal_Bool_4QNode_Bool_bufchan_d[0]) || lizzieLet0_4MQNode_4QVal_Bool_4QNode_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QVal_Bool_4QNode_Bool_bufchan_d <= {16'd0,
                                                              1'd0};
    else
      if (lizzieLet0_4MQNode_4QVal_Bool_4QNode_Bool_r)
        lizzieLet0_4MQNode_4QVal_Bool_4QNode_Bool_bufchan_d <= lizzieLet0_4MQNode_4QVal_Bool_4QNode_Bool_d;
  Pointer_CTf_t lizzieLet0_4MQNode_4QVal_Bool_4QNode_Bool_bufchan_buf;
  assign lizzieLet0_4MQNode_4QVal_Bool_4QNode_Bool_bufchan_r = (! lizzieLet0_4MQNode_4QVal_Bool_4QNode_Bool_bufchan_buf[0]);
  assign lizzieLet0_4MQNode_4QVal_Bool_4QNode_Bool_1_argbuf_d = (lizzieLet0_4MQNode_4QVal_Bool_4QNode_Bool_bufchan_buf[0] ? lizzieLet0_4MQNode_4QVal_Bool_4QNode_Bool_bufchan_buf :
                                                                 lizzieLet0_4MQNode_4QVal_Bool_4QNode_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QVal_Bool_4QNode_Bool_bufchan_buf <= {16'd0,
                                                                1'd0};
    else
      if ((lizzieLet0_4MQNode_4QVal_Bool_4QNode_Bool_1_argbuf_r && lizzieLet0_4MQNode_4QVal_Bool_4QNode_Bool_bufchan_buf[0]))
        lizzieLet0_4MQNode_4QVal_Bool_4QNode_Bool_bufchan_buf <= {16'd0,
                                                                  1'd0};
      else if (((! lizzieLet0_4MQNode_4QVal_Bool_4QNode_Bool_1_argbuf_r) && (! lizzieLet0_4MQNode_4QVal_Bool_4QNode_Bool_bufchan_buf[0])))
        lizzieLet0_4MQNode_4QVal_Bool_4QNode_Bool_bufchan_buf <= lizzieLet0_4MQNode_4QVal_Bool_4QNode_Bool_bufchan_d;
  
  /* buf (Ty Pointer_CTf) : (lizzieLet0_4MQNode_4QVal_Bool_4QNone_Bool,Pointer_CTf) > (lizzieLet0_4MQNode_4QVal_Bool_4QNone_Bool_1_argbuf,Pointer_CTf) */
  Pointer_CTf_t lizzieLet0_4MQNode_4QVal_Bool_4QNone_Bool_bufchan_d;
  logic lizzieLet0_4MQNode_4QVal_Bool_4QNone_Bool_bufchan_r;
  assign lizzieLet0_4MQNode_4QVal_Bool_4QNone_Bool_r = ((! lizzieLet0_4MQNode_4QVal_Bool_4QNone_Bool_bufchan_d[0]) || lizzieLet0_4MQNode_4QVal_Bool_4QNone_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QVal_Bool_4QNone_Bool_bufchan_d <= {16'd0,
                                                              1'd0};
    else
      if (lizzieLet0_4MQNode_4QVal_Bool_4QNone_Bool_r)
        lizzieLet0_4MQNode_4QVal_Bool_4QNone_Bool_bufchan_d <= lizzieLet0_4MQNode_4QVal_Bool_4QNone_Bool_d;
  Pointer_CTf_t lizzieLet0_4MQNode_4QVal_Bool_4QNone_Bool_bufchan_buf;
  assign lizzieLet0_4MQNode_4QVal_Bool_4QNone_Bool_bufchan_r = (! lizzieLet0_4MQNode_4QVal_Bool_4QNone_Bool_bufchan_buf[0]);
  assign lizzieLet0_4MQNode_4QVal_Bool_4QNone_Bool_1_argbuf_d = (lizzieLet0_4MQNode_4QVal_Bool_4QNone_Bool_bufchan_buf[0] ? lizzieLet0_4MQNode_4QVal_Bool_4QNone_Bool_bufchan_buf :
                                                                 lizzieLet0_4MQNode_4QVal_Bool_4QNone_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QVal_Bool_4QNone_Bool_bufchan_buf <= {16'd0,
                                                                1'd0};
    else
      if ((lizzieLet0_4MQNode_4QVal_Bool_4QNone_Bool_1_argbuf_r && lizzieLet0_4MQNode_4QVal_Bool_4QNone_Bool_bufchan_buf[0]))
        lizzieLet0_4MQNode_4QVal_Bool_4QNone_Bool_bufchan_buf <= {16'd0,
                                                                  1'd0};
      else if (((! lizzieLet0_4MQNode_4QVal_Bool_4QNone_Bool_1_argbuf_r) && (! lizzieLet0_4MQNode_4QVal_Bool_4QNone_Bool_bufchan_buf[0])))
        lizzieLet0_4MQNode_4QVal_Bool_4QNone_Bool_bufchan_buf <= lizzieLet0_4MQNode_4QVal_Bool_4QNone_Bool_bufchan_d;
  
  /* demux (Ty QTree_Bool,
       Ty MyBool) : (lizzieLet0_4MQNode_4QVal_Bool_5,QTree_Bool) (v1a8h_destruct,MyBool) > [(_81,MyBool),
                                                                                            (lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool,MyBool),
                                                                                            (_80,MyBool),
                                                                                            (_79,MyBool)] */
  logic [3:0] v1a8h_destruct_onehotd;
  always_comb
    if ((lizzieLet0_4MQNode_4QVal_Bool_5_d[0] && v1a8h_destruct_d[0]))
      unique case (lizzieLet0_4MQNode_4QVal_Bool_5_d[2:1])
        2'd0: v1a8h_destruct_onehotd = 4'd1;
        2'd1: v1a8h_destruct_onehotd = 4'd2;
        2'd2: v1a8h_destruct_onehotd = 4'd4;
        2'd3: v1a8h_destruct_onehotd = 4'd8;
        default: v1a8h_destruct_onehotd = 4'd0;
      endcase
    else v1a8h_destruct_onehotd = 4'd0;
  assign _81_d = {v1a8h_destruct_d[1:1], v1a8h_destruct_onehotd[0]};
  assign lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_d = {v1a8h_destruct_d[1:1],
                                                       v1a8h_destruct_onehotd[1]};
  assign _80_d = {v1a8h_destruct_d[1:1], v1a8h_destruct_onehotd[2]};
  assign _79_d = {v1a8h_destruct_d[1:1], v1a8h_destruct_onehotd[3]};
  assign v1a8h_destruct_r = (| (v1a8h_destruct_onehotd & {_79_r,
                                                          _80_r,
                                                          lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_r,
                                                          _81_r}));
  assign lizzieLet0_4MQNode_4QVal_Bool_5_r = v1a8h_destruct_r;
  
  /* fork (Ty MyBool) : (lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool,MyBool) > [(lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1,MyBool),
                                                                        (lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_2,MyBool),
                                                                        (lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3,MyBool)] */
  logic [2:0] lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_emitted;
  logic [2:0] lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_done;
  assign lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1_d = {lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_d[1:1],
                                                         (lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_d[0] && (! lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_emitted[0]))};
  assign lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_2_d = {lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_d[1:1],
                                                         (lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_d[0] && (! lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_emitted[1]))};
  assign lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3_d = {lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_d[1:1],
                                                         (lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_d[0] && (! lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_emitted[2]))};
  assign lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_done = (lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_emitted | ({lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3_d[0],
                                                                                                               lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_2_d[0],
                                                                                                               lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1_d[0]} & {lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3_r,
                                                                                                                                                                   lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_2_r,
                                                                                                                                                                   lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1_r}));
  assign lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_r = (& lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_emitted <= 3'd0;
    else
      lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_emitted <= (lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_r ? 3'd0 :
                                                           lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_done);
  
  /* demux (Ty MyBool,
       Ty Go) : (lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1,MyBool) (lizzieLet0_4MQNode_4QVal_Bool_3QVal_Bool,Go) > [(lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyFalse,Go),
                                                                                                                     (lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyTrue,Go)] */
  logic [1:0] lizzieLet0_4MQNode_4QVal_Bool_3QVal_Bool_onehotd;
  always_comb
    if ((lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1_d[0] && lizzieLet0_4MQNode_4QVal_Bool_3QVal_Bool_d[0]))
      unique case (lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1_d[1:1])
        1'd0: lizzieLet0_4MQNode_4QVal_Bool_3QVal_Bool_onehotd = 2'd1;
        1'd1: lizzieLet0_4MQNode_4QVal_Bool_3QVal_Bool_onehotd = 2'd2;
        default: lizzieLet0_4MQNode_4QVal_Bool_3QVal_Bool_onehotd = 2'd0;
      endcase
    else lizzieLet0_4MQNode_4QVal_Bool_3QVal_Bool_onehotd = 2'd0;
  assign lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyFalse_d = lizzieLet0_4MQNode_4QVal_Bool_3QVal_Bool_onehotd[0];
  assign lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyTrue_d = lizzieLet0_4MQNode_4QVal_Bool_3QVal_Bool_onehotd[1];
  assign lizzieLet0_4MQNode_4QVal_Bool_3QVal_Bool_r = (| (lizzieLet0_4MQNode_4QVal_Bool_3QVal_Bool_onehotd & {lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyTrue_r,
                                                                                                              lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyFalse_r}));
  assign lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1_r = lizzieLet0_4MQNode_4QVal_Bool_3QVal_Bool_r;
  
  /* fork (Ty Go) : (lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyTrue,Go) > [(lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyTrue_1,Go),
                                                                        (lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyTrue_2,Go)] */
  logic [1:0] lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyTrue_emitted;
  logic [1:0] lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyTrue_done;
  assign lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyTrue_1_d = (lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyTrue_d[0] && (! lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyTrue_emitted[0]));
  assign lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyTrue_2_d = (lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyTrue_d[0] && (! lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyTrue_emitted[1]));
  assign lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyTrue_done = (lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyTrue_emitted | ({lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyTrue_2_d[0],
                                                                                                                               lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyTrue_1_d[0]} & {lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyTrue_2_r,
                                                                                                                                                                                           lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyTrue_1_r}));
  assign lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyTrue_r = (& lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyTrue_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyTrue_emitted <= 2'd0;
    else
      lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyTrue_emitted <= (lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyTrue_r ? 2'd0 :
                                                                   lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyTrue_done);
  
  /* dcon (Ty QTree_Bool,
      Dcon QError_Bool) : [(lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyTrue_1,Go)] > (lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyTrue_1QError_Bool,QTree_Bool) */
  assign lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyTrue_1QError_Bool_d = QError_Bool_dc((& {lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyTrue_1_d[0]}), lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyTrue_1_d);
  assign {lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyTrue_1_r} = {1 {(lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyTrue_1QError_Bool_r && lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyTrue_1QError_Bool_d[0])}};
  
  /* buf (Ty QTree_Bool) : (lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyTrue_1QError_Bool,QTree_Bool) > (lizzieLet12_1_argbuf,QTree_Bool) */
  QTree_Bool_t lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyTrue_1QError_Bool_bufchan_d;
  logic lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyTrue_1QError_Bool_bufchan_r;
  assign lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyTrue_1QError_Bool_r = ((! lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyTrue_1QError_Bool_bufchan_d[0]) || lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyTrue_1QError_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyTrue_1QError_Bool_bufchan_d <= {66'd0,
                                                                                  1'd0};
    else
      if (lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyTrue_1QError_Bool_r)
        lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyTrue_1QError_Bool_bufchan_d <= lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyTrue_1QError_Bool_d;
  QTree_Bool_t lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyTrue_1QError_Bool_bufchan_buf;
  assign lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyTrue_1QError_Bool_bufchan_r = (! lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyTrue_1QError_Bool_bufchan_buf[0]);
  assign lizzieLet12_1_argbuf_d = (lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyTrue_1QError_Bool_bufchan_buf[0] ? lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyTrue_1QError_Bool_bufchan_buf :
                                   lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyTrue_1QError_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyTrue_1QError_Bool_bufchan_buf <= {66'd0,
                                                                                    1'd0};
    else
      if ((lizzieLet12_1_argbuf_r && lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyTrue_1QError_Bool_bufchan_buf[0]))
        lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyTrue_1QError_Bool_bufchan_buf <= {66'd0,
                                                                                      1'd0};
      else if (((! lizzieLet12_1_argbuf_r) && (! lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyTrue_1QError_Bool_bufchan_buf[0])))
        lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyTrue_1QError_Bool_bufchan_buf <= lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyTrue_1QError_Bool_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyTrue_2,Go) > (lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyTrue_2_argbuf,Go) */
  Go_t lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyTrue_2_bufchan_d;
  logic lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyTrue_2_bufchan_r;
  assign lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyTrue_2_r = ((! lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyTrue_2_bufchan_d[0]) || lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyTrue_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyTrue_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyTrue_2_r)
        lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyTrue_2_bufchan_d <= lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyTrue_2_d;
  Go_t lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyTrue_2_bufchan_buf;
  assign lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyTrue_2_bufchan_r = (! lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyTrue_2_bufchan_buf[0]);
  assign lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyTrue_2_argbuf_d = (lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyTrue_2_bufchan_buf[0] ? lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyTrue_2_bufchan_buf :
                                                                        lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyTrue_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyTrue_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyTrue_2_argbuf_r && lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyTrue_2_bufchan_buf[0]))
        lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyTrue_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyTrue_2_argbuf_r) && (! lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyTrue_2_bufchan_buf[0])))
        lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyTrue_2_bufchan_buf <= lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyTrue_2_bufchan_d;
  
  /* demux (Ty MyBool,
       Ty Pointer_CTf) : (lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_2,MyBool) (lizzieLet0_4MQNode_4QVal_Bool_4QVal_Bool,Pointer_CTf) > [(lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_2MyFalse,Pointer_CTf),
                                                                                                                                       (lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_2MyTrue,Pointer_CTf)] */
  logic [1:0] lizzieLet0_4MQNode_4QVal_Bool_4QVal_Bool_onehotd;
  always_comb
    if ((lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_2_d[0] && lizzieLet0_4MQNode_4QVal_Bool_4QVal_Bool_d[0]))
      unique case (lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_2_d[1:1])
        1'd0: lizzieLet0_4MQNode_4QVal_Bool_4QVal_Bool_onehotd = 2'd1;
        1'd1: lizzieLet0_4MQNode_4QVal_Bool_4QVal_Bool_onehotd = 2'd2;
        default: lizzieLet0_4MQNode_4QVal_Bool_4QVal_Bool_onehotd = 2'd0;
      endcase
    else lizzieLet0_4MQNode_4QVal_Bool_4QVal_Bool_onehotd = 2'd0;
  assign lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_2MyFalse_d = {lizzieLet0_4MQNode_4QVal_Bool_4QVal_Bool_d[16:1],
                                                                lizzieLet0_4MQNode_4QVal_Bool_4QVal_Bool_onehotd[0]};
  assign lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_2MyTrue_d = {lizzieLet0_4MQNode_4QVal_Bool_4QVal_Bool_d[16:1],
                                                               lizzieLet0_4MQNode_4QVal_Bool_4QVal_Bool_onehotd[1]};
  assign lizzieLet0_4MQNode_4QVal_Bool_4QVal_Bool_r = (| (lizzieLet0_4MQNode_4QVal_Bool_4QVal_Bool_onehotd & {lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_2MyTrue_r,
                                                                                                              lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_2MyFalse_r}));
  assign lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_2_r = lizzieLet0_4MQNode_4QVal_Bool_4QVal_Bool_r;
  
  /* buf (Ty Pointer_CTf) : (lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_2MyTrue,Pointer_CTf) > (lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_2MyTrue_1_argbuf,Pointer_CTf) */
  Pointer_CTf_t lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_2MyTrue_bufchan_d;
  logic lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_2MyTrue_bufchan_r;
  assign lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_2MyTrue_r = ((! lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_2MyTrue_bufchan_d[0]) || lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_2MyTrue_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_2MyTrue_bufchan_d <= {16'd0,
                                                                     1'd0};
    else
      if (lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_2MyTrue_r)
        lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_2MyTrue_bufchan_d <= lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_2MyTrue_d;
  Pointer_CTf_t lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_2MyTrue_bufchan_buf;
  assign lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_2MyTrue_bufchan_r = (! lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_2MyTrue_bufchan_buf[0]);
  assign lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_2MyTrue_1_argbuf_d = (lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_2MyTrue_bufchan_buf[0] ? lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_2MyTrue_bufchan_buf :
                                                                        lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_2MyTrue_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_2MyTrue_bufchan_buf <= {16'd0,
                                                                       1'd0};
    else
      if ((lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_2MyTrue_1_argbuf_r && lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_2MyTrue_bufchan_buf[0]))
        lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_2MyTrue_bufchan_buf <= {16'd0,
                                                                         1'd0};
      else if (((! lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_2MyTrue_1_argbuf_r) && (! lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_2MyTrue_bufchan_buf[0])))
        lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_2MyTrue_bufchan_buf <= lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_2MyTrue_bufchan_d;
  
  /* demux (Ty MyBool,
       Ty MyBool) : (lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3,MyBool) (va8i_destruct,MyBool) > [(lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse,MyBool),
                                                                                                  (_78,MyBool)] */
  logic [1:0] va8i_destruct_onehotd;
  always_comb
    if ((lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3_d[0] && va8i_destruct_d[0]))
      unique case (lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3_d[1:1])
        1'd0: va8i_destruct_onehotd = 2'd1;
        1'd1: va8i_destruct_onehotd = 2'd2;
        default: va8i_destruct_onehotd = 2'd0;
      endcase
    else va8i_destruct_onehotd = 2'd0;
  assign lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_d = {va8i_destruct_d[1:1],
                                                                va8i_destruct_onehotd[0]};
  assign _78_d = {va8i_destruct_d[1:1], va8i_destruct_onehotd[1]};
  assign va8i_destruct_r = (| (va8i_destruct_onehotd & {_78_r,
                                                        lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_r}));
  assign lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3_r = va8i_destruct_r;
  
  /* fork (Ty MyBool) : (lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse,MyBool) > [(lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1,MyBool),
                                                                                 (lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_2,MyBool)] */
  logic [1:0] lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_emitted;
  logic [1:0] lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_done;
  assign lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1_d = {lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_d[1:1],
                                                                  (lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_d[0] && (! lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_emitted[0]))};
  assign lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_2_d = {lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_d[1:1],
                                                                  (lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_d[0] && (! lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_emitted[1]))};
  assign lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_done = (lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_emitted | ({lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_2_d[0],
                                                                                                                                 lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1_d[0]} & {lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_2_r,
                                                                                                                                                                                              lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1_r}));
  assign lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_r = (& lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_emitted <= 2'd0;
    else
      lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_emitted <= (lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_r ? 2'd0 :
                                                                    lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_done);
  
  /* demux (Ty MyBool,
       Ty Go) : (lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1,MyBool) (lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyFalse,Go) > [(lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyFalse,Go),
                                                                                                                                       (lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyTrue,Go)] */
  logic [1:0] lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyFalse_onehotd;
  always_comb
    if ((lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1_d[0] && lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyFalse_d[0]))
      unique case (lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1_d[1:1])
        1'd0:
          lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyFalse_onehotd = 2'd1;
        1'd1:
          lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyFalse_onehotd = 2'd2;
        default:
          lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyFalse_onehotd = 2'd0;
      endcase
    else
      lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyFalse_onehotd = 2'd0;
  assign lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyFalse_d = lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyFalse_onehotd[0];
  assign lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyTrue_d = lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyFalse_onehotd[1];
  assign lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyFalse_r = (| (lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyFalse_onehotd & {lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyTrue_r,
                                                                                                                                lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyFalse_r}));
  assign lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1_r = lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_1MyFalse_r;
  
  /* fork (Ty Go) : (lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyFalse,Go) > [(lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyFalse_1,Go),
                                                                                  (lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyFalse_2,Go)] */
  logic [1:0] lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyFalse_emitted;
  logic [1:0] lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyFalse_done;
  assign lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyFalse_1_d = (lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyFalse_d[0] && (! lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyFalse_emitted[0]));
  assign lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyFalse_2_d = (lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyFalse_d[0] && (! lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyFalse_emitted[1]));
  assign lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyFalse_done = (lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyFalse_emitted | ({lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyFalse_2_d[0],
                                                                                                                                                   lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyFalse_1_d[0]} & {lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyFalse_2_r,
                                                                                                                                                                                                                         lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyFalse_1_r}));
  assign lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyFalse_r = (& lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyFalse_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyFalse_emitted <= 2'd0;
    else
      lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyFalse_emitted <= (lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyFalse_r ? 2'd0 :
                                                                             lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyFalse_done);
  
  /* dcon (Ty QTree_Bool,
      Dcon QNone_Bool) : [(lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyFalse_1,Go)] > (lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool,QTree_Bool) */
  assign lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_d = QNone_Bool_dc((& {lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyFalse_1_d[0]}), lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyFalse_1_d);
  assign {lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyFalse_1_r} = {1 {(lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_r && lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_d[0])}};
  
  /* buf (Ty QTree_Bool) : (lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool,QTree_Bool) > (lizzieLet10_1_argbuf,QTree_Bool) */
  QTree_Bool_t lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_bufchan_d;
  logic lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_bufchan_r;
  assign lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_r = ((! lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_bufchan_d[0]) || lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_bufchan_d <= {66'd0,
                                                                                           1'd0};
    else
      if (lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_r)
        lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_bufchan_d <= lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_d;
  QTree_Bool_t lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_bufchan_buf;
  assign lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_bufchan_r = (! lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_bufchan_buf[0]);
  assign lizzieLet10_1_argbuf_d = (lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_bufchan_buf[0] ? lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_bufchan_buf :
                                   lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_bufchan_buf <= {66'd0,
                                                                                             1'd0};
    else
      if ((lizzieLet10_1_argbuf_r && lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_bufchan_buf[0]))
        lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_bufchan_buf <= {66'd0,
                                                                                               1'd0};
      else if (((! lizzieLet10_1_argbuf_r) && (! lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_bufchan_buf[0])))
        lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_bufchan_buf <= lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyFalse_2,Go) > (lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyFalse_2_argbuf,Go) */
  Go_t lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyFalse_2_bufchan_d;
  logic lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyFalse_2_bufchan_r;
  assign lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyFalse_2_r = ((! lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyFalse_2_bufchan_d[0]) || lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyFalse_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyFalse_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyFalse_2_r)
        lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyFalse_2_bufchan_d <= lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyFalse_2_d;
  Go_t lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyFalse_2_bufchan_buf;
  assign lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyFalse_2_bufchan_r = (! lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyFalse_2_bufchan_buf[0]);
  assign lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyFalse_2_argbuf_d = (lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyFalse_2_bufchan_buf[0] ? lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyFalse_2_bufchan_buf :
                                                                                  lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyFalse_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyFalse_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyFalse_2_argbuf_r && lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyFalse_2_bufchan_buf[0]))
        lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyFalse_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyFalse_2_argbuf_r) && (! lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyFalse_2_bufchan_buf[0])))
        lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyFalse_2_bufchan_buf <= lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyFalse_2_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyTrue,Go) > [(lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyTrue_1,Go),
                                                                                 (lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyTrue_2,Go)] */
  logic [1:0] lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyTrue_emitted;
  logic [1:0] lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyTrue_done;
  assign lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyTrue_1_d = (lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyTrue_d[0] && (! lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyTrue_emitted[0]));
  assign lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyTrue_2_d = (lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyTrue_d[0] && (! lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyTrue_emitted[1]));
  assign lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyTrue_done = (lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyTrue_emitted | ({lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyTrue_2_d[0],
                                                                                                                                                 lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyTrue_1_d[0]} & {lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyTrue_2_r,
                                                                                                                                                                                                                      lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyTrue_1_r}));
  assign lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyTrue_r = (& lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyTrue_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyTrue_emitted <= 2'd0;
    else
      lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyTrue_emitted <= (lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyTrue_r ? 2'd0 :
                                                                            lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyTrue_done);
  
  /* dcon (Ty QTree_Bool,
      Dcon QError_Bool) : [(lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyTrue_1,Go)] > (lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyTrue_1QError_Bool,QTree_Bool) */
  assign lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyTrue_1QError_Bool_d = QError_Bool_dc((& {lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyTrue_1_d[0]}), lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyTrue_1_d);
  assign {lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyTrue_1_r} = {1 {(lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyTrue_1QError_Bool_r && lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyTrue_1QError_Bool_d[0])}};
  
  /* buf (Ty QTree_Bool) : (lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyTrue_1QError_Bool,QTree_Bool) > (lizzieLet11_1_argbuf,QTree_Bool) */
  QTree_Bool_t lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyTrue_1QError_Bool_bufchan_d;
  logic lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyTrue_1QError_Bool_bufchan_r;
  assign lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyTrue_1QError_Bool_r = ((! lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyTrue_1QError_Bool_bufchan_d[0]) || lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyTrue_1QError_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyTrue_1QError_Bool_bufchan_d <= {66'd0,
                                                                                           1'd0};
    else
      if (lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyTrue_1QError_Bool_r)
        lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyTrue_1QError_Bool_bufchan_d <= lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyTrue_1QError_Bool_d;
  QTree_Bool_t lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyTrue_1QError_Bool_bufchan_buf;
  assign lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyTrue_1QError_Bool_bufchan_r = (! lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyTrue_1QError_Bool_bufchan_buf[0]);
  assign lizzieLet11_1_argbuf_d = (lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyTrue_1QError_Bool_bufchan_buf[0] ? lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyTrue_1QError_Bool_bufchan_buf :
                                   lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyTrue_1QError_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyTrue_1QError_Bool_bufchan_buf <= {66'd0,
                                                                                             1'd0};
    else
      if ((lizzieLet11_1_argbuf_r && lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyTrue_1QError_Bool_bufchan_buf[0]))
        lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyTrue_1QError_Bool_bufchan_buf <= {66'd0,
                                                                                               1'd0};
      else if (((! lizzieLet11_1_argbuf_r) && (! lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyTrue_1QError_Bool_bufchan_buf[0])))
        lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyTrue_1QError_Bool_bufchan_buf <= lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyTrue_1QError_Bool_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyTrue_2,Go) > (lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyTrue_2_argbuf,Go) */
  Go_t lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyTrue_2_bufchan_d;
  logic lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyTrue_2_bufchan_r;
  assign lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyTrue_2_r = ((! lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyTrue_2_bufchan_d[0]) || lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyTrue_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyTrue_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyTrue_2_r)
        lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyTrue_2_bufchan_d <= lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyTrue_2_d;
  Go_t lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyTrue_2_bufchan_buf;
  assign lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyTrue_2_bufchan_r = (! lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyTrue_2_bufchan_buf[0]);
  assign lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyTrue_2_argbuf_d = (lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyTrue_2_bufchan_buf[0] ? lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyTrue_2_bufchan_buf :
                                                                                 lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyTrue_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyTrue_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyTrue_2_argbuf_r && lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyTrue_2_bufchan_buf[0]))
        lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyTrue_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyTrue_2_argbuf_r) && (! lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyTrue_2_bufchan_buf[0])))
        lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyTrue_2_bufchan_buf <= lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_1MyTrue_2_bufchan_d;
  
  /* demux (Ty MyBool,
       Ty Pointer_CTf) : (lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_2,MyBool) (lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_2MyFalse,Pointer_CTf) > [(lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_2MyFalse,Pointer_CTf),
                                                                                                                                                         (lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_2MyTrue,Pointer_CTf)] */
  logic [1:0] lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_2MyFalse_onehotd;
  always_comb
    if ((lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_2_d[0] && lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_2MyFalse_d[0]))
      unique case (lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_2_d[1:1])
        1'd0:
          lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_2MyFalse_onehotd = 2'd1;
        1'd1:
          lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_2MyFalse_onehotd = 2'd2;
        default:
          lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_2MyFalse_onehotd = 2'd0;
      endcase
    else
      lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_2MyFalse_onehotd = 2'd0;
  assign lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_2MyFalse_d = {lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_2MyFalse_d[16:1],
                                                                         lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_2MyFalse_onehotd[0]};
  assign lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_2MyTrue_d = {lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_2MyFalse_d[16:1],
                                                                        lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_2MyFalse_onehotd[1]};
  assign lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_2MyFalse_r = (| (lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_2MyFalse_onehotd & {lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_2MyTrue_r,
                                                                                                                                lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_2MyFalse_r}));
  assign lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_2_r = lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_2MyFalse_r;
  
  /* buf (Ty Pointer_CTf) : (lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_2MyFalse,Pointer_CTf) > (lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_2MyFalse_1_argbuf,Pointer_CTf) */
  Pointer_CTf_t lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_2MyFalse_bufchan_d;
  logic lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_2MyFalse_bufchan_r;
  assign lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_2MyFalse_r = ((! lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_2MyFalse_bufchan_d[0]) || lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_2MyFalse_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_2MyFalse_bufchan_d <= {16'd0,
                                                                               1'd0};
    else
      if (lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_2MyFalse_r)
        lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_2MyFalse_bufchan_d <= lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_2MyFalse_d;
  Pointer_CTf_t lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_2MyFalse_bufchan_buf;
  assign lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_2MyFalse_bufchan_r = (! lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_2MyFalse_bufchan_buf[0]);
  assign lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_2MyFalse_1_argbuf_d = (lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_2MyFalse_bufchan_buf[0] ? lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_2MyFalse_bufchan_buf :
                                                                                  lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_2MyFalse_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_2MyFalse_bufchan_buf <= {16'd0,
                                                                                 1'd0};
    else
      if ((lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_2MyFalse_1_argbuf_r && lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_2MyFalse_bufchan_buf[0]))
        lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_2MyFalse_bufchan_buf <= {16'd0,
                                                                                   1'd0};
      else if (((! lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_2MyFalse_1_argbuf_r) && (! lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_2MyFalse_bufchan_buf[0])))
        lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_2MyFalse_bufchan_buf <= lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_2MyFalse_bufchan_d;
  
  /* buf (Ty Pointer_CTf) : (lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_2MyTrue,Pointer_CTf) > (lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_2MyTrue_1_argbuf,Pointer_CTf) */
  Pointer_CTf_t lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_2MyTrue_bufchan_d;
  logic lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_2MyTrue_bufchan_r;
  assign lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_2MyTrue_r = ((! lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_2MyTrue_bufchan_d[0]) || lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_2MyTrue_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_2MyTrue_bufchan_d <= {16'd0,
                                                                              1'd0};
    else
      if (lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_2MyTrue_r)
        lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_2MyTrue_bufchan_d <= lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_2MyTrue_d;
  Pointer_CTf_t lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_2MyTrue_bufchan_buf;
  assign lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_2MyTrue_bufchan_r = (! lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_2MyTrue_bufchan_buf[0]);
  assign lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_2MyTrue_1_argbuf_d = (lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_2MyTrue_bufchan_buf[0] ? lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_2MyTrue_bufchan_buf :
                                                                                 lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_2MyTrue_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_2MyTrue_bufchan_buf <= {16'd0,
                                                                                1'd0};
    else
      if ((lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_2MyTrue_1_argbuf_r && lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_2MyTrue_bufchan_buf[0]))
        lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_2MyTrue_bufchan_buf <= {16'd0,
                                                                                  1'd0};
      else if (((! lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_2MyTrue_1_argbuf_r) && (! lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_2MyTrue_bufchan_buf[0])))
        lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_2MyTrue_bufchan_buf <= lizzieLet0_4MQNode_4QVal_Bool_5QVal_Bool_3MyFalse_2MyTrue_bufchan_d;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_CTf) : (lizzieLet0_4MQNode_5,QTree_Bool) (lizzieLet0_8MQNode,Pointer_CTf) > [(lizzieLet0_4MQNode_5QNone_Bool,Pointer_CTf),
                                                                                               (lizzieLet0_4MQNode_5QVal_Bool,Pointer_CTf),
                                                                                               (lizzieLet0_4MQNode_5QNode_Bool,Pointer_CTf),
                                                                                               (lizzieLet0_4MQNode_5QError_Bool,Pointer_CTf)] */
  logic [3:0] lizzieLet0_8MQNode_onehotd;
  always_comb
    if ((lizzieLet0_4MQNode_5_d[0] && lizzieLet0_8MQNode_d[0]))
      unique case (lizzieLet0_4MQNode_5_d[2:1])
        2'd0: lizzieLet0_8MQNode_onehotd = 4'd1;
        2'd1: lizzieLet0_8MQNode_onehotd = 4'd2;
        2'd2: lizzieLet0_8MQNode_onehotd = 4'd4;
        2'd3: lizzieLet0_8MQNode_onehotd = 4'd8;
        default: lizzieLet0_8MQNode_onehotd = 4'd0;
      endcase
    else lizzieLet0_8MQNode_onehotd = 4'd0;
  assign lizzieLet0_4MQNode_5QNone_Bool_d = {lizzieLet0_8MQNode_d[16:1],
                                             lizzieLet0_8MQNode_onehotd[0]};
  assign lizzieLet0_4MQNode_5QVal_Bool_d = {lizzieLet0_8MQNode_d[16:1],
                                            lizzieLet0_8MQNode_onehotd[1]};
  assign lizzieLet0_4MQNode_5QNode_Bool_d = {lizzieLet0_8MQNode_d[16:1],
                                             lizzieLet0_8MQNode_onehotd[2]};
  assign lizzieLet0_4MQNode_5QError_Bool_d = {lizzieLet0_8MQNode_d[16:1],
                                              lizzieLet0_8MQNode_onehotd[3]};
  assign lizzieLet0_8MQNode_r = (| (lizzieLet0_8MQNode_onehotd & {lizzieLet0_4MQNode_5QError_Bool_r,
                                                                  lizzieLet0_4MQNode_5QNode_Bool_r,
                                                                  lizzieLet0_4MQNode_5QVal_Bool_r,
                                                                  lizzieLet0_4MQNode_5QNone_Bool_r}));
  assign lizzieLet0_4MQNode_5_r = lizzieLet0_8MQNode_r;
  
  /* buf (Ty Pointer_CTf) : (lizzieLet0_4MQNode_5QError_Bool,Pointer_CTf) > (lizzieLet0_4MQNode_5QError_Bool_1_argbuf,Pointer_CTf) */
  Pointer_CTf_t lizzieLet0_4MQNode_5QError_Bool_bufchan_d;
  logic lizzieLet0_4MQNode_5QError_Bool_bufchan_r;
  assign lizzieLet0_4MQNode_5QError_Bool_r = ((! lizzieLet0_4MQNode_5QError_Bool_bufchan_d[0]) || lizzieLet0_4MQNode_5QError_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_5QError_Bool_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet0_4MQNode_5QError_Bool_r)
        lizzieLet0_4MQNode_5QError_Bool_bufchan_d <= lizzieLet0_4MQNode_5QError_Bool_d;
  Pointer_CTf_t lizzieLet0_4MQNode_5QError_Bool_bufchan_buf;
  assign lizzieLet0_4MQNode_5QError_Bool_bufchan_r = (! lizzieLet0_4MQNode_5QError_Bool_bufchan_buf[0]);
  assign lizzieLet0_4MQNode_5QError_Bool_1_argbuf_d = (lizzieLet0_4MQNode_5QError_Bool_bufchan_buf[0] ? lizzieLet0_4MQNode_5QError_Bool_bufchan_buf :
                                                       lizzieLet0_4MQNode_5QError_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4MQNode_5QError_Bool_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet0_4MQNode_5QError_Bool_1_argbuf_r && lizzieLet0_4MQNode_5QError_Bool_bufchan_buf[0]))
        lizzieLet0_4MQNode_5QError_Bool_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet0_4MQNode_5QError_Bool_1_argbuf_r) && (! lizzieLet0_4MQNode_5QError_Bool_bufchan_buf[0])))
        lizzieLet0_4MQNode_5QError_Bool_bufchan_buf <= lizzieLet0_4MQNode_5QError_Bool_bufchan_d;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_MaskQTree) : (lizzieLet0_4MQNode_6,QTree_Bool) (q1a88_destruct,Pointer_MaskQTree) > [(lizzieLet0_4MQNode_6QNone_Bool,Pointer_MaskQTree),
                                                                                                       (_77,Pointer_MaskQTree),
                                                                                                       (lizzieLet0_4MQNode_6QNode_Bool,Pointer_MaskQTree),
                                                                                                       (_76,Pointer_MaskQTree)] */
  logic [3:0] q1a88_destruct_onehotd;
  always_comb
    if ((lizzieLet0_4MQNode_6_d[0] && q1a88_destruct_d[0]))
      unique case (lizzieLet0_4MQNode_6_d[2:1])
        2'd0: q1a88_destruct_onehotd = 4'd1;
        2'd1: q1a88_destruct_onehotd = 4'd2;
        2'd2: q1a88_destruct_onehotd = 4'd4;
        2'd3: q1a88_destruct_onehotd = 4'd8;
        default: q1a88_destruct_onehotd = 4'd0;
      endcase
    else q1a88_destruct_onehotd = 4'd0;
  assign lizzieLet0_4MQNode_6QNone_Bool_d = {q1a88_destruct_d[16:1],
                                             q1a88_destruct_onehotd[0]};
  assign _77_d = {q1a88_destruct_d[16:1], q1a88_destruct_onehotd[1]};
  assign lizzieLet0_4MQNode_6QNode_Bool_d = {q1a88_destruct_d[16:1],
                                             q1a88_destruct_onehotd[2]};
  assign _76_d = {q1a88_destruct_d[16:1], q1a88_destruct_onehotd[3]};
  assign q1a88_destruct_r = (| (q1a88_destruct_onehotd & {_76_r,
                                                          lizzieLet0_4MQNode_6QNode_Bool_r,
                                                          _77_r,
                                                          lizzieLet0_4MQNode_6QNone_Bool_r}));
  assign lizzieLet0_4MQNode_6_r = q1a88_destruct_r;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_MaskQTree) : (lizzieLet0_4MQNode_7,QTree_Bool) (q2a89_destruct,Pointer_MaskQTree) > [(lizzieLet0_4MQNode_7QNone_Bool,Pointer_MaskQTree),
                                                                                                       (_75,Pointer_MaskQTree),
                                                                                                       (lizzieLet0_4MQNode_7QNode_Bool,Pointer_MaskQTree),
                                                                                                       (_74,Pointer_MaskQTree)] */
  logic [3:0] q2a89_destruct_onehotd;
  always_comb
    if ((lizzieLet0_4MQNode_7_d[0] && q2a89_destruct_d[0]))
      unique case (lizzieLet0_4MQNode_7_d[2:1])
        2'd0: q2a89_destruct_onehotd = 4'd1;
        2'd1: q2a89_destruct_onehotd = 4'd2;
        2'd2: q2a89_destruct_onehotd = 4'd4;
        2'd3: q2a89_destruct_onehotd = 4'd8;
        default: q2a89_destruct_onehotd = 4'd0;
      endcase
    else q2a89_destruct_onehotd = 4'd0;
  assign lizzieLet0_4MQNode_7QNone_Bool_d = {q2a89_destruct_d[16:1],
                                             q2a89_destruct_onehotd[0]};
  assign _75_d = {q2a89_destruct_d[16:1], q2a89_destruct_onehotd[1]};
  assign lizzieLet0_4MQNode_7QNode_Bool_d = {q2a89_destruct_d[16:1],
                                             q2a89_destruct_onehotd[2]};
  assign _74_d = {q2a89_destruct_d[16:1], q2a89_destruct_onehotd[3]};
  assign q2a89_destruct_r = (| (q2a89_destruct_onehotd & {_74_r,
                                                          lizzieLet0_4MQNode_7QNode_Bool_r,
                                                          _75_r,
                                                          lizzieLet0_4MQNode_7QNone_Bool_r}));
  assign lizzieLet0_4MQNode_7_r = q2a89_destruct_r;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_MaskQTree) : (lizzieLet0_4MQNode_8,QTree_Bool) (q3a8a_destruct,Pointer_MaskQTree) > [(lizzieLet0_4MQNode_8QNone_Bool,Pointer_MaskQTree),
                                                                                                       (_73,Pointer_MaskQTree),
                                                                                                       (lizzieLet0_4MQNode_8QNode_Bool,Pointer_MaskQTree),
                                                                                                       (_72,Pointer_MaskQTree)] */
  logic [3:0] q3a8a_destruct_onehotd;
  always_comb
    if ((lizzieLet0_4MQNode_8_d[0] && q3a8a_destruct_d[0]))
      unique case (lizzieLet0_4MQNode_8_d[2:1])
        2'd0: q3a8a_destruct_onehotd = 4'd1;
        2'd1: q3a8a_destruct_onehotd = 4'd2;
        2'd2: q3a8a_destruct_onehotd = 4'd4;
        2'd3: q3a8a_destruct_onehotd = 4'd8;
        default: q3a8a_destruct_onehotd = 4'd0;
      endcase
    else q3a8a_destruct_onehotd = 4'd0;
  assign lizzieLet0_4MQNode_8QNone_Bool_d = {q3a8a_destruct_d[16:1],
                                             q3a8a_destruct_onehotd[0]};
  assign _73_d = {q3a8a_destruct_d[16:1], q3a8a_destruct_onehotd[1]};
  assign lizzieLet0_4MQNode_8QNode_Bool_d = {q3a8a_destruct_d[16:1],
                                             q3a8a_destruct_onehotd[2]};
  assign _72_d = {q3a8a_destruct_d[16:1], q3a8a_destruct_onehotd[3]};
  assign q3a8a_destruct_r = (| (q3a8a_destruct_onehotd & {_72_r,
                                                          lizzieLet0_4MQNode_8QNode_Bool_r,
                                                          _73_r,
                                                          lizzieLet0_4MQNode_8QNone_Bool_r}));
  assign lizzieLet0_4MQNode_8_r = q3a8a_destruct_r;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_MaskQTree) : (lizzieLet0_4MQNode_9,QTree_Bool) (q4a8b_destruct,Pointer_MaskQTree) > [(lizzieLet0_4MQNode_9QNone_Bool,Pointer_MaskQTree),
                                                                                                       (_71,Pointer_MaskQTree),
                                                                                                       (lizzieLet0_4MQNode_9QNode_Bool,Pointer_MaskQTree),
                                                                                                       (_70,Pointer_MaskQTree)] */
  logic [3:0] q4a8b_destruct_onehotd;
  always_comb
    if ((lizzieLet0_4MQNode_9_d[0] && q4a8b_destruct_d[0]))
      unique case (lizzieLet0_4MQNode_9_d[2:1])
        2'd0: q4a8b_destruct_onehotd = 4'd1;
        2'd1: q4a8b_destruct_onehotd = 4'd2;
        2'd2: q4a8b_destruct_onehotd = 4'd4;
        2'd3: q4a8b_destruct_onehotd = 4'd8;
        default: q4a8b_destruct_onehotd = 4'd0;
      endcase
    else q4a8b_destruct_onehotd = 4'd0;
  assign lizzieLet0_4MQNode_9QNone_Bool_d = {q4a8b_destruct_d[16:1],
                                             q4a8b_destruct_onehotd[0]};
  assign _71_d = {q4a8b_destruct_d[16:1], q4a8b_destruct_onehotd[1]};
  assign lizzieLet0_4MQNode_9QNode_Bool_d = {q4a8b_destruct_d[16:1],
                                             q4a8b_destruct_onehotd[2]};
  assign _70_d = {q4a8b_destruct_d[16:1], q4a8b_destruct_onehotd[3]};
  assign q4a8b_destruct_r = (| (q4a8b_destruct_onehotd & {_70_r,
                                                          lizzieLet0_4MQNode_9QNode_Bool_r,
                                                          _71_r,
                                                          lizzieLet0_4MQNode_9QNone_Bool_r}));
  assign lizzieLet0_4MQNode_9_r = q4a8b_destruct_r;
  
  /* demux (Ty MaskQTree,
       Ty QTree_Bool) : (lizzieLet0_5,MaskQTree) (readPointer_QTree_Boolm3a87_1_argbuf_rwb,QTree_Bool) > [(_69,QTree_Bool),
                                                                                                          (_68,QTree_Bool),
                                                                                                          (lizzieLet0_5MQNode,QTree_Bool)] */
  logic [2:0] readPointer_QTree_Boolm3a87_1_argbuf_rwb_onehotd;
  always_comb
    if ((lizzieLet0_5_d[0] && readPointer_QTree_Boolm3a87_1_argbuf_rwb_d[0]))
      unique case (lizzieLet0_5_d[2:1])
        2'd0: readPointer_QTree_Boolm3a87_1_argbuf_rwb_onehotd = 3'd1;
        2'd1: readPointer_QTree_Boolm3a87_1_argbuf_rwb_onehotd = 3'd2;
        2'd2: readPointer_QTree_Boolm3a87_1_argbuf_rwb_onehotd = 3'd4;
        default: readPointer_QTree_Boolm3a87_1_argbuf_rwb_onehotd = 3'd0;
      endcase
    else readPointer_QTree_Boolm3a87_1_argbuf_rwb_onehotd = 3'd0;
  assign _69_d = {readPointer_QTree_Boolm3a87_1_argbuf_rwb_d[66:1],
                  readPointer_QTree_Boolm3a87_1_argbuf_rwb_onehotd[0]};
  assign _68_d = {readPointer_QTree_Boolm3a87_1_argbuf_rwb_d[66:1],
                  readPointer_QTree_Boolm3a87_1_argbuf_rwb_onehotd[1]};
  assign lizzieLet0_5MQNode_d = {readPointer_QTree_Boolm3a87_1_argbuf_rwb_d[66:1],
                                 readPointer_QTree_Boolm3a87_1_argbuf_rwb_onehotd[2]};
  assign readPointer_QTree_Boolm3a87_1_argbuf_rwb_r = (| (readPointer_QTree_Boolm3a87_1_argbuf_rwb_onehotd & {lizzieLet0_5MQNode_r,
                                                                                                              _68_r,
                                                                                                              _69_r}));
  assign lizzieLet0_5_r = readPointer_QTree_Boolm3a87_1_argbuf_rwb_r;
  
  /* demux (Ty MaskQTree,
       Ty Pointer_QTree_Bool) : (lizzieLet0_6,MaskQTree) (m2a86_2,Pointer_QTree_Bool) > [(_67,Pointer_QTree_Bool),
                                                                                         (lizzieLet0_6MQVal,Pointer_QTree_Bool),
                                                                                         (_66,Pointer_QTree_Bool)] */
  logic [2:0] m2a86_2_onehotd;
  always_comb
    if ((lizzieLet0_6_d[0] && m2a86_2_d[0]))
      unique case (lizzieLet0_6_d[2:1])
        2'd0: m2a86_2_onehotd = 3'd1;
        2'd1: m2a86_2_onehotd = 3'd2;
        2'd2: m2a86_2_onehotd = 3'd4;
        default: m2a86_2_onehotd = 3'd0;
      endcase
    else m2a86_2_onehotd = 3'd0;
  assign _67_d = {m2a86_2_d[16:1], m2a86_2_onehotd[0]};
  assign lizzieLet0_6MQVal_d = {m2a86_2_d[16:1], m2a86_2_onehotd[1]};
  assign _66_d = {m2a86_2_d[16:1], m2a86_2_onehotd[2]};
  assign m2a86_2_r = (| (m2a86_2_onehotd & {_66_r,
                                            lizzieLet0_6MQVal_r,
                                            _67_r}));
  assign lizzieLet0_6_r = m2a86_2_r;
  
  /* buf (Ty Pointer_QTree_Bool) : (lizzieLet0_6MQVal,Pointer_QTree_Bool) > (lizzieLet0_6MQVal_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t lizzieLet0_6MQVal_bufchan_d;
  logic lizzieLet0_6MQVal_bufchan_r;
  assign lizzieLet0_6MQVal_r = ((! lizzieLet0_6MQVal_bufchan_d[0]) || lizzieLet0_6MQVal_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet0_6MQVal_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet0_6MQVal_r)
        lizzieLet0_6MQVal_bufchan_d <= lizzieLet0_6MQVal_d;
  Pointer_QTree_Bool_t lizzieLet0_6MQVal_bufchan_buf;
  assign lizzieLet0_6MQVal_bufchan_r = (! lizzieLet0_6MQVal_bufchan_buf[0]);
  assign lizzieLet0_6MQVal_1_argbuf_d = (lizzieLet0_6MQVal_bufchan_buf[0] ? lizzieLet0_6MQVal_bufchan_buf :
                                         lizzieLet0_6MQVal_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_6MQVal_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet0_6MQVal_1_argbuf_r && lizzieLet0_6MQVal_bufchan_buf[0]))
        lizzieLet0_6MQVal_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet0_6MQVal_1_argbuf_r) && (! lizzieLet0_6MQVal_bufchan_buf[0])))
        lizzieLet0_6MQVal_bufchan_buf <= lizzieLet0_6MQVal_bufchan_d;
  
  /* demux (Ty MaskQTree,
       Ty Pointer_QTree_Bool) : (lizzieLet0_7,MaskQTree) (m3a87_2,Pointer_QTree_Bool) > [(_65,Pointer_QTree_Bool),
                                                                                         (lizzieLet0_7MQVal,Pointer_QTree_Bool),
                                                                                         (_64,Pointer_QTree_Bool)] */
  logic [2:0] m3a87_2_onehotd;
  always_comb
    if ((lizzieLet0_7_d[0] && m3a87_2_d[0]))
      unique case (lizzieLet0_7_d[2:1])
        2'd0: m3a87_2_onehotd = 3'd1;
        2'd1: m3a87_2_onehotd = 3'd2;
        2'd2: m3a87_2_onehotd = 3'd4;
        default: m3a87_2_onehotd = 3'd0;
      endcase
    else m3a87_2_onehotd = 3'd0;
  assign _65_d = {m3a87_2_d[16:1], m3a87_2_onehotd[0]};
  assign lizzieLet0_7MQVal_d = {m3a87_2_d[16:1], m3a87_2_onehotd[1]};
  assign _64_d = {m3a87_2_d[16:1], m3a87_2_onehotd[2]};
  assign m3a87_2_r = (| (m3a87_2_onehotd & {_64_r,
                                            lizzieLet0_7MQVal_r,
                                            _65_r}));
  assign lizzieLet0_7_r = m3a87_2_r;
  
  /* buf (Ty Pointer_QTree_Bool) : (lizzieLet0_7MQVal,Pointer_QTree_Bool) > (lizzieLet0_7MQVal_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t lizzieLet0_7MQVal_bufchan_d;
  logic lizzieLet0_7MQVal_bufchan_r;
  assign lizzieLet0_7MQVal_r = ((! lizzieLet0_7MQVal_bufchan_d[0]) || lizzieLet0_7MQVal_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet0_7MQVal_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet0_7MQVal_r)
        lizzieLet0_7MQVal_bufchan_d <= lizzieLet0_7MQVal_d;
  Pointer_QTree_Bool_t lizzieLet0_7MQVal_bufchan_buf;
  assign lizzieLet0_7MQVal_bufchan_r = (! lizzieLet0_7MQVal_bufchan_buf[0]);
  assign lizzieLet0_7MQVal_1_argbuf_d = (lizzieLet0_7MQVal_bufchan_buf[0] ? lizzieLet0_7MQVal_bufchan_buf :
                                         lizzieLet0_7MQVal_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_7MQVal_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet0_7MQVal_1_argbuf_r && lizzieLet0_7MQVal_bufchan_buf[0]))
        lizzieLet0_7MQVal_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet0_7MQVal_1_argbuf_r) && (! lizzieLet0_7MQVal_bufchan_buf[0])))
        lizzieLet0_7MQVal_bufchan_buf <= lizzieLet0_7MQVal_bufchan_d;
  
  /* demux (Ty MaskQTree,
       Ty Pointer_CTf) : (lizzieLet0_8,MaskQTree) (sc_0_goMux_mux,Pointer_CTf) > [(lizzieLet0_8MQNone,Pointer_CTf),
                                                                                  (lizzieLet0_8MQVal,Pointer_CTf),
                                                                                  (lizzieLet0_8MQNode,Pointer_CTf)] */
  logic [2:0] sc_0_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet0_8_d[0] && sc_0_goMux_mux_d[0]))
      unique case (lizzieLet0_8_d[2:1])
        2'd0: sc_0_goMux_mux_onehotd = 3'd1;
        2'd1: sc_0_goMux_mux_onehotd = 3'd2;
        2'd2: sc_0_goMux_mux_onehotd = 3'd4;
        default: sc_0_goMux_mux_onehotd = 3'd0;
      endcase
    else sc_0_goMux_mux_onehotd = 3'd0;
  assign lizzieLet0_8MQNone_d = {sc_0_goMux_mux_d[16:1],
                                 sc_0_goMux_mux_onehotd[0]};
  assign lizzieLet0_8MQVal_d = {sc_0_goMux_mux_d[16:1],
                                sc_0_goMux_mux_onehotd[1]};
  assign lizzieLet0_8MQNode_d = {sc_0_goMux_mux_d[16:1],
                                 sc_0_goMux_mux_onehotd[2]};
  assign sc_0_goMux_mux_r = (| (sc_0_goMux_mux_onehotd & {lizzieLet0_8MQNode_r,
                                                          lizzieLet0_8MQVal_r,
                                                          lizzieLet0_8MQNone_r}));
  assign lizzieLet0_8_r = sc_0_goMux_mux_r;
  
  /* buf (Ty Pointer_CTf) : (lizzieLet0_8MQNone,Pointer_CTf) > (lizzieLet0_8MQNone_1_argbuf,Pointer_CTf) */
  Pointer_CTf_t lizzieLet0_8MQNone_bufchan_d;
  logic lizzieLet0_8MQNone_bufchan_r;
  assign lizzieLet0_8MQNone_r = ((! lizzieLet0_8MQNone_bufchan_d[0]) || lizzieLet0_8MQNone_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet0_8MQNone_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet0_8MQNone_r)
        lizzieLet0_8MQNone_bufchan_d <= lizzieLet0_8MQNone_d;
  Pointer_CTf_t lizzieLet0_8MQNone_bufchan_buf;
  assign lizzieLet0_8MQNone_bufchan_r = (! lizzieLet0_8MQNone_bufchan_buf[0]);
  assign lizzieLet0_8MQNone_1_argbuf_d = (lizzieLet0_8MQNone_bufchan_buf[0] ? lizzieLet0_8MQNone_bufchan_buf :
                                          lizzieLet0_8MQNone_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_8MQNone_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet0_8MQNone_1_argbuf_r && lizzieLet0_8MQNone_bufchan_buf[0]))
        lizzieLet0_8MQNone_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet0_8MQNone_1_argbuf_r) && (! lizzieLet0_8MQNone_bufchan_buf[0])))
        lizzieLet0_8MQNone_bufchan_buf <= lizzieLet0_8MQNone_bufchan_d;
  
  /* buf (Ty Pointer_CTf) : (lizzieLet0_8MQVal,Pointer_CTf) > (lizzieLet0_8MQVal_1_argbuf,Pointer_CTf) */
  Pointer_CTf_t lizzieLet0_8MQVal_bufchan_d;
  logic lizzieLet0_8MQVal_bufchan_r;
  assign lizzieLet0_8MQVal_r = ((! lizzieLet0_8MQVal_bufchan_d[0]) || lizzieLet0_8MQVal_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet0_8MQVal_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet0_8MQVal_r)
        lizzieLet0_8MQVal_bufchan_d <= lizzieLet0_8MQVal_d;
  Pointer_CTf_t lizzieLet0_8MQVal_bufchan_buf;
  assign lizzieLet0_8MQVal_bufchan_r = (! lizzieLet0_8MQVal_bufchan_buf[0]);
  assign lizzieLet0_8MQVal_1_argbuf_d = (lizzieLet0_8MQVal_bufchan_buf[0] ? lizzieLet0_8MQVal_bufchan_buf :
                                         lizzieLet0_8MQVal_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_8MQVal_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet0_8MQVal_1_argbuf_r && lizzieLet0_8MQVal_bufchan_buf[0]))
        lizzieLet0_8MQVal_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet0_8MQVal_1_argbuf_r) && (! lizzieLet0_8MQVal_bufchan_buf[0])))
        lizzieLet0_8MQVal_bufchan_buf <= lizzieLet0_8MQVal_bufchan_d;
  
  /* destruct (Ty QTree_Bool,
          Dcon QNode_Bool) : (lizzieLet20_1_1QNode_Bool,QTree_Bool) > [(q1a8P_destruct,Pointer_QTree_Bool),
                                                                       (q2a8Q_destruct,Pointer_QTree_Bool),
                                                                       (q3a8R_destruct,Pointer_QTree_Bool),
                                                                       (q4a8S_destruct,Pointer_QTree_Bool)] */
  logic [3:0] lizzieLet20_1_1QNode_Bool_emitted;
  logic [3:0] lizzieLet20_1_1QNode_Bool_done;
  assign q1a8P_destruct_d = {lizzieLet20_1_1QNode_Bool_d[18:3],
                             (lizzieLet20_1_1QNode_Bool_d[0] && (! lizzieLet20_1_1QNode_Bool_emitted[0]))};
  assign q2a8Q_destruct_d = {lizzieLet20_1_1QNode_Bool_d[34:19],
                             (lizzieLet20_1_1QNode_Bool_d[0] && (! lizzieLet20_1_1QNode_Bool_emitted[1]))};
  assign q3a8R_destruct_d = {lizzieLet20_1_1QNode_Bool_d[50:35],
                             (lizzieLet20_1_1QNode_Bool_d[0] && (! lizzieLet20_1_1QNode_Bool_emitted[2]))};
  assign q4a8S_destruct_d = {lizzieLet20_1_1QNode_Bool_d[66:51],
                             (lizzieLet20_1_1QNode_Bool_d[0] && (! lizzieLet20_1_1QNode_Bool_emitted[3]))};
  assign lizzieLet20_1_1QNode_Bool_done = (lizzieLet20_1_1QNode_Bool_emitted | ({q4a8S_destruct_d[0],
                                                                                 q3a8R_destruct_d[0],
                                                                                 q2a8Q_destruct_d[0],
                                                                                 q1a8P_destruct_d[0]} & {q4a8S_destruct_r,
                                                                                                         q3a8R_destruct_r,
                                                                                                         q2a8Q_destruct_r,
                                                                                                         q1a8P_destruct_r}));
  assign lizzieLet20_1_1QNode_Bool_r = (& lizzieLet20_1_1QNode_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet20_1_1QNode_Bool_emitted <= 4'd0;
    else
      lizzieLet20_1_1QNode_Bool_emitted <= (lizzieLet20_1_1QNode_Bool_r ? 4'd0 :
                                            lizzieLet20_1_1QNode_Bool_done);
  
  /* destruct (Ty QTree_Bool,
          Dcon QVal_Bool) : (lizzieLet20_1_1QVal_Bool,QTree_Bool) > [(v1a8J_destruct,MyBool)] */
  assign v1a8J_destruct_d = {lizzieLet20_1_1QVal_Bool_d[3:3],
                             lizzieLet20_1_1QVal_Bool_d[0]};
  assign lizzieLet20_1_1QVal_Bool_r = v1a8J_destruct_r;
  
  /* demux (Ty QTree_Bool,
       Ty QTree_Bool) : (lizzieLet20_1_2,QTree_Bool) (lizzieLet20_1_1,QTree_Bool) > [(_63,QTree_Bool),
                                                                                     (lizzieLet20_1_1QVal_Bool,QTree_Bool),
                                                                                     (lizzieLet20_1_1QNode_Bool,QTree_Bool),
                                                                                     (_62,QTree_Bool)] */
  logic [3:0] lizzieLet20_1_1_onehotd;
  always_comb
    if ((lizzieLet20_1_2_d[0] && lizzieLet20_1_1_d[0]))
      unique case (lizzieLet20_1_2_d[2:1])
        2'd0: lizzieLet20_1_1_onehotd = 4'd1;
        2'd1: lizzieLet20_1_1_onehotd = 4'd2;
        2'd2: lizzieLet20_1_1_onehotd = 4'd4;
        2'd3: lizzieLet20_1_1_onehotd = 4'd8;
        default: lizzieLet20_1_1_onehotd = 4'd0;
      endcase
    else lizzieLet20_1_1_onehotd = 4'd0;
  assign _63_d = {lizzieLet20_1_1_d[66:1],
                  lizzieLet20_1_1_onehotd[0]};
  assign lizzieLet20_1_1QVal_Bool_d = {lizzieLet20_1_1_d[66:1],
                                       lizzieLet20_1_1_onehotd[1]};
  assign lizzieLet20_1_1QNode_Bool_d = {lizzieLet20_1_1_d[66:1],
                                        lizzieLet20_1_1_onehotd[2]};
  assign _62_d = {lizzieLet20_1_1_d[66:1],
                  lizzieLet20_1_1_onehotd[3]};
  assign lizzieLet20_1_1_r = (| (lizzieLet20_1_1_onehotd & {_62_r,
                                                            lizzieLet20_1_1QNode_Bool_r,
                                                            lizzieLet20_1_1QVal_Bool_r,
                                                            _63_r}));
  assign lizzieLet20_1_2_r = lizzieLet20_1_1_r;
  
  /* demux (Ty QTree_Bool,
       Ty Go) : (lizzieLet20_1_3,QTree_Bool) (go_3_goMux_data,Go) > [(lizzieLet20_1_3QNone_Bool,Go),
                                                                     (lizzieLet20_1_3QVal_Bool,Go),
                                                                     (lizzieLet20_1_3QNode_Bool,Go),
                                                                     (lizzieLet20_1_3QError_Bool,Go)] */
  logic [3:0] go_3_goMux_data_onehotd;
  always_comb
    if ((lizzieLet20_1_3_d[0] && go_3_goMux_data_d[0]))
      unique case (lizzieLet20_1_3_d[2:1])
        2'd0: go_3_goMux_data_onehotd = 4'd1;
        2'd1: go_3_goMux_data_onehotd = 4'd2;
        2'd2: go_3_goMux_data_onehotd = 4'd4;
        2'd3: go_3_goMux_data_onehotd = 4'd8;
        default: go_3_goMux_data_onehotd = 4'd0;
      endcase
    else go_3_goMux_data_onehotd = 4'd0;
  assign lizzieLet20_1_3QNone_Bool_d = go_3_goMux_data_onehotd[0];
  assign lizzieLet20_1_3QVal_Bool_d = go_3_goMux_data_onehotd[1];
  assign lizzieLet20_1_3QNode_Bool_d = go_3_goMux_data_onehotd[2];
  assign lizzieLet20_1_3QError_Bool_d = go_3_goMux_data_onehotd[3];
  assign go_3_goMux_data_r = (| (go_3_goMux_data_onehotd & {lizzieLet20_1_3QError_Bool_r,
                                                            lizzieLet20_1_3QNode_Bool_r,
                                                            lizzieLet20_1_3QVal_Bool_r,
                                                            lizzieLet20_1_3QNone_Bool_r}));
  assign lizzieLet20_1_3_r = go_3_goMux_data_r;
  
  /* fork (Ty Go) : (lizzieLet20_1_3QError_Bool,Go) > [(lizzieLet20_1_3QError_Bool_1,Go),
                                                  (lizzieLet20_1_3QError_Bool_2,Go)] */
  logic [1:0] lizzieLet20_1_3QError_Bool_emitted;
  logic [1:0] lizzieLet20_1_3QError_Bool_done;
  assign lizzieLet20_1_3QError_Bool_1_d = (lizzieLet20_1_3QError_Bool_d[0] && (! lizzieLet20_1_3QError_Bool_emitted[0]));
  assign lizzieLet20_1_3QError_Bool_2_d = (lizzieLet20_1_3QError_Bool_d[0] && (! lizzieLet20_1_3QError_Bool_emitted[1]));
  assign lizzieLet20_1_3QError_Bool_done = (lizzieLet20_1_3QError_Bool_emitted | ({lizzieLet20_1_3QError_Bool_2_d[0],
                                                                                   lizzieLet20_1_3QError_Bool_1_d[0]} & {lizzieLet20_1_3QError_Bool_2_r,
                                                                                                                         lizzieLet20_1_3QError_Bool_1_r}));
  assign lizzieLet20_1_3QError_Bool_r = (& lizzieLet20_1_3QError_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet20_1_3QError_Bool_emitted <= 2'd0;
    else
      lizzieLet20_1_3QError_Bool_emitted <= (lizzieLet20_1_3QError_Bool_r ? 2'd0 :
                                             lizzieLet20_1_3QError_Bool_done);
  
  /* dcon (Ty QTree_Bool,
      Dcon QError_Bool) : [(lizzieLet20_1_3QError_Bool_1,Go)] > (lizzieLet20_1_3QError_Bool_1QError_Bool,QTree_Bool) */
  assign lizzieLet20_1_3QError_Bool_1QError_Bool_d = QError_Bool_dc((& {lizzieLet20_1_3QError_Bool_1_d[0]}), lizzieLet20_1_3QError_Bool_1_d);
  assign {lizzieLet20_1_3QError_Bool_1_r} = {1 {(lizzieLet20_1_3QError_Bool_1QError_Bool_r && lizzieLet20_1_3QError_Bool_1QError_Bool_d[0])}};
  
  /* buf (Ty QTree_Bool) : (lizzieLet20_1_3QError_Bool_1QError_Bool,QTree_Bool) > (lizzieLet31_1_argbuf,QTree_Bool) */
  QTree_Bool_t lizzieLet20_1_3QError_Bool_1QError_Bool_bufchan_d;
  logic lizzieLet20_1_3QError_Bool_1QError_Bool_bufchan_r;
  assign lizzieLet20_1_3QError_Bool_1QError_Bool_r = ((! lizzieLet20_1_3QError_Bool_1QError_Bool_bufchan_d[0]) || lizzieLet20_1_3QError_Bool_1QError_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet20_1_3QError_Bool_1QError_Bool_bufchan_d <= {66'd0, 1'd0};
    else
      if (lizzieLet20_1_3QError_Bool_1QError_Bool_r)
        lizzieLet20_1_3QError_Bool_1QError_Bool_bufchan_d <= lizzieLet20_1_3QError_Bool_1QError_Bool_d;
  QTree_Bool_t lizzieLet20_1_3QError_Bool_1QError_Bool_bufchan_buf;
  assign lizzieLet20_1_3QError_Bool_1QError_Bool_bufchan_r = (! lizzieLet20_1_3QError_Bool_1QError_Bool_bufchan_buf[0]);
  assign lizzieLet31_1_argbuf_d = (lizzieLet20_1_3QError_Bool_1QError_Bool_bufchan_buf[0] ? lizzieLet20_1_3QError_Bool_1QError_Bool_bufchan_buf :
                                   lizzieLet20_1_3QError_Bool_1QError_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet20_1_3QError_Bool_1QError_Bool_bufchan_buf <= {66'd0,
                                                              1'd0};
    else
      if ((lizzieLet31_1_argbuf_r && lizzieLet20_1_3QError_Bool_1QError_Bool_bufchan_buf[0]))
        lizzieLet20_1_3QError_Bool_1QError_Bool_bufchan_buf <= {66'd0,
                                                                1'd0};
      else if (((! lizzieLet31_1_argbuf_r) && (! lizzieLet20_1_3QError_Bool_1QError_Bool_bufchan_buf[0])))
        lizzieLet20_1_3QError_Bool_1QError_Bool_bufchan_buf <= lizzieLet20_1_3QError_Bool_1QError_Bool_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet20_1_3QError_Bool_2,Go) > (lizzieLet20_1_3QError_Bool_2_argbuf,Go) */
  Go_t lizzieLet20_1_3QError_Bool_2_bufchan_d;
  logic lizzieLet20_1_3QError_Bool_2_bufchan_r;
  assign lizzieLet20_1_3QError_Bool_2_r = ((! lizzieLet20_1_3QError_Bool_2_bufchan_d[0]) || lizzieLet20_1_3QError_Bool_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet20_1_3QError_Bool_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet20_1_3QError_Bool_2_r)
        lizzieLet20_1_3QError_Bool_2_bufchan_d <= lizzieLet20_1_3QError_Bool_2_d;
  Go_t lizzieLet20_1_3QError_Bool_2_bufchan_buf;
  assign lizzieLet20_1_3QError_Bool_2_bufchan_r = (! lizzieLet20_1_3QError_Bool_2_bufchan_buf[0]);
  assign lizzieLet20_1_3QError_Bool_2_argbuf_d = (lizzieLet20_1_3QError_Bool_2_bufchan_buf[0] ? lizzieLet20_1_3QError_Bool_2_bufchan_buf :
                                                  lizzieLet20_1_3QError_Bool_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet20_1_3QError_Bool_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet20_1_3QError_Bool_2_argbuf_r && lizzieLet20_1_3QError_Bool_2_bufchan_buf[0]))
        lizzieLet20_1_3QError_Bool_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet20_1_3QError_Bool_2_argbuf_r) && (! lizzieLet20_1_3QError_Bool_2_bufchan_buf[0])))
        lizzieLet20_1_3QError_Bool_2_bufchan_buf <= lizzieLet20_1_3QError_Bool_2_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet20_1_3QNone_Bool,Go) > (lizzieLet20_1_3QNone_Bool_1_argbuf,Go) */
  Go_t lizzieLet20_1_3QNone_Bool_bufchan_d;
  logic lizzieLet20_1_3QNone_Bool_bufchan_r;
  assign lizzieLet20_1_3QNone_Bool_r = ((! lizzieLet20_1_3QNone_Bool_bufchan_d[0]) || lizzieLet20_1_3QNone_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet20_1_3QNone_Bool_bufchan_d <= 1'd0;
    else
      if (lizzieLet20_1_3QNone_Bool_r)
        lizzieLet20_1_3QNone_Bool_bufchan_d <= lizzieLet20_1_3QNone_Bool_d;
  Go_t lizzieLet20_1_3QNone_Bool_bufchan_buf;
  assign lizzieLet20_1_3QNone_Bool_bufchan_r = (! lizzieLet20_1_3QNone_Bool_bufchan_buf[0]);
  assign lizzieLet20_1_3QNone_Bool_1_argbuf_d = (lizzieLet20_1_3QNone_Bool_bufchan_buf[0] ? lizzieLet20_1_3QNone_Bool_bufchan_buf :
                                                 lizzieLet20_1_3QNone_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet20_1_3QNone_Bool_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet20_1_3QNone_Bool_1_argbuf_r && lizzieLet20_1_3QNone_Bool_bufchan_buf[0]))
        lizzieLet20_1_3QNone_Bool_bufchan_buf <= 1'd0;
      else if (((! lizzieLet20_1_3QNone_Bool_1_argbuf_r) && (! lizzieLet20_1_3QNone_Bool_bufchan_buf[0])))
        lizzieLet20_1_3QNone_Bool_bufchan_buf <= lizzieLet20_1_3QNone_Bool_bufchan_d;
  
  /* mergectrl (Ty C12,
           Ty Go) : [(lizzieLet20_1_3QNone_Bool_1_argbuf,Go),
                     (lizzieLet48_3Lcall_f'0_1_argbuf,Go),
                     (lizzieLet20_1_4QVal_Bool_3QNone_Bool_1_argbuf,Go),
                     (lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_argbuf,Go),
                     (lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_argbuf,Go),
                     (lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyTrue_2_argbuf,Go),
                     (lizzieLet20_1_4QVal_Bool_3QNode_Bool_2_argbuf,Go),
                     (lizzieLet20_1_4QVal_Bool_3QError_Bool_2_argbuf,Go),
                     (lizzieLet20_1_4QNode_Bool_3QNone_Bool_1_argbuf,Go),
                     (lizzieLet20_1_4QNode_Bool_3QVal_Bool_2_argbuf,Go),
                     (lizzieLet20_1_4QNode_Bool_3QError_Bool_2_argbuf,Go),
                     (lizzieLet20_1_3QError_Bool_2_argbuf,Go)] > (go_10_goMux_choice,C12) (go_10_goMux_data,Go) */
  logic [11:0] lizzieLet20_1_3QNone_Bool_1_argbuf_select_d;
  assign lizzieLet20_1_3QNone_Bool_1_argbuf_select_d = ((| lizzieLet20_1_3QNone_Bool_1_argbuf_select_q) ? lizzieLet20_1_3QNone_Bool_1_argbuf_select_q :
                                                        (lizzieLet20_1_3QNone_Bool_1_argbuf_d[0] ? 12'd1 :
                                                         (\lizzieLet48_3Lcall_f'0_1_argbuf_d [0] ? 12'd2 :
                                                          (lizzieLet20_1_4QVal_Bool_3QNone_Bool_1_argbuf_d[0] ? 12'd4 :
                                                           (lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_argbuf_d[0] ? 12'd8 :
                                                            (lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_argbuf_d[0] ? 12'd16 :
                                                             (lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyTrue_2_argbuf_d[0] ? 12'd32 :
                                                              (lizzieLet20_1_4QVal_Bool_3QNode_Bool_2_argbuf_d[0] ? 12'd64 :
                                                               (lizzieLet20_1_4QVal_Bool_3QError_Bool_2_argbuf_d[0] ? 12'd128 :
                                                                (lizzieLet20_1_4QNode_Bool_3QNone_Bool_1_argbuf_d[0] ? 12'd256 :
                                                                 (lizzieLet20_1_4QNode_Bool_3QVal_Bool_2_argbuf_d[0] ? 12'd512 :
                                                                  (lizzieLet20_1_4QNode_Bool_3QError_Bool_2_argbuf_d[0] ? 12'd1024 :
                                                                   (lizzieLet20_1_3QError_Bool_2_argbuf_d[0] ? 12'd2048 :
                                                                    12'd0)))))))))))));
  logic [11:0] lizzieLet20_1_3QNone_Bool_1_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet20_1_3QNone_Bool_1_argbuf_select_q <= 12'd0;
    else
      lizzieLet20_1_3QNone_Bool_1_argbuf_select_q <= (lizzieLet20_1_3QNone_Bool_1_argbuf_done ? 12'd0 :
                                                      lizzieLet20_1_3QNone_Bool_1_argbuf_select_d);
  logic [1:0] lizzieLet20_1_3QNone_Bool_1_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet20_1_3QNone_Bool_1_argbuf_emit_q <= 2'd0;
    else
      lizzieLet20_1_3QNone_Bool_1_argbuf_emit_q <= (lizzieLet20_1_3QNone_Bool_1_argbuf_done ? 2'd0 :
                                                    lizzieLet20_1_3QNone_Bool_1_argbuf_emit_d);
  logic [1:0] lizzieLet20_1_3QNone_Bool_1_argbuf_emit_d;
  assign lizzieLet20_1_3QNone_Bool_1_argbuf_emit_d = (lizzieLet20_1_3QNone_Bool_1_argbuf_emit_q | ({go_10_goMux_choice_d[0],
                                                                                                    go_10_goMux_data_d[0]} & {go_10_goMux_choice_r,
                                                                                                                              go_10_goMux_data_r}));
  logic lizzieLet20_1_3QNone_Bool_1_argbuf_done;
  assign lizzieLet20_1_3QNone_Bool_1_argbuf_done = (& lizzieLet20_1_3QNone_Bool_1_argbuf_emit_d);
  assign {lizzieLet20_1_3QError_Bool_2_argbuf_r,
          lizzieLet20_1_4QNode_Bool_3QError_Bool_2_argbuf_r,
          lizzieLet20_1_4QNode_Bool_3QVal_Bool_2_argbuf_r,
          lizzieLet20_1_4QNode_Bool_3QNone_Bool_1_argbuf_r,
          lizzieLet20_1_4QVal_Bool_3QError_Bool_2_argbuf_r,
          lizzieLet20_1_4QVal_Bool_3QNode_Bool_2_argbuf_r,
          lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyTrue_2_argbuf_r,
          lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_argbuf_r,
          lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_argbuf_r,
          lizzieLet20_1_4QVal_Bool_3QNone_Bool_1_argbuf_r,
          \lizzieLet48_3Lcall_f'0_1_argbuf_r ,
          lizzieLet20_1_3QNone_Bool_1_argbuf_r} = (lizzieLet20_1_3QNone_Bool_1_argbuf_done ? lizzieLet20_1_3QNone_Bool_1_argbuf_select_d :
                                                   12'd0);
  assign go_10_goMux_data_d = ((lizzieLet20_1_3QNone_Bool_1_argbuf_select_d[0] && (! lizzieLet20_1_3QNone_Bool_1_argbuf_emit_q[0])) ? lizzieLet20_1_3QNone_Bool_1_argbuf_d :
                               ((lizzieLet20_1_3QNone_Bool_1_argbuf_select_d[1] && (! lizzieLet20_1_3QNone_Bool_1_argbuf_emit_q[0])) ? \lizzieLet48_3Lcall_f'0_1_argbuf_d  :
                                ((lizzieLet20_1_3QNone_Bool_1_argbuf_select_d[2] && (! lizzieLet20_1_3QNone_Bool_1_argbuf_emit_q[0])) ? lizzieLet20_1_4QVal_Bool_3QNone_Bool_1_argbuf_d :
                                 ((lizzieLet20_1_3QNone_Bool_1_argbuf_select_d[3] && (! lizzieLet20_1_3QNone_Bool_1_argbuf_emit_q[0])) ? lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_argbuf_d :
                                  ((lizzieLet20_1_3QNone_Bool_1_argbuf_select_d[4] && (! lizzieLet20_1_3QNone_Bool_1_argbuf_emit_q[0])) ? lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_argbuf_d :
                                   ((lizzieLet20_1_3QNone_Bool_1_argbuf_select_d[5] && (! lizzieLet20_1_3QNone_Bool_1_argbuf_emit_q[0])) ? lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyTrue_2_argbuf_d :
                                    ((lizzieLet20_1_3QNone_Bool_1_argbuf_select_d[6] && (! lizzieLet20_1_3QNone_Bool_1_argbuf_emit_q[0])) ? lizzieLet20_1_4QVal_Bool_3QNode_Bool_2_argbuf_d :
                                     ((lizzieLet20_1_3QNone_Bool_1_argbuf_select_d[7] && (! lizzieLet20_1_3QNone_Bool_1_argbuf_emit_q[0])) ? lizzieLet20_1_4QVal_Bool_3QError_Bool_2_argbuf_d :
                                      ((lizzieLet20_1_3QNone_Bool_1_argbuf_select_d[8] && (! lizzieLet20_1_3QNone_Bool_1_argbuf_emit_q[0])) ? lizzieLet20_1_4QNode_Bool_3QNone_Bool_1_argbuf_d :
                                       ((lizzieLet20_1_3QNone_Bool_1_argbuf_select_d[9] && (! lizzieLet20_1_3QNone_Bool_1_argbuf_emit_q[0])) ? lizzieLet20_1_4QNode_Bool_3QVal_Bool_2_argbuf_d :
                                        ((lizzieLet20_1_3QNone_Bool_1_argbuf_select_d[10] && (! lizzieLet20_1_3QNone_Bool_1_argbuf_emit_q[0])) ? lizzieLet20_1_4QNode_Bool_3QError_Bool_2_argbuf_d :
                                         ((lizzieLet20_1_3QNone_Bool_1_argbuf_select_d[11] && (! lizzieLet20_1_3QNone_Bool_1_argbuf_emit_q[0])) ? lizzieLet20_1_3QError_Bool_2_argbuf_d :
                                          1'd0))))))))))));
  assign go_10_goMux_choice_d = ((lizzieLet20_1_3QNone_Bool_1_argbuf_select_d[0] && (! lizzieLet20_1_3QNone_Bool_1_argbuf_emit_q[1])) ? C1_12_dc(1'd1) :
                                 ((lizzieLet20_1_3QNone_Bool_1_argbuf_select_d[1] && (! lizzieLet20_1_3QNone_Bool_1_argbuf_emit_q[1])) ? C2_12_dc(1'd1) :
                                  ((lizzieLet20_1_3QNone_Bool_1_argbuf_select_d[2] && (! lizzieLet20_1_3QNone_Bool_1_argbuf_emit_q[1])) ? C3_12_dc(1'd1) :
                                   ((lizzieLet20_1_3QNone_Bool_1_argbuf_select_d[3] && (! lizzieLet20_1_3QNone_Bool_1_argbuf_emit_q[1])) ? C4_12_dc(1'd1) :
                                    ((lizzieLet20_1_3QNone_Bool_1_argbuf_select_d[4] && (! lizzieLet20_1_3QNone_Bool_1_argbuf_emit_q[1])) ? C5_12_dc(1'd1) :
                                     ((lizzieLet20_1_3QNone_Bool_1_argbuf_select_d[5] && (! lizzieLet20_1_3QNone_Bool_1_argbuf_emit_q[1])) ? C6_12_dc(1'd1) :
                                      ((lizzieLet20_1_3QNone_Bool_1_argbuf_select_d[6] && (! lizzieLet20_1_3QNone_Bool_1_argbuf_emit_q[1])) ? C7_12_dc(1'd1) :
                                       ((lizzieLet20_1_3QNone_Bool_1_argbuf_select_d[7] && (! lizzieLet20_1_3QNone_Bool_1_argbuf_emit_q[1])) ? C8_12_dc(1'd1) :
                                        ((lizzieLet20_1_3QNone_Bool_1_argbuf_select_d[8] && (! lizzieLet20_1_3QNone_Bool_1_argbuf_emit_q[1])) ? C9_12_dc(1'd1) :
                                         ((lizzieLet20_1_3QNone_Bool_1_argbuf_select_d[9] && (! lizzieLet20_1_3QNone_Bool_1_argbuf_emit_q[1])) ? C10_12_dc(1'd1) :
                                          ((lizzieLet20_1_3QNone_Bool_1_argbuf_select_d[10] && (! lizzieLet20_1_3QNone_Bool_1_argbuf_emit_q[1])) ? C11_12_dc(1'd1) :
                                           ((lizzieLet20_1_3QNone_Bool_1_argbuf_select_d[11] && (! lizzieLet20_1_3QNone_Bool_1_argbuf_emit_q[1])) ? C12_12_dc(1'd1) :
                                            {4'd0, 1'd0}))))))))))));
  
  /* demux (Ty QTree_Bool,
       Ty QTree_Bool) : (lizzieLet20_1_4,QTree_Bool) (readPointer_QTree_Boolm3a8I_1_argbuf_rwb,QTree_Bool) > [(_61,QTree_Bool),
                                                                                                              (lizzieLet20_1_4QVal_Bool,QTree_Bool),
                                                                                                              (lizzieLet20_1_4QNode_Bool,QTree_Bool),
                                                                                                              (_60,QTree_Bool)] */
  logic [3:0] readPointer_QTree_Boolm3a8I_1_argbuf_rwb_onehotd;
  always_comb
    if ((lizzieLet20_1_4_d[0] && readPointer_QTree_Boolm3a8I_1_argbuf_rwb_d[0]))
      unique case (lizzieLet20_1_4_d[2:1])
        2'd0: readPointer_QTree_Boolm3a8I_1_argbuf_rwb_onehotd = 4'd1;
        2'd1: readPointer_QTree_Boolm3a8I_1_argbuf_rwb_onehotd = 4'd2;
        2'd2: readPointer_QTree_Boolm3a8I_1_argbuf_rwb_onehotd = 4'd4;
        2'd3: readPointer_QTree_Boolm3a8I_1_argbuf_rwb_onehotd = 4'd8;
        default: readPointer_QTree_Boolm3a8I_1_argbuf_rwb_onehotd = 4'd0;
      endcase
    else readPointer_QTree_Boolm3a8I_1_argbuf_rwb_onehotd = 4'd0;
  assign _61_d = {readPointer_QTree_Boolm3a8I_1_argbuf_rwb_d[66:1],
                  readPointer_QTree_Boolm3a8I_1_argbuf_rwb_onehotd[0]};
  assign lizzieLet20_1_4QVal_Bool_d = {readPointer_QTree_Boolm3a8I_1_argbuf_rwb_d[66:1],
                                       readPointer_QTree_Boolm3a8I_1_argbuf_rwb_onehotd[1]};
  assign lizzieLet20_1_4QNode_Bool_d = {readPointer_QTree_Boolm3a8I_1_argbuf_rwb_d[66:1],
                                        readPointer_QTree_Boolm3a8I_1_argbuf_rwb_onehotd[2]};
  assign _60_d = {readPointer_QTree_Boolm3a8I_1_argbuf_rwb_d[66:1],
                  readPointer_QTree_Boolm3a8I_1_argbuf_rwb_onehotd[3]};
  assign readPointer_QTree_Boolm3a8I_1_argbuf_rwb_r = (| (readPointer_QTree_Boolm3a8I_1_argbuf_rwb_onehotd & {_60_r,
                                                                                                              lizzieLet20_1_4QNode_Bool_r,
                                                                                                              lizzieLet20_1_4QVal_Bool_r,
                                                                                                              _61_r}));
  assign lizzieLet20_1_4_r = readPointer_QTree_Boolm3a8I_1_argbuf_rwb_r;
  
  /* fork (Ty QTree_Bool) : (lizzieLet20_1_4QNode_Bool,QTree_Bool) > [(lizzieLet20_1_4QNode_Bool_1,QTree_Bool),
                                                                 (lizzieLet20_1_4QNode_Bool_2,QTree_Bool),
                                                                 (lizzieLet20_1_4QNode_Bool_3,QTree_Bool),
                                                                 (lizzieLet20_1_4QNode_Bool_4,QTree_Bool),
                                                                 (lizzieLet20_1_4QNode_Bool_5,QTree_Bool),
                                                                 (lizzieLet20_1_4QNode_Bool_6,QTree_Bool),
                                                                 (lizzieLet20_1_4QNode_Bool_7,QTree_Bool),
                                                                 (lizzieLet20_1_4QNode_Bool_8,QTree_Bool),
                                                                 (lizzieLet20_1_4QNode_Bool_9,QTree_Bool)] */
  logic [8:0] lizzieLet20_1_4QNode_Bool_emitted;
  logic [8:0] lizzieLet20_1_4QNode_Bool_done;
  assign lizzieLet20_1_4QNode_Bool_1_d = {lizzieLet20_1_4QNode_Bool_d[66:1],
                                          (lizzieLet20_1_4QNode_Bool_d[0] && (! lizzieLet20_1_4QNode_Bool_emitted[0]))};
  assign lizzieLet20_1_4QNode_Bool_2_d = {lizzieLet20_1_4QNode_Bool_d[66:1],
                                          (lizzieLet20_1_4QNode_Bool_d[0] && (! lizzieLet20_1_4QNode_Bool_emitted[1]))};
  assign lizzieLet20_1_4QNode_Bool_3_d = {lizzieLet20_1_4QNode_Bool_d[66:1],
                                          (lizzieLet20_1_4QNode_Bool_d[0] && (! lizzieLet20_1_4QNode_Bool_emitted[2]))};
  assign lizzieLet20_1_4QNode_Bool_4_d = {lizzieLet20_1_4QNode_Bool_d[66:1],
                                          (lizzieLet20_1_4QNode_Bool_d[0] && (! lizzieLet20_1_4QNode_Bool_emitted[3]))};
  assign lizzieLet20_1_4QNode_Bool_5_d = {lizzieLet20_1_4QNode_Bool_d[66:1],
                                          (lizzieLet20_1_4QNode_Bool_d[0] && (! lizzieLet20_1_4QNode_Bool_emitted[4]))};
  assign lizzieLet20_1_4QNode_Bool_6_d = {lizzieLet20_1_4QNode_Bool_d[66:1],
                                          (lizzieLet20_1_4QNode_Bool_d[0] && (! lizzieLet20_1_4QNode_Bool_emitted[5]))};
  assign lizzieLet20_1_4QNode_Bool_7_d = {lizzieLet20_1_4QNode_Bool_d[66:1],
                                          (lizzieLet20_1_4QNode_Bool_d[0] && (! lizzieLet20_1_4QNode_Bool_emitted[6]))};
  assign lizzieLet20_1_4QNode_Bool_8_d = {lizzieLet20_1_4QNode_Bool_d[66:1],
                                          (lizzieLet20_1_4QNode_Bool_d[0] && (! lizzieLet20_1_4QNode_Bool_emitted[7]))};
  assign lizzieLet20_1_4QNode_Bool_9_d = {lizzieLet20_1_4QNode_Bool_d[66:1],
                                          (lizzieLet20_1_4QNode_Bool_d[0] && (! lizzieLet20_1_4QNode_Bool_emitted[8]))};
  assign lizzieLet20_1_4QNode_Bool_done = (lizzieLet20_1_4QNode_Bool_emitted | ({lizzieLet20_1_4QNode_Bool_9_d[0],
                                                                                 lizzieLet20_1_4QNode_Bool_8_d[0],
                                                                                 lizzieLet20_1_4QNode_Bool_7_d[0],
                                                                                 lizzieLet20_1_4QNode_Bool_6_d[0],
                                                                                 lizzieLet20_1_4QNode_Bool_5_d[0],
                                                                                 lizzieLet20_1_4QNode_Bool_4_d[0],
                                                                                 lizzieLet20_1_4QNode_Bool_3_d[0],
                                                                                 lizzieLet20_1_4QNode_Bool_2_d[0],
                                                                                 lizzieLet20_1_4QNode_Bool_1_d[0]} & {lizzieLet20_1_4QNode_Bool_9_r,
                                                                                                                      lizzieLet20_1_4QNode_Bool_8_r,
                                                                                                                      lizzieLet20_1_4QNode_Bool_7_r,
                                                                                                                      lizzieLet20_1_4QNode_Bool_6_r,
                                                                                                                      lizzieLet20_1_4QNode_Bool_5_r,
                                                                                                                      lizzieLet20_1_4QNode_Bool_4_r,
                                                                                                                      lizzieLet20_1_4QNode_Bool_3_r,
                                                                                                                      lizzieLet20_1_4QNode_Bool_2_r,
                                                                                                                      lizzieLet20_1_4QNode_Bool_1_r}));
  assign lizzieLet20_1_4QNode_Bool_r = (& lizzieLet20_1_4QNode_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet20_1_4QNode_Bool_emitted <= 9'd0;
    else
      lizzieLet20_1_4QNode_Bool_emitted <= (lizzieLet20_1_4QNode_Bool_r ? 9'd0 :
                                            lizzieLet20_1_4QNode_Bool_done);
  
  /* destruct (Ty QTree_Bool,
          Dcon QNode_Bool) : (lizzieLet20_1_4QNode_Bool_1QNode_Bool,QTree_Bool) > [(t1a8U_destruct,Pointer_QTree_Bool),
                                                                                   (t2a8V_destruct,Pointer_QTree_Bool),
                                                                                   (t3a8W_destruct,Pointer_QTree_Bool),
                                                                                   (t4a8X_destruct,Pointer_QTree_Bool)] */
  logic [3:0] lizzieLet20_1_4QNode_Bool_1QNode_Bool_emitted;
  logic [3:0] lizzieLet20_1_4QNode_Bool_1QNode_Bool_done;
  assign t1a8U_destruct_d = {lizzieLet20_1_4QNode_Bool_1QNode_Bool_d[18:3],
                             (lizzieLet20_1_4QNode_Bool_1QNode_Bool_d[0] && (! lizzieLet20_1_4QNode_Bool_1QNode_Bool_emitted[0]))};
  assign t2a8V_destruct_d = {lizzieLet20_1_4QNode_Bool_1QNode_Bool_d[34:19],
                             (lizzieLet20_1_4QNode_Bool_1QNode_Bool_d[0] && (! lizzieLet20_1_4QNode_Bool_1QNode_Bool_emitted[1]))};
  assign t3a8W_destruct_d = {lizzieLet20_1_4QNode_Bool_1QNode_Bool_d[50:35],
                             (lizzieLet20_1_4QNode_Bool_1QNode_Bool_d[0] && (! lizzieLet20_1_4QNode_Bool_1QNode_Bool_emitted[2]))};
  assign t4a8X_destruct_d = {lizzieLet20_1_4QNode_Bool_1QNode_Bool_d[66:51],
                             (lizzieLet20_1_4QNode_Bool_1QNode_Bool_d[0] && (! lizzieLet20_1_4QNode_Bool_1QNode_Bool_emitted[3]))};
  assign lizzieLet20_1_4QNode_Bool_1QNode_Bool_done = (lizzieLet20_1_4QNode_Bool_1QNode_Bool_emitted | ({t4a8X_destruct_d[0],
                                                                                                         t3a8W_destruct_d[0],
                                                                                                         t2a8V_destruct_d[0],
                                                                                                         t1a8U_destruct_d[0]} & {t4a8X_destruct_r,
                                                                                                                                 t3a8W_destruct_r,
                                                                                                                                 t2a8V_destruct_r,
                                                                                                                                 t1a8U_destruct_r}));
  assign lizzieLet20_1_4QNode_Bool_1QNode_Bool_r = (& lizzieLet20_1_4QNode_Bool_1QNode_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet20_1_4QNode_Bool_1QNode_Bool_emitted <= 4'd0;
    else
      lizzieLet20_1_4QNode_Bool_1QNode_Bool_emitted <= (lizzieLet20_1_4QNode_Bool_1QNode_Bool_r ? 4'd0 :
                                                        lizzieLet20_1_4QNode_Bool_1QNode_Bool_done);
  
  /* demux (Ty QTree_Bool,
       Ty QTree_Bool) : (lizzieLet20_1_4QNode_Bool_2,QTree_Bool) (lizzieLet20_1_4QNode_Bool_1,QTree_Bool) > [(_59,QTree_Bool),
                                                                                                             (_58,QTree_Bool),
                                                                                                             (lizzieLet20_1_4QNode_Bool_1QNode_Bool,QTree_Bool),
                                                                                                             (_57,QTree_Bool)] */
  logic [3:0] lizzieLet20_1_4QNode_Bool_1_onehotd;
  always_comb
    if ((lizzieLet20_1_4QNode_Bool_2_d[0] && lizzieLet20_1_4QNode_Bool_1_d[0]))
      unique case (lizzieLet20_1_4QNode_Bool_2_d[2:1])
        2'd0: lizzieLet20_1_4QNode_Bool_1_onehotd = 4'd1;
        2'd1: lizzieLet20_1_4QNode_Bool_1_onehotd = 4'd2;
        2'd2: lizzieLet20_1_4QNode_Bool_1_onehotd = 4'd4;
        2'd3: lizzieLet20_1_4QNode_Bool_1_onehotd = 4'd8;
        default: lizzieLet20_1_4QNode_Bool_1_onehotd = 4'd0;
      endcase
    else lizzieLet20_1_4QNode_Bool_1_onehotd = 4'd0;
  assign _59_d = {lizzieLet20_1_4QNode_Bool_1_d[66:1],
                  lizzieLet20_1_4QNode_Bool_1_onehotd[0]};
  assign _58_d = {lizzieLet20_1_4QNode_Bool_1_d[66:1],
                  lizzieLet20_1_4QNode_Bool_1_onehotd[1]};
  assign lizzieLet20_1_4QNode_Bool_1QNode_Bool_d = {lizzieLet20_1_4QNode_Bool_1_d[66:1],
                                                    lizzieLet20_1_4QNode_Bool_1_onehotd[2]};
  assign _57_d = {lizzieLet20_1_4QNode_Bool_1_d[66:1],
                  lizzieLet20_1_4QNode_Bool_1_onehotd[3]};
  assign lizzieLet20_1_4QNode_Bool_1_r = (| (lizzieLet20_1_4QNode_Bool_1_onehotd & {_57_r,
                                                                                    lizzieLet20_1_4QNode_Bool_1QNode_Bool_r,
                                                                                    _58_r,
                                                                                    _59_r}));
  assign lizzieLet20_1_4QNode_Bool_2_r = lizzieLet20_1_4QNode_Bool_1_r;
  
  /* demux (Ty QTree_Bool,
       Ty Go) : (lizzieLet20_1_4QNode_Bool_3,QTree_Bool) (lizzieLet20_1_3QNode_Bool,Go) > [(lizzieLet20_1_4QNode_Bool_3QNone_Bool,Go),
                                                                                           (lizzieLet20_1_4QNode_Bool_3QVal_Bool,Go),
                                                                                           (lizzieLet20_1_4QNode_Bool_3QNode_Bool,Go),
                                                                                           (lizzieLet20_1_4QNode_Bool_3QError_Bool,Go)] */
  logic [3:0] lizzieLet20_1_3QNode_Bool_onehotd;
  always_comb
    if ((lizzieLet20_1_4QNode_Bool_3_d[0] && lizzieLet20_1_3QNode_Bool_d[0]))
      unique case (lizzieLet20_1_4QNode_Bool_3_d[2:1])
        2'd0: lizzieLet20_1_3QNode_Bool_onehotd = 4'd1;
        2'd1: lizzieLet20_1_3QNode_Bool_onehotd = 4'd2;
        2'd2: lizzieLet20_1_3QNode_Bool_onehotd = 4'd4;
        2'd3: lizzieLet20_1_3QNode_Bool_onehotd = 4'd8;
        default: lizzieLet20_1_3QNode_Bool_onehotd = 4'd0;
      endcase
    else lizzieLet20_1_3QNode_Bool_onehotd = 4'd0;
  assign lizzieLet20_1_4QNode_Bool_3QNone_Bool_d = lizzieLet20_1_3QNode_Bool_onehotd[0];
  assign lizzieLet20_1_4QNode_Bool_3QVal_Bool_d = lizzieLet20_1_3QNode_Bool_onehotd[1];
  assign lizzieLet20_1_4QNode_Bool_3QNode_Bool_d = lizzieLet20_1_3QNode_Bool_onehotd[2];
  assign lizzieLet20_1_4QNode_Bool_3QError_Bool_d = lizzieLet20_1_3QNode_Bool_onehotd[3];
  assign lizzieLet20_1_3QNode_Bool_r = (| (lizzieLet20_1_3QNode_Bool_onehotd & {lizzieLet20_1_4QNode_Bool_3QError_Bool_r,
                                                                                lizzieLet20_1_4QNode_Bool_3QNode_Bool_r,
                                                                                lizzieLet20_1_4QNode_Bool_3QVal_Bool_r,
                                                                                lizzieLet20_1_4QNode_Bool_3QNone_Bool_r}));
  assign lizzieLet20_1_4QNode_Bool_3_r = lizzieLet20_1_3QNode_Bool_r;
  
  /* fork (Ty Go) : (lizzieLet20_1_4QNode_Bool_3QError_Bool,Go) > [(lizzieLet20_1_4QNode_Bool_3QError_Bool_1,Go),
                                                              (lizzieLet20_1_4QNode_Bool_3QError_Bool_2,Go)] */
  logic [1:0] lizzieLet20_1_4QNode_Bool_3QError_Bool_emitted;
  logic [1:0] lizzieLet20_1_4QNode_Bool_3QError_Bool_done;
  assign lizzieLet20_1_4QNode_Bool_3QError_Bool_1_d = (lizzieLet20_1_4QNode_Bool_3QError_Bool_d[0] && (! lizzieLet20_1_4QNode_Bool_3QError_Bool_emitted[0]));
  assign lizzieLet20_1_4QNode_Bool_3QError_Bool_2_d = (lizzieLet20_1_4QNode_Bool_3QError_Bool_d[0] && (! lizzieLet20_1_4QNode_Bool_3QError_Bool_emitted[1]));
  assign lizzieLet20_1_4QNode_Bool_3QError_Bool_done = (lizzieLet20_1_4QNode_Bool_3QError_Bool_emitted | ({lizzieLet20_1_4QNode_Bool_3QError_Bool_2_d[0],
                                                                                                           lizzieLet20_1_4QNode_Bool_3QError_Bool_1_d[0]} & {lizzieLet20_1_4QNode_Bool_3QError_Bool_2_r,
                                                                                                                                                             lizzieLet20_1_4QNode_Bool_3QError_Bool_1_r}));
  assign lizzieLet20_1_4QNode_Bool_3QError_Bool_r = (& lizzieLet20_1_4QNode_Bool_3QError_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet20_1_4QNode_Bool_3QError_Bool_emitted <= 2'd0;
    else
      lizzieLet20_1_4QNode_Bool_3QError_Bool_emitted <= (lizzieLet20_1_4QNode_Bool_3QError_Bool_r ? 2'd0 :
                                                         lizzieLet20_1_4QNode_Bool_3QError_Bool_done);
  
  /* dcon (Ty QTree_Bool,
      Dcon QError_Bool) : [(lizzieLet20_1_4QNode_Bool_3QError_Bool_1,Go)] > (lizzieLet20_1_4QNode_Bool_3QError_Bool_1QError_Bool,QTree_Bool) */
  assign lizzieLet20_1_4QNode_Bool_3QError_Bool_1QError_Bool_d = QError_Bool_dc((& {lizzieLet20_1_4QNode_Bool_3QError_Bool_1_d[0]}), lizzieLet20_1_4QNode_Bool_3QError_Bool_1_d);
  assign {lizzieLet20_1_4QNode_Bool_3QError_Bool_1_r} = {1 {(lizzieLet20_1_4QNode_Bool_3QError_Bool_1QError_Bool_r && lizzieLet20_1_4QNode_Bool_3QError_Bool_1QError_Bool_d[0])}};
  
  /* buf (Ty QTree_Bool) : (lizzieLet20_1_4QNode_Bool_3QError_Bool_1QError_Bool,QTree_Bool) > (lizzieLet30_1_argbuf,QTree_Bool) */
  QTree_Bool_t lizzieLet20_1_4QNode_Bool_3QError_Bool_1QError_Bool_bufchan_d;
  logic lizzieLet20_1_4QNode_Bool_3QError_Bool_1QError_Bool_bufchan_r;
  assign lizzieLet20_1_4QNode_Bool_3QError_Bool_1QError_Bool_r = ((! lizzieLet20_1_4QNode_Bool_3QError_Bool_1QError_Bool_bufchan_d[0]) || lizzieLet20_1_4QNode_Bool_3QError_Bool_1QError_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet20_1_4QNode_Bool_3QError_Bool_1QError_Bool_bufchan_d <= {66'd0,
                                                                        1'd0};
    else
      if (lizzieLet20_1_4QNode_Bool_3QError_Bool_1QError_Bool_r)
        lizzieLet20_1_4QNode_Bool_3QError_Bool_1QError_Bool_bufchan_d <= lizzieLet20_1_4QNode_Bool_3QError_Bool_1QError_Bool_d;
  QTree_Bool_t lizzieLet20_1_4QNode_Bool_3QError_Bool_1QError_Bool_bufchan_buf;
  assign lizzieLet20_1_4QNode_Bool_3QError_Bool_1QError_Bool_bufchan_r = (! lizzieLet20_1_4QNode_Bool_3QError_Bool_1QError_Bool_bufchan_buf[0]);
  assign lizzieLet30_1_argbuf_d = (lizzieLet20_1_4QNode_Bool_3QError_Bool_1QError_Bool_bufchan_buf[0] ? lizzieLet20_1_4QNode_Bool_3QError_Bool_1QError_Bool_bufchan_buf :
                                   lizzieLet20_1_4QNode_Bool_3QError_Bool_1QError_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet20_1_4QNode_Bool_3QError_Bool_1QError_Bool_bufchan_buf <= {66'd0,
                                                                          1'd0};
    else
      if ((lizzieLet30_1_argbuf_r && lizzieLet20_1_4QNode_Bool_3QError_Bool_1QError_Bool_bufchan_buf[0]))
        lizzieLet20_1_4QNode_Bool_3QError_Bool_1QError_Bool_bufchan_buf <= {66'd0,
                                                                            1'd0};
      else if (((! lizzieLet30_1_argbuf_r) && (! lizzieLet20_1_4QNode_Bool_3QError_Bool_1QError_Bool_bufchan_buf[0])))
        lizzieLet20_1_4QNode_Bool_3QError_Bool_1QError_Bool_bufchan_buf <= lizzieLet20_1_4QNode_Bool_3QError_Bool_1QError_Bool_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet20_1_4QNode_Bool_3QError_Bool_2,Go) > (lizzieLet20_1_4QNode_Bool_3QError_Bool_2_argbuf,Go) */
  Go_t lizzieLet20_1_4QNode_Bool_3QError_Bool_2_bufchan_d;
  logic lizzieLet20_1_4QNode_Bool_3QError_Bool_2_bufchan_r;
  assign lizzieLet20_1_4QNode_Bool_3QError_Bool_2_r = ((! lizzieLet20_1_4QNode_Bool_3QError_Bool_2_bufchan_d[0]) || lizzieLet20_1_4QNode_Bool_3QError_Bool_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet20_1_4QNode_Bool_3QError_Bool_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet20_1_4QNode_Bool_3QError_Bool_2_r)
        lizzieLet20_1_4QNode_Bool_3QError_Bool_2_bufchan_d <= lizzieLet20_1_4QNode_Bool_3QError_Bool_2_d;
  Go_t lizzieLet20_1_4QNode_Bool_3QError_Bool_2_bufchan_buf;
  assign lizzieLet20_1_4QNode_Bool_3QError_Bool_2_bufchan_r = (! lizzieLet20_1_4QNode_Bool_3QError_Bool_2_bufchan_buf[0]);
  assign lizzieLet20_1_4QNode_Bool_3QError_Bool_2_argbuf_d = (lizzieLet20_1_4QNode_Bool_3QError_Bool_2_bufchan_buf[0] ? lizzieLet20_1_4QNode_Bool_3QError_Bool_2_bufchan_buf :
                                                              lizzieLet20_1_4QNode_Bool_3QError_Bool_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet20_1_4QNode_Bool_3QError_Bool_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet20_1_4QNode_Bool_3QError_Bool_2_argbuf_r && lizzieLet20_1_4QNode_Bool_3QError_Bool_2_bufchan_buf[0]))
        lizzieLet20_1_4QNode_Bool_3QError_Bool_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet20_1_4QNode_Bool_3QError_Bool_2_argbuf_r) && (! lizzieLet20_1_4QNode_Bool_3QError_Bool_2_bufchan_buf[0])))
        lizzieLet20_1_4QNode_Bool_3QError_Bool_2_bufchan_buf <= lizzieLet20_1_4QNode_Bool_3QError_Bool_2_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet20_1_4QNode_Bool_3QNode_Bool,Go) > (lizzieLet20_1_4QNode_Bool_3QNode_Bool_1_argbuf,Go) */
  Go_t lizzieLet20_1_4QNode_Bool_3QNode_Bool_bufchan_d;
  logic lizzieLet20_1_4QNode_Bool_3QNode_Bool_bufchan_r;
  assign lizzieLet20_1_4QNode_Bool_3QNode_Bool_r = ((! lizzieLet20_1_4QNode_Bool_3QNode_Bool_bufchan_d[0]) || lizzieLet20_1_4QNode_Bool_3QNode_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet20_1_4QNode_Bool_3QNode_Bool_bufchan_d <= 1'd0;
    else
      if (lizzieLet20_1_4QNode_Bool_3QNode_Bool_r)
        lizzieLet20_1_4QNode_Bool_3QNode_Bool_bufchan_d <= lizzieLet20_1_4QNode_Bool_3QNode_Bool_d;
  Go_t lizzieLet20_1_4QNode_Bool_3QNode_Bool_bufchan_buf;
  assign lizzieLet20_1_4QNode_Bool_3QNode_Bool_bufchan_r = (! lizzieLet20_1_4QNode_Bool_3QNode_Bool_bufchan_buf[0]);
  assign lizzieLet20_1_4QNode_Bool_3QNode_Bool_1_argbuf_d = (lizzieLet20_1_4QNode_Bool_3QNode_Bool_bufchan_buf[0] ? lizzieLet20_1_4QNode_Bool_3QNode_Bool_bufchan_buf :
                                                             lizzieLet20_1_4QNode_Bool_3QNode_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet20_1_4QNode_Bool_3QNode_Bool_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet20_1_4QNode_Bool_3QNode_Bool_1_argbuf_r && lizzieLet20_1_4QNode_Bool_3QNode_Bool_bufchan_buf[0]))
        lizzieLet20_1_4QNode_Bool_3QNode_Bool_bufchan_buf <= 1'd0;
      else if (((! lizzieLet20_1_4QNode_Bool_3QNode_Bool_1_argbuf_r) && (! lizzieLet20_1_4QNode_Bool_3QNode_Bool_bufchan_buf[0])))
        lizzieLet20_1_4QNode_Bool_3QNode_Bool_bufchan_buf <= lizzieLet20_1_4QNode_Bool_3QNode_Bool_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet20_1_4QNode_Bool_3QNone_Bool,Go) > (lizzieLet20_1_4QNode_Bool_3QNone_Bool_1_argbuf,Go) */
  Go_t lizzieLet20_1_4QNode_Bool_3QNone_Bool_bufchan_d;
  logic lizzieLet20_1_4QNode_Bool_3QNone_Bool_bufchan_r;
  assign lizzieLet20_1_4QNode_Bool_3QNone_Bool_r = ((! lizzieLet20_1_4QNode_Bool_3QNone_Bool_bufchan_d[0]) || lizzieLet20_1_4QNode_Bool_3QNone_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet20_1_4QNode_Bool_3QNone_Bool_bufchan_d <= 1'd0;
    else
      if (lizzieLet20_1_4QNode_Bool_3QNone_Bool_r)
        lizzieLet20_1_4QNode_Bool_3QNone_Bool_bufchan_d <= lizzieLet20_1_4QNode_Bool_3QNone_Bool_d;
  Go_t lizzieLet20_1_4QNode_Bool_3QNone_Bool_bufchan_buf;
  assign lizzieLet20_1_4QNode_Bool_3QNone_Bool_bufchan_r = (! lizzieLet20_1_4QNode_Bool_3QNone_Bool_bufchan_buf[0]);
  assign lizzieLet20_1_4QNode_Bool_3QNone_Bool_1_argbuf_d = (lizzieLet20_1_4QNode_Bool_3QNone_Bool_bufchan_buf[0] ? lizzieLet20_1_4QNode_Bool_3QNone_Bool_bufchan_buf :
                                                             lizzieLet20_1_4QNode_Bool_3QNone_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet20_1_4QNode_Bool_3QNone_Bool_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet20_1_4QNode_Bool_3QNone_Bool_1_argbuf_r && lizzieLet20_1_4QNode_Bool_3QNone_Bool_bufchan_buf[0]))
        lizzieLet20_1_4QNode_Bool_3QNone_Bool_bufchan_buf <= 1'd0;
      else if (((! lizzieLet20_1_4QNode_Bool_3QNone_Bool_1_argbuf_r) && (! lizzieLet20_1_4QNode_Bool_3QNone_Bool_bufchan_buf[0])))
        lizzieLet20_1_4QNode_Bool_3QNone_Bool_bufchan_buf <= lizzieLet20_1_4QNode_Bool_3QNone_Bool_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet20_1_4QNode_Bool_3QVal_Bool,Go) > [(lizzieLet20_1_4QNode_Bool_3QVal_Bool_1,Go),
                                                            (lizzieLet20_1_4QNode_Bool_3QVal_Bool_2,Go)] */
  logic [1:0] lizzieLet20_1_4QNode_Bool_3QVal_Bool_emitted;
  logic [1:0] lizzieLet20_1_4QNode_Bool_3QVal_Bool_done;
  assign lizzieLet20_1_4QNode_Bool_3QVal_Bool_1_d = (lizzieLet20_1_4QNode_Bool_3QVal_Bool_d[0] && (! lizzieLet20_1_4QNode_Bool_3QVal_Bool_emitted[0]));
  assign lizzieLet20_1_4QNode_Bool_3QVal_Bool_2_d = (lizzieLet20_1_4QNode_Bool_3QVal_Bool_d[0] && (! lizzieLet20_1_4QNode_Bool_3QVal_Bool_emitted[1]));
  assign lizzieLet20_1_4QNode_Bool_3QVal_Bool_done = (lizzieLet20_1_4QNode_Bool_3QVal_Bool_emitted | ({lizzieLet20_1_4QNode_Bool_3QVal_Bool_2_d[0],
                                                                                                       lizzieLet20_1_4QNode_Bool_3QVal_Bool_1_d[0]} & {lizzieLet20_1_4QNode_Bool_3QVal_Bool_2_r,
                                                                                                                                                       lizzieLet20_1_4QNode_Bool_3QVal_Bool_1_r}));
  assign lizzieLet20_1_4QNode_Bool_3QVal_Bool_r = (& lizzieLet20_1_4QNode_Bool_3QVal_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet20_1_4QNode_Bool_3QVal_Bool_emitted <= 2'd0;
    else
      lizzieLet20_1_4QNode_Bool_3QVal_Bool_emitted <= (lizzieLet20_1_4QNode_Bool_3QVal_Bool_r ? 2'd0 :
                                                       lizzieLet20_1_4QNode_Bool_3QVal_Bool_done);
  
  /* dcon (Ty QTree_Bool,
      Dcon QError_Bool) : [(lizzieLet20_1_4QNode_Bool_3QVal_Bool_1,Go)] > (lizzieLet20_1_4QNode_Bool_3QVal_Bool_1QError_Bool,QTree_Bool) */
  assign lizzieLet20_1_4QNode_Bool_3QVal_Bool_1QError_Bool_d = QError_Bool_dc((& {lizzieLet20_1_4QNode_Bool_3QVal_Bool_1_d[0]}), lizzieLet20_1_4QNode_Bool_3QVal_Bool_1_d);
  assign {lizzieLet20_1_4QNode_Bool_3QVal_Bool_1_r} = {1 {(lizzieLet20_1_4QNode_Bool_3QVal_Bool_1QError_Bool_r && lizzieLet20_1_4QNode_Bool_3QVal_Bool_1QError_Bool_d[0])}};
  
  /* buf (Ty QTree_Bool) : (lizzieLet20_1_4QNode_Bool_3QVal_Bool_1QError_Bool,QTree_Bool) > (lizzieLet28_1_argbuf,QTree_Bool) */
  QTree_Bool_t lizzieLet20_1_4QNode_Bool_3QVal_Bool_1QError_Bool_bufchan_d;
  logic lizzieLet20_1_4QNode_Bool_3QVal_Bool_1QError_Bool_bufchan_r;
  assign lizzieLet20_1_4QNode_Bool_3QVal_Bool_1QError_Bool_r = ((! lizzieLet20_1_4QNode_Bool_3QVal_Bool_1QError_Bool_bufchan_d[0]) || lizzieLet20_1_4QNode_Bool_3QVal_Bool_1QError_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet20_1_4QNode_Bool_3QVal_Bool_1QError_Bool_bufchan_d <= {66'd0,
                                                                      1'd0};
    else
      if (lizzieLet20_1_4QNode_Bool_3QVal_Bool_1QError_Bool_r)
        lizzieLet20_1_4QNode_Bool_3QVal_Bool_1QError_Bool_bufchan_d <= lizzieLet20_1_4QNode_Bool_3QVal_Bool_1QError_Bool_d;
  QTree_Bool_t lizzieLet20_1_4QNode_Bool_3QVal_Bool_1QError_Bool_bufchan_buf;
  assign lizzieLet20_1_4QNode_Bool_3QVal_Bool_1QError_Bool_bufchan_r = (! lizzieLet20_1_4QNode_Bool_3QVal_Bool_1QError_Bool_bufchan_buf[0]);
  assign lizzieLet28_1_argbuf_d = (lizzieLet20_1_4QNode_Bool_3QVal_Bool_1QError_Bool_bufchan_buf[0] ? lizzieLet20_1_4QNode_Bool_3QVal_Bool_1QError_Bool_bufchan_buf :
                                   lizzieLet20_1_4QNode_Bool_3QVal_Bool_1QError_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet20_1_4QNode_Bool_3QVal_Bool_1QError_Bool_bufchan_buf <= {66'd0,
                                                                        1'd0};
    else
      if ((lizzieLet28_1_argbuf_r && lizzieLet20_1_4QNode_Bool_3QVal_Bool_1QError_Bool_bufchan_buf[0]))
        lizzieLet20_1_4QNode_Bool_3QVal_Bool_1QError_Bool_bufchan_buf <= {66'd0,
                                                                          1'd0};
      else if (((! lizzieLet28_1_argbuf_r) && (! lizzieLet20_1_4QNode_Bool_3QVal_Bool_1QError_Bool_bufchan_buf[0])))
        lizzieLet20_1_4QNode_Bool_3QVal_Bool_1QError_Bool_bufchan_buf <= lizzieLet20_1_4QNode_Bool_3QVal_Bool_1QError_Bool_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet20_1_4QNode_Bool_3QVal_Bool_2,Go) > (lizzieLet20_1_4QNode_Bool_3QVal_Bool_2_argbuf,Go) */
  Go_t lizzieLet20_1_4QNode_Bool_3QVal_Bool_2_bufchan_d;
  logic lizzieLet20_1_4QNode_Bool_3QVal_Bool_2_bufchan_r;
  assign lizzieLet20_1_4QNode_Bool_3QVal_Bool_2_r = ((! lizzieLet20_1_4QNode_Bool_3QVal_Bool_2_bufchan_d[0]) || lizzieLet20_1_4QNode_Bool_3QVal_Bool_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet20_1_4QNode_Bool_3QVal_Bool_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet20_1_4QNode_Bool_3QVal_Bool_2_r)
        lizzieLet20_1_4QNode_Bool_3QVal_Bool_2_bufchan_d <= lizzieLet20_1_4QNode_Bool_3QVal_Bool_2_d;
  Go_t lizzieLet20_1_4QNode_Bool_3QVal_Bool_2_bufchan_buf;
  assign lizzieLet20_1_4QNode_Bool_3QVal_Bool_2_bufchan_r = (! lizzieLet20_1_4QNode_Bool_3QVal_Bool_2_bufchan_buf[0]);
  assign lizzieLet20_1_4QNode_Bool_3QVal_Bool_2_argbuf_d = (lizzieLet20_1_4QNode_Bool_3QVal_Bool_2_bufchan_buf[0] ? lizzieLet20_1_4QNode_Bool_3QVal_Bool_2_bufchan_buf :
                                                            lizzieLet20_1_4QNode_Bool_3QVal_Bool_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet20_1_4QNode_Bool_3QVal_Bool_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet20_1_4QNode_Bool_3QVal_Bool_2_argbuf_r && lizzieLet20_1_4QNode_Bool_3QVal_Bool_2_bufchan_buf[0]))
        lizzieLet20_1_4QNode_Bool_3QVal_Bool_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet20_1_4QNode_Bool_3QVal_Bool_2_argbuf_r) && (! lizzieLet20_1_4QNode_Bool_3QVal_Bool_2_bufchan_buf[0])))
        lizzieLet20_1_4QNode_Bool_3QVal_Bool_2_bufchan_buf <= lizzieLet20_1_4QNode_Bool_3QVal_Bool_2_bufchan_d;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_QTree_Bool) : (lizzieLet20_1_4QNode_Bool_4,QTree_Bool) (lizzieLet20_1_5QNode_Bool,Pointer_QTree_Bool) > [(lizzieLet20_1_4QNode_Bool_4QNone_Bool,Pointer_QTree_Bool),
                                                                                                                           (_56,Pointer_QTree_Bool),
                                                                                                                           (_55,Pointer_QTree_Bool),
                                                                                                                           (_54,Pointer_QTree_Bool)] */
  logic [3:0] lizzieLet20_1_5QNode_Bool_onehotd;
  always_comb
    if ((lizzieLet20_1_4QNode_Bool_4_d[0] && lizzieLet20_1_5QNode_Bool_d[0]))
      unique case (lizzieLet20_1_4QNode_Bool_4_d[2:1])
        2'd0: lizzieLet20_1_5QNode_Bool_onehotd = 4'd1;
        2'd1: lizzieLet20_1_5QNode_Bool_onehotd = 4'd2;
        2'd2: lizzieLet20_1_5QNode_Bool_onehotd = 4'd4;
        2'd3: lizzieLet20_1_5QNode_Bool_onehotd = 4'd8;
        default: lizzieLet20_1_5QNode_Bool_onehotd = 4'd0;
      endcase
    else lizzieLet20_1_5QNode_Bool_onehotd = 4'd0;
  assign lizzieLet20_1_4QNode_Bool_4QNone_Bool_d = {lizzieLet20_1_5QNode_Bool_d[16:1],
                                                    lizzieLet20_1_5QNode_Bool_onehotd[0]};
  assign _56_d = {lizzieLet20_1_5QNode_Bool_d[16:1],
                  lizzieLet20_1_5QNode_Bool_onehotd[1]};
  assign _55_d = {lizzieLet20_1_5QNode_Bool_d[16:1],
                  lizzieLet20_1_5QNode_Bool_onehotd[2]};
  assign _54_d = {lizzieLet20_1_5QNode_Bool_d[16:1],
                  lizzieLet20_1_5QNode_Bool_onehotd[3]};
  assign lizzieLet20_1_5QNode_Bool_r = (| (lizzieLet20_1_5QNode_Bool_onehotd & {_54_r,
                                                                                _55_r,
                                                                                _56_r,
                                                                                lizzieLet20_1_4QNode_Bool_4QNone_Bool_r}));
  assign lizzieLet20_1_4QNode_Bool_4_r = lizzieLet20_1_5QNode_Bool_r;
  
  /* buf (Ty Pointer_QTree_Bool) : (lizzieLet20_1_4QNode_Bool_4QNone_Bool,Pointer_QTree_Bool) > (lizzieLet20_1_4QNode_Bool_4QNone_Bool_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t lizzieLet20_1_4QNode_Bool_4QNone_Bool_bufchan_d;
  logic lizzieLet20_1_4QNode_Bool_4QNone_Bool_bufchan_r;
  assign lizzieLet20_1_4QNode_Bool_4QNone_Bool_r = ((! lizzieLet20_1_4QNode_Bool_4QNone_Bool_bufchan_d[0]) || lizzieLet20_1_4QNode_Bool_4QNone_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet20_1_4QNode_Bool_4QNone_Bool_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet20_1_4QNode_Bool_4QNone_Bool_r)
        lizzieLet20_1_4QNode_Bool_4QNone_Bool_bufchan_d <= lizzieLet20_1_4QNode_Bool_4QNone_Bool_d;
  Pointer_QTree_Bool_t lizzieLet20_1_4QNode_Bool_4QNone_Bool_bufchan_buf;
  assign lizzieLet20_1_4QNode_Bool_4QNone_Bool_bufchan_r = (! lizzieLet20_1_4QNode_Bool_4QNone_Bool_bufchan_buf[0]);
  assign lizzieLet20_1_4QNode_Bool_4QNone_Bool_1_argbuf_d = (lizzieLet20_1_4QNode_Bool_4QNone_Bool_bufchan_buf[0] ? lizzieLet20_1_4QNode_Bool_4QNone_Bool_bufchan_buf :
                                                             lizzieLet20_1_4QNode_Bool_4QNone_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet20_1_4QNode_Bool_4QNone_Bool_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet20_1_4QNode_Bool_4QNone_Bool_1_argbuf_r && lizzieLet20_1_4QNode_Bool_4QNone_Bool_bufchan_buf[0]))
        lizzieLet20_1_4QNode_Bool_4QNone_Bool_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet20_1_4QNode_Bool_4QNone_Bool_1_argbuf_r) && (! lizzieLet20_1_4QNode_Bool_4QNone_Bool_bufchan_buf[0])))
        lizzieLet20_1_4QNode_Bool_4QNone_Bool_bufchan_buf <= lizzieLet20_1_4QNode_Bool_4QNone_Bool_bufchan_d;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_CTf') : (lizzieLet20_1_4QNode_Bool_5,QTree_Bool) (lizzieLet20_1_7QNode_Bool,Pointer_CTf') > [(lizzieLet20_1_4QNode_Bool_5QNone_Bool,Pointer_CTf'),
                                                                                                               (lizzieLet20_1_4QNode_Bool_5QVal_Bool,Pointer_CTf'),
                                                                                                               (lizzieLet20_1_4QNode_Bool_5QNode_Bool,Pointer_CTf'),
                                                                                                               (lizzieLet20_1_4QNode_Bool_5QError_Bool,Pointer_CTf')] */
  logic [3:0] lizzieLet20_1_7QNode_Bool_onehotd;
  always_comb
    if ((lizzieLet20_1_4QNode_Bool_5_d[0] && lizzieLet20_1_7QNode_Bool_d[0]))
      unique case (lizzieLet20_1_4QNode_Bool_5_d[2:1])
        2'd0: lizzieLet20_1_7QNode_Bool_onehotd = 4'd1;
        2'd1: lizzieLet20_1_7QNode_Bool_onehotd = 4'd2;
        2'd2: lizzieLet20_1_7QNode_Bool_onehotd = 4'd4;
        2'd3: lizzieLet20_1_7QNode_Bool_onehotd = 4'd8;
        default: lizzieLet20_1_7QNode_Bool_onehotd = 4'd0;
      endcase
    else lizzieLet20_1_7QNode_Bool_onehotd = 4'd0;
  assign lizzieLet20_1_4QNode_Bool_5QNone_Bool_d = {lizzieLet20_1_7QNode_Bool_d[16:1],
                                                    lizzieLet20_1_7QNode_Bool_onehotd[0]};
  assign lizzieLet20_1_4QNode_Bool_5QVal_Bool_d = {lizzieLet20_1_7QNode_Bool_d[16:1],
                                                   lizzieLet20_1_7QNode_Bool_onehotd[1]};
  assign lizzieLet20_1_4QNode_Bool_5QNode_Bool_d = {lizzieLet20_1_7QNode_Bool_d[16:1],
                                                    lizzieLet20_1_7QNode_Bool_onehotd[2]};
  assign lizzieLet20_1_4QNode_Bool_5QError_Bool_d = {lizzieLet20_1_7QNode_Bool_d[16:1],
                                                     lizzieLet20_1_7QNode_Bool_onehotd[3]};
  assign lizzieLet20_1_7QNode_Bool_r = (| (lizzieLet20_1_7QNode_Bool_onehotd & {lizzieLet20_1_4QNode_Bool_5QError_Bool_r,
                                                                                lizzieLet20_1_4QNode_Bool_5QNode_Bool_r,
                                                                                lizzieLet20_1_4QNode_Bool_5QVal_Bool_r,
                                                                                lizzieLet20_1_4QNode_Bool_5QNone_Bool_r}));
  assign lizzieLet20_1_4QNode_Bool_5_r = lizzieLet20_1_7QNode_Bool_r;
  
  /* buf (Ty Pointer_CTf') : (lizzieLet20_1_4QNode_Bool_5QError_Bool,Pointer_CTf') > (lizzieLet20_1_4QNode_Bool_5QError_Bool_1_argbuf,Pointer_CTf') */
  \Pointer_CTf'_t  lizzieLet20_1_4QNode_Bool_5QError_Bool_bufchan_d;
  logic lizzieLet20_1_4QNode_Bool_5QError_Bool_bufchan_r;
  assign lizzieLet20_1_4QNode_Bool_5QError_Bool_r = ((! lizzieLet20_1_4QNode_Bool_5QError_Bool_bufchan_d[0]) || lizzieLet20_1_4QNode_Bool_5QError_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet20_1_4QNode_Bool_5QError_Bool_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet20_1_4QNode_Bool_5QError_Bool_r)
        lizzieLet20_1_4QNode_Bool_5QError_Bool_bufchan_d <= lizzieLet20_1_4QNode_Bool_5QError_Bool_d;
  \Pointer_CTf'_t  lizzieLet20_1_4QNode_Bool_5QError_Bool_bufchan_buf;
  assign lizzieLet20_1_4QNode_Bool_5QError_Bool_bufchan_r = (! lizzieLet20_1_4QNode_Bool_5QError_Bool_bufchan_buf[0]);
  assign lizzieLet20_1_4QNode_Bool_5QError_Bool_1_argbuf_d = (lizzieLet20_1_4QNode_Bool_5QError_Bool_bufchan_buf[0] ? lizzieLet20_1_4QNode_Bool_5QError_Bool_bufchan_buf :
                                                              lizzieLet20_1_4QNode_Bool_5QError_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet20_1_4QNode_Bool_5QError_Bool_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((lizzieLet20_1_4QNode_Bool_5QError_Bool_1_argbuf_r && lizzieLet20_1_4QNode_Bool_5QError_Bool_bufchan_buf[0]))
        lizzieLet20_1_4QNode_Bool_5QError_Bool_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! lizzieLet20_1_4QNode_Bool_5QError_Bool_1_argbuf_r) && (! lizzieLet20_1_4QNode_Bool_5QError_Bool_bufchan_buf[0])))
        lizzieLet20_1_4QNode_Bool_5QError_Bool_bufchan_buf <= lizzieLet20_1_4QNode_Bool_5QError_Bool_bufchan_d;
  
  /* dcon (Ty CTf',
      Dcon Lcall_f'3) : [(lizzieLet20_1_4QNode_Bool_5QNode_Bool,Pointer_CTf'),
                         (lizzieLet20_1_4QNode_Bool_6QNode_Bool,Pointer_QTree_Bool),
                         (t1a8U_destruct,Pointer_QTree_Bool),
                         (lizzieLet20_1_4QNode_Bool_7QNode_Bool,Pointer_QTree_Bool),
                         (t2a8V_destruct,Pointer_QTree_Bool),
                         (lizzieLet20_1_4QNode_Bool_8QNode_Bool,Pointer_QTree_Bool),
                         (t3a8W_destruct,Pointer_QTree_Bool)] > (lizzieLet20_1_4QNode_Bool_5QNode_Bool_1lizzieLet20_1_4QNode_Bool_6QNode_Bool_1t1a8U_1lizzieLet20_1_4QNode_Bool_7QNode_Bool_1t2a8V_1lizzieLet20_1_4QNode_Bool_8QNode_Bool_1t3a8W_1Lcall_f'3,CTf') */
  assign \lizzieLet20_1_4QNode_Bool_5QNode_Bool_1lizzieLet20_1_4QNode_Bool_6QNode_Bool_1t1a8U_1lizzieLet20_1_4QNode_Bool_7QNode_Bool_1t2a8V_1lizzieLet20_1_4QNode_Bool_8QNode_Bool_1t3a8W_1Lcall_f'3_d  = \Lcall_f'3_dc ((& {lizzieLet20_1_4QNode_Bool_5QNode_Bool_d[0],
                                                                                                                                                                                                                             lizzieLet20_1_4QNode_Bool_6QNode_Bool_d[0],
                                                                                                                                                                                                                             t1a8U_destruct_d[0],
                                                                                                                                                                                                                             lizzieLet20_1_4QNode_Bool_7QNode_Bool_d[0],
                                                                                                                                                                                                                             t2a8V_destruct_d[0],
                                                                                                                                                                                                                             lizzieLet20_1_4QNode_Bool_8QNode_Bool_d[0],
                                                                                                                                                                                                                             t3a8W_destruct_d[0]}), lizzieLet20_1_4QNode_Bool_5QNode_Bool_d, lizzieLet20_1_4QNode_Bool_6QNode_Bool_d, t1a8U_destruct_d, lizzieLet20_1_4QNode_Bool_7QNode_Bool_d, t2a8V_destruct_d, lizzieLet20_1_4QNode_Bool_8QNode_Bool_d, t3a8W_destruct_d);
  assign {lizzieLet20_1_4QNode_Bool_5QNode_Bool_r,
          lizzieLet20_1_4QNode_Bool_6QNode_Bool_r,
          t1a8U_destruct_r,
          lizzieLet20_1_4QNode_Bool_7QNode_Bool_r,
          t2a8V_destruct_r,
          lizzieLet20_1_4QNode_Bool_8QNode_Bool_r,
          t3a8W_destruct_r} = {7 {(\lizzieLet20_1_4QNode_Bool_5QNode_Bool_1lizzieLet20_1_4QNode_Bool_6QNode_Bool_1t1a8U_1lizzieLet20_1_4QNode_Bool_7QNode_Bool_1t2a8V_1lizzieLet20_1_4QNode_Bool_8QNode_Bool_1t3a8W_1Lcall_f'3_r  && \lizzieLet20_1_4QNode_Bool_5QNode_Bool_1lizzieLet20_1_4QNode_Bool_6QNode_Bool_1t1a8U_1lizzieLet20_1_4QNode_Bool_7QNode_Bool_1t2a8V_1lizzieLet20_1_4QNode_Bool_8QNode_Bool_1t3a8W_1Lcall_f'3_d [0])}};
  
  /* buf (Ty CTf') : (lizzieLet20_1_4QNode_Bool_5QNode_Bool_1lizzieLet20_1_4QNode_Bool_6QNode_Bool_1t1a8U_1lizzieLet20_1_4QNode_Bool_7QNode_Bool_1t2a8V_1lizzieLet20_1_4QNode_Bool_8QNode_Bool_1t3a8W_1Lcall_f'3,CTf') > (lizzieLet29_1_argbuf,CTf') */
  \CTf'_t  \lizzieLet20_1_4QNode_Bool_5QNode_Bool_1lizzieLet20_1_4QNode_Bool_6QNode_Bool_1t1a8U_1lizzieLet20_1_4QNode_Bool_7QNode_Bool_1t2a8V_1lizzieLet20_1_4QNode_Bool_8QNode_Bool_1t3a8W_1Lcall_f'3_bufchan_d ;
  logic \lizzieLet20_1_4QNode_Bool_5QNode_Bool_1lizzieLet20_1_4QNode_Bool_6QNode_Bool_1t1a8U_1lizzieLet20_1_4QNode_Bool_7QNode_Bool_1t2a8V_1lizzieLet20_1_4QNode_Bool_8QNode_Bool_1t3a8W_1Lcall_f'3_bufchan_r ;
  assign \lizzieLet20_1_4QNode_Bool_5QNode_Bool_1lizzieLet20_1_4QNode_Bool_6QNode_Bool_1t1a8U_1lizzieLet20_1_4QNode_Bool_7QNode_Bool_1t2a8V_1lizzieLet20_1_4QNode_Bool_8QNode_Bool_1t3a8W_1Lcall_f'3_r  = ((! \lizzieLet20_1_4QNode_Bool_5QNode_Bool_1lizzieLet20_1_4QNode_Bool_6QNode_Bool_1t1a8U_1lizzieLet20_1_4QNode_Bool_7QNode_Bool_1t2a8V_1lizzieLet20_1_4QNode_Bool_8QNode_Bool_1t3a8W_1Lcall_f'3_bufchan_d [0]) || \lizzieLet20_1_4QNode_Bool_5QNode_Bool_1lizzieLet20_1_4QNode_Bool_6QNode_Bool_1t1a8U_1lizzieLet20_1_4QNode_Bool_7QNode_Bool_1t2a8V_1lizzieLet20_1_4QNode_Bool_8QNode_Bool_1t3a8W_1Lcall_f'3_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet20_1_4QNode_Bool_5QNode_Bool_1lizzieLet20_1_4QNode_Bool_6QNode_Bool_1t1a8U_1lizzieLet20_1_4QNode_Bool_7QNode_Bool_1t2a8V_1lizzieLet20_1_4QNode_Bool_8QNode_Bool_1t3a8W_1Lcall_f'3_bufchan_d  <= {115'd0,
                                                                                                                                                                                                                 1'd0};
    else
      if (\lizzieLet20_1_4QNode_Bool_5QNode_Bool_1lizzieLet20_1_4QNode_Bool_6QNode_Bool_1t1a8U_1lizzieLet20_1_4QNode_Bool_7QNode_Bool_1t2a8V_1lizzieLet20_1_4QNode_Bool_8QNode_Bool_1t3a8W_1Lcall_f'3_r )
        \lizzieLet20_1_4QNode_Bool_5QNode_Bool_1lizzieLet20_1_4QNode_Bool_6QNode_Bool_1t1a8U_1lizzieLet20_1_4QNode_Bool_7QNode_Bool_1t2a8V_1lizzieLet20_1_4QNode_Bool_8QNode_Bool_1t3a8W_1Lcall_f'3_bufchan_d  <= \lizzieLet20_1_4QNode_Bool_5QNode_Bool_1lizzieLet20_1_4QNode_Bool_6QNode_Bool_1t1a8U_1lizzieLet20_1_4QNode_Bool_7QNode_Bool_1t2a8V_1lizzieLet20_1_4QNode_Bool_8QNode_Bool_1t3a8W_1Lcall_f'3_d ;
  \CTf'_t  \lizzieLet20_1_4QNode_Bool_5QNode_Bool_1lizzieLet20_1_4QNode_Bool_6QNode_Bool_1t1a8U_1lizzieLet20_1_4QNode_Bool_7QNode_Bool_1t2a8V_1lizzieLet20_1_4QNode_Bool_8QNode_Bool_1t3a8W_1Lcall_f'3_bufchan_buf ;
  assign \lizzieLet20_1_4QNode_Bool_5QNode_Bool_1lizzieLet20_1_4QNode_Bool_6QNode_Bool_1t1a8U_1lizzieLet20_1_4QNode_Bool_7QNode_Bool_1t2a8V_1lizzieLet20_1_4QNode_Bool_8QNode_Bool_1t3a8W_1Lcall_f'3_bufchan_r  = (! \lizzieLet20_1_4QNode_Bool_5QNode_Bool_1lizzieLet20_1_4QNode_Bool_6QNode_Bool_1t1a8U_1lizzieLet20_1_4QNode_Bool_7QNode_Bool_1t2a8V_1lizzieLet20_1_4QNode_Bool_8QNode_Bool_1t3a8W_1Lcall_f'3_bufchan_buf [0]);
  assign lizzieLet29_1_argbuf_d = (\lizzieLet20_1_4QNode_Bool_5QNode_Bool_1lizzieLet20_1_4QNode_Bool_6QNode_Bool_1t1a8U_1lizzieLet20_1_4QNode_Bool_7QNode_Bool_1t2a8V_1lizzieLet20_1_4QNode_Bool_8QNode_Bool_1t3a8W_1Lcall_f'3_bufchan_buf [0] ? \lizzieLet20_1_4QNode_Bool_5QNode_Bool_1lizzieLet20_1_4QNode_Bool_6QNode_Bool_1t1a8U_1lizzieLet20_1_4QNode_Bool_7QNode_Bool_1t2a8V_1lizzieLet20_1_4QNode_Bool_8QNode_Bool_1t3a8W_1Lcall_f'3_bufchan_buf  :
                                   \lizzieLet20_1_4QNode_Bool_5QNode_Bool_1lizzieLet20_1_4QNode_Bool_6QNode_Bool_1t1a8U_1lizzieLet20_1_4QNode_Bool_7QNode_Bool_1t2a8V_1lizzieLet20_1_4QNode_Bool_8QNode_Bool_1t3a8W_1Lcall_f'3_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet20_1_4QNode_Bool_5QNode_Bool_1lizzieLet20_1_4QNode_Bool_6QNode_Bool_1t1a8U_1lizzieLet20_1_4QNode_Bool_7QNode_Bool_1t2a8V_1lizzieLet20_1_4QNode_Bool_8QNode_Bool_1t3a8W_1Lcall_f'3_bufchan_buf  <= {115'd0,
                                                                                                                                                                                                                   1'd0};
    else
      if ((lizzieLet29_1_argbuf_r && \lizzieLet20_1_4QNode_Bool_5QNode_Bool_1lizzieLet20_1_4QNode_Bool_6QNode_Bool_1t1a8U_1lizzieLet20_1_4QNode_Bool_7QNode_Bool_1t2a8V_1lizzieLet20_1_4QNode_Bool_8QNode_Bool_1t3a8W_1Lcall_f'3_bufchan_buf [0]))
        \lizzieLet20_1_4QNode_Bool_5QNode_Bool_1lizzieLet20_1_4QNode_Bool_6QNode_Bool_1t1a8U_1lizzieLet20_1_4QNode_Bool_7QNode_Bool_1t2a8V_1lizzieLet20_1_4QNode_Bool_8QNode_Bool_1t3a8W_1Lcall_f'3_bufchan_buf  <= {115'd0,
                                                                                                                                                                                                                     1'd0};
      else if (((! lizzieLet29_1_argbuf_r) && (! \lizzieLet20_1_4QNode_Bool_5QNode_Bool_1lizzieLet20_1_4QNode_Bool_6QNode_Bool_1t1a8U_1lizzieLet20_1_4QNode_Bool_7QNode_Bool_1t2a8V_1lizzieLet20_1_4QNode_Bool_8QNode_Bool_1t3a8W_1Lcall_f'3_bufchan_buf [0])))
        \lizzieLet20_1_4QNode_Bool_5QNode_Bool_1lizzieLet20_1_4QNode_Bool_6QNode_Bool_1t1a8U_1lizzieLet20_1_4QNode_Bool_7QNode_Bool_1t2a8V_1lizzieLet20_1_4QNode_Bool_8QNode_Bool_1t3a8W_1Lcall_f'3_bufchan_buf  <= \lizzieLet20_1_4QNode_Bool_5QNode_Bool_1lizzieLet20_1_4QNode_Bool_6QNode_Bool_1t1a8U_1lizzieLet20_1_4QNode_Bool_7QNode_Bool_1t2a8V_1lizzieLet20_1_4QNode_Bool_8QNode_Bool_1t3a8W_1Lcall_f'3_bufchan_d ;
  
  /* buf (Ty Pointer_CTf') : (lizzieLet20_1_4QNode_Bool_5QNone_Bool,Pointer_CTf') > (lizzieLet20_1_4QNode_Bool_5QNone_Bool_1_argbuf,Pointer_CTf') */
  \Pointer_CTf'_t  lizzieLet20_1_4QNode_Bool_5QNone_Bool_bufchan_d;
  logic lizzieLet20_1_4QNode_Bool_5QNone_Bool_bufchan_r;
  assign lizzieLet20_1_4QNode_Bool_5QNone_Bool_r = ((! lizzieLet20_1_4QNode_Bool_5QNone_Bool_bufchan_d[0]) || lizzieLet20_1_4QNode_Bool_5QNone_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet20_1_4QNode_Bool_5QNone_Bool_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet20_1_4QNode_Bool_5QNone_Bool_r)
        lizzieLet20_1_4QNode_Bool_5QNone_Bool_bufchan_d <= lizzieLet20_1_4QNode_Bool_5QNone_Bool_d;
  \Pointer_CTf'_t  lizzieLet20_1_4QNode_Bool_5QNone_Bool_bufchan_buf;
  assign lizzieLet20_1_4QNode_Bool_5QNone_Bool_bufchan_r = (! lizzieLet20_1_4QNode_Bool_5QNone_Bool_bufchan_buf[0]);
  assign lizzieLet20_1_4QNode_Bool_5QNone_Bool_1_argbuf_d = (lizzieLet20_1_4QNode_Bool_5QNone_Bool_bufchan_buf[0] ? lizzieLet20_1_4QNode_Bool_5QNone_Bool_bufchan_buf :
                                                             lizzieLet20_1_4QNode_Bool_5QNone_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet20_1_4QNode_Bool_5QNone_Bool_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet20_1_4QNode_Bool_5QNone_Bool_1_argbuf_r && lizzieLet20_1_4QNode_Bool_5QNone_Bool_bufchan_buf[0]))
        lizzieLet20_1_4QNode_Bool_5QNone_Bool_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet20_1_4QNode_Bool_5QNone_Bool_1_argbuf_r) && (! lizzieLet20_1_4QNode_Bool_5QNone_Bool_bufchan_buf[0])))
        lizzieLet20_1_4QNode_Bool_5QNone_Bool_bufchan_buf <= lizzieLet20_1_4QNode_Bool_5QNone_Bool_bufchan_d;
  
  /* buf (Ty Pointer_CTf') : (lizzieLet20_1_4QNode_Bool_5QVal_Bool,Pointer_CTf') > (lizzieLet20_1_4QNode_Bool_5QVal_Bool_1_argbuf,Pointer_CTf') */
  \Pointer_CTf'_t  lizzieLet20_1_4QNode_Bool_5QVal_Bool_bufchan_d;
  logic lizzieLet20_1_4QNode_Bool_5QVal_Bool_bufchan_r;
  assign lizzieLet20_1_4QNode_Bool_5QVal_Bool_r = ((! lizzieLet20_1_4QNode_Bool_5QVal_Bool_bufchan_d[0]) || lizzieLet20_1_4QNode_Bool_5QVal_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet20_1_4QNode_Bool_5QVal_Bool_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet20_1_4QNode_Bool_5QVal_Bool_r)
        lizzieLet20_1_4QNode_Bool_5QVal_Bool_bufchan_d <= lizzieLet20_1_4QNode_Bool_5QVal_Bool_d;
  \Pointer_CTf'_t  lizzieLet20_1_4QNode_Bool_5QVal_Bool_bufchan_buf;
  assign lizzieLet20_1_4QNode_Bool_5QVal_Bool_bufchan_r = (! lizzieLet20_1_4QNode_Bool_5QVal_Bool_bufchan_buf[0]);
  assign lizzieLet20_1_4QNode_Bool_5QVal_Bool_1_argbuf_d = (lizzieLet20_1_4QNode_Bool_5QVal_Bool_bufchan_buf[0] ? lizzieLet20_1_4QNode_Bool_5QVal_Bool_bufchan_buf :
                                                            lizzieLet20_1_4QNode_Bool_5QVal_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet20_1_4QNode_Bool_5QVal_Bool_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet20_1_4QNode_Bool_5QVal_Bool_1_argbuf_r && lizzieLet20_1_4QNode_Bool_5QVal_Bool_bufchan_buf[0]))
        lizzieLet20_1_4QNode_Bool_5QVal_Bool_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet20_1_4QNode_Bool_5QVal_Bool_1_argbuf_r) && (! lizzieLet20_1_4QNode_Bool_5QVal_Bool_bufchan_buf[0])))
        lizzieLet20_1_4QNode_Bool_5QVal_Bool_bufchan_buf <= lizzieLet20_1_4QNode_Bool_5QVal_Bool_bufchan_d;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_QTree_Bool) : (lizzieLet20_1_4QNode_Bool_6,QTree_Bool) (q1a8P_destruct,Pointer_QTree_Bool) > [(_53,Pointer_QTree_Bool),
                                                                                                                (_52,Pointer_QTree_Bool),
                                                                                                                (lizzieLet20_1_4QNode_Bool_6QNode_Bool,Pointer_QTree_Bool),
                                                                                                                (_51,Pointer_QTree_Bool)] */
  logic [3:0] q1a8P_destruct_onehotd;
  always_comb
    if ((lizzieLet20_1_4QNode_Bool_6_d[0] && q1a8P_destruct_d[0]))
      unique case (lizzieLet20_1_4QNode_Bool_6_d[2:1])
        2'd0: q1a8P_destruct_onehotd = 4'd1;
        2'd1: q1a8P_destruct_onehotd = 4'd2;
        2'd2: q1a8P_destruct_onehotd = 4'd4;
        2'd3: q1a8P_destruct_onehotd = 4'd8;
        default: q1a8P_destruct_onehotd = 4'd0;
      endcase
    else q1a8P_destruct_onehotd = 4'd0;
  assign _53_d = {q1a8P_destruct_d[16:1], q1a8P_destruct_onehotd[0]};
  assign _52_d = {q1a8P_destruct_d[16:1], q1a8P_destruct_onehotd[1]};
  assign lizzieLet20_1_4QNode_Bool_6QNode_Bool_d = {q1a8P_destruct_d[16:1],
                                                    q1a8P_destruct_onehotd[2]};
  assign _51_d = {q1a8P_destruct_d[16:1], q1a8P_destruct_onehotd[3]};
  assign q1a8P_destruct_r = (| (q1a8P_destruct_onehotd & {_51_r,
                                                          lizzieLet20_1_4QNode_Bool_6QNode_Bool_r,
                                                          _52_r,
                                                          _53_r}));
  assign lizzieLet20_1_4QNode_Bool_6_r = q1a8P_destruct_r;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_QTree_Bool) : (lizzieLet20_1_4QNode_Bool_7,QTree_Bool) (q2a8Q_destruct,Pointer_QTree_Bool) > [(_50,Pointer_QTree_Bool),
                                                                                                                (_49,Pointer_QTree_Bool),
                                                                                                                (lizzieLet20_1_4QNode_Bool_7QNode_Bool,Pointer_QTree_Bool),
                                                                                                                (_48,Pointer_QTree_Bool)] */
  logic [3:0] q2a8Q_destruct_onehotd;
  always_comb
    if ((lizzieLet20_1_4QNode_Bool_7_d[0] && q2a8Q_destruct_d[0]))
      unique case (lizzieLet20_1_4QNode_Bool_7_d[2:1])
        2'd0: q2a8Q_destruct_onehotd = 4'd1;
        2'd1: q2a8Q_destruct_onehotd = 4'd2;
        2'd2: q2a8Q_destruct_onehotd = 4'd4;
        2'd3: q2a8Q_destruct_onehotd = 4'd8;
        default: q2a8Q_destruct_onehotd = 4'd0;
      endcase
    else q2a8Q_destruct_onehotd = 4'd0;
  assign _50_d = {q2a8Q_destruct_d[16:1], q2a8Q_destruct_onehotd[0]};
  assign _49_d = {q2a8Q_destruct_d[16:1], q2a8Q_destruct_onehotd[1]};
  assign lizzieLet20_1_4QNode_Bool_7QNode_Bool_d = {q2a8Q_destruct_d[16:1],
                                                    q2a8Q_destruct_onehotd[2]};
  assign _48_d = {q2a8Q_destruct_d[16:1], q2a8Q_destruct_onehotd[3]};
  assign q2a8Q_destruct_r = (| (q2a8Q_destruct_onehotd & {_48_r,
                                                          lizzieLet20_1_4QNode_Bool_7QNode_Bool_r,
                                                          _49_r,
                                                          _50_r}));
  assign lizzieLet20_1_4QNode_Bool_7_r = q2a8Q_destruct_r;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_QTree_Bool) : (lizzieLet20_1_4QNode_Bool_8,QTree_Bool) (q3a8R_destruct,Pointer_QTree_Bool) > [(_47,Pointer_QTree_Bool),
                                                                                                                (_46,Pointer_QTree_Bool),
                                                                                                                (lizzieLet20_1_4QNode_Bool_8QNode_Bool,Pointer_QTree_Bool),
                                                                                                                (_45,Pointer_QTree_Bool)] */
  logic [3:0] q3a8R_destruct_onehotd;
  always_comb
    if ((lizzieLet20_1_4QNode_Bool_8_d[0] && q3a8R_destruct_d[0]))
      unique case (lizzieLet20_1_4QNode_Bool_8_d[2:1])
        2'd0: q3a8R_destruct_onehotd = 4'd1;
        2'd1: q3a8R_destruct_onehotd = 4'd2;
        2'd2: q3a8R_destruct_onehotd = 4'd4;
        2'd3: q3a8R_destruct_onehotd = 4'd8;
        default: q3a8R_destruct_onehotd = 4'd0;
      endcase
    else q3a8R_destruct_onehotd = 4'd0;
  assign _47_d = {q3a8R_destruct_d[16:1], q3a8R_destruct_onehotd[0]};
  assign _46_d = {q3a8R_destruct_d[16:1], q3a8R_destruct_onehotd[1]};
  assign lizzieLet20_1_4QNode_Bool_8QNode_Bool_d = {q3a8R_destruct_d[16:1],
                                                    q3a8R_destruct_onehotd[2]};
  assign _45_d = {q3a8R_destruct_d[16:1], q3a8R_destruct_onehotd[3]};
  assign q3a8R_destruct_r = (| (q3a8R_destruct_onehotd & {_45_r,
                                                          lizzieLet20_1_4QNode_Bool_8QNode_Bool_r,
                                                          _46_r,
                                                          _47_r}));
  assign lizzieLet20_1_4QNode_Bool_8_r = q3a8R_destruct_r;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_QTree_Bool) : (lizzieLet20_1_4QNode_Bool_9,QTree_Bool) (q4a8S_destruct,Pointer_QTree_Bool) > [(_44,Pointer_QTree_Bool),
                                                                                                                (_43,Pointer_QTree_Bool),
                                                                                                                (lizzieLet20_1_4QNode_Bool_9QNode_Bool,Pointer_QTree_Bool),
                                                                                                                (_42,Pointer_QTree_Bool)] */
  logic [3:0] q4a8S_destruct_onehotd;
  always_comb
    if ((lizzieLet20_1_4QNode_Bool_9_d[0] && q4a8S_destruct_d[0]))
      unique case (lizzieLet20_1_4QNode_Bool_9_d[2:1])
        2'd0: q4a8S_destruct_onehotd = 4'd1;
        2'd1: q4a8S_destruct_onehotd = 4'd2;
        2'd2: q4a8S_destruct_onehotd = 4'd4;
        2'd3: q4a8S_destruct_onehotd = 4'd8;
        default: q4a8S_destruct_onehotd = 4'd0;
      endcase
    else q4a8S_destruct_onehotd = 4'd0;
  assign _44_d = {q4a8S_destruct_d[16:1], q4a8S_destruct_onehotd[0]};
  assign _43_d = {q4a8S_destruct_d[16:1], q4a8S_destruct_onehotd[1]};
  assign lizzieLet20_1_4QNode_Bool_9QNode_Bool_d = {q4a8S_destruct_d[16:1],
                                                    q4a8S_destruct_onehotd[2]};
  assign _42_d = {q4a8S_destruct_d[16:1], q4a8S_destruct_onehotd[3]};
  assign q4a8S_destruct_r = (| (q4a8S_destruct_onehotd & {_42_r,
                                                          lizzieLet20_1_4QNode_Bool_9QNode_Bool_r,
                                                          _43_r,
                                                          _44_r}));
  assign lizzieLet20_1_4QNode_Bool_9_r = q4a8S_destruct_r;
  
  /* buf (Ty Pointer_QTree_Bool) : (lizzieLet20_1_4QNode_Bool_9QNode_Bool,Pointer_QTree_Bool) > (lizzieLet20_1_4QNode_Bool_9QNode_Bool_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t lizzieLet20_1_4QNode_Bool_9QNode_Bool_bufchan_d;
  logic lizzieLet20_1_4QNode_Bool_9QNode_Bool_bufchan_r;
  assign lizzieLet20_1_4QNode_Bool_9QNode_Bool_r = ((! lizzieLet20_1_4QNode_Bool_9QNode_Bool_bufchan_d[0]) || lizzieLet20_1_4QNode_Bool_9QNode_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet20_1_4QNode_Bool_9QNode_Bool_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet20_1_4QNode_Bool_9QNode_Bool_r)
        lizzieLet20_1_4QNode_Bool_9QNode_Bool_bufchan_d <= lizzieLet20_1_4QNode_Bool_9QNode_Bool_d;
  Pointer_QTree_Bool_t lizzieLet20_1_4QNode_Bool_9QNode_Bool_bufchan_buf;
  assign lizzieLet20_1_4QNode_Bool_9QNode_Bool_bufchan_r = (! lizzieLet20_1_4QNode_Bool_9QNode_Bool_bufchan_buf[0]);
  assign lizzieLet20_1_4QNode_Bool_9QNode_Bool_1_argbuf_d = (lizzieLet20_1_4QNode_Bool_9QNode_Bool_bufchan_buf[0] ? lizzieLet20_1_4QNode_Bool_9QNode_Bool_bufchan_buf :
                                                             lizzieLet20_1_4QNode_Bool_9QNode_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet20_1_4QNode_Bool_9QNode_Bool_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet20_1_4QNode_Bool_9QNode_Bool_1_argbuf_r && lizzieLet20_1_4QNode_Bool_9QNode_Bool_bufchan_buf[0]))
        lizzieLet20_1_4QNode_Bool_9QNode_Bool_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet20_1_4QNode_Bool_9QNode_Bool_1_argbuf_r) && (! lizzieLet20_1_4QNode_Bool_9QNode_Bool_bufchan_buf[0])))
        lizzieLet20_1_4QNode_Bool_9QNode_Bool_bufchan_buf <= lizzieLet20_1_4QNode_Bool_9QNode_Bool_bufchan_d;
  
  /* fork (Ty QTree_Bool) : (lizzieLet20_1_4QVal_Bool,QTree_Bool) > [(lizzieLet20_1_4QVal_Bool_1,QTree_Bool),
                                                                (lizzieLet20_1_4QVal_Bool_2,QTree_Bool),
                                                                (lizzieLet20_1_4QVal_Bool_3,QTree_Bool),
                                                                (lizzieLet20_1_4QVal_Bool_4,QTree_Bool),
                                                                (lizzieLet20_1_4QVal_Bool_5,QTree_Bool),
                                                                (lizzieLet20_1_4QVal_Bool_6,QTree_Bool)] */
  logic [5:0] lizzieLet20_1_4QVal_Bool_emitted;
  logic [5:0] lizzieLet20_1_4QVal_Bool_done;
  assign lizzieLet20_1_4QVal_Bool_1_d = {lizzieLet20_1_4QVal_Bool_d[66:1],
                                         (lizzieLet20_1_4QVal_Bool_d[0] && (! lizzieLet20_1_4QVal_Bool_emitted[0]))};
  assign lizzieLet20_1_4QVal_Bool_2_d = {lizzieLet20_1_4QVal_Bool_d[66:1],
                                         (lizzieLet20_1_4QVal_Bool_d[0] && (! lizzieLet20_1_4QVal_Bool_emitted[1]))};
  assign lizzieLet20_1_4QVal_Bool_3_d = {lizzieLet20_1_4QVal_Bool_d[66:1],
                                         (lizzieLet20_1_4QVal_Bool_d[0] && (! lizzieLet20_1_4QVal_Bool_emitted[2]))};
  assign lizzieLet20_1_4QVal_Bool_4_d = {lizzieLet20_1_4QVal_Bool_d[66:1],
                                         (lizzieLet20_1_4QVal_Bool_d[0] && (! lizzieLet20_1_4QVal_Bool_emitted[3]))};
  assign lizzieLet20_1_4QVal_Bool_5_d = {lizzieLet20_1_4QVal_Bool_d[66:1],
                                         (lizzieLet20_1_4QVal_Bool_d[0] && (! lizzieLet20_1_4QVal_Bool_emitted[4]))};
  assign lizzieLet20_1_4QVal_Bool_6_d = {lizzieLet20_1_4QVal_Bool_d[66:1],
                                         (lizzieLet20_1_4QVal_Bool_d[0] && (! lizzieLet20_1_4QVal_Bool_emitted[5]))};
  assign lizzieLet20_1_4QVal_Bool_done = (lizzieLet20_1_4QVal_Bool_emitted | ({lizzieLet20_1_4QVal_Bool_6_d[0],
                                                                               lizzieLet20_1_4QVal_Bool_5_d[0],
                                                                               lizzieLet20_1_4QVal_Bool_4_d[0],
                                                                               lizzieLet20_1_4QVal_Bool_3_d[0],
                                                                               lizzieLet20_1_4QVal_Bool_2_d[0],
                                                                               lizzieLet20_1_4QVal_Bool_1_d[0]} & {lizzieLet20_1_4QVal_Bool_6_r,
                                                                                                                   lizzieLet20_1_4QVal_Bool_5_r,
                                                                                                                   lizzieLet20_1_4QVal_Bool_4_r,
                                                                                                                   lizzieLet20_1_4QVal_Bool_3_r,
                                                                                                                   lizzieLet20_1_4QVal_Bool_2_r,
                                                                                                                   lizzieLet20_1_4QVal_Bool_1_r}));
  assign lizzieLet20_1_4QVal_Bool_r = (& lizzieLet20_1_4QVal_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet20_1_4QVal_Bool_emitted <= 6'd0;
    else
      lizzieLet20_1_4QVal_Bool_emitted <= (lizzieLet20_1_4QVal_Bool_r ? 6'd0 :
                                           lizzieLet20_1_4QVal_Bool_done);
  
  /* destruct (Ty QTree_Bool,
          Dcon QVal_Bool) : (lizzieLet20_1_4QVal_Bool_1QVal_Bool,QTree_Bool) > [(va8K_destruct,MyBool)] */
  assign va8K_destruct_d = {lizzieLet20_1_4QVal_Bool_1QVal_Bool_d[3:3],
                            lizzieLet20_1_4QVal_Bool_1QVal_Bool_d[0]};
  assign lizzieLet20_1_4QVal_Bool_1QVal_Bool_r = va8K_destruct_r;
  
  /* demux (Ty QTree_Bool,
       Ty QTree_Bool) : (lizzieLet20_1_4QVal_Bool_2,QTree_Bool) (lizzieLet20_1_4QVal_Bool_1,QTree_Bool) > [(_41,QTree_Bool),
                                                                                                           (lizzieLet20_1_4QVal_Bool_1QVal_Bool,QTree_Bool),
                                                                                                           (_40,QTree_Bool),
                                                                                                           (_39,QTree_Bool)] */
  logic [3:0] lizzieLet20_1_4QVal_Bool_1_onehotd;
  always_comb
    if ((lizzieLet20_1_4QVal_Bool_2_d[0] && lizzieLet20_1_4QVal_Bool_1_d[0]))
      unique case (lizzieLet20_1_4QVal_Bool_2_d[2:1])
        2'd0: lizzieLet20_1_4QVal_Bool_1_onehotd = 4'd1;
        2'd1: lizzieLet20_1_4QVal_Bool_1_onehotd = 4'd2;
        2'd2: lizzieLet20_1_4QVal_Bool_1_onehotd = 4'd4;
        2'd3: lizzieLet20_1_4QVal_Bool_1_onehotd = 4'd8;
        default: lizzieLet20_1_4QVal_Bool_1_onehotd = 4'd0;
      endcase
    else lizzieLet20_1_4QVal_Bool_1_onehotd = 4'd0;
  assign _41_d = {lizzieLet20_1_4QVal_Bool_1_d[66:1],
                  lizzieLet20_1_4QVal_Bool_1_onehotd[0]};
  assign lizzieLet20_1_4QVal_Bool_1QVal_Bool_d = {lizzieLet20_1_4QVal_Bool_1_d[66:1],
                                                  lizzieLet20_1_4QVal_Bool_1_onehotd[1]};
  assign _40_d = {lizzieLet20_1_4QVal_Bool_1_d[66:1],
                  lizzieLet20_1_4QVal_Bool_1_onehotd[2]};
  assign _39_d = {lizzieLet20_1_4QVal_Bool_1_d[66:1],
                  lizzieLet20_1_4QVal_Bool_1_onehotd[3]};
  assign lizzieLet20_1_4QVal_Bool_1_r = (| (lizzieLet20_1_4QVal_Bool_1_onehotd & {_39_r,
                                                                                  _40_r,
                                                                                  lizzieLet20_1_4QVal_Bool_1QVal_Bool_r,
                                                                                  _41_r}));
  assign lizzieLet20_1_4QVal_Bool_2_r = lizzieLet20_1_4QVal_Bool_1_r;
  
  /* demux (Ty QTree_Bool,
       Ty Go) : (lizzieLet20_1_4QVal_Bool_3,QTree_Bool) (lizzieLet20_1_3QVal_Bool,Go) > [(lizzieLet20_1_4QVal_Bool_3QNone_Bool,Go),
                                                                                         (lizzieLet20_1_4QVal_Bool_3QVal_Bool,Go),
                                                                                         (lizzieLet20_1_4QVal_Bool_3QNode_Bool,Go),
                                                                                         (lizzieLet20_1_4QVal_Bool_3QError_Bool,Go)] */
  logic [3:0] lizzieLet20_1_3QVal_Bool_onehotd;
  always_comb
    if ((lizzieLet20_1_4QVal_Bool_3_d[0] && lizzieLet20_1_3QVal_Bool_d[0]))
      unique case (lizzieLet20_1_4QVal_Bool_3_d[2:1])
        2'd0: lizzieLet20_1_3QVal_Bool_onehotd = 4'd1;
        2'd1: lizzieLet20_1_3QVal_Bool_onehotd = 4'd2;
        2'd2: lizzieLet20_1_3QVal_Bool_onehotd = 4'd4;
        2'd3: lizzieLet20_1_3QVal_Bool_onehotd = 4'd8;
        default: lizzieLet20_1_3QVal_Bool_onehotd = 4'd0;
      endcase
    else lizzieLet20_1_3QVal_Bool_onehotd = 4'd0;
  assign lizzieLet20_1_4QVal_Bool_3QNone_Bool_d = lizzieLet20_1_3QVal_Bool_onehotd[0];
  assign lizzieLet20_1_4QVal_Bool_3QVal_Bool_d = lizzieLet20_1_3QVal_Bool_onehotd[1];
  assign lizzieLet20_1_4QVal_Bool_3QNode_Bool_d = lizzieLet20_1_3QVal_Bool_onehotd[2];
  assign lizzieLet20_1_4QVal_Bool_3QError_Bool_d = lizzieLet20_1_3QVal_Bool_onehotd[3];
  assign lizzieLet20_1_3QVal_Bool_r = (| (lizzieLet20_1_3QVal_Bool_onehotd & {lizzieLet20_1_4QVal_Bool_3QError_Bool_r,
                                                                              lizzieLet20_1_4QVal_Bool_3QNode_Bool_r,
                                                                              lizzieLet20_1_4QVal_Bool_3QVal_Bool_r,
                                                                              lizzieLet20_1_4QVal_Bool_3QNone_Bool_r}));
  assign lizzieLet20_1_4QVal_Bool_3_r = lizzieLet20_1_3QVal_Bool_r;
  
  /* fork (Ty Go) : (lizzieLet20_1_4QVal_Bool_3QError_Bool,Go) > [(lizzieLet20_1_4QVal_Bool_3QError_Bool_1,Go),
                                                             (lizzieLet20_1_4QVal_Bool_3QError_Bool_2,Go)] */
  logic [1:0] lizzieLet20_1_4QVal_Bool_3QError_Bool_emitted;
  logic [1:0] lizzieLet20_1_4QVal_Bool_3QError_Bool_done;
  assign lizzieLet20_1_4QVal_Bool_3QError_Bool_1_d = (lizzieLet20_1_4QVal_Bool_3QError_Bool_d[0] && (! lizzieLet20_1_4QVal_Bool_3QError_Bool_emitted[0]));
  assign lizzieLet20_1_4QVal_Bool_3QError_Bool_2_d = (lizzieLet20_1_4QVal_Bool_3QError_Bool_d[0] && (! lizzieLet20_1_4QVal_Bool_3QError_Bool_emitted[1]));
  assign lizzieLet20_1_4QVal_Bool_3QError_Bool_done = (lizzieLet20_1_4QVal_Bool_3QError_Bool_emitted | ({lizzieLet20_1_4QVal_Bool_3QError_Bool_2_d[0],
                                                                                                         lizzieLet20_1_4QVal_Bool_3QError_Bool_1_d[0]} & {lizzieLet20_1_4QVal_Bool_3QError_Bool_2_r,
                                                                                                                                                          lizzieLet20_1_4QVal_Bool_3QError_Bool_1_r}));
  assign lizzieLet20_1_4QVal_Bool_3QError_Bool_r = (& lizzieLet20_1_4QVal_Bool_3QError_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet20_1_4QVal_Bool_3QError_Bool_emitted <= 2'd0;
    else
      lizzieLet20_1_4QVal_Bool_3QError_Bool_emitted <= (lizzieLet20_1_4QVal_Bool_3QError_Bool_r ? 2'd0 :
                                                        lizzieLet20_1_4QVal_Bool_3QError_Bool_done);
  
  /* dcon (Ty QTree_Bool,
      Dcon QError_Bool) : [(lizzieLet20_1_4QVal_Bool_3QError_Bool_1,Go)] > (lizzieLet20_1_4QVal_Bool_3QError_Bool_1QError_Bool,QTree_Bool) */
  assign lizzieLet20_1_4QVal_Bool_3QError_Bool_1QError_Bool_d = QError_Bool_dc((& {lizzieLet20_1_4QVal_Bool_3QError_Bool_1_d[0]}), lizzieLet20_1_4QVal_Bool_3QError_Bool_1_d);
  assign {lizzieLet20_1_4QVal_Bool_3QError_Bool_1_r} = {1 {(lizzieLet20_1_4QVal_Bool_3QError_Bool_1QError_Bool_r && lizzieLet20_1_4QVal_Bool_3QError_Bool_1QError_Bool_d[0])}};
  
  /* buf (Ty QTree_Bool) : (lizzieLet20_1_4QVal_Bool_3QError_Bool_1QError_Bool,QTree_Bool) > (lizzieLet26_1_1_argbuf,QTree_Bool) */
  QTree_Bool_t lizzieLet20_1_4QVal_Bool_3QError_Bool_1QError_Bool_bufchan_d;
  logic lizzieLet20_1_4QVal_Bool_3QError_Bool_1QError_Bool_bufchan_r;
  assign lizzieLet20_1_4QVal_Bool_3QError_Bool_1QError_Bool_r = ((! lizzieLet20_1_4QVal_Bool_3QError_Bool_1QError_Bool_bufchan_d[0]) || lizzieLet20_1_4QVal_Bool_3QError_Bool_1QError_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet20_1_4QVal_Bool_3QError_Bool_1QError_Bool_bufchan_d <= {66'd0,
                                                                       1'd0};
    else
      if (lizzieLet20_1_4QVal_Bool_3QError_Bool_1QError_Bool_r)
        lizzieLet20_1_4QVal_Bool_3QError_Bool_1QError_Bool_bufchan_d <= lizzieLet20_1_4QVal_Bool_3QError_Bool_1QError_Bool_d;
  QTree_Bool_t lizzieLet20_1_4QVal_Bool_3QError_Bool_1QError_Bool_bufchan_buf;
  assign lizzieLet20_1_4QVal_Bool_3QError_Bool_1QError_Bool_bufchan_r = (! lizzieLet20_1_4QVal_Bool_3QError_Bool_1QError_Bool_bufchan_buf[0]);
  assign lizzieLet26_1_1_argbuf_d = (lizzieLet20_1_4QVal_Bool_3QError_Bool_1QError_Bool_bufchan_buf[0] ? lizzieLet20_1_4QVal_Bool_3QError_Bool_1QError_Bool_bufchan_buf :
                                     lizzieLet20_1_4QVal_Bool_3QError_Bool_1QError_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet20_1_4QVal_Bool_3QError_Bool_1QError_Bool_bufchan_buf <= {66'd0,
                                                                         1'd0};
    else
      if ((lizzieLet26_1_1_argbuf_r && lizzieLet20_1_4QVal_Bool_3QError_Bool_1QError_Bool_bufchan_buf[0]))
        lizzieLet20_1_4QVal_Bool_3QError_Bool_1QError_Bool_bufchan_buf <= {66'd0,
                                                                           1'd0};
      else if (((! lizzieLet26_1_1_argbuf_r) && (! lizzieLet20_1_4QVal_Bool_3QError_Bool_1QError_Bool_bufchan_buf[0])))
        lizzieLet20_1_4QVal_Bool_3QError_Bool_1QError_Bool_bufchan_buf <= lizzieLet20_1_4QVal_Bool_3QError_Bool_1QError_Bool_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet20_1_4QVal_Bool_3QError_Bool_2,Go) > (lizzieLet20_1_4QVal_Bool_3QError_Bool_2_argbuf,Go) */
  Go_t lizzieLet20_1_4QVal_Bool_3QError_Bool_2_bufchan_d;
  logic lizzieLet20_1_4QVal_Bool_3QError_Bool_2_bufchan_r;
  assign lizzieLet20_1_4QVal_Bool_3QError_Bool_2_r = ((! lizzieLet20_1_4QVal_Bool_3QError_Bool_2_bufchan_d[0]) || lizzieLet20_1_4QVal_Bool_3QError_Bool_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet20_1_4QVal_Bool_3QError_Bool_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet20_1_4QVal_Bool_3QError_Bool_2_r)
        lizzieLet20_1_4QVal_Bool_3QError_Bool_2_bufchan_d <= lizzieLet20_1_4QVal_Bool_3QError_Bool_2_d;
  Go_t lizzieLet20_1_4QVal_Bool_3QError_Bool_2_bufchan_buf;
  assign lizzieLet20_1_4QVal_Bool_3QError_Bool_2_bufchan_r = (! lizzieLet20_1_4QVal_Bool_3QError_Bool_2_bufchan_buf[0]);
  assign lizzieLet20_1_4QVal_Bool_3QError_Bool_2_argbuf_d = (lizzieLet20_1_4QVal_Bool_3QError_Bool_2_bufchan_buf[0] ? lizzieLet20_1_4QVal_Bool_3QError_Bool_2_bufchan_buf :
                                                             lizzieLet20_1_4QVal_Bool_3QError_Bool_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet20_1_4QVal_Bool_3QError_Bool_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet20_1_4QVal_Bool_3QError_Bool_2_argbuf_r && lizzieLet20_1_4QVal_Bool_3QError_Bool_2_bufchan_buf[0]))
        lizzieLet20_1_4QVal_Bool_3QError_Bool_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet20_1_4QVal_Bool_3QError_Bool_2_argbuf_r) && (! lizzieLet20_1_4QVal_Bool_3QError_Bool_2_bufchan_buf[0])))
        lizzieLet20_1_4QVal_Bool_3QError_Bool_2_bufchan_buf <= lizzieLet20_1_4QVal_Bool_3QError_Bool_2_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet20_1_4QVal_Bool_3QNode_Bool,Go) > [(lizzieLet20_1_4QVal_Bool_3QNode_Bool_1,Go),
                                                            (lizzieLet20_1_4QVal_Bool_3QNode_Bool_2,Go)] */
  logic [1:0] lizzieLet20_1_4QVal_Bool_3QNode_Bool_emitted;
  logic [1:0] lizzieLet20_1_4QVal_Bool_3QNode_Bool_done;
  assign lizzieLet20_1_4QVal_Bool_3QNode_Bool_1_d = (lizzieLet20_1_4QVal_Bool_3QNode_Bool_d[0] && (! lizzieLet20_1_4QVal_Bool_3QNode_Bool_emitted[0]));
  assign lizzieLet20_1_4QVal_Bool_3QNode_Bool_2_d = (lizzieLet20_1_4QVal_Bool_3QNode_Bool_d[0] && (! lizzieLet20_1_4QVal_Bool_3QNode_Bool_emitted[1]));
  assign lizzieLet20_1_4QVal_Bool_3QNode_Bool_done = (lizzieLet20_1_4QVal_Bool_3QNode_Bool_emitted | ({lizzieLet20_1_4QVal_Bool_3QNode_Bool_2_d[0],
                                                                                                       lizzieLet20_1_4QVal_Bool_3QNode_Bool_1_d[0]} & {lizzieLet20_1_4QVal_Bool_3QNode_Bool_2_r,
                                                                                                                                                       lizzieLet20_1_4QVal_Bool_3QNode_Bool_1_r}));
  assign lizzieLet20_1_4QVal_Bool_3QNode_Bool_r = (& lizzieLet20_1_4QVal_Bool_3QNode_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet20_1_4QVal_Bool_3QNode_Bool_emitted <= 2'd0;
    else
      lizzieLet20_1_4QVal_Bool_3QNode_Bool_emitted <= (lizzieLet20_1_4QVal_Bool_3QNode_Bool_r ? 2'd0 :
                                                       lizzieLet20_1_4QVal_Bool_3QNode_Bool_done);
  
  /* dcon (Ty QTree_Bool,
      Dcon QError_Bool) : [(lizzieLet20_1_4QVal_Bool_3QNode_Bool_1,Go)] > (lizzieLet20_1_4QVal_Bool_3QNode_Bool_1QError_Bool,QTree_Bool) */
  assign lizzieLet20_1_4QVal_Bool_3QNode_Bool_1QError_Bool_d = QError_Bool_dc((& {lizzieLet20_1_4QVal_Bool_3QNode_Bool_1_d[0]}), lizzieLet20_1_4QVal_Bool_3QNode_Bool_1_d);
  assign {lizzieLet20_1_4QVal_Bool_3QNode_Bool_1_r} = {1 {(lizzieLet20_1_4QVal_Bool_3QNode_Bool_1QError_Bool_r && lizzieLet20_1_4QVal_Bool_3QNode_Bool_1QError_Bool_d[0])}};
  
  /* buf (Ty QTree_Bool) : (lizzieLet20_1_4QVal_Bool_3QNode_Bool_1QError_Bool,QTree_Bool) > (lizzieLet25_1_1_argbuf,QTree_Bool) */
  QTree_Bool_t lizzieLet20_1_4QVal_Bool_3QNode_Bool_1QError_Bool_bufchan_d;
  logic lizzieLet20_1_4QVal_Bool_3QNode_Bool_1QError_Bool_bufchan_r;
  assign lizzieLet20_1_4QVal_Bool_3QNode_Bool_1QError_Bool_r = ((! lizzieLet20_1_4QVal_Bool_3QNode_Bool_1QError_Bool_bufchan_d[0]) || lizzieLet20_1_4QVal_Bool_3QNode_Bool_1QError_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet20_1_4QVal_Bool_3QNode_Bool_1QError_Bool_bufchan_d <= {66'd0,
                                                                      1'd0};
    else
      if (lizzieLet20_1_4QVal_Bool_3QNode_Bool_1QError_Bool_r)
        lizzieLet20_1_4QVal_Bool_3QNode_Bool_1QError_Bool_bufchan_d <= lizzieLet20_1_4QVal_Bool_3QNode_Bool_1QError_Bool_d;
  QTree_Bool_t lizzieLet20_1_4QVal_Bool_3QNode_Bool_1QError_Bool_bufchan_buf;
  assign lizzieLet20_1_4QVal_Bool_3QNode_Bool_1QError_Bool_bufchan_r = (! lizzieLet20_1_4QVal_Bool_3QNode_Bool_1QError_Bool_bufchan_buf[0]);
  assign lizzieLet25_1_1_argbuf_d = (lizzieLet20_1_4QVal_Bool_3QNode_Bool_1QError_Bool_bufchan_buf[0] ? lizzieLet20_1_4QVal_Bool_3QNode_Bool_1QError_Bool_bufchan_buf :
                                     lizzieLet20_1_4QVal_Bool_3QNode_Bool_1QError_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet20_1_4QVal_Bool_3QNode_Bool_1QError_Bool_bufchan_buf <= {66'd0,
                                                                        1'd0};
    else
      if ((lizzieLet25_1_1_argbuf_r && lizzieLet20_1_4QVal_Bool_3QNode_Bool_1QError_Bool_bufchan_buf[0]))
        lizzieLet20_1_4QVal_Bool_3QNode_Bool_1QError_Bool_bufchan_buf <= {66'd0,
                                                                          1'd0};
      else if (((! lizzieLet25_1_1_argbuf_r) && (! lizzieLet20_1_4QVal_Bool_3QNode_Bool_1QError_Bool_bufchan_buf[0])))
        lizzieLet20_1_4QVal_Bool_3QNode_Bool_1QError_Bool_bufchan_buf <= lizzieLet20_1_4QVal_Bool_3QNode_Bool_1QError_Bool_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet20_1_4QVal_Bool_3QNode_Bool_2,Go) > (lizzieLet20_1_4QVal_Bool_3QNode_Bool_2_argbuf,Go) */
  Go_t lizzieLet20_1_4QVal_Bool_3QNode_Bool_2_bufchan_d;
  logic lizzieLet20_1_4QVal_Bool_3QNode_Bool_2_bufchan_r;
  assign lizzieLet20_1_4QVal_Bool_3QNode_Bool_2_r = ((! lizzieLet20_1_4QVal_Bool_3QNode_Bool_2_bufchan_d[0]) || lizzieLet20_1_4QVal_Bool_3QNode_Bool_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet20_1_4QVal_Bool_3QNode_Bool_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet20_1_4QVal_Bool_3QNode_Bool_2_r)
        lizzieLet20_1_4QVal_Bool_3QNode_Bool_2_bufchan_d <= lizzieLet20_1_4QVal_Bool_3QNode_Bool_2_d;
  Go_t lizzieLet20_1_4QVal_Bool_3QNode_Bool_2_bufchan_buf;
  assign lizzieLet20_1_4QVal_Bool_3QNode_Bool_2_bufchan_r = (! lizzieLet20_1_4QVal_Bool_3QNode_Bool_2_bufchan_buf[0]);
  assign lizzieLet20_1_4QVal_Bool_3QNode_Bool_2_argbuf_d = (lizzieLet20_1_4QVal_Bool_3QNode_Bool_2_bufchan_buf[0] ? lizzieLet20_1_4QVal_Bool_3QNode_Bool_2_bufchan_buf :
                                                            lizzieLet20_1_4QVal_Bool_3QNode_Bool_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet20_1_4QVal_Bool_3QNode_Bool_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet20_1_4QVal_Bool_3QNode_Bool_2_argbuf_r && lizzieLet20_1_4QVal_Bool_3QNode_Bool_2_bufchan_buf[0]))
        lizzieLet20_1_4QVal_Bool_3QNode_Bool_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet20_1_4QVal_Bool_3QNode_Bool_2_argbuf_r) && (! lizzieLet20_1_4QVal_Bool_3QNode_Bool_2_bufchan_buf[0])))
        lizzieLet20_1_4QVal_Bool_3QNode_Bool_2_bufchan_buf <= lizzieLet20_1_4QVal_Bool_3QNode_Bool_2_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet20_1_4QVal_Bool_3QNone_Bool,Go) > (lizzieLet20_1_4QVal_Bool_3QNone_Bool_1_argbuf,Go) */
  Go_t lizzieLet20_1_4QVal_Bool_3QNone_Bool_bufchan_d;
  logic lizzieLet20_1_4QVal_Bool_3QNone_Bool_bufchan_r;
  assign lizzieLet20_1_4QVal_Bool_3QNone_Bool_r = ((! lizzieLet20_1_4QVal_Bool_3QNone_Bool_bufchan_d[0]) || lizzieLet20_1_4QVal_Bool_3QNone_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet20_1_4QVal_Bool_3QNone_Bool_bufchan_d <= 1'd0;
    else
      if (lizzieLet20_1_4QVal_Bool_3QNone_Bool_r)
        lizzieLet20_1_4QVal_Bool_3QNone_Bool_bufchan_d <= lizzieLet20_1_4QVal_Bool_3QNone_Bool_d;
  Go_t lizzieLet20_1_4QVal_Bool_3QNone_Bool_bufchan_buf;
  assign lizzieLet20_1_4QVal_Bool_3QNone_Bool_bufchan_r = (! lizzieLet20_1_4QVal_Bool_3QNone_Bool_bufchan_buf[0]);
  assign lizzieLet20_1_4QVal_Bool_3QNone_Bool_1_argbuf_d = (lizzieLet20_1_4QVal_Bool_3QNone_Bool_bufchan_buf[0] ? lizzieLet20_1_4QVal_Bool_3QNone_Bool_bufchan_buf :
                                                            lizzieLet20_1_4QVal_Bool_3QNone_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet20_1_4QVal_Bool_3QNone_Bool_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet20_1_4QVal_Bool_3QNone_Bool_1_argbuf_r && lizzieLet20_1_4QVal_Bool_3QNone_Bool_bufchan_buf[0]))
        lizzieLet20_1_4QVal_Bool_3QNone_Bool_bufchan_buf <= 1'd0;
      else if (((! lizzieLet20_1_4QVal_Bool_3QNone_Bool_1_argbuf_r) && (! lizzieLet20_1_4QVal_Bool_3QNone_Bool_bufchan_buf[0])))
        lizzieLet20_1_4QVal_Bool_3QNone_Bool_bufchan_buf <= lizzieLet20_1_4QVal_Bool_3QNone_Bool_bufchan_d;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_QTree_Bool) : (lizzieLet20_1_4QVal_Bool_4,QTree_Bool) (lizzieLet20_1_5QVal_Bool,Pointer_QTree_Bool) > [(lizzieLet20_1_4QVal_Bool_4QNone_Bool,Pointer_QTree_Bool),
                                                                                                                         (_38,Pointer_QTree_Bool),
                                                                                                                         (_37,Pointer_QTree_Bool),
                                                                                                                         (_36,Pointer_QTree_Bool)] */
  logic [3:0] lizzieLet20_1_5QVal_Bool_onehotd;
  always_comb
    if ((lizzieLet20_1_4QVal_Bool_4_d[0] && lizzieLet20_1_5QVal_Bool_d[0]))
      unique case (lizzieLet20_1_4QVal_Bool_4_d[2:1])
        2'd0: lizzieLet20_1_5QVal_Bool_onehotd = 4'd1;
        2'd1: lizzieLet20_1_5QVal_Bool_onehotd = 4'd2;
        2'd2: lizzieLet20_1_5QVal_Bool_onehotd = 4'd4;
        2'd3: lizzieLet20_1_5QVal_Bool_onehotd = 4'd8;
        default: lizzieLet20_1_5QVal_Bool_onehotd = 4'd0;
      endcase
    else lizzieLet20_1_5QVal_Bool_onehotd = 4'd0;
  assign lizzieLet20_1_4QVal_Bool_4QNone_Bool_d = {lizzieLet20_1_5QVal_Bool_d[16:1],
                                                   lizzieLet20_1_5QVal_Bool_onehotd[0]};
  assign _38_d = {lizzieLet20_1_5QVal_Bool_d[16:1],
                  lizzieLet20_1_5QVal_Bool_onehotd[1]};
  assign _37_d = {lizzieLet20_1_5QVal_Bool_d[16:1],
                  lizzieLet20_1_5QVal_Bool_onehotd[2]};
  assign _36_d = {lizzieLet20_1_5QVal_Bool_d[16:1],
                  lizzieLet20_1_5QVal_Bool_onehotd[3]};
  assign lizzieLet20_1_5QVal_Bool_r = (| (lizzieLet20_1_5QVal_Bool_onehotd & {_36_r,
                                                                              _37_r,
                                                                              _38_r,
                                                                              lizzieLet20_1_4QVal_Bool_4QNone_Bool_r}));
  assign lizzieLet20_1_4QVal_Bool_4_r = lizzieLet20_1_5QVal_Bool_r;
  
  /* buf (Ty Pointer_QTree_Bool) : (lizzieLet20_1_4QVal_Bool_4QNone_Bool,Pointer_QTree_Bool) > (lizzieLet20_1_4QVal_Bool_4QNone_Bool_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t lizzieLet20_1_4QVal_Bool_4QNone_Bool_bufchan_d;
  logic lizzieLet20_1_4QVal_Bool_4QNone_Bool_bufchan_r;
  assign lizzieLet20_1_4QVal_Bool_4QNone_Bool_r = ((! lizzieLet20_1_4QVal_Bool_4QNone_Bool_bufchan_d[0]) || lizzieLet20_1_4QVal_Bool_4QNone_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet20_1_4QVal_Bool_4QNone_Bool_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet20_1_4QVal_Bool_4QNone_Bool_r)
        lizzieLet20_1_4QVal_Bool_4QNone_Bool_bufchan_d <= lizzieLet20_1_4QVal_Bool_4QNone_Bool_d;
  Pointer_QTree_Bool_t lizzieLet20_1_4QVal_Bool_4QNone_Bool_bufchan_buf;
  assign lizzieLet20_1_4QVal_Bool_4QNone_Bool_bufchan_r = (! lizzieLet20_1_4QVal_Bool_4QNone_Bool_bufchan_buf[0]);
  assign lizzieLet20_1_4QVal_Bool_4QNone_Bool_1_argbuf_d = (lizzieLet20_1_4QVal_Bool_4QNone_Bool_bufchan_buf[0] ? lizzieLet20_1_4QVal_Bool_4QNone_Bool_bufchan_buf :
                                                            lizzieLet20_1_4QVal_Bool_4QNone_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet20_1_4QVal_Bool_4QNone_Bool_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet20_1_4QVal_Bool_4QNone_Bool_1_argbuf_r && lizzieLet20_1_4QVal_Bool_4QNone_Bool_bufchan_buf[0]))
        lizzieLet20_1_4QVal_Bool_4QNone_Bool_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet20_1_4QVal_Bool_4QNone_Bool_1_argbuf_r) && (! lizzieLet20_1_4QVal_Bool_4QNone_Bool_bufchan_buf[0])))
        lizzieLet20_1_4QVal_Bool_4QNone_Bool_bufchan_buf <= lizzieLet20_1_4QVal_Bool_4QNone_Bool_bufchan_d;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_CTf') : (lizzieLet20_1_4QVal_Bool_5,QTree_Bool) (lizzieLet20_1_7QVal_Bool,Pointer_CTf') > [(lizzieLet20_1_4QVal_Bool_5QNone_Bool,Pointer_CTf'),
                                                                                                             (lizzieLet20_1_4QVal_Bool_5QVal_Bool,Pointer_CTf'),
                                                                                                             (lizzieLet20_1_4QVal_Bool_5QNode_Bool,Pointer_CTf'),
                                                                                                             (lizzieLet20_1_4QVal_Bool_5QError_Bool,Pointer_CTf')] */
  logic [3:0] lizzieLet20_1_7QVal_Bool_onehotd;
  always_comb
    if ((lizzieLet20_1_4QVal_Bool_5_d[0] && lizzieLet20_1_7QVal_Bool_d[0]))
      unique case (lizzieLet20_1_4QVal_Bool_5_d[2:1])
        2'd0: lizzieLet20_1_7QVal_Bool_onehotd = 4'd1;
        2'd1: lizzieLet20_1_7QVal_Bool_onehotd = 4'd2;
        2'd2: lizzieLet20_1_7QVal_Bool_onehotd = 4'd4;
        2'd3: lizzieLet20_1_7QVal_Bool_onehotd = 4'd8;
        default: lizzieLet20_1_7QVal_Bool_onehotd = 4'd0;
      endcase
    else lizzieLet20_1_7QVal_Bool_onehotd = 4'd0;
  assign lizzieLet20_1_4QVal_Bool_5QNone_Bool_d = {lizzieLet20_1_7QVal_Bool_d[16:1],
                                                   lizzieLet20_1_7QVal_Bool_onehotd[0]};
  assign lizzieLet20_1_4QVal_Bool_5QVal_Bool_d = {lizzieLet20_1_7QVal_Bool_d[16:1],
                                                  lizzieLet20_1_7QVal_Bool_onehotd[1]};
  assign lizzieLet20_1_4QVal_Bool_5QNode_Bool_d = {lizzieLet20_1_7QVal_Bool_d[16:1],
                                                   lizzieLet20_1_7QVal_Bool_onehotd[2]};
  assign lizzieLet20_1_4QVal_Bool_5QError_Bool_d = {lizzieLet20_1_7QVal_Bool_d[16:1],
                                                    lizzieLet20_1_7QVal_Bool_onehotd[3]};
  assign lizzieLet20_1_7QVal_Bool_r = (| (lizzieLet20_1_7QVal_Bool_onehotd & {lizzieLet20_1_4QVal_Bool_5QError_Bool_r,
                                                                              lizzieLet20_1_4QVal_Bool_5QNode_Bool_r,
                                                                              lizzieLet20_1_4QVal_Bool_5QVal_Bool_r,
                                                                              lizzieLet20_1_4QVal_Bool_5QNone_Bool_r}));
  assign lizzieLet20_1_4QVal_Bool_5_r = lizzieLet20_1_7QVal_Bool_r;
  
  /* buf (Ty Pointer_CTf') : (lizzieLet20_1_4QVal_Bool_5QError_Bool,Pointer_CTf') > (lizzieLet20_1_4QVal_Bool_5QError_Bool_1_argbuf,Pointer_CTf') */
  \Pointer_CTf'_t  lizzieLet20_1_4QVal_Bool_5QError_Bool_bufchan_d;
  logic lizzieLet20_1_4QVal_Bool_5QError_Bool_bufchan_r;
  assign lizzieLet20_1_4QVal_Bool_5QError_Bool_r = ((! lizzieLet20_1_4QVal_Bool_5QError_Bool_bufchan_d[0]) || lizzieLet20_1_4QVal_Bool_5QError_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet20_1_4QVal_Bool_5QError_Bool_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet20_1_4QVal_Bool_5QError_Bool_r)
        lizzieLet20_1_4QVal_Bool_5QError_Bool_bufchan_d <= lizzieLet20_1_4QVal_Bool_5QError_Bool_d;
  \Pointer_CTf'_t  lizzieLet20_1_4QVal_Bool_5QError_Bool_bufchan_buf;
  assign lizzieLet20_1_4QVal_Bool_5QError_Bool_bufchan_r = (! lizzieLet20_1_4QVal_Bool_5QError_Bool_bufchan_buf[0]);
  assign lizzieLet20_1_4QVal_Bool_5QError_Bool_1_argbuf_d = (lizzieLet20_1_4QVal_Bool_5QError_Bool_bufchan_buf[0] ? lizzieLet20_1_4QVal_Bool_5QError_Bool_bufchan_buf :
                                                             lizzieLet20_1_4QVal_Bool_5QError_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet20_1_4QVal_Bool_5QError_Bool_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet20_1_4QVal_Bool_5QError_Bool_1_argbuf_r && lizzieLet20_1_4QVal_Bool_5QError_Bool_bufchan_buf[0]))
        lizzieLet20_1_4QVal_Bool_5QError_Bool_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet20_1_4QVal_Bool_5QError_Bool_1_argbuf_r) && (! lizzieLet20_1_4QVal_Bool_5QError_Bool_bufchan_buf[0])))
        lizzieLet20_1_4QVal_Bool_5QError_Bool_bufchan_buf <= lizzieLet20_1_4QVal_Bool_5QError_Bool_bufchan_d;
  
  /* buf (Ty Pointer_CTf') : (lizzieLet20_1_4QVal_Bool_5QNode_Bool,Pointer_CTf') > (lizzieLet20_1_4QVal_Bool_5QNode_Bool_1_argbuf,Pointer_CTf') */
  \Pointer_CTf'_t  lizzieLet20_1_4QVal_Bool_5QNode_Bool_bufchan_d;
  logic lizzieLet20_1_4QVal_Bool_5QNode_Bool_bufchan_r;
  assign lizzieLet20_1_4QVal_Bool_5QNode_Bool_r = ((! lizzieLet20_1_4QVal_Bool_5QNode_Bool_bufchan_d[0]) || lizzieLet20_1_4QVal_Bool_5QNode_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet20_1_4QVal_Bool_5QNode_Bool_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet20_1_4QVal_Bool_5QNode_Bool_r)
        lizzieLet20_1_4QVal_Bool_5QNode_Bool_bufchan_d <= lizzieLet20_1_4QVal_Bool_5QNode_Bool_d;
  \Pointer_CTf'_t  lizzieLet20_1_4QVal_Bool_5QNode_Bool_bufchan_buf;
  assign lizzieLet20_1_4QVal_Bool_5QNode_Bool_bufchan_r = (! lizzieLet20_1_4QVal_Bool_5QNode_Bool_bufchan_buf[0]);
  assign lizzieLet20_1_4QVal_Bool_5QNode_Bool_1_argbuf_d = (lizzieLet20_1_4QVal_Bool_5QNode_Bool_bufchan_buf[0] ? lizzieLet20_1_4QVal_Bool_5QNode_Bool_bufchan_buf :
                                                            lizzieLet20_1_4QVal_Bool_5QNode_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet20_1_4QVal_Bool_5QNode_Bool_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet20_1_4QVal_Bool_5QNode_Bool_1_argbuf_r && lizzieLet20_1_4QVal_Bool_5QNode_Bool_bufchan_buf[0]))
        lizzieLet20_1_4QVal_Bool_5QNode_Bool_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet20_1_4QVal_Bool_5QNode_Bool_1_argbuf_r) && (! lizzieLet20_1_4QVal_Bool_5QNode_Bool_bufchan_buf[0])))
        lizzieLet20_1_4QVal_Bool_5QNode_Bool_bufchan_buf <= lizzieLet20_1_4QVal_Bool_5QNode_Bool_bufchan_d;
  
  /* buf (Ty Pointer_CTf') : (lizzieLet20_1_4QVal_Bool_5QNone_Bool,Pointer_CTf') > (lizzieLet20_1_4QVal_Bool_5QNone_Bool_1_argbuf,Pointer_CTf') */
  \Pointer_CTf'_t  lizzieLet20_1_4QVal_Bool_5QNone_Bool_bufchan_d;
  logic lizzieLet20_1_4QVal_Bool_5QNone_Bool_bufchan_r;
  assign lizzieLet20_1_4QVal_Bool_5QNone_Bool_r = ((! lizzieLet20_1_4QVal_Bool_5QNone_Bool_bufchan_d[0]) || lizzieLet20_1_4QVal_Bool_5QNone_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet20_1_4QVal_Bool_5QNone_Bool_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet20_1_4QVal_Bool_5QNone_Bool_r)
        lizzieLet20_1_4QVal_Bool_5QNone_Bool_bufchan_d <= lizzieLet20_1_4QVal_Bool_5QNone_Bool_d;
  \Pointer_CTf'_t  lizzieLet20_1_4QVal_Bool_5QNone_Bool_bufchan_buf;
  assign lizzieLet20_1_4QVal_Bool_5QNone_Bool_bufchan_r = (! lizzieLet20_1_4QVal_Bool_5QNone_Bool_bufchan_buf[0]);
  assign lizzieLet20_1_4QVal_Bool_5QNone_Bool_1_argbuf_d = (lizzieLet20_1_4QVal_Bool_5QNone_Bool_bufchan_buf[0] ? lizzieLet20_1_4QVal_Bool_5QNone_Bool_bufchan_buf :
                                                            lizzieLet20_1_4QVal_Bool_5QNone_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet20_1_4QVal_Bool_5QNone_Bool_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet20_1_4QVal_Bool_5QNone_Bool_1_argbuf_r && lizzieLet20_1_4QVal_Bool_5QNone_Bool_bufchan_buf[0]))
        lizzieLet20_1_4QVal_Bool_5QNone_Bool_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet20_1_4QVal_Bool_5QNone_Bool_1_argbuf_r) && (! lizzieLet20_1_4QVal_Bool_5QNone_Bool_bufchan_buf[0])))
        lizzieLet20_1_4QVal_Bool_5QNone_Bool_bufchan_buf <= lizzieLet20_1_4QVal_Bool_5QNone_Bool_bufchan_d;
  
  /* demux (Ty QTree_Bool,
       Ty MyBool) : (lizzieLet20_1_4QVal_Bool_6,QTree_Bool) (v1a8J_destruct,MyBool) > [(_35,MyBool),
                                                                                       (lizzieLet20_1_4QVal_Bool_6QVal_Bool,MyBool),
                                                                                       (_34,MyBool),
                                                                                       (_33,MyBool)] */
  logic [3:0] v1a8J_destruct_onehotd;
  always_comb
    if ((lizzieLet20_1_4QVal_Bool_6_d[0] && v1a8J_destruct_d[0]))
      unique case (lizzieLet20_1_4QVal_Bool_6_d[2:1])
        2'd0: v1a8J_destruct_onehotd = 4'd1;
        2'd1: v1a8J_destruct_onehotd = 4'd2;
        2'd2: v1a8J_destruct_onehotd = 4'd4;
        2'd3: v1a8J_destruct_onehotd = 4'd8;
        default: v1a8J_destruct_onehotd = 4'd0;
      endcase
    else v1a8J_destruct_onehotd = 4'd0;
  assign _35_d = {v1a8J_destruct_d[1:1], v1a8J_destruct_onehotd[0]};
  assign lizzieLet20_1_4QVal_Bool_6QVal_Bool_d = {v1a8J_destruct_d[1:1],
                                                  v1a8J_destruct_onehotd[1]};
  assign _34_d = {v1a8J_destruct_d[1:1], v1a8J_destruct_onehotd[2]};
  assign _33_d = {v1a8J_destruct_d[1:1], v1a8J_destruct_onehotd[3]};
  assign v1a8J_destruct_r = (| (v1a8J_destruct_onehotd & {_33_r,
                                                          _34_r,
                                                          lizzieLet20_1_4QVal_Bool_6QVal_Bool_r,
                                                          _35_r}));
  assign lizzieLet20_1_4QVal_Bool_6_r = v1a8J_destruct_r;
  
  /* fork (Ty MyBool) : (lizzieLet20_1_4QVal_Bool_6QVal_Bool,MyBool) > [(lizzieLet20_1_4QVal_Bool_6QVal_Bool_1,MyBool),
                                                                   (lizzieLet20_1_4QVal_Bool_6QVal_Bool_2,MyBool),
                                                                   (lizzieLet20_1_4QVal_Bool_6QVal_Bool_3,MyBool)] */
  logic [2:0] lizzieLet20_1_4QVal_Bool_6QVal_Bool_emitted;
  logic [2:0] lizzieLet20_1_4QVal_Bool_6QVal_Bool_done;
  assign lizzieLet20_1_4QVal_Bool_6QVal_Bool_1_d = {lizzieLet20_1_4QVal_Bool_6QVal_Bool_d[1:1],
                                                    (lizzieLet20_1_4QVal_Bool_6QVal_Bool_d[0] && (! lizzieLet20_1_4QVal_Bool_6QVal_Bool_emitted[0]))};
  assign lizzieLet20_1_4QVal_Bool_6QVal_Bool_2_d = {lizzieLet20_1_4QVal_Bool_6QVal_Bool_d[1:1],
                                                    (lizzieLet20_1_4QVal_Bool_6QVal_Bool_d[0] && (! lizzieLet20_1_4QVal_Bool_6QVal_Bool_emitted[1]))};
  assign lizzieLet20_1_4QVal_Bool_6QVal_Bool_3_d = {lizzieLet20_1_4QVal_Bool_6QVal_Bool_d[1:1],
                                                    (lizzieLet20_1_4QVal_Bool_6QVal_Bool_d[0] && (! lizzieLet20_1_4QVal_Bool_6QVal_Bool_emitted[2]))};
  assign lizzieLet20_1_4QVal_Bool_6QVal_Bool_done = (lizzieLet20_1_4QVal_Bool_6QVal_Bool_emitted | ({lizzieLet20_1_4QVal_Bool_6QVal_Bool_3_d[0],
                                                                                                     lizzieLet20_1_4QVal_Bool_6QVal_Bool_2_d[0],
                                                                                                     lizzieLet20_1_4QVal_Bool_6QVal_Bool_1_d[0]} & {lizzieLet20_1_4QVal_Bool_6QVal_Bool_3_r,
                                                                                                                                                    lizzieLet20_1_4QVal_Bool_6QVal_Bool_2_r,
                                                                                                                                                    lizzieLet20_1_4QVal_Bool_6QVal_Bool_1_r}));
  assign lizzieLet20_1_4QVal_Bool_6QVal_Bool_r = (& lizzieLet20_1_4QVal_Bool_6QVal_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet20_1_4QVal_Bool_6QVal_Bool_emitted <= 3'd0;
    else
      lizzieLet20_1_4QVal_Bool_6QVal_Bool_emitted <= (lizzieLet20_1_4QVal_Bool_6QVal_Bool_r ? 3'd0 :
                                                      lizzieLet20_1_4QVal_Bool_6QVal_Bool_done);
  
  /* demux (Ty MyBool,
       Ty Go) : (lizzieLet20_1_4QVal_Bool_6QVal_Bool_1,MyBool) (lizzieLet20_1_4QVal_Bool_3QVal_Bool,Go) > [(lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyFalse,Go),
                                                                                                           (lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyTrue,Go)] */
  logic [1:0] lizzieLet20_1_4QVal_Bool_3QVal_Bool_onehotd;
  always_comb
    if ((lizzieLet20_1_4QVal_Bool_6QVal_Bool_1_d[0] && lizzieLet20_1_4QVal_Bool_3QVal_Bool_d[0]))
      unique case (lizzieLet20_1_4QVal_Bool_6QVal_Bool_1_d[1:1])
        1'd0: lizzieLet20_1_4QVal_Bool_3QVal_Bool_onehotd = 2'd1;
        1'd1: lizzieLet20_1_4QVal_Bool_3QVal_Bool_onehotd = 2'd2;
        default: lizzieLet20_1_4QVal_Bool_3QVal_Bool_onehotd = 2'd0;
      endcase
    else lizzieLet20_1_4QVal_Bool_3QVal_Bool_onehotd = 2'd0;
  assign lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyFalse_d = lizzieLet20_1_4QVal_Bool_3QVal_Bool_onehotd[0];
  assign lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyTrue_d = lizzieLet20_1_4QVal_Bool_3QVal_Bool_onehotd[1];
  assign lizzieLet20_1_4QVal_Bool_3QVal_Bool_r = (| (lizzieLet20_1_4QVal_Bool_3QVal_Bool_onehotd & {lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyTrue_r,
                                                                                                    lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyFalse_r}));
  assign lizzieLet20_1_4QVal_Bool_6QVal_Bool_1_r = lizzieLet20_1_4QVal_Bool_3QVal_Bool_r;
  
  /* fork (Ty Go) : (lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyTrue,Go) > [(lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyTrue_1,Go),
                                                                   (lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyTrue_2,Go)] */
  logic [1:0] lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyTrue_emitted;
  logic [1:0] lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyTrue_done;
  assign lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyTrue_1_d = (lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyTrue_d[0] && (! lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyTrue_emitted[0]));
  assign lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyTrue_2_d = (lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyTrue_d[0] && (! lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyTrue_emitted[1]));
  assign lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyTrue_done = (lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyTrue_emitted | ({lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyTrue_2_d[0],
                                                                                                                     lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyTrue_1_d[0]} & {lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyTrue_2_r,
                                                                                                                                                                            lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyTrue_1_r}));
  assign lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyTrue_r = (& lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyTrue_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyTrue_emitted <= 2'd0;
    else
      lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyTrue_emitted <= (lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyTrue_r ? 2'd0 :
                                                              lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyTrue_done);
  
  /* buf (Ty Go) : (lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyTrue_1,Go) > (lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyTrue_1_argbuf,Go) */
  Go_t lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyTrue_1_bufchan_d;
  logic lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyTrue_1_bufchan_r;
  assign lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyTrue_1_r = ((! lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyTrue_1_bufchan_d[0]) || lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyTrue_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyTrue_1_bufchan_d <= 1'd0;
    else
      if (lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyTrue_1_r)
        lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyTrue_1_bufchan_d <= lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyTrue_1_d;
  Go_t lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyTrue_1_bufchan_buf;
  assign lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyTrue_1_bufchan_r = (! lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyTrue_1_bufchan_buf[0]);
  assign lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyTrue_1_argbuf_d = (lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyTrue_1_bufchan_buf[0] ? lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyTrue_1_bufchan_buf :
                                                                   lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyTrue_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyTrue_1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyTrue_1_argbuf_r && lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyTrue_1_bufchan_buf[0]))
        lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyTrue_1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyTrue_1_argbuf_r) && (! lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyTrue_1_bufchan_buf[0])))
        lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyTrue_1_bufchan_buf <= lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyTrue_1_bufchan_d;
  
  /* dcon (Ty TupGo,
      Dcon TupGo) : [(lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyTrue_1_argbuf,Go)] > (lvlrcX-0TupGo2,TupGo) */
  assign \lvlrcX-0TupGo2_d  = TupGo_dc((& {lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyTrue_1_argbuf_d[0]}), lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyTrue_1_argbuf_d);
  assign {lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyTrue_1_argbuf_r} = {1 {(\lvlrcX-0TupGo2_r  && \lvlrcX-0TupGo2_d [0])}};
  
  /* buf (Ty Go) : (lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyTrue_2,Go) > (lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyTrue_2_argbuf,Go) */
  Go_t lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyTrue_2_bufchan_d;
  logic lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyTrue_2_bufchan_r;
  assign lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyTrue_2_r = ((! lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyTrue_2_bufchan_d[0]) || lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyTrue_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyTrue_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyTrue_2_r)
        lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyTrue_2_bufchan_d <= lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyTrue_2_d;
  Go_t lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyTrue_2_bufchan_buf;
  assign lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyTrue_2_bufchan_r = (! lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyTrue_2_bufchan_buf[0]);
  assign lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyTrue_2_argbuf_d = (lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyTrue_2_bufchan_buf[0] ? lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyTrue_2_bufchan_buf :
                                                                   lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyTrue_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyTrue_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyTrue_2_argbuf_r && lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyTrue_2_bufchan_buf[0]))
        lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyTrue_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyTrue_2_argbuf_r) && (! lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyTrue_2_bufchan_buf[0])))
        lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyTrue_2_bufchan_buf <= lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyTrue_2_bufchan_d;
  
  /* demux (Ty MyBool,
       Ty Pointer_CTf') : (lizzieLet20_1_4QVal_Bool_6QVal_Bool_2,MyBool) (lizzieLet20_1_4QVal_Bool_5QVal_Bool,Pointer_CTf') > [(lizzieLet20_1_4QVal_Bool_6QVal_Bool_2MyFalse,Pointer_CTf'),
                                                                                                                               (lizzieLet20_1_4QVal_Bool_6QVal_Bool_2MyTrue,Pointer_CTf')] */
  logic [1:0] lizzieLet20_1_4QVal_Bool_5QVal_Bool_onehotd;
  always_comb
    if ((lizzieLet20_1_4QVal_Bool_6QVal_Bool_2_d[0] && lizzieLet20_1_4QVal_Bool_5QVal_Bool_d[0]))
      unique case (lizzieLet20_1_4QVal_Bool_6QVal_Bool_2_d[1:1])
        1'd0: lizzieLet20_1_4QVal_Bool_5QVal_Bool_onehotd = 2'd1;
        1'd1: lizzieLet20_1_4QVal_Bool_5QVal_Bool_onehotd = 2'd2;
        default: lizzieLet20_1_4QVal_Bool_5QVal_Bool_onehotd = 2'd0;
      endcase
    else lizzieLet20_1_4QVal_Bool_5QVal_Bool_onehotd = 2'd0;
  assign lizzieLet20_1_4QVal_Bool_6QVal_Bool_2MyFalse_d = {lizzieLet20_1_4QVal_Bool_5QVal_Bool_d[16:1],
                                                           lizzieLet20_1_4QVal_Bool_5QVal_Bool_onehotd[0]};
  assign lizzieLet20_1_4QVal_Bool_6QVal_Bool_2MyTrue_d = {lizzieLet20_1_4QVal_Bool_5QVal_Bool_d[16:1],
                                                          lizzieLet20_1_4QVal_Bool_5QVal_Bool_onehotd[1]};
  assign lizzieLet20_1_4QVal_Bool_5QVal_Bool_r = (| (lizzieLet20_1_4QVal_Bool_5QVal_Bool_onehotd & {lizzieLet20_1_4QVal_Bool_6QVal_Bool_2MyTrue_r,
                                                                                                    lizzieLet20_1_4QVal_Bool_6QVal_Bool_2MyFalse_r}));
  assign lizzieLet20_1_4QVal_Bool_6QVal_Bool_2_r = lizzieLet20_1_4QVal_Bool_5QVal_Bool_r;
  
  /* buf (Ty Pointer_CTf') : (lizzieLet20_1_4QVal_Bool_6QVal_Bool_2MyTrue,Pointer_CTf') > (lizzieLet20_1_4QVal_Bool_6QVal_Bool_2MyTrue_1_argbuf,Pointer_CTf') */
  \Pointer_CTf'_t  lizzieLet20_1_4QVal_Bool_6QVal_Bool_2MyTrue_bufchan_d;
  logic lizzieLet20_1_4QVal_Bool_6QVal_Bool_2MyTrue_bufchan_r;
  assign lizzieLet20_1_4QVal_Bool_6QVal_Bool_2MyTrue_r = ((! lizzieLet20_1_4QVal_Bool_6QVal_Bool_2MyTrue_bufchan_d[0]) || lizzieLet20_1_4QVal_Bool_6QVal_Bool_2MyTrue_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet20_1_4QVal_Bool_6QVal_Bool_2MyTrue_bufchan_d <= {16'd0,
                                                                1'd0};
    else
      if (lizzieLet20_1_4QVal_Bool_6QVal_Bool_2MyTrue_r)
        lizzieLet20_1_4QVal_Bool_6QVal_Bool_2MyTrue_bufchan_d <= lizzieLet20_1_4QVal_Bool_6QVal_Bool_2MyTrue_d;
  \Pointer_CTf'_t  lizzieLet20_1_4QVal_Bool_6QVal_Bool_2MyTrue_bufchan_buf;
  assign lizzieLet20_1_4QVal_Bool_6QVal_Bool_2MyTrue_bufchan_r = (! lizzieLet20_1_4QVal_Bool_6QVal_Bool_2MyTrue_bufchan_buf[0]);
  assign lizzieLet20_1_4QVal_Bool_6QVal_Bool_2MyTrue_1_argbuf_d = (lizzieLet20_1_4QVal_Bool_6QVal_Bool_2MyTrue_bufchan_buf[0] ? lizzieLet20_1_4QVal_Bool_6QVal_Bool_2MyTrue_bufchan_buf :
                                                                   lizzieLet20_1_4QVal_Bool_6QVal_Bool_2MyTrue_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet20_1_4QVal_Bool_6QVal_Bool_2MyTrue_bufchan_buf <= {16'd0,
                                                                  1'd0};
    else
      if ((lizzieLet20_1_4QVal_Bool_6QVal_Bool_2MyTrue_1_argbuf_r && lizzieLet20_1_4QVal_Bool_6QVal_Bool_2MyTrue_bufchan_buf[0]))
        lizzieLet20_1_4QVal_Bool_6QVal_Bool_2MyTrue_bufchan_buf <= {16'd0,
                                                                    1'd0};
      else if (((! lizzieLet20_1_4QVal_Bool_6QVal_Bool_2MyTrue_1_argbuf_r) && (! lizzieLet20_1_4QVal_Bool_6QVal_Bool_2MyTrue_bufchan_buf[0])))
        lizzieLet20_1_4QVal_Bool_6QVal_Bool_2MyTrue_bufchan_buf <= lizzieLet20_1_4QVal_Bool_6QVal_Bool_2MyTrue_bufchan_d;
  
  /* demux (Ty MyBool,
       Ty MyBool) : (lizzieLet20_1_4QVal_Bool_6QVal_Bool_3,MyBool) (va8K_destruct,MyBool) > [(lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse,MyBool),
                                                                                             (_32,MyBool)] */
  logic [1:0] va8K_destruct_onehotd;
  always_comb
    if ((lizzieLet20_1_4QVal_Bool_6QVal_Bool_3_d[0] && va8K_destruct_d[0]))
      unique case (lizzieLet20_1_4QVal_Bool_6QVal_Bool_3_d[1:1])
        1'd0: va8K_destruct_onehotd = 2'd1;
        1'd1: va8K_destruct_onehotd = 2'd2;
        default: va8K_destruct_onehotd = 2'd0;
      endcase
    else va8K_destruct_onehotd = 2'd0;
  assign lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_d = {va8K_destruct_d[1:1],
                                                           va8K_destruct_onehotd[0]};
  assign _32_d = {va8K_destruct_d[1:1], va8K_destruct_onehotd[1]};
  assign va8K_destruct_r = (| (va8K_destruct_onehotd & {_32_r,
                                                        lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_r}));
  assign lizzieLet20_1_4QVal_Bool_6QVal_Bool_3_r = va8K_destruct_r;
  
  /* fork (Ty MyBool) : (lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse,MyBool) > [(lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1,MyBool),
                                                                            (lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_2,MyBool)] */
  logic [1:0] lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_emitted;
  logic [1:0] lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_done;
  assign lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1_d = {lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_d[1:1],
                                                             (lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_d[0] && (! lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_emitted[0]))};
  assign lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_2_d = {lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_d[1:1],
                                                             (lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_d[0] && (! lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_emitted[1]))};
  assign lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_done = (lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_emitted | ({lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_2_d[0],
                                                                                                                       lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1_d[0]} & {lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_2_r,
                                                                                                                                                                               lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1_r}));
  assign lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_r = (& lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_emitted <= 2'd0;
    else
      lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_emitted <= (lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_r ? 2'd0 :
                                                               lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_done);
  
  /* demux (Ty MyBool,
       Ty Go) : (lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1,MyBool) (lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyFalse,Go) > [(lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse,Go),
                                                                                                                             (lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue,Go)] */
  logic [1:0] lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyFalse_onehotd;
  always_comb
    if ((lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1_d[0] && lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyFalse_d[0]))
      unique case (lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1_d[1:1])
        1'd0: lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyFalse_onehotd = 2'd1;
        1'd1: lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyFalse_onehotd = 2'd2;
        default:
          lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyFalse_onehotd = 2'd0;
      endcase
    else lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyFalse_onehotd = 2'd0;
  assign lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_d = lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyFalse_onehotd[0];
  assign lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_d = lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyFalse_onehotd[1];
  assign lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyFalse_r = (| (lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyFalse_onehotd & {lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_r,
                                                                                                                      lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_r}));
  assign lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1_r = lizzieLet20_1_4QVal_Bool_6QVal_Bool_1MyFalse_r;
  
  /* fork (Ty Go) : (lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse,Go) > [(lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1,Go),
                                                                             (lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2,Go)] */
  logic [1:0] lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_emitted;
  logic [1:0] lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_done;
  assign lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1_d = (lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_d[0] && (! lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_emitted[0]));
  assign lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_d = (lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_d[0] && (! lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_emitted[1]));
  assign lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_done = (lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_emitted | ({lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_d[0],
                                                                                                                                         lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1_d[0]} & {lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_r,
                                                                                                                                                                                                          lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1_r}));
  assign lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_r = (& lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_emitted <= 2'd0;
    else
      lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_emitted <= (lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_r ? 2'd0 :
                                                                        lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_done);
  
  /* dcon (Ty QTree_Bool,
      Dcon QNone_Bool) : [(lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1,Go)] > (lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool,QTree_Bool) */
  assign lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_d = QNone_Bool_dc((& {lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1_d[0]}), lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1_d);
  assign {lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1_r} = {1 {(lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_r && lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_d[0])}};
  
  /* buf (Ty QTree_Bool) : (lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool,QTree_Bool) > (lizzieLet22_1_1_argbuf,QTree_Bool) */
  QTree_Bool_t lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_bufchan_d;
  logic lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_bufchan_r;
  assign lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_r = ((! lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_bufchan_d[0]) || lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_bufchan_d <= {66'd0,
                                                                                      1'd0};
    else
      if (lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_r)
        lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_bufchan_d <= lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_d;
  QTree_Bool_t lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_bufchan_buf;
  assign lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_bufchan_r = (! lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_bufchan_buf[0]);
  assign lizzieLet22_1_1_argbuf_d = (lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_bufchan_buf[0] ? lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_bufchan_buf :
                                     lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_bufchan_buf <= {66'd0,
                                                                                        1'd0};
    else
      if ((lizzieLet22_1_1_argbuf_r && lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_bufchan_buf[0]))
        lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_bufchan_buf <= {66'd0,
                                                                                          1'd0};
      else if (((! lizzieLet22_1_1_argbuf_r) && (! lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_bufchan_buf[0])))
        lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_bufchan_buf <= lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_1QNone_Bool_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2,Go) > (lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_argbuf,Go) */
  Go_t lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_bufchan_d;
  logic lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_bufchan_r;
  assign lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_r = ((! lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_bufchan_d[0]) || lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_r)
        lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_bufchan_d <= lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_d;
  Go_t lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_bufchan_buf;
  assign lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_bufchan_r = (! lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_bufchan_buf[0]);
  assign lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_argbuf_d = (lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_bufchan_buf[0] ? lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_bufchan_buf :
                                                                             lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_argbuf_r && lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_bufchan_buf[0]))
        lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_argbuf_r) && (! lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_bufchan_buf[0])))
        lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_bufchan_buf <= lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyFalse_2_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue,Go) > [(lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1,Go),
                                                                            (lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2,Go)] */
  logic [1:0] lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_emitted;
  logic [1:0] lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_done;
  assign lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_d = (lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_d[0] && (! lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_emitted[0]));
  assign lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_d = (lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_d[0] && (! lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_emitted[1]));
  assign lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_done = (lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_emitted | ({lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_d[0],
                                                                                                                                       lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_d[0]} & {lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_r,
                                                                                                                                                                                                       lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_r}));
  assign lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_r = (& lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_emitted <= 2'd0;
    else
      lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_emitted <= (lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_r ? 2'd0 :
                                                                       lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_done);
  
  /* buf (Ty Go) : (lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1,Go) > (lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_argbuf,Go) */
  Go_t lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_bufchan_d;
  logic lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_bufchan_r;
  assign lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_r = ((! lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_bufchan_d[0]) || lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_bufchan_d <= 1'd0;
    else
      if (lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_r)
        lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_bufchan_d <= lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_d;
  Go_t lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_bufchan_buf;
  assign lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_bufchan_r = (! lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_bufchan_buf[0]);
  assign lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_argbuf_d = (lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_bufchan_buf[0] ? lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_bufchan_buf :
                                                                            lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_argbuf_r && lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_bufchan_buf[0]))
        lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_argbuf_r) && (! lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_bufchan_buf[0])))
        lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_bufchan_buf <= lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_bufchan_d;
  
  /* dcon (Ty TupGo,
      Dcon TupGo) : [(lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_argbuf,Go)] > (lvlrcX-0TupGo_1,TupGo) */
  assign \lvlrcX-0TupGo_1_d  = TupGo_dc((& {lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_argbuf_d[0]}), lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_argbuf_d);
  assign {lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_1_argbuf_r} = {1 {(\lvlrcX-0TupGo_1_r  && \lvlrcX-0TupGo_1_d [0])}};
  
  /* buf (Ty Go) : (lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2,Go) > (lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_argbuf,Go) */
  Go_t lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_bufchan_d;
  logic lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_bufchan_r;
  assign lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_r = ((! lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_bufchan_d[0]) || lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_r)
        lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_bufchan_d <= lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_d;
  Go_t lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_bufchan_buf;
  assign lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_bufchan_r = (! lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_bufchan_buf[0]);
  assign lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_argbuf_d = (lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_bufchan_buf[0] ? lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_bufchan_buf :
                                                                            lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_argbuf_r && lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_bufchan_buf[0]))
        lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_argbuf_r) && (! lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_bufchan_buf[0])))
        lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_bufchan_buf <= lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_1MyTrue_2_bufchan_d;
  
  /* demux (Ty MyBool,
       Ty Pointer_CTf') : (lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_2,MyBool) (lizzieLet20_1_4QVal_Bool_6QVal_Bool_2MyFalse,Pointer_CTf') > [(lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_2MyFalse,Pointer_CTf'),
                                                                                                                                                 (lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_2MyTrue,Pointer_CTf')] */
  logic [1:0] lizzieLet20_1_4QVal_Bool_6QVal_Bool_2MyFalse_onehotd;
  always_comb
    if ((lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_2_d[0] && lizzieLet20_1_4QVal_Bool_6QVal_Bool_2MyFalse_d[0]))
      unique case (lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_2_d[1:1])
        1'd0: lizzieLet20_1_4QVal_Bool_6QVal_Bool_2MyFalse_onehotd = 2'd1;
        1'd1: lizzieLet20_1_4QVal_Bool_6QVal_Bool_2MyFalse_onehotd = 2'd2;
        default:
          lizzieLet20_1_4QVal_Bool_6QVal_Bool_2MyFalse_onehotd = 2'd0;
      endcase
    else lizzieLet20_1_4QVal_Bool_6QVal_Bool_2MyFalse_onehotd = 2'd0;
  assign lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_2MyFalse_d = {lizzieLet20_1_4QVal_Bool_6QVal_Bool_2MyFalse_d[16:1],
                                                                    lizzieLet20_1_4QVal_Bool_6QVal_Bool_2MyFalse_onehotd[0]};
  assign lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_2MyTrue_d = {lizzieLet20_1_4QVal_Bool_6QVal_Bool_2MyFalse_d[16:1],
                                                                   lizzieLet20_1_4QVal_Bool_6QVal_Bool_2MyFalse_onehotd[1]};
  assign lizzieLet20_1_4QVal_Bool_6QVal_Bool_2MyFalse_r = (| (lizzieLet20_1_4QVal_Bool_6QVal_Bool_2MyFalse_onehotd & {lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_2MyTrue_r,
                                                                                                                      lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_2MyFalse_r}));
  assign lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_2_r = lizzieLet20_1_4QVal_Bool_6QVal_Bool_2MyFalse_r;
  
  /* buf (Ty Pointer_CTf') : (lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_2MyFalse,Pointer_CTf') > (lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_2MyFalse_1_argbuf,Pointer_CTf') */
  \Pointer_CTf'_t  lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_2MyFalse_bufchan_d;
  logic lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_2MyFalse_bufchan_r;
  assign lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_2MyFalse_r = ((! lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_2MyFalse_bufchan_d[0]) || lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_2MyFalse_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_2MyFalse_bufchan_d <= {16'd0,
                                                                          1'd0};
    else
      if (lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_2MyFalse_r)
        lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_2MyFalse_bufchan_d <= lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_2MyFalse_d;
  \Pointer_CTf'_t  lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_2MyFalse_bufchan_buf;
  assign lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_2MyFalse_bufchan_r = (! lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_2MyFalse_bufchan_buf[0]);
  assign lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_2MyFalse_1_argbuf_d = (lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_2MyFalse_bufchan_buf[0] ? lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_2MyFalse_bufchan_buf :
                                                                             lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_2MyFalse_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_2MyFalse_bufchan_buf <= {16'd0,
                                                                            1'd0};
    else
      if ((lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_2MyFalse_1_argbuf_r && lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_2MyFalse_bufchan_buf[0]))
        lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_2MyFalse_bufchan_buf <= {16'd0,
                                                                              1'd0};
      else if (((! lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_2MyFalse_1_argbuf_r) && (! lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_2MyFalse_bufchan_buf[0])))
        lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_2MyFalse_bufchan_buf <= lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_2MyFalse_bufchan_d;
  
  /* buf (Ty Pointer_CTf') : (lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_2MyTrue,Pointer_CTf') > (lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_2MyTrue_1_argbuf,Pointer_CTf') */
  \Pointer_CTf'_t  lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_2MyTrue_bufchan_d;
  logic lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_2MyTrue_bufchan_r;
  assign lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_2MyTrue_r = ((! lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_2MyTrue_bufchan_d[0]) || lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_2MyTrue_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_2MyTrue_bufchan_d <= {16'd0,
                                                                         1'd0};
    else
      if (lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_2MyTrue_r)
        lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_2MyTrue_bufchan_d <= lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_2MyTrue_d;
  \Pointer_CTf'_t  lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_2MyTrue_bufchan_buf;
  assign lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_2MyTrue_bufchan_r = (! lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_2MyTrue_bufchan_buf[0]);
  assign lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_2MyTrue_1_argbuf_d = (lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_2MyTrue_bufchan_buf[0] ? lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_2MyTrue_bufchan_buf :
                                                                            lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_2MyTrue_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_2MyTrue_bufchan_buf <= {16'd0,
                                                                           1'd0};
    else
      if ((lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_2MyTrue_1_argbuf_r && lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_2MyTrue_bufchan_buf[0]))
        lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_2MyTrue_bufchan_buf <= {16'd0,
                                                                             1'd0};
      else if (((! lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_2MyTrue_1_argbuf_r) && (! lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_2MyTrue_bufchan_buf[0])))
        lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_2MyTrue_bufchan_buf <= lizzieLet20_1_4QVal_Bool_6QVal_Bool_3MyFalse_2MyTrue_bufchan_d;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_QTree_Bool) : (lizzieLet20_1_5,QTree_Bool) (m2a8H_2,Pointer_QTree_Bool) > [(_31,Pointer_QTree_Bool),
                                                                                             (lizzieLet20_1_5QVal_Bool,Pointer_QTree_Bool),
                                                                                             (lizzieLet20_1_5QNode_Bool,Pointer_QTree_Bool),
                                                                                             (_30,Pointer_QTree_Bool)] */
  logic [3:0] m2a8H_2_onehotd;
  always_comb
    if ((lizzieLet20_1_5_d[0] && m2a8H_2_d[0]))
      unique case (lizzieLet20_1_5_d[2:1])
        2'd0: m2a8H_2_onehotd = 4'd1;
        2'd1: m2a8H_2_onehotd = 4'd2;
        2'd2: m2a8H_2_onehotd = 4'd4;
        2'd3: m2a8H_2_onehotd = 4'd8;
        default: m2a8H_2_onehotd = 4'd0;
      endcase
    else m2a8H_2_onehotd = 4'd0;
  assign _31_d = {m2a8H_2_d[16:1], m2a8H_2_onehotd[0]};
  assign lizzieLet20_1_5QVal_Bool_d = {m2a8H_2_d[16:1],
                                       m2a8H_2_onehotd[1]};
  assign lizzieLet20_1_5QNode_Bool_d = {m2a8H_2_d[16:1],
                                        m2a8H_2_onehotd[2]};
  assign _30_d = {m2a8H_2_d[16:1], m2a8H_2_onehotd[3]};
  assign m2a8H_2_r = (| (m2a8H_2_onehotd & {_30_r,
                                            lizzieLet20_1_5QNode_Bool_r,
                                            lizzieLet20_1_5QVal_Bool_r,
                                            _31_r}));
  assign lizzieLet20_1_5_r = m2a8H_2_r;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_QTree_Bool) : (lizzieLet20_1_6,QTree_Bool) (m3a8I_2,Pointer_QTree_Bool) > [(lizzieLet20_1_6QNone_Bool,Pointer_QTree_Bool),
                                                                                             (_29,Pointer_QTree_Bool),
                                                                                             (_28,Pointer_QTree_Bool),
                                                                                             (_27,Pointer_QTree_Bool)] */
  logic [3:0] m3a8I_2_onehotd;
  always_comb
    if ((lizzieLet20_1_6_d[0] && m3a8I_2_d[0]))
      unique case (lizzieLet20_1_6_d[2:1])
        2'd0: m3a8I_2_onehotd = 4'd1;
        2'd1: m3a8I_2_onehotd = 4'd2;
        2'd2: m3a8I_2_onehotd = 4'd4;
        2'd3: m3a8I_2_onehotd = 4'd8;
        default: m3a8I_2_onehotd = 4'd0;
      endcase
    else m3a8I_2_onehotd = 4'd0;
  assign lizzieLet20_1_6QNone_Bool_d = {m3a8I_2_d[16:1],
                                        m3a8I_2_onehotd[0]};
  assign _29_d = {m3a8I_2_d[16:1], m3a8I_2_onehotd[1]};
  assign _28_d = {m3a8I_2_d[16:1], m3a8I_2_onehotd[2]};
  assign _27_d = {m3a8I_2_d[16:1], m3a8I_2_onehotd[3]};
  assign m3a8I_2_r = (| (m3a8I_2_onehotd & {_27_r,
                                            _28_r,
                                            _29_r,
                                            lizzieLet20_1_6QNone_Bool_r}));
  assign lizzieLet20_1_6_r = m3a8I_2_r;
  
  /* buf (Ty Pointer_QTree_Bool) : (lizzieLet20_1_6QNone_Bool,Pointer_QTree_Bool) > (lizzieLet20_1_6QNone_Bool_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t lizzieLet20_1_6QNone_Bool_bufchan_d;
  logic lizzieLet20_1_6QNone_Bool_bufchan_r;
  assign lizzieLet20_1_6QNone_Bool_r = ((! lizzieLet20_1_6QNone_Bool_bufchan_d[0]) || lizzieLet20_1_6QNone_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet20_1_6QNone_Bool_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet20_1_6QNone_Bool_r)
        lizzieLet20_1_6QNone_Bool_bufchan_d <= lizzieLet20_1_6QNone_Bool_d;
  Pointer_QTree_Bool_t lizzieLet20_1_6QNone_Bool_bufchan_buf;
  assign lizzieLet20_1_6QNone_Bool_bufchan_r = (! lizzieLet20_1_6QNone_Bool_bufchan_buf[0]);
  assign lizzieLet20_1_6QNone_Bool_1_argbuf_d = (lizzieLet20_1_6QNone_Bool_bufchan_buf[0] ? lizzieLet20_1_6QNone_Bool_bufchan_buf :
                                                 lizzieLet20_1_6QNone_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet20_1_6QNone_Bool_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet20_1_6QNone_Bool_1_argbuf_r && lizzieLet20_1_6QNone_Bool_bufchan_buf[0]))
        lizzieLet20_1_6QNone_Bool_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet20_1_6QNone_Bool_1_argbuf_r) && (! lizzieLet20_1_6QNone_Bool_bufchan_buf[0])))
        lizzieLet20_1_6QNone_Bool_bufchan_buf <= lizzieLet20_1_6QNone_Bool_bufchan_d;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_CTf') : (lizzieLet20_1_7,QTree_Bool) (sc_0_1_goMux_mux,Pointer_CTf') > [(lizzieLet20_1_7QNone_Bool,Pointer_CTf'),
                                                                                          (lizzieLet20_1_7QVal_Bool,Pointer_CTf'),
                                                                                          (lizzieLet20_1_7QNode_Bool,Pointer_CTf'),
                                                                                          (lizzieLet20_1_7QError_Bool,Pointer_CTf')] */
  logic [3:0] sc_0_1_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet20_1_7_d[0] && sc_0_1_goMux_mux_d[0]))
      unique case (lizzieLet20_1_7_d[2:1])
        2'd0: sc_0_1_goMux_mux_onehotd = 4'd1;
        2'd1: sc_0_1_goMux_mux_onehotd = 4'd2;
        2'd2: sc_0_1_goMux_mux_onehotd = 4'd4;
        2'd3: sc_0_1_goMux_mux_onehotd = 4'd8;
        default: sc_0_1_goMux_mux_onehotd = 4'd0;
      endcase
    else sc_0_1_goMux_mux_onehotd = 4'd0;
  assign lizzieLet20_1_7QNone_Bool_d = {sc_0_1_goMux_mux_d[16:1],
                                        sc_0_1_goMux_mux_onehotd[0]};
  assign lizzieLet20_1_7QVal_Bool_d = {sc_0_1_goMux_mux_d[16:1],
                                       sc_0_1_goMux_mux_onehotd[1]};
  assign lizzieLet20_1_7QNode_Bool_d = {sc_0_1_goMux_mux_d[16:1],
                                        sc_0_1_goMux_mux_onehotd[2]};
  assign lizzieLet20_1_7QError_Bool_d = {sc_0_1_goMux_mux_d[16:1],
                                         sc_0_1_goMux_mux_onehotd[3]};
  assign sc_0_1_goMux_mux_r = (| (sc_0_1_goMux_mux_onehotd & {lizzieLet20_1_7QError_Bool_r,
                                                              lizzieLet20_1_7QNode_Bool_r,
                                                              lizzieLet20_1_7QVal_Bool_r,
                                                              lizzieLet20_1_7QNone_Bool_r}));
  assign lizzieLet20_1_7_r = sc_0_1_goMux_mux_r;
  
  /* buf (Ty Pointer_CTf') : (lizzieLet20_1_7QError_Bool,Pointer_CTf') > (lizzieLet20_1_7QError_Bool_1_argbuf,Pointer_CTf') */
  \Pointer_CTf'_t  lizzieLet20_1_7QError_Bool_bufchan_d;
  logic lizzieLet20_1_7QError_Bool_bufchan_r;
  assign lizzieLet20_1_7QError_Bool_r = ((! lizzieLet20_1_7QError_Bool_bufchan_d[0]) || lizzieLet20_1_7QError_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet20_1_7QError_Bool_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet20_1_7QError_Bool_r)
        lizzieLet20_1_7QError_Bool_bufchan_d <= lizzieLet20_1_7QError_Bool_d;
  \Pointer_CTf'_t  lizzieLet20_1_7QError_Bool_bufchan_buf;
  assign lizzieLet20_1_7QError_Bool_bufchan_r = (! lizzieLet20_1_7QError_Bool_bufchan_buf[0]);
  assign lizzieLet20_1_7QError_Bool_1_argbuf_d = (lizzieLet20_1_7QError_Bool_bufchan_buf[0] ? lizzieLet20_1_7QError_Bool_bufchan_buf :
                                                  lizzieLet20_1_7QError_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet20_1_7QError_Bool_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet20_1_7QError_Bool_1_argbuf_r && lizzieLet20_1_7QError_Bool_bufchan_buf[0]))
        lizzieLet20_1_7QError_Bool_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet20_1_7QError_Bool_1_argbuf_r) && (! lizzieLet20_1_7QError_Bool_bufchan_buf[0])))
        lizzieLet20_1_7QError_Bool_bufchan_buf <= lizzieLet20_1_7QError_Bool_bufchan_d;
  
  /* buf (Ty Pointer_CTf') : (lizzieLet20_1_7QNone_Bool,Pointer_CTf') > (lizzieLet20_1_7QNone_Bool_1_argbuf,Pointer_CTf') */
  \Pointer_CTf'_t  lizzieLet20_1_7QNone_Bool_bufchan_d;
  logic lizzieLet20_1_7QNone_Bool_bufchan_r;
  assign lizzieLet20_1_7QNone_Bool_r = ((! lizzieLet20_1_7QNone_Bool_bufchan_d[0]) || lizzieLet20_1_7QNone_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet20_1_7QNone_Bool_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet20_1_7QNone_Bool_r)
        lizzieLet20_1_7QNone_Bool_bufchan_d <= lizzieLet20_1_7QNone_Bool_d;
  \Pointer_CTf'_t  lizzieLet20_1_7QNone_Bool_bufchan_buf;
  assign lizzieLet20_1_7QNone_Bool_bufchan_r = (! lizzieLet20_1_7QNone_Bool_bufchan_buf[0]);
  assign lizzieLet20_1_7QNone_Bool_1_argbuf_d = (lizzieLet20_1_7QNone_Bool_bufchan_buf[0] ? lizzieLet20_1_7QNone_Bool_bufchan_buf :
                                                 lizzieLet20_1_7QNone_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet20_1_7QNone_Bool_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet20_1_7QNone_Bool_1_argbuf_r && lizzieLet20_1_7QNone_Bool_bufchan_buf[0]))
        lizzieLet20_1_7QNone_Bool_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet20_1_7QNone_Bool_1_argbuf_r) && (! lizzieLet20_1_7QNone_Bool_bufchan_buf[0])))
        lizzieLet20_1_7QNone_Bool_bufchan_buf <= lizzieLet20_1_7QNone_Bool_bufchan_d;
  
  /* destruct (Ty MaskQTree,
          Dcon MQNode) : (lizzieLet32_1MQNode,MaskQTree) > [(q1a8y_destruct,Pointer_MaskQTree),
                                                            (q2a8z_destruct,Pointer_MaskQTree),
                                                            (q3a8A_destruct,Pointer_MaskQTree),
                                                            (q5a8B_destruct,Pointer_MaskQTree)] */
  logic [3:0] lizzieLet32_1MQNode_emitted;
  logic [3:0] lizzieLet32_1MQNode_done;
  assign q1a8y_destruct_d = {lizzieLet32_1MQNode_d[18:3],
                             (lizzieLet32_1MQNode_d[0] && (! lizzieLet32_1MQNode_emitted[0]))};
  assign q2a8z_destruct_d = {lizzieLet32_1MQNode_d[34:19],
                             (lizzieLet32_1MQNode_d[0] && (! lizzieLet32_1MQNode_emitted[1]))};
  assign q3a8A_destruct_d = {lizzieLet32_1MQNode_d[50:35],
                             (lizzieLet32_1MQNode_d[0] && (! lizzieLet32_1MQNode_emitted[2]))};
  assign q5a8B_destruct_d = {lizzieLet32_1MQNode_d[66:51],
                             (lizzieLet32_1MQNode_d[0] && (! lizzieLet32_1MQNode_emitted[3]))};
  assign lizzieLet32_1MQNode_done = (lizzieLet32_1MQNode_emitted | ({q5a8B_destruct_d[0],
                                                                     q3a8A_destruct_d[0],
                                                                     q2a8z_destruct_d[0],
                                                                     q1a8y_destruct_d[0]} & {q5a8B_destruct_r,
                                                                                             q3a8A_destruct_r,
                                                                                             q2a8z_destruct_r,
                                                                                             q1a8y_destruct_r}));
  assign lizzieLet32_1MQNode_r = (& lizzieLet32_1MQNode_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet32_1MQNode_emitted <= 4'd0;
    else
      lizzieLet32_1MQNode_emitted <= (lizzieLet32_1MQNode_r ? 4'd0 :
                                      lizzieLet32_1MQNode_done);
  
  /* demux (Ty MaskQTree,
       Ty MaskQTree) : (lizzieLet32_2,MaskQTree) (lizzieLet32_1,MaskQTree) > [(_26,MaskQTree),
                                                                              (_25,MaskQTree),
                                                                              (lizzieLet32_1MQNode,MaskQTree)] */
  logic [2:0] lizzieLet32_1_onehotd;
  always_comb
    if ((lizzieLet32_2_d[0] && lizzieLet32_1_d[0]))
      unique case (lizzieLet32_2_d[2:1])
        2'd0: lizzieLet32_1_onehotd = 3'd1;
        2'd1: lizzieLet32_1_onehotd = 3'd2;
        2'd2: lizzieLet32_1_onehotd = 3'd4;
        default: lizzieLet32_1_onehotd = 3'd0;
      endcase
    else lizzieLet32_1_onehotd = 3'd0;
  assign _26_d = {lizzieLet32_1_d[66:1], lizzieLet32_1_onehotd[0]};
  assign _25_d = {lizzieLet32_1_d[66:1], lizzieLet32_1_onehotd[1]};
  assign lizzieLet32_1MQNode_d = {lizzieLet32_1_d[66:1],
                                  lizzieLet32_1_onehotd[2]};
  assign lizzieLet32_1_r = (| (lizzieLet32_1_onehotd & {lizzieLet32_1MQNode_r,
                                                        _25_r,
                                                        _26_r}));
  assign lizzieLet32_2_r = lizzieLet32_1_r;
  
  /* demux (Ty MaskQTree,
       Ty Go) : (lizzieLet32_3,MaskQTree) (go_4_goMux_data,Go) > [(lizzieLet32_3MQNone,Go),
                                                                  (lizzieLet32_3MQVal,Go),
                                                                  (lizzieLet32_3MQNode,Go)] */
  logic [2:0] go_4_goMux_data_onehotd;
  always_comb
    if ((lizzieLet32_3_d[0] && go_4_goMux_data_d[0]))
      unique case (lizzieLet32_3_d[2:1])
        2'd0: go_4_goMux_data_onehotd = 3'd1;
        2'd1: go_4_goMux_data_onehotd = 3'd2;
        2'd2: go_4_goMux_data_onehotd = 3'd4;
        default: go_4_goMux_data_onehotd = 3'd0;
      endcase
    else go_4_goMux_data_onehotd = 3'd0;
  assign lizzieLet32_3MQNone_d = go_4_goMux_data_onehotd[0];
  assign lizzieLet32_3MQVal_d = go_4_goMux_data_onehotd[1];
  assign lizzieLet32_3MQNode_d = go_4_goMux_data_onehotd[2];
  assign go_4_goMux_data_r = (| (go_4_goMux_data_onehotd & {lizzieLet32_3MQNode_r,
                                                            lizzieLet32_3MQVal_r,
                                                            lizzieLet32_3MQNone_r}));
  assign lizzieLet32_3_r = go_4_goMux_data_r;
  
  /* fork (Ty Go) : (lizzieLet32_3MQNone,Go) > [(lizzieLet32_3MQNone_1,Go),
                                           (lizzieLet32_3MQNone_2,Go)] */
  logic [1:0] lizzieLet32_3MQNone_emitted;
  logic [1:0] lizzieLet32_3MQNone_done;
  assign lizzieLet32_3MQNone_1_d = (lizzieLet32_3MQNone_d[0] && (! lizzieLet32_3MQNone_emitted[0]));
  assign lizzieLet32_3MQNone_2_d = (lizzieLet32_3MQNone_d[0] && (! lizzieLet32_3MQNone_emitted[1]));
  assign lizzieLet32_3MQNone_done = (lizzieLet32_3MQNone_emitted | ({lizzieLet32_3MQNone_2_d[0],
                                                                     lizzieLet32_3MQNone_1_d[0]} & {lizzieLet32_3MQNone_2_r,
                                                                                                    lizzieLet32_3MQNone_1_r}));
  assign lizzieLet32_3MQNone_r = (& lizzieLet32_3MQNone_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet32_3MQNone_emitted <= 2'd0;
    else
      lizzieLet32_3MQNone_emitted <= (lizzieLet32_3MQNone_r ? 2'd0 :
                                      lizzieLet32_3MQNone_done);
  
  /* dcon (Ty QTree_Bool,
      Dcon QNone_Bool) : [(lizzieLet32_3MQNone_1,Go)] > (lizzieLet32_3MQNone_1QNone_Bool,QTree_Bool) */
  assign lizzieLet32_3MQNone_1QNone_Bool_d = QNone_Bool_dc((& {lizzieLet32_3MQNone_1_d[0]}), lizzieLet32_3MQNone_1_d);
  assign {lizzieLet32_3MQNone_1_r} = {1 {(lizzieLet32_3MQNone_1QNone_Bool_r && lizzieLet32_3MQNone_1QNone_Bool_d[0])}};
  
  /* buf (Ty QTree_Bool) : (lizzieLet32_3MQNone_1QNone_Bool,QTree_Bool) > (lizzieLet33_1_argbuf,QTree_Bool) */
  QTree_Bool_t lizzieLet32_3MQNone_1QNone_Bool_bufchan_d;
  logic lizzieLet32_3MQNone_1QNone_Bool_bufchan_r;
  assign lizzieLet32_3MQNone_1QNone_Bool_r = ((! lizzieLet32_3MQNone_1QNone_Bool_bufchan_d[0]) || lizzieLet32_3MQNone_1QNone_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet32_3MQNone_1QNone_Bool_bufchan_d <= {66'd0, 1'd0};
    else
      if (lizzieLet32_3MQNone_1QNone_Bool_r)
        lizzieLet32_3MQNone_1QNone_Bool_bufchan_d <= lizzieLet32_3MQNone_1QNone_Bool_d;
  QTree_Bool_t lizzieLet32_3MQNone_1QNone_Bool_bufchan_buf;
  assign lizzieLet32_3MQNone_1QNone_Bool_bufchan_r = (! lizzieLet32_3MQNone_1QNone_Bool_bufchan_buf[0]);
  assign lizzieLet33_1_argbuf_d = (lizzieLet32_3MQNone_1QNone_Bool_bufchan_buf[0] ? lizzieLet32_3MQNone_1QNone_Bool_bufchan_buf :
                                   lizzieLet32_3MQNone_1QNone_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet32_3MQNone_1QNone_Bool_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((lizzieLet33_1_argbuf_r && lizzieLet32_3MQNone_1QNone_Bool_bufchan_buf[0]))
        lizzieLet32_3MQNone_1QNone_Bool_bufchan_buf <= {66'd0, 1'd0};
      else if (((! lizzieLet33_1_argbuf_r) && (! lizzieLet32_3MQNone_1QNone_Bool_bufchan_buf[0])))
        lizzieLet32_3MQNone_1QNone_Bool_bufchan_buf <= lizzieLet32_3MQNone_1QNone_Bool_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet32_3MQNone_2,Go) > (lizzieLet32_3MQNone_2_argbuf,Go) */
  Go_t lizzieLet32_3MQNone_2_bufchan_d;
  logic lizzieLet32_3MQNone_2_bufchan_r;
  assign lizzieLet32_3MQNone_2_r = ((! lizzieLet32_3MQNone_2_bufchan_d[0]) || lizzieLet32_3MQNone_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet32_3MQNone_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet32_3MQNone_2_r)
        lizzieLet32_3MQNone_2_bufchan_d <= lizzieLet32_3MQNone_2_d;
  Go_t lizzieLet32_3MQNone_2_bufchan_buf;
  assign lizzieLet32_3MQNone_2_bufchan_r = (! lizzieLet32_3MQNone_2_bufchan_buf[0]);
  assign lizzieLet32_3MQNone_2_argbuf_d = (lizzieLet32_3MQNone_2_bufchan_buf[0] ? lizzieLet32_3MQNone_2_bufchan_buf :
                                           lizzieLet32_3MQNone_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet32_3MQNone_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet32_3MQNone_2_argbuf_r && lizzieLet32_3MQNone_2_bufchan_buf[0]))
        lizzieLet32_3MQNone_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet32_3MQNone_2_argbuf_r) && (! lizzieLet32_3MQNone_2_bufchan_buf[0])))
        lizzieLet32_3MQNone_2_bufchan_buf <= lizzieLet32_3MQNone_2_bufchan_d;
  
  /* mergectrl (Ty C6,Ty Go) : [(lizzieLet32_3MQNone_2_argbuf,Go),
                           (lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool0_1_argbuf,Go),
                           (lizzieLet32_3MQVal_1_argbuf,Go),
                           (lizzieLet32_4MQNode_3QNone_Bool_2_argbuf,Go),
                           (lizzieLet32_4MQNode_3QVal_Bool_2_argbuf,Go),
                           (lizzieLet32_4MQNode_3QError_Bool_2_argbuf,Go)] > (go_11_goMux_choice,C6) (go_11_goMux_data,Go) */
  logic [5:0] lizzieLet32_3MQNone_2_argbuf_select_d;
  assign lizzieLet32_3MQNone_2_argbuf_select_d = ((| lizzieLet32_3MQNone_2_argbuf_select_q) ? lizzieLet32_3MQNone_2_argbuf_select_q :
                                                  (lizzieLet32_3MQNone_2_argbuf_d[0] ? 6'd1 :
                                                   (\lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool0_1_argbuf_d [0] ? 6'd2 :
                                                    (lizzieLet32_3MQVal_1_argbuf_d[0] ? 6'd4 :
                                                     (lizzieLet32_4MQNode_3QNone_Bool_2_argbuf_d[0] ? 6'd8 :
                                                      (lizzieLet32_4MQNode_3QVal_Bool_2_argbuf_d[0] ? 6'd16 :
                                                       (lizzieLet32_4MQNode_3QError_Bool_2_argbuf_d[0] ? 6'd32 :
                                                        6'd0)))))));
  logic [5:0] lizzieLet32_3MQNone_2_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet32_3MQNone_2_argbuf_select_q <= 6'd0;
    else
      lizzieLet32_3MQNone_2_argbuf_select_q <= (lizzieLet32_3MQNone_2_argbuf_done ? 6'd0 :
                                                lizzieLet32_3MQNone_2_argbuf_select_d);
  logic [1:0] lizzieLet32_3MQNone_2_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet32_3MQNone_2_argbuf_emit_q <= 2'd0;
    else
      lizzieLet32_3MQNone_2_argbuf_emit_q <= (lizzieLet32_3MQNone_2_argbuf_done ? 2'd0 :
                                              lizzieLet32_3MQNone_2_argbuf_emit_d);
  logic [1:0] lizzieLet32_3MQNone_2_argbuf_emit_d;
  assign lizzieLet32_3MQNone_2_argbuf_emit_d = (lizzieLet32_3MQNone_2_argbuf_emit_q | ({go_11_goMux_choice_d[0],
                                                                                        go_11_goMux_data_d[0]} & {go_11_goMux_choice_r,
                                                                                                                  go_11_goMux_data_r}));
  logic lizzieLet32_3MQNone_2_argbuf_done;
  assign lizzieLet32_3MQNone_2_argbuf_done = (& lizzieLet32_3MQNone_2_argbuf_emit_d);
  assign {lizzieLet32_4MQNode_3QError_Bool_2_argbuf_r,
          lizzieLet32_4MQNode_3QVal_Bool_2_argbuf_r,
          lizzieLet32_4MQNode_3QNone_Bool_2_argbuf_r,
          lizzieLet32_3MQVal_1_argbuf_r,
          \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool0_1_argbuf_r ,
          lizzieLet32_3MQNone_2_argbuf_r} = (lizzieLet32_3MQNone_2_argbuf_done ? lizzieLet32_3MQNone_2_argbuf_select_d :
                                             6'd0);
  assign go_11_goMux_data_d = ((lizzieLet32_3MQNone_2_argbuf_select_d[0] && (! lizzieLet32_3MQNone_2_argbuf_emit_q[0])) ? lizzieLet32_3MQNone_2_argbuf_d :
                               ((lizzieLet32_3MQNone_2_argbuf_select_d[1] && (! lizzieLet32_3MQNone_2_argbuf_emit_q[0])) ? \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool0_1_argbuf_d  :
                                ((lizzieLet32_3MQNone_2_argbuf_select_d[2] && (! lizzieLet32_3MQNone_2_argbuf_emit_q[0])) ? lizzieLet32_3MQVal_1_argbuf_d :
                                 ((lizzieLet32_3MQNone_2_argbuf_select_d[3] && (! lizzieLet32_3MQNone_2_argbuf_emit_q[0])) ? lizzieLet32_4MQNode_3QNone_Bool_2_argbuf_d :
                                  ((lizzieLet32_3MQNone_2_argbuf_select_d[4] && (! lizzieLet32_3MQNone_2_argbuf_emit_q[0])) ? lizzieLet32_4MQNode_3QVal_Bool_2_argbuf_d :
                                   ((lizzieLet32_3MQNone_2_argbuf_select_d[5] && (! lizzieLet32_3MQNone_2_argbuf_emit_q[0])) ? lizzieLet32_4MQNode_3QError_Bool_2_argbuf_d :
                                    1'd0))))));
  assign go_11_goMux_choice_d = ((lizzieLet32_3MQNone_2_argbuf_select_d[0] && (! lizzieLet32_3MQNone_2_argbuf_emit_q[1])) ? C1_6_dc(1'd1) :
                                 ((lizzieLet32_3MQNone_2_argbuf_select_d[1] && (! lizzieLet32_3MQNone_2_argbuf_emit_q[1])) ? C2_6_dc(1'd1) :
                                  ((lizzieLet32_3MQNone_2_argbuf_select_d[2] && (! lizzieLet32_3MQNone_2_argbuf_emit_q[1])) ? C3_6_dc(1'd1) :
                                   ((lizzieLet32_3MQNone_2_argbuf_select_d[3] && (! lizzieLet32_3MQNone_2_argbuf_emit_q[1])) ? C4_6_dc(1'd1) :
                                    ((lizzieLet32_3MQNone_2_argbuf_select_d[4] && (! lizzieLet32_3MQNone_2_argbuf_emit_q[1])) ? C5_6_dc(1'd1) :
                                     ((lizzieLet32_3MQNone_2_argbuf_select_d[5] && (! lizzieLet32_3MQNone_2_argbuf_emit_q[1])) ? C6_6_dc(1'd1) :
                                      {3'd0, 1'd0}))))));
  
  /* buf (Ty Go) : (lizzieLet32_3MQVal,Go) > (lizzieLet32_3MQVal_1_argbuf,Go) */
  Go_t lizzieLet32_3MQVal_bufchan_d;
  logic lizzieLet32_3MQVal_bufchan_r;
  assign lizzieLet32_3MQVal_r = ((! lizzieLet32_3MQVal_bufchan_d[0]) || lizzieLet32_3MQVal_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet32_3MQVal_bufchan_d <= 1'd0;
    else
      if (lizzieLet32_3MQVal_r)
        lizzieLet32_3MQVal_bufchan_d <= lizzieLet32_3MQVal_d;
  Go_t lizzieLet32_3MQVal_bufchan_buf;
  assign lizzieLet32_3MQVal_bufchan_r = (! lizzieLet32_3MQVal_bufchan_buf[0]);
  assign lizzieLet32_3MQVal_1_argbuf_d = (lizzieLet32_3MQVal_bufchan_buf[0] ? lizzieLet32_3MQVal_bufchan_buf :
                                          lizzieLet32_3MQVal_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet32_3MQVal_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet32_3MQVal_1_argbuf_r && lizzieLet32_3MQVal_bufchan_buf[0]))
        lizzieLet32_3MQVal_bufchan_buf <= 1'd0;
      else if (((! lizzieLet32_3MQVal_1_argbuf_r) && (! lizzieLet32_3MQVal_bufchan_buf[0])))
        lizzieLet32_3MQVal_bufchan_buf <= lizzieLet32_3MQVal_bufchan_d;
  
  /* demux (Ty MaskQTree,
       Ty QTree_Bool) : (lizzieLet32_4,MaskQTree) (readPointer_QTree_Boolq4'a8x_1_argbuf_rwb,QTree_Bool) > [(_24,QTree_Bool),
                                                                                                            (_23,QTree_Bool),
                                                                                                            (lizzieLet32_4MQNode,QTree_Bool)] */
  logic [2:0] \readPointer_QTree_Boolq4'a8x_1_argbuf_rwb_onehotd ;
  always_comb
    if ((lizzieLet32_4_d[0] && \readPointer_QTree_Boolq4'a8x_1_argbuf_rwb_d [0]))
      unique case (lizzieLet32_4_d[2:1])
        2'd0: \readPointer_QTree_Boolq4'a8x_1_argbuf_rwb_onehotd  = 3'd1;
        2'd1: \readPointer_QTree_Boolq4'a8x_1_argbuf_rwb_onehotd  = 3'd2;
        2'd2: \readPointer_QTree_Boolq4'a8x_1_argbuf_rwb_onehotd  = 3'd4;
        default:
          \readPointer_QTree_Boolq4'a8x_1_argbuf_rwb_onehotd  = 3'd0;
      endcase
    else \readPointer_QTree_Boolq4'a8x_1_argbuf_rwb_onehotd  = 3'd0;
  assign _24_d = {\readPointer_QTree_Boolq4'a8x_1_argbuf_rwb_d [66:1],
                  \readPointer_QTree_Boolq4'a8x_1_argbuf_rwb_onehotd [0]};
  assign _23_d = {\readPointer_QTree_Boolq4'a8x_1_argbuf_rwb_d [66:1],
                  \readPointer_QTree_Boolq4'a8x_1_argbuf_rwb_onehotd [1]};
  assign lizzieLet32_4MQNode_d = {\readPointer_QTree_Boolq4'a8x_1_argbuf_rwb_d [66:1],
                                  \readPointer_QTree_Boolq4'a8x_1_argbuf_rwb_onehotd [2]};
  assign \readPointer_QTree_Boolq4'a8x_1_argbuf_rwb_r  = (| (\readPointer_QTree_Boolq4'a8x_1_argbuf_rwb_onehotd  & {lizzieLet32_4MQNode_r,
                                                                                                                    _23_r,
                                                                                                                    _24_r}));
  assign lizzieLet32_4_r = \readPointer_QTree_Boolq4'a8x_1_argbuf_rwb_r ;
  
  /* fork (Ty QTree_Bool) : (lizzieLet32_4MQNode,QTree_Bool) > [(lizzieLet32_4MQNode_1,QTree_Bool),
                                                           (lizzieLet32_4MQNode_2,QTree_Bool),
                                                           (lizzieLet32_4MQNode_3,QTree_Bool),
                                                           (lizzieLet32_4MQNode_4,QTree_Bool),
                                                           (lizzieLet32_4MQNode_5,QTree_Bool),
                                                           (lizzieLet32_4MQNode_6,QTree_Bool),
                                                           (lizzieLet32_4MQNode_7,QTree_Bool),
                                                           (lizzieLet32_4MQNode_8,QTree_Bool)] */
  logic [7:0] lizzieLet32_4MQNode_emitted;
  logic [7:0] lizzieLet32_4MQNode_done;
  assign lizzieLet32_4MQNode_1_d = {lizzieLet32_4MQNode_d[66:1],
                                    (lizzieLet32_4MQNode_d[0] && (! lizzieLet32_4MQNode_emitted[0]))};
  assign lizzieLet32_4MQNode_2_d = {lizzieLet32_4MQNode_d[66:1],
                                    (lizzieLet32_4MQNode_d[0] && (! lizzieLet32_4MQNode_emitted[1]))};
  assign lizzieLet32_4MQNode_3_d = {lizzieLet32_4MQNode_d[66:1],
                                    (lizzieLet32_4MQNode_d[0] && (! lizzieLet32_4MQNode_emitted[2]))};
  assign lizzieLet32_4MQNode_4_d = {lizzieLet32_4MQNode_d[66:1],
                                    (lizzieLet32_4MQNode_d[0] && (! lizzieLet32_4MQNode_emitted[3]))};
  assign lizzieLet32_4MQNode_5_d = {lizzieLet32_4MQNode_d[66:1],
                                    (lizzieLet32_4MQNode_d[0] && (! lizzieLet32_4MQNode_emitted[4]))};
  assign lizzieLet32_4MQNode_6_d = {lizzieLet32_4MQNode_d[66:1],
                                    (lizzieLet32_4MQNode_d[0] && (! lizzieLet32_4MQNode_emitted[5]))};
  assign lizzieLet32_4MQNode_7_d = {lizzieLet32_4MQNode_d[66:1],
                                    (lizzieLet32_4MQNode_d[0] && (! lizzieLet32_4MQNode_emitted[6]))};
  assign lizzieLet32_4MQNode_8_d = {lizzieLet32_4MQNode_d[66:1],
                                    (lizzieLet32_4MQNode_d[0] && (! lizzieLet32_4MQNode_emitted[7]))};
  assign lizzieLet32_4MQNode_done = (lizzieLet32_4MQNode_emitted | ({lizzieLet32_4MQNode_8_d[0],
                                                                     lizzieLet32_4MQNode_7_d[0],
                                                                     lizzieLet32_4MQNode_6_d[0],
                                                                     lizzieLet32_4MQNode_5_d[0],
                                                                     lizzieLet32_4MQNode_4_d[0],
                                                                     lizzieLet32_4MQNode_3_d[0],
                                                                     lizzieLet32_4MQNode_2_d[0],
                                                                     lizzieLet32_4MQNode_1_d[0]} & {lizzieLet32_4MQNode_8_r,
                                                                                                    lizzieLet32_4MQNode_7_r,
                                                                                                    lizzieLet32_4MQNode_6_r,
                                                                                                    lizzieLet32_4MQNode_5_r,
                                                                                                    lizzieLet32_4MQNode_4_r,
                                                                                                    lizzieLet32_4MQNode_3_r,
                                                                                                    lizzieLet32_4MQNode_2_r,
                                                                                                    lizzieLet32_4MQNode_1_r}));
  assign lizzieLet32_4MQNode_r = (& lizzieLet32_4MQNode_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet32_4MQNode_emitted <= 8'd0;
    else
      lizzieLet32_4MQNode_emitted <= (lizzieLet32_4MQNode_r ? 8'd0 :
                                      lizzieLet32_4MQNode_done);
  
  /* destruct (Ty QTree_Bool,
          Dcon QNode_Bool) : (lizzieLet32_4MQNode_1QNode_Bool,QTree_Bool) > [(t1a8D_destruct,Pointer_QTree_Bool),
                                                                             (t2a8E_destruct,Pointer_QTree_Bool),
                                                                             (t3a8F_destruct,Pointer_QTree_Bool),
                                                                             (t4a8G_destruct,Pointer_QTree_Bool)] */
  logic [3:0] lizzieLet32_4MQNode_1QNode_Bool_emitted;
  logic [3:0] lizzieLet32_4MQNode_1QNode_Bool_done;
  assign t1a8D_destruct_d = {lizzieLet32_4MQNode_1QNode_Bool_d[18:3],
                             (lizzieLet32_4MQNode_1QNode_Bool_d[0] && (! lizzieLet32_4MQNode_1QNode_Bool_emitted[0]))};
  assign t2a8E_destruct_d = {lizzieLet32_4MQNode_1QNode_Bool_d[34:19],
                             (lizzieLet32_4MQNode_1QNode_Bool_d[0] && (! lizzieLet32_4MQNode_1QNode_Bool_emitted[1]))};
  assign t3a8F_destruct_d = {lizzieLet32_4MQNode_1QNode_Bool_d[50:35],
                             (lizzieLet32_4MQNode_1QNode_Bool_d[0] && (! lizzieLet32_4MQNode_1QNode_Bool_emitted[2]))};
  assign t4a8G_destruct_d = {lizzieLet32_4MQNode_1QNode_Bool_d[66:51],
                             (lizzieLet32_4MQNode_1QNode_Bool_d[0] && (! lizzieLet32_4MQNode_1QNode_Bool_emitted[3]))};
  assign lizzieLet32_4MQNode_1QNode_Bool_done = (lizzieLet32_4MQNode_1QNode_Bool_emitted | ({t4a8G_destruct_d[0],
                                                                                             t3a8F_destruct_d[0],
                                                                                             t2a8E_destruct_d[0],
                                                                                             t1a8D_destruct_d[0]} & {t4a8G_destruct_r,
                                                                                                                     t3a8F_destruct_r,
                                                                                                                     t2a8E_destruct_r,
                                                                                                                     t1a8D_destruct_r}));
  assign lizzieLet32_4MQNode_1QNode_Bool_r = (& lizzieLet32_4MQNode_1QNode_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet32_4MQNode_1QNode_Bool_emitted <= 4'd0;
    else
      lizzieLet32_4MQNode_1QNode_Bool_emitted <= (lizzieLet32_4MQNode_1QNode_Bool_r ? 4'd0 :
                                                  lizzieLet32_4MQNode_1QNode_Bool_done);
  
  /* demux (Ty QTree_Bool,
       Ty QTree_Bool) : (lizzieLet32_4MQNode_2,QTree_Bool) (lizzieLet32_4MQNode_1,QTree_Bool) > [(_22,QTree_Bool),
                                                                                                 (_21,QTree_Bool),
                                                                                                 (lizzieLet32_4MQNode_1QNode_Bool,QTree_Bool),
                                                                                                 (_20,QTree_Bool)] */
  logic [3:0] lizzieLet32_4MQNode_1_onehotd;
  always_comb
    if ((lizzieLet32_4MQNode_2_d[0] && lizzieLet32_4MQNode_1_d[0]))
      unique case (lizzieLet32_4MQNode_2_d[2:1])
        2'd0: lizzieLet32_4MQNode_1_onehotd = 4'd1;
        2'd1: lizzieLet32_4MQNode_1_onehotd = 4'd2;
        2'd2: lizzieLet32_4MQNode_1_onehotd = 4'd4;
        2'd3: lizzieLet32_4MQNode_1_onehotd = 4'd8;
        default: lizzieLet32_4MQNode_1_onehotd = 4'd0;
      endcase
    else lizzieLet32_4MQNode_1_onehotd = 4'd0;
  assign _22_d = {lizzieLet32_4MQNode_1_d[66:1],
                  lizzieLet32_4MQNode_1_onehotd[0]};
  assign _21_d = {lizzieLet32_4MQNode_1_d[66:1],
                  lizzieLet32_4MQNode_1_onehotd[1]};
  assign lizzieLet32_4MQNode_1QNode_Bool_d = {lizzieLet32_4MQNode_1_d[66:1],
                                              lizzieLet32_4MQNode_1_onehotd[2]};
  assign _20_d = {lizzieLet32_4MQNode_1_d[66:1],
                  lizzieLet32_4MQNode_1_onehotd[3]};
  assign lizzieLet32_4MQNode_1_r = (| (lizzieLet32_4MQNode_1_onehotd & {_20_r,
                                                                        lizzieLet32_4MQNode_1QNode_Bool_r,
                                                                        _21_r,
                                                                        _22_r}));
  assign lizzieLet32_4MQNode_2_r = lizzieLet32_4MQNode_1_r;
  
  /* demux (Ty QTree_Bool,
       Ty Go) : (lizzieLet32_4MQNode_3,QTree_Bool) (lizzieLet32_3MQNode,Go) > [(lizzieLet32_4MQNode_3QNone_Bool,Go),
                                                                               (lizzieLet32_4MQNode_3QVal_Bool,Go),
                                                                               (lizzieLet32_4MQNode_3QNode_Bool,Go),
                                                                               (lizzieLet32_4MQNode_3QError_Bool,Go)] */
  logic [3:0] lizzieLet32_3MQNode_onehotd;
  always_comb
    if ((lizzieLet32_4MQNode_3_d[0] && lizzieLet32_3MQNode_d[0]))
      unique case (lizzieLet32_4MQNode_3_d[2:1])
        2'd0: lizzieLet32_3MQNode_onehotd = 4'd1;
        2'd1: lizzieLet32_3MQNode_onehotd = 4'd2;
        2'd2: lizzieLet32_3MQNode_onehotd = 4'd4;
        2'd3: lizzieLet32_3MQNode_onehotd = 4'd8;
        default: lizzieLet32_3MQNode_onehotd = 4'd0;
      endcase
    else lizzieLet32_3MQNode_onehotd = 4'd0;
  assign lizzieLet32_4MQNode_3QNone_Bool_d = lizzieLet32_3MQNode_onehotd[0];
  assign lizzieLet32_4MQNode_3QVal_Bool_d = lizzieLet32_3MQNode_onehotd[1];
  assign lizzieLet32_4MQNode_3QNode_Bool_d = lizzieLet32_3MQNode_onehotd[2];
  assign lizzieLet32_4MQNode_3QError_Bool_d = lizzieLet32_3MQNode_onehotd[3];
  assign lizzieLet32_3MQNode_r = (| (lizzieLet32_3MQNode_onehotd & {lizzieLet32_4MQNode_3QError_Bool_r,
                                                                    lizzieLet32_4MQNode_3QNode_Bool_r,
                                                                    lizzieLet32_4MQNode_3QVal_Bool_r,
                                                                    lizzieLet32_4MQNode_3QNone_Bool_r}));
  assign lizzieLet32_4MQNode_3_r = lizzieLet32_3MQNode_r;
  
  /* fork (Ty Go) : (lizzieLet32_4MQNode_3QError_Bool,Go) > [(lizzieLet32_4MQNode_3QError_Bool_1,Go),
                                                        (lizzieLet32_4MQNode_3QError_Bool_2,Go)] */
  logic [1:0] lizzieLet32_4MQNode_3QError_Bool_emitted;
  logic [1:0] lizzieLet32_4MQNode_3QError_Bool_done;
  assign lizzieLet32_4MQNode_3QError_Bool_1_d = (lizzieLet32_4MQNode_3QError_Bool_d[0] && (! lizzieLet32_4MQNode_3QError_Bool_emitted[0]));
  assign lizzieLet32_4MQNode_3QError_Bool_2_d = (lizzieLet32_4MQNode_3QError_Bool_d[0] && (! lizzieLet32_4MQNode_3QError_Bool_emitted[1]));
  assign lizzieLet32_4MQNode_3QError_Bool_done = (lizzieLet32_4MQNode_3QError_Bool_emitted | ({lizzieLet32_4MQNode_3QError_Bool_2_d[0],
                                                                                               lizzieLet32_4MQNode_3QError_Bool_1_d[0]} & {lizzieLet32_4MQNode_3QError_Bool_2_r,
                                                                                                                                           lizzieLet32_4MQNode_3QError_Bool_1_r}));
  assign lizzieLet32_4MQNode_3QError_Bool_r = (& lizzieLet32_4MQNode_3QError_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet32_4MQNode_3QError_Bool_emitted <= 2'd0;
    else
      lizzieLet32_4MQNode_3QError_Bool_emitted <= (lizzieLet32_4MQNode_3QError_Bool_r ? 2'd0 :
                                                   lizzieLet32_4MQNode_3QError_Bool_done);
  
  /* dcon (Ty QTree_Bool,
      Dcon QError_Bool) : [(lizzieLet32_4MQNode_3QError_Bool_1,Go)] > (lizzieLet32_4MQNode_3QError_Bool_1QError_Bool,QTree_Bool) */
  assign lizzieLet32_4MQNode_3QError_Bool_1QError_Bool_d = QError_Bool_dc((& {lizzieLet32_4MQNode_3QError_Bool_1_d[0]}), lizzieLet32_4MQNode_3QError_Bool_1_d);
  assign {lizzieLet32_4MQNode_3QError_Bool_1_r} = {1 {(lizzieLet32_4MQNode_3QError_Bool_1QError_Bool_r && lizzieLet32_4MQNode_3QError_Bool_1QError_Bool_d[0])}};
  
  /* buf (Ty QTree_Bool) : (lizzieLet32_4MQNode_3QError_Bool_1QError_Bool,QTree_Bool) > (lizzieLet38_1_argbuf,QTree_Bool) */
  QTree_Bool_t lizzieLet32_4MQNode_3QError_Bool_1QError_Bool_bufchan_d;
  logic lizzieLet32_4MQNode_3QError_Bool_1QError_Bool_bufchan_r;
  assign lizzieLet32_4MQNode_3QError_Bool_1QError_Bool_r = ((! lizzieLet32_4MQNode_3QError_Bool_1QError_Bool_bufchan_d[0]) || lizzieLet32_4MQNode_3QError_Bool_1QError_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet32_4MQNode_3QError_Bool_1QError_Bool_bufchan_d <= {66'd0,
                                                                  1'd0};
    else
      if (lizzieLet32_4MQNode_3QError_Bool_1QError_Bool_r)
        lizzieLet32_4MQNode_3QError_Bool_1QError_Bool_bufchan_d <= lizzieLet32_4MQNode_3QError_Bool_1QError_Bool_d;
  QTree_Bool_t lizzieLet32_4MQNode_3QError_Bool_1QError_Bool_bufchan_buf;
  assign lizzieLet32_4MQNode_3QError_Bool_1QError_Bool_bufchan_r = (! lizzieLet32_4MQNode_3QError_Bool_1QError_Bool_bufchan_buf[0]);
  assign lizzieLet38_1_argbuf_d = (lizzieLet32_4MQNode_3QError_Bool_1QError_Bool_bufchan_buf[0] ? lizzieLet32_4MQNode_3QError_Bool_1QError_Bool_bufchan_buf :
                                   lizzieLet32_4MQNode_3QError_Bool_1QError_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet32_4MQNode_3QError_Bool_1QError_Bool_bufchan_buf <= {66'd0,
                                                                    1'd0};
    else
      if ((lizzieLet38_1_argbuf_r && lizzieLet32_4MQNode_3QError_Bool_1QError_Bool_bufchan_buf[0]))
        lizzieLet32_4MQNode_3QError_Bool_1QError_Bool_bufchan_buf <= {66'd0,
                                                                      1'd0};
      else if (((! lizzieLet38_1_argbuf_r) && (! lizzieLet32_4MQNode_3QError_Bool_1QError_Bool_bufchan_buf[0])))
        lizzieLet32_4MQNode_3QError_Bool_1QError_Bool_bufchan_buf <= lizzieLet32_4MQNode_3QError_Bool_1QError_Bool_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet32_4MQNode_3QError_Bool_2,Go) > (lizzieLet32_4MQNode_3QError_Bool_2_argbuf,Go) */
  Go_t lizzieLet32_4MQNode_3QError_Bool_2_bufchan_d;
  logic lizzieLet32_4MQNode_3QError_Bool_2_bufchan_r;
  assign lizzieLet32_4MQNode_3QError_Bool_2_r = ((! lizzieLet32_4MQNode_3QError_Bool_2_bufchan_d[0]) || lizzieLet32_4MQNode_3QError_Bool_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet32_4MQNode_3QError_Bool_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet32_4MQNode_3QError_Bool_2_r)
        lizzieLet32_4MQNode_3QError_Bool_2_bufchan_d <= lizzieLet32_4MQNode_3QError_Bool_2_d;
  Go_t lizzieLet32_4MQNode_3QError_Bool_2_bufchan_buf;
  assign lizzieLet32_4MQNode_3QError_Bool_2_bufchan_r = (! lizzieLet32_4MQNode_3QError_Bool_2_bufchan_buf[0]);
  assign lizzieLet32_4MQNode_3QError_Bool_2_argbuf_d = (lizzieLet32_4MQNode_3QError_Bool_2_bufchan_buf[0] ? lizzieLet32_4MQNode_3QError_Bool_2_bufchan_buf :
                                                        lizzieLet32_4MQNode_3QError_Bool_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet32_4MQNode_3QError_Bool_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet32_4MQNode_3QError_Bool_2_argbuf_r && lizzieLet32_4MQNode_3QError_Bool_2_bufchan_buf[0]))
        lizzieLet32_4MQNode_3QError_Bool_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet32_4MQNode_3QError_Bool_2_argbuf_r) && (! lizzieLet32_4MQNode_3QError_Bool_2_bufchan_buf[0])))
        lizzieLet32_4MQNode_3QError_Bool_2_bufchan_buf <= lizzieLet32_4MQNode_3QError_Bool_2_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet32_4MQNode_3QNode_Bool,Go) > (lizzieLet32_4MQNode_3QNode_Bool_1_argbuf,Go) */
  Go_t lizzieLet32_4MQNode_3QNode_Bool_bufchan_d;
  logic lizzieLet32_4MQNode_3QNode_Bool_bufchan_r;
  assign lizzieLet32_4MQNode_3QNode_Bool_r = ((! lizzieLet32_4MQNode_3QNode_Bool_bufchan_d[0]) || lizzieLet32_4MQNode_3QNode_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet32_4MQNode_3QNode_Bool_bufchan_d <= 1'd0;
    else
      if (lizzieLet32_4MQNode_3QNode_Bool_r)
        lizzieLet32_4MQNode_3QNode_Bool_bufchan_d <= lizzieLet32_4MQNode_3QNode_Bool_d;
  Go_t lizzieLet32_4MQNode_3QNode_Bool_bufchan_buf;
  assign lizzieLet32_4MQNode_3QNode_Bool_bufchan_r = (! lizzieLet32_4MQNode_3QNode_Bool_bufchan_buf[0]);
  assign lizzieLet32_4MQNode_3QNode_Bool_1_argbuf_d = (lizzieLet32_4MQNode_3QNode_Bool_bufchan_buf[0] ? lizzieLet32_4MQNode_3QNode_Bool_bufchan_buf :
                                                       lizzieLet32_4MQNode_3QNode_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet32_4MQNode_3QNode_Bool_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet32_4MQNode_3QNode_Bool_1_argbuf_r && lizzieLet32_4MQNode_3QNode_Bool_bufchan_buf[0]))
        lizzieLet32_4MQNode_3QNode_Bool_bufchan_buf <= 1'd0;
      else if (((! lizzieLet32_4MQNode_3QNode_Bool_1_argbuf_r) && (! lizzieLet32_4MQNode_3QNode_Bool_bufchan_buf[0])))
        lizzieLet32_4MQNode_3QNode_Bool_bufchan_buf <= lizzieLet32_4MQNode_3QNode_Bool_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet32_4MQNode_3QNone_Bool,Go) > [(lizzieLet32_4MQNode_3QNone_Bool_1,Go),
                                                       (lizzieLet32_4MQNode_3QNone_Bool_2,Go)] */
  logic [1:0] lizzieLet32_4MQNode_3QNone_Bool_emitted;
  logic [1:0] lizzieLet32_4MQNode_3QNone_Bool_done;
  assign lizzieLet32_4MQNode_3QNone_Bool_1_d = (lizzieLet32_4MQNode_3QNone_Bool_d[0] && (! lizzieLet32_4MQNode_3QNone_Bool_emitted[0]));
  assign lizzieLet32_4MQNode_3QNone_Bool_2_d = (lizzieLet32_4MQNode_3QNone_Bool_d[0] && (! lizzieLet32_4MQNode_3QNone_Bool_emitted[1]));
  assign lizzieLet32_4MQNode_3QNone_Bool_done = (lizzieLet32_4MQNode_3QNone_Bool_emitted | ({lizzieLet32_4MQNode_3QNone_Bool_2_d[0],
                                                                                             lizzieLet32_4MQNode_3QNone_Bool_1_d[0]} & {lizzieLet32_4MQNode_3QNone_Bool_2_r,
                                                                                                                                        lizzieLet32_4MQNode_3QNone_Bool_1_r}));
  assign lizzieLet32_4MQNode_3QNone_Bool_r = (& lizzieLet32_4MQNode_3QNone_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet32_4MQNode_3QNone_Bool_emitted <= 2'd0;
    else
      lizzieLet32_4MQNode_3QNone_Bool_emitted <= (lizzieLet32_4MQNode_3QNone_Bool_r ? 2'd0 :
                                                  lizzieLet32_4MQNode_3QNone_Bool_done);
  
  /* dcon (Ty QTree_Bool,
      Dcon QNone_Bool) : [(lizzieLet32_4MQNode_3QNone_Bool_1,Go)] > (lizzieLet32_4MQNode_3QNone_Bool_1QNone_Bool,QTree_Bool) */
  assign lizzieLet32_4MQNode_3QNone_Bool_1QNone_Bool_d = QNone_Bool_dc((& {lizzieLet32_4MQNode_3QNone_Bool_1_d[0]}), lizzieLet32_4MQNode_3QNone_Bool_1_d);
  assign {lizzieLet32_4MQNode_3QNone_Bool_1_r} = {1 {(lizzieLet32_4MQNode_3QNone_Bool_1QNone_Bool_r && lizzieLet32_4MQNode_3QNone_Bool_1QNone_Bool_d[0])}};
  
  /* buf (Ty QTree_Bool) : (lizzieLet32_4MQNode_3QNone_Bool_1QNone_Bool,QTree_Bool) > (lizzieLet35_1_argbuf,QTree_Bool) */
  QTree_Bool_t lizzieLet32_4MQNode_3QNone_Bool_1QNone_Bool_bufchan_d;
  logic lizzieLet32_4MQNode_3QNone_Bool_1QNone_Bool_bufchan_r;
  assign lizzieLet32_4MQNode_3QNone_Bool_1QNone_Bool_r = ((! lizzieLet32_4MQNode_3QNone_Bool_1QNone_Bool_bufchan_d[0]) || lizzieLet32_4MQNode_3QNone_Bool_1QNone_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet32_4MQNode_3QNone_Bool_1QNone_Bool_bufchan_d <= {66'd0,
                                                                1'd0};
    else
      if (lizzieLet32_4MQNode_3QNone_Bool_1QNone_Bool_r)
        lizzieLet32_4MQNode_3QNone_Bool_1QNone_Bool_bufchan_d <= lizzieLet32_4MQNode_3QNone_Bool_1QNone_Bool_d;
  QTree_Bool_t lizzieLet32_4MQNode_3QNone_Bool_1QNone_Bool_bufchan_buf;
  assign lizzieLet32_4MQNode_3QNone_Bool_1QNone_Bool_bufchan_r = (! lizzieLet32_4MQNode_3QNone_Bool_1QNone_Bool_bufchan_buf[0]);
  assign lizzieLet35_1_argbuf_d = (lizzieLet32_4MQNode_3QNone_Bool_1QNone_Bool_bufchan_buf[0] ? lizzieLet32_4MQNode_3QNone_Bool_1QNone_Bool_bufchan_buf :
                                   lizzieLet32_4MQNode_3QNone_Bool_1QNone_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet32_4MQNode_3QNone_Bool_1QNone_Bool_bufchan_buf <= {66'd0,
                                                                  1'd0};
    else
      if ((lizzieLet35_1_argbuf_r && lizzieLet32_4MQNode_3QNone_Bool_1QNone_Bool_bufchan_buf[0]))
        lizzieLet32_4MQNode_3QNone_Bool_1QNone_Bool_bufchan_buf <= {66'd0,
                                                                    1'd0};
      else if (((! lizzieLet35_1_argbuf_r) && (! lizzieLet32_4MQNode_3QNone_Bool_1QNone_Bool_bufchan_buf[0])))
        lizzieLet32_4MQNode_3QNone_Bool_1QNone_Bool_bufchan_buf <= lizzieLet32_4MQNode_3QNone_Bool_1QNone_Bool_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet32_4MQNode_3QNone_Bool_2,Go) > (lizzieLet32_4MQNode_3QNone_Bool_2_argbuf,Go) */
  Go_t lizzieLet32_4MQNode_3QNone_Bool_2_bufchan_d;
  logic lizzieLet32_4MQNode_3QNone_Bool_2_bufchan_r;
  assign lizzieLet32_4MQNode_3QNone_Bool_2_r = ((! lizzieLet32_4MQNode_3QNone_Bool_2_bufchan_d[0]) || lizzieLet32_4MQNode_3QNone_Bool_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet32_4MQNode_3QNone_Bool_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet32_4MQNode_3QNone_Bool_2_r)
        lizzieLet32_4MQNode_3QNone_Bool_2_bufchan_d <= lizzieLet32_4MQNode_3QNone_Bool_2_d;
  Go_t lizzieLet32_4MQNode_3QNone_Bool_2_bufchan_buf;
  assign lizzieLet32_4MQNode_3QNone_Bool_2_bufchan_r = (! lizzieLet32_4MQNode_3QNone_Bool_2_bufchan_buf[0]);
  assign lizzieLet32_4MQNode_3QNone_Bool_2_argbuf_d = (lizzieLet32_4MQNode_3QNone_Bool_2_bufchan_buf[0] ? lizzieLet32_4MQNode_3QNone_Bool_2_bufchan_buf :
                                                       lizzieLet32_4MQNode_3QNone_Bool_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet32_4MQNode_3QNone_Bool_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet32_4MQNode_3QNone_Bool_2_argbuf_r && lizzieLet32_4MQNode_3QNone_Bool_2_bufchan_buf[0]))
        lizzieLet32_4MQNode_3QNone_Bool_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet32_4MQNode_3QNone_Bool_2_argbuf_r) && (! lizzieLet32_4MQNode_3QNone_Bool_2_bufchan_buf[0])))
        lizzieLet32_4MQNode_3QNone_Bool_2_bufchan_buf <= lizzieLet32_4MQNode_3QNone_Bool_2_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet32_4MQNode_3QVal_Bool,Go) > [(lizzieLet32_4MQNode_3QVal_Bool_1,Go),
                                                      (lizzieLet32_4MQNode_3QVal_Bool_2,Go)] */
  logic [1:0] lizzieLet32_4MQNode_3QVal_Bool_emitted;
  logic [1:0] lizzieLet32_4MQNode_3QVal_Bool_done;
  assign lizzieLet32_4MQNode_3QVal_Bool_1_d = (lizzieLet32_4MQNode_3QVal_Bool_d[0] && (! lizzieLet32_4MQNode_3QVal_Bool_emitted[0]));
  assign lizzieLet32_4MQNode_3QVal_Bool_2_d = (lizzieLet32_4MQNode_3QVal_Bool_d[0] && (! lizzieLet32_4MQNode_3QVal_Bool_emitted[1]));
  assign lizzieLet32_4MQNode_3QVal_Bool_done = (lizzieLet32_4MQNode_3QVal_Bool_emitted | ({lizzieLet32_4MQNode_3QVal_Bool_2_d[0],
                                                                                           lizzieLet32_4MQNode_3QVal_Bool_1_d[0]} & {lizzieLet32_4MQNode_3QVal_Bool_2_r,
                                                                                                                                     lizzieLet32_4MQNode_3QVal_Bool_1_r}));
  assign lizzieLet32_4MQNode_3QVal_Bool_r = (& lizzieLet32_4MQNode_3QVal_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet32_4MQNode_3QVal_Bool_emitted <= 2'd0;
    else
      lizzieLet32_4MQNode_3QVal_Bool_emitted <= (lizzieLet32_4MQNode_3QVal_Bool_r ? 2'd0 :
                                                 lizzieLet32_4MQNode_3QVal_Bool_done);
  
  /* dcon (Ty QTree_Bool,
      Dcon QError_Bool) : [(lizzieLet32_4MQNode_3QVal_Bool_1,Go)] > (lizzieLet32_4MQNode_3QVal_Bool_1QError_Bool,QTree_Bool) */
  assign lizzieLet32_4MQNode_3QVal_Bool_1QError_Bool_d = QError_Bool_dc((& {lizzieLet32_4MQNode_3QVal_Bool_1_d[0]}), lizzieLet32_4MQNode_3QVal_Bool_1_d);
  assign {lizzieLet32_4MQNode_3QVal_Bool_1_r} = {1 {(lizzieLet32_4MQNode_3QVal_Bool_1QError_Bool_r && lizzieLet32_4MQNode_3QVal_Bool_1QError_Bool_d[0])}};
  
  /* buf (Ty QTree_Bool) : (lizzieLet32_4MQNode_3QVal_Bool_1QError_Bool,QTree_Bool) > (lizzieLet36_1_argbuf,QTree_Bool) */
  QTree_Bool_t lizzieLet32_4MQNode_3QVal_Bool_1QError_Bool_bufchan_d;
  logic lizzieLet32_4MQNode_3QVal_Bool_1QError_Bool_bufchan_r;
  assign lizzieLet32_4MQNode_3QVal_Bool_1QError_Bool_r = ((! lizzieLet32_4MQNode_3QVal_Bool_1QError_Bool_bufchan_d[0]) || lizzieLet32_4MQNode_3QVal_Bool_1QError_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet32_4MQNode_3QVal_Bool_1QError_Bool_bufchan_d <= {66'd0,
                                                                1'd0};
    else
      if (lizzieLet32_4MQNode_3QVal_Bool_1QError_Bool_r)
        lizzieLet32_4MQNode_3QVal_Bool_1QError_Bool_bufchan_d <= lizzieLet32_4MQNode_3QVal_Bool_1QError_Bool_d;
  QTree_Bool_t lizzieLet32_4MQNode_3QVal_Bool_1QError_Bool_bufchan_buf;
  assign lizzieLet32_4MQNode_3QVal_Bool_1QError_Bool_bufchan_r = (! lizzieLet32_4MQNode_3QVal_Bool_1QError_Bool_bufchan_buf[0]);
  assign lizzieLet36_1_argbuf_d = (lizzieLet32_4MQNode_3QVal_Bool_1QError_Bool_bufchan_buf[0] ? lizzieLet32_4MQNode_3QVal_Bool_1QError_Bool_bufchan_buf :
                                   lizzieLet32_4MQNode_3QVal_Bool_1QError_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet32_4MQNode_3QVal_Bool_1QError_Bool_bufchan_buf <= {66'd0,
                                                                  1'd0};
    else
      if ((lizzieLet36_1_argbuf_r && lizzieLet32_4MQNode_3QVal_Bool_1QError_Bool_bufchan_buf[0]))
        lizzieLet32_4MQNode_3QVal_Bool_1QError_Bool_bufchan_buf <= {66'd0,
                                                                    1'd0};
      else if (((! lizzieLet36_1_argbuf_r) && (! lizzieLet32_4MQNode_3QVal_Bool_1QError_Bool_bufchan_buf[0])))
        lizzieLet32_4MQNode_3QVal_Bool_1QError_Bool_bufchan_buf <= lizzieLet32_4MQNode_3QVal_Bool_1QError_Bool_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet32_4MQNode_3QVal_Bool_2,Go) > (lizzieLet32_4MQNode_3QVal_Bool_2_argbuf,Go) */
  Go_t lizzieLet32_4MQNode_3QVal_Bool_2_bufchan_d;
  logic lizzieLet32_4MQNode_3QVal_Bool_2_bufchan_r;
  assign lizzieLet32_4MQNode_3QVal_Bool_2_r = ((! lizzieLet32_4MQNode_3QVal_Bool_2_bufchan_d[0]) || lizzieLet32_4MQNode_3QVal_Bool_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet32_4MQNode_3QVal_Bool_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet32_4MQNode_3QVal_Bool_2_r)
        lizzieLet32_4MQNode_3QVal_Bool_2_bufchan_d <= lizzieLet32_4MQNode_3QVal_Bool_2_d;
  Go_t lizzieLet32_4MQNode_3QVal_Bool_2_bufchan_buf;
  assign lizzieLet32_4MQNode_3QVal_Bool_2_bufchan_r = (! lizzieLet32_4MQNode_3QVal_Bool_2_bufchan_buf[0]);
  assign lizzieLet32_4MQNode_3QVal_Bool_2_argbuf_d = (lizzieLet32_4MQNode_3QVal_Bool_2_bufchan_buf[0] ? lizzieLet32_4MQNode_3QVal_Bool_2_bufchan_buf :
                                                      lizzieLet32_4MQNode_3QVal_Bool_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet32_4MQNode_3QVal_Bool_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet32_4MQNode_3QVal_Bool_2_argbuf_r && lizzieLet32_4MQNode_3QVal_Bool_2_bufchan_buf[0]))
        lizzieLet32_4MQNode_3QVal_Bool_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet32_4MQNode_3QVal_Bool_2_argbuf_r) && (! lizzieLet32_4MQNode_3QVal_Bool_2_bufchan_buf[0])))
        lizzieLet32_4MQNode_3QVal_Bool_2_bufchan_buf <= lizzieLet32_4MQNode_3QVal_Bool_2_bufchan_d;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_CTf'''''''''_f'''''''''_Bool) : (lizzieLet32_4MQNode_4,QTree_Bool) (lizzieLet32_6MQNode,Pointer_CTf'''''''''_f'''''''''_Bool) > [(lizzieLet32_4MQNode_4QNone_Bool,Pointer_CTf'''''''''_f'''''''''_Bool),
                                                                                                                                                   (lizzieLet32_4MQNode_4QVal_Bool,Pointer_CTf'''''''''_f'''''''''_Bool),
                                                                                                                                                   (lizzieLet32_4MQNode_4QNode_Bool,Pointer_CTf'''''''''_f'''''''''_Bool),
                                                                                                                                                   (lizzieLet32_4MQNode_4QError_Bool,Pointer_CTf'''''''''_f'''''''''_Bool)] */
  logic [3:0] lizzieLet32_6MQNode_onehotd;
  always_comb
    if ((lizzieLet32_4MQNode_4_d[0] && lizzieLet32_6MQNode_d[0]))
      unique case (lizzieLet32_4MQNode_4_d[2:1])
        2'd0: lizzieLet32_6MQNode_onehotd = 4'd1;
        2'd1: lizzieLet32_6MQNode_onehotd = 4'd2;
        2'd2: lizzieLet32_6MQNode_onehotd = 4'd4;
        2'd3: lizzieLet32_6MQNode_onehotd = 4'd8;
        default: lizzieLet32_6MQNode_onehotd = 4'd0;
      endcase
    else lizzieLet32_6MQNode_onehotd = 4'd0;
  assign lizzieLet32_4MQNode_4QNone_Bool_d = {lizzieLet32_6MQNode_d[16:1],
                                              lizzieLet32_6MQNode_onehotd[0]};
  assign lizzieLet32_4MQNode_4QVal_Bool_d = {lizzieLet32_6MQNode_d[16:1],
                                             lizzieLet32_6MQNode_onehotd[1]};
  assign lizzieLet32_4MQNode_4QNode_Bool_d = {lizzieLet32_6MQNode_d[16:1],
                                              lizzieLet32_6MQNode_onehotd[2]};
  assign lizzieLet32_4MQNode_4QError_Bool_d = {lizzieLet32_6MQNode_d[16:1],
                                               lizzieLet32_6MQNode_onehotd[3]};
  assign lizzieLet32_6MQNode_r = (| (lizzieLet32_6MQNode_onehotd & {lizzieLet32_4MQNode_4QError_Bool_r,
                                                                    lizzieLet32_4MQNode_4QNode_Bool_r,
                                                                    lizzieLet32_4MQNode_4QVal_Bool_r,
                                                                    lizzieLet32_4MQNode_4QNone_Bool_r}));
  assign lizzieLet32_4MQNode_4_r = lizzieLet32_6MQNode_r;
  
  /* buf (Ty Pointer_CTf'''''''''_f'''''''''_Bool) : (lizzieLet32_4MQNode_4QError_Bool,Pointer_CTf'''''''''_f'''''''''_Bool) > (lizzieLet32_4MQNode_4QError_Bool_1_argbuf,Pointer_CTf'''''''''_f'''''''''_Bool) */
  \Pointer_CTf'''''''''_f'''''''''_Bool_t  lizzieLet32_4MQNode_4QError_Bool_bufchan_d;
  logic lizzieLet32_4MQNode_4QError_Bool_bufchan_r;
  assign lizzieLet32_4MQNode_4QError_Bool_r = ((! lizzieLet32_4MQNode_4QError_Bool_bufchan_d[0]) || lizzieLet32_4MQNode_4QError_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet32_4MQNode_4QError_Bool_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet32_4MQNode_4QError_Bool_r)
        lizzieLet32_4MQNode_4QError_Bool_bufchan_d <= lizzieLet32_4MQNode_4QError_Bool_d;
  \Pointer_CTf'''''''''_f'''''''''_Bool_t  lizzieLet32_4MQNode_4QError_Bool_bufchan_buf;
  assign lizzieLet32_4MQNode_4QError_Bool_bufchan_r = (! lizzieLet32_4MQNode_4QError_Bool_bufchan_buf[0]);
  assign lizzieLet32_4MQNode_4QError_Bool_1_argbuf_d = (lizzieLet32_4MQNode_4QError_Bool_bufchan_buf[0] ? lizzieLet32_4MQNode_4QError_Bool_bufchan_buf :
                                                        lizzieLet32_4MQNode_4QError_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet32_4MQNode_4QError_Bool_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet32_4MQNode_4QError_Bool_1_argbuf_r && lizzieLet32_4MQNode_4QError_Bool_bufchan_buf[0]))
        lizzieLet32_4MQNode_4QError_Bool_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet32_4MQNode_4QError_Bool_1_argbuf_r) && (! lizzieLet32_4MQNode_4QError_Bool_bufchan_buf[0])))
        lizzieLet32_4MQNode_4QError_Bool_bufchan_buf <= lizzieLet32_4MQNode_4QError_Bool_bufchan_d;
  
  /* dcon (Ty CTf'''''''''_f'''''''''_Bool,
      Dcon Lcall_f'''''''''_f'''''''''_Bool3) : [(lizzieLet32_4MQNode_4QNode_Bool,Pointer_CTf'''''''''_f'''''''''_Bool),
                                                 (lizzieLet32_4MQNode_5QNode_Bool,Pointer_MaskQTree),
                                                 (t1a8D_destruct,Pointer_QTree_Bool),
                                                 (lizzieLet32_4MQNode_6QNode_Bool,Pointer_MaskQTree),
                                                 (t2a8E_destruct,Pointer_QTree_Bool),
                                                 (lizzieLet32_4MQNode_7QNode_Bool,Pointer_MaskQTree),
                                                 (t3a8F_destruct,Pointer_QTree_Bool)] > (lizzieLet32_4MQNode_4QNode_Bool_1lizzieLet32_4MQNode_5QNode_Bool_1t1a8D_1lizzieLet32_4MQNode_6QNode_Bool_1t2a8E_1lizzieLet32_4MQNode_7QNode_Bool_1t3a8F_1Lcall_f'''''''''_f'''''''''_Bool3,CTf'''''''''_f'''''''''_Bool) */
  assign \lizzieLet32_4MQNode_4QNode_Bool_1lizzieLet32_4MQNode_5QNode_Bool_1t1a8D_1lizzieLet32_4MQNode_6QNode_Bool_1t2a8E_1lizzieLet32_4MQNode_7QNode_Bool_1t3a8F_1Lcall_f'''''''''_f'''''''''_Bool3_d  = \Lcall_f'''''''''_f'''''''''_Bool3_dc ((& {lizzieLet32_4MQNode_4QNode_Bool_d[0],
                                                                                                                                                                                                                                                     lizzieLet32_4MQNode_5QNode_Bool_d[0],
                                                                                                                                                                                                                                                     t1a8D_destruct_d[0],
                                                                                                                                                                                                                                                     lizzieLet32_4MQNode_6QNode_Bool_d[0],
                                                                                                                                                                                                                                                     t2a8E_destruct_d[0],
                                                                                                                                                                                                                                                     lizzieLet32_4MQNode_7QNode_Bool_d[0],
                                                                                                                                                                                                                                                     t3a8F_destruct_d[0]}), lizzieLet32_4MQNode_4QNode_Bool_d, lizzieLet32_4MQNode_5QNode_Bool_d, t1a8D_destruct_d, lizzieLet32_4MQNode_6QNode_Bool_d, t2a8E_destruct_d, lizzieLet32_4MQNode_7QNode_Bool_d, t3a8F_destruct_d);
  assign {lizzieLet32_4MQNode_4QNode_Bool_r,
          lizzieLet32_4MQNode_5QNode_Bool_r,
          t1a8D_destruct_r,
          lizzieLet32_4MQNode_6QNode_Bool_r,
          t2a8E_destruct_r,
          lizzieLet32_4MQNode_7QNode_Bool_r,
          t3a8F_destruct_r} = {7 {(\lizzieLet32_4MQNode_4QNode_Bool_1lizzieLet32_4MQNode_5QNode_Bool_1t1a8D_1lizzieLet32_4MQNode_6QNode_Bool_1t2a8E_1lizzieLet32_4MQNode_7QNode_Bool_1t3a8F_1Lcall_f'''''''''_f'''''''''_Bool3_r  && \lizzieLet32_4MQNode_4QNode_Bool_1lizzieLet32_4MQNode_5QNode_Bool_1t1a8D_1lizzieLet32_4MQNode_6QNode_Bool_1t2a8E_1lizzieLet32_4MQNode_7QNode_Bool_1t3a8F_1Lcall_f'''''''''_f'''''''''_Bool3_d [0])}};
  
  /* buf (Ty CTf'''''''''_f'''''''''_Bool) : (lizzieLet32_4MQNode_4QNode_Bool_1lizzieLet32_4MQNode_5QNode_Bool_1t1a8D_1lizzieLet32_4MQNode_6QNode_Bool_1t2a8E_1lizzieLet32_4MQNode_7QNode_Bool_1t3a8F_1Lcall_f'''''''''_f'''''''''_Bool3,CTf'''''''''_f'''''''''_Bool) > (lizzieLet37_1_argbuf,CTf'''''''''_f'''''''''_Bool) */
  \CTf'''''''''_f'''''''''_Bool_t  \lizzieLet32_4MQNode_4QNode_Bool_1lizzieLet32_4MQNode_5QNode_Bool_1t1a8D_1lizzieLet32_4MQNode_6QNode_Bool_1t2a8E_1lizzieLet32_4MQNode_7QNode_Bool_1t3a8F_1Lcall_f'''''''''_f'''''''''_Bool3_bufchan_d ;
  logic \lizzieLet32_4MQNode_4QNode_Bool_1lizzieLet32_4MQNode_5QNode_Bool_1t1a8D_1lizzieLet32_4MQNode_6QNode_Bool_1t2a8E_1lizzieLet32_4MQNode_7QNode_Bool_1t3a8F_1Lcall_f'''''''''_f'''''''''_Bool3_bufchan_r ;
  assign \lizzieLet32_4MQNode_4QNode_Bool_1lizzieLet32_4MQNode_5QNode_Bool_1t1a8D_1lizzieLet32_4MQNode_6QNode_Bool_1t2a8E_1lizzieLet32_4MQNode_7QNode_Bool_1t3a8F_1Lcall_f'''''''''_f'''''''''_Bool3_r  = ((! \lizzieLet32_4MQNode_4QNode_Bool_1lizzieLet32_4MQNode_5QNode_Bool_1t1a8D_1lizzieLet32_4MQNode_6QNode_Bool_1t2a8E_1lizzieLet32_4MQNode_7QNode_Bool_1t3a8F_1Lcall_f'''''''''_f'''''''''_Bool3_bufchan_d [0]) || \lizzieLet32_4MQNode_4QNode_Bool_1lizzieLet32_4MQNode_5QNode_Bool_1t1a8D_1lizzieLet32_4MQNode_6QNode_Bool_1t2a8E_1lizzieLet32_4MQNode_7QNode_Bool_1t3a8F_1Lcall_f'''''''''_f'''''''''_Bool3_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet32_4MQNode_4QNode_Bool_1lizzieLet32_4MQNode_5QNode_Bool_1t1a8D_1lizzieLet32_4MQNode_6QNode_Bool_1t2a8E_1lizzieLet32_4MQNode_7QNode_Bool_1t3a8F_1Lcall_f'''''''''_f'''''''''_Bool3_bufchan_d  <= {115'd0,
                                                                                                                                                                                                                 1'd0};
    else
      if (\lizzieLet32_4MQNode_4QNode_Bool_1lizzieLet32_4MQNode_5QNode_Bool_1t1a8D_1lizzieLet32_4MQNode_6QNode_Bool_1t2a8E_1lizzieLet32_4MQNode_7QNode_Bool_1t3a8F_1Lcall_f'''''''''_f'''''''''_Bool3_r )
        \lizzieLet32_4MQNode_4QNode_Bool_1lizzieLet32_4MQNode_5QNode_Bool_1t1a8D_1lizzieLet32_4MQNode_6QNode_Bool_1t2a8E_1lizzieLet32_4MQNode_7QNode_Bool_1t3a8F_1Lcall_f'''''''''_f'''''''''_Bool3_bufchan_d  <= \lizzieLet32_4MQNode_4QNode_Bool_1lizzieLet32_4MQNode_5QNode_Bool_1t1a8D_1lizzieLet32_4MQNode_6QNode_Bool_1t2a8E_1lizzieLet32_4MQNode_7QNode_Bool_1t3a8F_1Lcall_f'''''''''_f'''''''''_Bool3_d ;
  \CTf'''''''''_f'''''''''_Bool_t  \lizzieLet32_4MQNode_4QNode_Bool_1lizzieLet32_4MQNode_5QNode_Bool_1t1a8D_1lizzieLet32_4MQNode_6QNode_Bool_1t2a8E_1lizzieLet32_4MQNode_7QNode_Bool_1t3a8F_1Lcall_f'''''''''_f'''''''''_Bool3_bufchan_buf ;
  assign \lizzieLet32_4MQNode_4QNode_Bool_1lizzieLet32_4MQNode_5QNode_Bool_1t1a8D_1lizzieLet32_4MQNode_6QNode_Bool_1t2a8E_1lizzieLet32_4MQNode_7QNode_Bool_1t3a8F_1Lcall_f'''''''''_f'''''''''_Bool3_bufchan_r  = (! \lizzieLet32_4MQNode_4QNode_Bool_1lizzieLet32_4MQNode_5QNode_Bool_1t1a8D_1lizzieLet32_4MQNode_6QNode_Bool_1t2a8E_1lizzieLet32_4MQNode_7QNode_Bool_1t3a8F_1Lcall_f'''''''''_f'''''''''_Bool3_bufchan_buf [0]);
  assign lizzieLet37_1_argbuf_d = (\lizzieLet32_4MQNode_4QNode_Bool_1lizzieLet32_4MQNode_5QNode_Bool_1t1a8D_1lizzieLet32_4MQNode_6QNode_Bool_1t2a8E_1lizzieLet32_4MQNode_7QNode_Bool_1t3a8F_1Lcall_f'''''''''_f'''''''''_Bool3_bufchan_buf [0] ? \lizzieLet32_4MQNode_4QNode_Bool_1lizzieLet32_4MQNode_5QNode_Bool_1t1a8D_1lizzieLet32_4MQNode_6QNode_Bool_1t2a8E_1lizzieLet32_4MQNode_7QNode_Bool_1t3a8F_1Lcall_f'''''''''_f'''''''''_Bool3_bufchan_buf  :
                                   \lizzieLet32_4MQNode_4QNode_Bool_1lizzieLet32_4MQNode_5QNode_Bool_1t1a8D_1lizzieLet32_4MQNode_6QNode_Bool_1t2a8E_1lizzieLet32_4MQNode_7QNode_Bool_1t3a8F_1Lcall_f'''''''''_f'''''''''_Bool3_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet32_4MQNode_4QNode_Bool_1lizzieLet32_4MQNode_5QNode_Bool_1t1a8D_1lizzieLet32_4MQNode_6QNode_Bool_1t2a8E_1lizzieLet32_4MQNode_7QNode_Bool_1t3a8F_1Lcall_f'''''''''_f'''''''''_Bool3_bufchan_buf  <= {115'd0,
                                                                                                                                                                                                                   1'd0};
    else
      if ((lizzieLet37_1_argbuf_r && \lizzieLet32_4MQNode_4QNode_Bool_1lizzieLet32_4MQNode_5QNode_Bool_1t1a8D_1lizzieLet32_4MQNode_6QNode_Bool_1t2a8E_1lizzieLet32_4MQNode_7QNode_Bool_1t3a8F_1Lcall_f'''''''''_f'''''''''_Bool3_bufchan_buf [0]))
        \lizzieLet32_4MQNode_4QNode_Bool_1lizzieLet32_4MQNode_5QNode_Bool_1t1a8D_1lizzieLet32_4MQNode_6QNode_Bool_1t2a8E_1lizzieLet32_4MQNode_7QNode_Bool_1t3a8F_1Lcall_f'''''''''_f'''''''''_Bool3_bufchan_buf  <= {115'd0,
                                                                                                                                                                                                                     1'd0};
      else if (((! lizzieLet37_1_argbuf_r) && (! \lizzieLet32_4MQNode_4QNode_Bool_1lizzieLet32_4MQNode_5QNode_Bool_1t1a8D_1lizzieLet32_4MQNode_6QNode_Bool_1t2a8E_1lizzieLet32_4MQNode_7QNode_Bool_1t3a8F_1Lcall_f'''''''''_f'''''''''_Bool3_bufchan_buf [0])))
        \lizzieLet32_4MQNode_4QNode_Bool_1lizzieLet32_4MQNode_5QNode_Bool_1t1a8D_1lizzieLet32_4MQNode_6QNode_Bool_1t2a8E_1lizzieLet32_4MQNode_7QNode_Bool_1t3a8F_1Lcall_f'''''''''_f'''''''''_Bool3_bufchan_buf  <= \lizzieLet32_4MQNode_4QNode_Bool_1lizzieLet32_4MQNode_5QNode_Bool_1t1a8D_1lizzieLet32_4MQNode_6QNode_Bool_1t2a8E_1lizzieLet32_4MQNode_7QNode_Bool_1t3a8F_1Lcall_f'''''''''_f'''''''''_Bool3_bufchan_d ;
  
  /* buf (Ty Pointer_CTf'''''''''_f'''''''''_Bool) : (lizzieLet32_4MQNode_4QNone_Bool,Pointer_CTf'''''''''_f'''''''''_Bool) > (lizzieLet32_4MQNode_4QNone_Bool_1_argbuf,Pointer_CTf'''''''''_f'''''''''_Bool) */
  \Pointer_CTf'''''''''_f'''''''''_Bool_t  lizzieLet32_4MQNode_4QNone_Bool_bufchan_d;
  logic lizzieLet32_4MQNode_4QNone_Bool_bufchan_r;
  assign lizzieLet32_4MQNode_4QNone_Bool_r = ((! lizzieLet32_4MQNode_4QNone_Bool_bufchan_d[0]) || lizzieLet32_4MQNode_4QNone_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet32_4MQNode_4QNone_Bool_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet32_4MQNode_4QNone_Bool_r)
        lizzieLet32_4MQNode_4QNone_Bool_bufchan_d <= lizzieLet32_4MQNode_4QNone_Bool_d;
  \Pointer_CTf'''''''''_f'''''''''_Bool_t  lizzieLet32_4MQNode_4QNone_Bool_bufchan_buf;
  assign lizzieLet32_4MQNode_4QNone_Bool_bufchan_r = (! lizzieLet32_4MQNode_4QNone_Bool_bufchan_buf[0]);
  assign lizzieLet32_4MQNode_4QNone_Bool_1_argbuf_d = (lizzieLet32_4MQNode_4QNone_Bool_bufchan_buf[0] ? lizzieLet32_4MQNode_4QNone_Bool_bufchan_buf :
                                                       lizzieLet32_4MQNode_4QNone_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet32_4MQNode_4QNone_Bool_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet32_4MQNode_4QNone_Bool_1_argbuf_r && lizzieLet32_4MQNode_4QNone_Bool_bufchan_buf[0]))
        lizzieLet32_4MQNode_4QNone_Bool_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet32_4MQNode_4QNone_Bool_1_argbuf_r) && (! lizzieLet32_4MQNode_4QNone_Bool_bufchan_buf[0])))
        lizzieLet32_4MQNode_4QNone_Bool_bufchan_buf <= lizzieLet32_4MQNode_4QNone_Bool_bufchan_d;
  
  /* buf (Ty Pointer_CTf'''''''''_f'''''''''_Bool) : (lizzieLet32_4MQNode_4QVal_Bool,Pointer_CTf'''''''''_f'''''''''_Bool) > (lizzieLet32_4MQNode_4QVal_Bool_1_argbuf,Pointer_CTf'''''''''_f'''''''''_Bool) */
  \Pointer_CTf'''''''''_f'''''''''_Bool_t  lizzieLet32_4MQNode_4QVal_Bool_bufchan_d;
  logic lizzieLet32_4MQNode_4QVal_Bool_bufchan_r;
  assign lizzieLet32_4MQNode_4QVal_Bool_r = ((! lizzieLet32_4MQNode_4QVal_Bool_bufchan_d[0]) || lizzieLet32_4MQNode_4QVal_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet32_4MQNode_4QVal_Bool_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet32_4MQNode_4QVal_Bool_r)
        lizzieLet32_4MQNode_4QVal_Bool_bufchan_d <= lizzieLet32_4MQNode_4QVal_Bool_d;
  \Pointer_CTf'''''''''_f'''''''''_Bool_t  lizzieLet32_4MQNode_4QVal_Bool_bufchan_buf;
  assign lizzieLet32_4MQNode_4QVal_Bool_bufchan_r = (! lizzieLet32_4MQNode_4QVal_Bool_bufchan_buf[0]);
  assign lizzieLet32_4MQNode_4QVal_Bool_1_argbuf_d = (lizzieLet32_4MQNode_4QVal_Bool_bufchan_buf[0] ? lizzieLet32_4MQNode_4QVal_Bool_bufchan_buf :
                                                      lizzieLet32_4MQNode_4QVal_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet32_4MQNode_4QVal_Bool_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet32_4MQNode_4QVal_Bool_1_argbuf_r && lizzieLet32_4MQNode_4QVal_Bool_bufchan_buf[0]))
        lizzieLet32_4MQNode_4QVal_Bool_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet32_4MQNode_4QVal_Bool_1_argbuf_r) && (! lizzieLet32_4MQNode_4QVal_Bool_bufchan_buf[0])))
        lizzieLet32_4MQNode_4QVal_Bool_bufchan_buf <= lizzieLet32_4MQNode_4QVal_Bool_bufchan_d;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_MaskQTree) : (lizzieLet32_4MQNode_5,QTree_Bool) (q1a8y_destruct,Pointer_MaskQTree) > [(_19,Pointer_MaskQTree),
                                                                                                        (_18,Pointer_MaskQTree),
                                                                                                        (lizzieLet32_4MQNode_5QNode_Bool,Pointer_MaskQTree),
                                                                                                        (_17,Pointer_MaskQTree)] */
  logic [3:0] q1a8y_destruct_onehotd;
  always_comb
    if ((lizzieLet32_4MQNode_5_d[0] && q1a8y_destruct_d[0]))
      unique case (lizzieLet32_4MQNode_5_d[2:1])
        2'd0: q1a8y_destruct_onehotd = 4'd1;
        2'd1: q1a8y_destruct_onehotd = 4'd2;
        2'd2: q1a8y_destruct_onehotd = 4'd4;
        2'd3: q1a8y_destruct_onehotd = 4'd8;
        default: q1a8y_destruct_onehotd = 4'd0;
      endcase
    else q1a8y_destruct_onehotd = 4'd0;
  assign _19_d = {q1a8y_destruct_d[16:1], q1a8y_destruct_onehotd[0]};
  assign _18_d = {q1a8y_destruct_d[16:1], q1a8y_destruct_onehotd[1]};
  assign lizzieLet32_4MQNode_5QNode_Bool_d = {q1a8y_destruct_d[16:1],
                                              q1a8y_destruct_onehotd[2]};
  assign _17_d = {q1a8y_destruct_d[16:1], q1a8y_destruct_onehotd[3]};
  assign q1a8y_destruct_r = (| (q1a8y_destruct_onehotd & {_17_r,
                                                          lizzieLet32_4MQNode_5QNode_Bool_r,
                                                          _18_r,
                                                          _19_r}));
  assign lizzieLet32_4MQNode_5_r = q1a8y_destruct_r;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_MaskQTree) : (lizzieLet32_4MQNode_6,QTree_Bool) (q2a8z_destruct,Pointer_MaskQTree) > [(_16,Pointer_MaskQTree),
                                                                                                        (_15,Pointer_MaskQTree),
                                                                                                        (lizzieLet32_4MQNode_6QNode_Bool,Pointer_MaskQTree),
                                                                                                        (_14,Pointer_MaskQTree)] */
  logic [3:0] q2a8z_destruct_onehotd;
  always_comb
    if ((lizzieLet32_4MQNode_6_d[0] && q2a8z_destruct_d[0]))
      unique case (lizzieLet32_4MQNode_6_d[2:1])
        2'd0: q2a8z_destruct_onehotd = 4'd1;
        2'd1: q2a8z_destruct_onehotd = 4'd2;
        2'd2: q2a8z_destruct_onehotd = 4'd4;
        2'd3: q2a8z_destruct_onehotd = 4'd8;
        default: q2a8z_destruct_onehotd = 4'd0;
      endcase
    else q2a8z_destruct_onehotd = 4'd0;
  assign _16_d = {q2a8z_destruct_d[16:1], q2a8z_destruct_onehotd[0]};
  assign _15_d = {q2a8z_destruct_d[16:1], q2a8z_destruct_onehotd[1]};
  assign lizzieLet32_4MQNode_6QNode_Bool_d = {q2a8z_destruct_d[16:1],
                                              q2a8z_destruct_onehotd[2]};
  assign _14_d = {q2a8z_destruct_d[16:1], q2a8z_destruct_onehotd[3]};
  assign q2a8z_destruct_r = (| (q2a8z_destruct_onehotd & {_14_r,
                                                          lizzieLet32_4MQNode_6QNode_Bool_r,
                                                          _15_r,
                                                          _16_r}));
  assign lizzieLet32_4MQNode_6_r = q2a8z_destruct_r;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_MaskQTree) : (lizzieLet32_4MQNode_7,QTree_Bool) (q3a8A_destruct,Pointer_MaskQTree) > [(_13,Pointer_MaskQTree),
                                                                                                        (_12,Pointer_MaskQTree),
                                                                                                        (lizzieLet32_4MQNode_7QNode_Bool,Pointer_MaskQTree),
                                                                                                        (_11,Pointer_MaskQTree)] */
  logic [3:0] q3a8A_destruct_onehotd;
  always_comb
    if ((lizzieLet32_4MQNode_7_d[0] && q3a8A_destruct_d[0]))
      unique case (lizzieLet32_4MQNode_7_d[2:1])
        2'd0: q3a8A_destruct_onehotd = 4'd1;
        2'd1: q3a8A_destruct_onehotd = 4'd2;
        2'd2: q3a8A_destruct_onehotd = 4'd4;
        2'd3: q3a8A_destruct_onehotd = 4'd8;
        default: q3a8A_destruct_onehotd = 4'd0;
      endcase
    else q3a8A_destruct_onehotd = 4'd0;
  assign _13_d = {q3a8A_destruct_d[16:1], q3a8A_destruct_onehotd[0]};
  assign _12_d = {q3a8A_destruct_d[16:1], q3a8A_destruct_onehotd[1]};
  assign lizzieLet32_4MQNode_7QNode_Bool_d = {q3a8A_destruct_d[16:1],
                                              q3a8A_destruct_onehotd[2]};
  assign _11_d = {q3a8A_destruct_d[16:1], q3a8A_destruct_onehotd[3]};
  assign q3a8A_destruct_r = (| (q3a8A_destruct_onehotd & {_11_r,
                                                          lizzieLet32_4MQNode_7QNode_Bool_r,
                                                          _12_r,
                                                          _13_r}));
  assign lizzieLet32_4MQNode_7_r = q3a8A_destruct_r;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_MaskQTree) : (lizzieLet32_4MQNode_8,QTree_Bool) (q5a8B_destruct,Pointer_MaskQTree) > [(_10,Pointer_MaskQTree),
                                                                                                        (_9,Pointer_MaskQTree),
                                                                                                        (lizzieLet32_4MQNode_8QNode_Bool,Pointer_MaskQTree),
                                                                                                        (_8,Pointer_MaskQTree)] */
  logic [3:0] q5a8B_destruct_onehotd;
  always_comb
    if ((lizzieLet32_4MQNode_8_d[0] && q5a8B_destruct_d[0]))
      unique case (lizzieLet32_4MQNode_8_d[2:1])
        2'd0: q5a8B_destruct_onehotd = 4'd1;
        2'd1: q5a8B_destruct_onehotd = 4'd2;
        2'd2: q5a8B_destruct_onehotd = 4'd4;
        2'd3: q5a8B_destruct_onehotd = 4'd8;
        default: q5a8B_destruct_onehotd = 4'd0;
      endcase
    else q5a8B_destruct_onehotd = 4'd0;
  assign _10_d = {q5a8B_destruct_d[16:1], q5a8B_destruct_onehotd[0]};
  assign _9_d = {q5a8B_destruct_d[16:1], q5a8B_destruct_onehotd[1]};
  assign lizzieLet32_4MQNode_8QNode_Bool_d = {q5a8B_destruct_d[16:1],
                                              q5a8B_destruct_onehotd[2]};
  assign _8_d = {q5a8B_destruct_d[16:1], q5a8B_destruct_onehotd[3]};
  assign q5a8B_destruct_r = (| (q5a8B_destruct_onehotd & {_8_r,
                                                          lizzieLet32_4MQNode_8QNode_Bool_r,
                                                          _9_r,
                                                          _10_r}));
  assign lizzieLet32_4MQNode_8_r = q5a8B_destruct_r;
  
  /* buf (Ty Pointer_MaskQTree) : (lizzieLet32_4MQNode_8QNode_Bool,Pointer_MaskQTree) > (lizzieLet32_4MQNode_8QNode_Bool_1_argbuf,Pointer_MaskQTree) */
  Pointer_MaskQTree_t lizzieLet32_4MQNode_8QNode_Bool_bufchan_d;
  logic lizzieLet32_4MQNode_8QNode_Bool_bufchan_r;
  assign lizzieLet32_4MQNode_8QNode_Bool_r = ((! lizzieLet32_4MQNode_8QNode_Bool_bufchan_d[0]) || lizzieLet32_4MQNode_8QNode_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet32_4MQNode_8QNode_Bool_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet32_4MQNode_8QNode_Bool_r)
        lizzieLet32_4MQNode_8QNode_Bool_bufchan_d <= lizzieLet32_4MQNode_8QNode_Bool_d;
  Pointer_MaskQTree_t lizzieLet32_4MQNode_8QNode_Bool_bufchan_buf;
  assign lizzieLet32_4MQNode_8QNode_Bool_bufchan_r = (! lizzieLet32_4MQNode_8QNode_Bool_bufchan_buf[0]);
  assign lizzieLet32_4MQNode_8QNode_Bool_1_argbuf_d = (lizzieLet32_4MQNode_8QNode_Bool_bufchan_buf[0] ? lizzieLet32_4MQNode_8QNode_Bool_bufchan_buf :
                                                       lizzieLet32_4MQNode_8QNode_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet32_4MQNode_8QNode_Bool_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet32_4MQNode_8QNode_Bool_1_argbuf_r && lizzieLet32_4MQNode_8QNode_Bool_bufchan_buf[0]))
        lizzieLet32_4MQNode_8QNode_Bool_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet32_4MQNode_8QNode_Bool_1_argbuf_r) && (! lizzieLet32_4MQNode_8QNode_Bool_bufchan_buf[0])))
        lizzieLet32_4MQNode_8QNode_Bool_bufchan_buf <= lizzieLet32_4MQNode_8QNode_Bool_bufchan_d;
  
  /* demux (Ty MaskQTree,
       Ty Pointer_QTree_Bool) : (lizzieLet32_5,MaskQTree) (q4'a8x_2,Pointer_QTree_Bool) > [(_7,Pointer_QTree_Bool),
                                                                                           (lizzieLet32_5MQVal,Pointer_QTree_Bool),
                                                                                           (_6,Pointer_QTree_Bool)] */
  logic [2:0] \q4'a8x_2_onehotd ;
  always_comb
    if ((lizzieLet32_5_d[0] && \q4'a8x_2_d [0]))
      unique case (lizzieLet32_5_d[2:1])
        2'd0: \q4'a8x_2_onehotd  = 3'd1;
        2'd1: \q4'a8x_2_onehotd  = 3'd2;
        2'd2: \q4'a8x_2_onehotd  = 3'd4;
        default: \q4'a8x_2_onehotd  = 3'd0;
      endcase
    else \q4'a8x_2_onehotd  = 3'd0;
  assign _7_d = {\q4'a8x_2_d [16:1], \q4'a8x_2_onehotd [0]};
  assign lizzieLet32_5MQVal_d = {\q4'a8x_2_d [16:1],
                                 \q4'a8x_2_onehotd [1]};
  assign _6_d = {\q4'a8x_2_d [16:1], \q4'a8x_2_onehotd [2]};
  assign \q4'a8x_2_r  = (| (\q4'a8x_2_onehotd  & {_6_r,
                                                  lizzieLet32_5MQVal_r,
                                                  _7_r}));
  assign lizzieLet32_5_r = \q4'a8x_2_r ;
  
  /* buf (Ty Pointer_QTree_Bool) : (lizzieLet32_5MQVal,Pointer_QTree_Bool) > (lizzieLet32_5MQVal_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t lizzieLet32_5MQVal_bufchan_d;
  logic lizzieLet32_5MQVal_bufchan_r;
  assign lizzieLet32_5MQVal_r = ((! lizzieLet32_5MQVal_bufchan_d[0]) || lizzieLet32_5MQVal_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet32_5MQVal_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet32_5MQVal_r)
        lizzieLet32_5MQVal_bufchan_d <= lizzieLet32_5MQVal_d;
  Pointer_QTree_Bool_t lizzieLet32_5MQVal_bufchan_buf;
  assign lizzieLet32_5MQVal_bufchan_r = (! lizzieLet32_5MQVal_bufchan_buf[0]);
  assign lizzieLet32_5MQVal_1_argbuf_d = (lizzieLet32_5MQVal_bufchan_buf[0] ? lizzieLet32_5MQVal_bufchan_buf :
                                          lizzieLet32_5MQVal_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet32_5MQVal_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet32_5MQVal_1_argbuf_r && lizzieLet32_5MQVal_bufchan_buf[0]))
        lizzieLet32_5MQVal_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet32_5MQVal_1_argbuf_r) && (! lizzieLet32_5MQVal_bufchan_buf[0])))
        lizzieLet32_5MQVal_bufchan_buf <= lizzieLet32_5MQVal_bufchan_d;
  
  /* demux (Ty MaskQTree,
       Ty Pointer_CTf'''''''''_f'''''''''_Bool) : (lizzieLet32_6,MaskQTree) (sc_0_2_goMux_mux,Pointer_CTf'''''''''_f'''''''''_Bool) > [(lizzieLet32_6MQNone,Pointer_CTf'''''''''_f'''''''''_Bool),
                                                                                                                                       (lizzieLet32_6MQVal,Pointer_CTf'''''''''_f'''''''''_Bool),
                                                                                                                                       (lizzieLet32_6MQNode,Pointer_CTf'''''''''_f'''''''''_Bool)] */
  logic [2:0] sc_0_2_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet32_6_d[0] && sc_0_2_goMux_mux_d[0]))
      unique case (lizzieLet32_6_d[2:1])
        2'd0: sc_0_2_goMux_mux_onehotd = 3'd1;
        2'd1: sc_0_2_goMux_mux_onehotd = 3'd2;
        2'd2: sc_0_2_goMux_mux_onehotd = 3'd4;
        default: sc_0_2_goMux_mux_onehotd = 3'd0;
      endcase
    else sc_0_2_goMux_mux_onehotd = 3'd0;
  assign lizzieLet32_6MQNone_d = {sc_0_2_goMux_mux_d[16:1],
                                  sc_0_2_goMux_mux_onehotd[0]};
  assign lizzieLet32_6MQVal_d = {sc_0_2_goMux_mux_d[16:1],
                                 sc_0_2_goMux_mux_onehotd[1]};
  assign lizzieLet32_6MQNode_d = {sc_0_2_goMux_mux_d[16:1],
                                  sc_0_2_goMux_mux_onehotd[2]};
  assign sc_0_2_goMux_mux_r = (| (sc_0_2_goMux_mux_onehotd & {lizzieLet32_6MQNode_r,
                                                              lizzieLet32_6MQVal_r,
                                                              lizzieLet32_6MQNone_r}));
  assign lizzieLet32_6_r = sc_0_2_goMux_mux_r;
  
  /* buf (Ty Pointer_CTf'''''''''_f'''''''''_Bool) : (lizzieLet32_6MQNone,Pointer_CTf'''''''''_f'''''''''_Bool) > (lizzieLet32_6MQNone_1_argbuf,Pointer_CTf'''''''''_f'''''''''_Bool) */
  \Pointer_CTf'''''''''_f'''''''''_Bool_t  lizzieLet32_6MQNone_bufchan_d;
  logic lizzieLet32_6MQNone_bufchan_r;
  assign lizzieLet32_6MQNone_r = ((! lizzieLet32_6MQNone_bufchan_d[0]) || lizzieLet32_6MQNone_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet32_6MQNone_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet32_6MQNone_r)
        lizzieLet32_6MQNone_bufchan_d <= lizzieLet32_6MQNone_d;
  \Pointer_CTf'''''''''_f'''''''''_Bool_t  lizzieLet32_6MQNone_bufchan_buf;
  assign lizzieLet32_6MQNone_bufchan_r = (! lizzieLet32_6MQNone_bufchan_buf[0]);
  assign lizzieLet32_6MQNone_1_argbuf_d = (lizzieLet32_6MQNone_bufchan_buf[0] ? lizzieLet32_6MQNone_bufchan_buf :
                                           lizzieLet32_6MQNone_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet32_6MQNone_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet32_6MQNone_1_argbuf_r && lizzieLet32_6MQNone_bufchan_buf[0]))
        lizzieLet32_6MQNone_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet32_6MQNone_1_argbuf_r) && (! lizzieLet32_6MQNone_bufchan_buf[0])))
        lizzieLet32_6MQNone_bufchan_buf <= lizzieLet32_6MQNone_bufchan_d;
  
  /* buf (Ty Pointer_CTf'''''''''_f'''''''''_Bool) : (lizzieLet32_6MQVal,Pointer_CTf'''''''''_f'''''''''_Bool) > (lizzieLet32_6MQVal_1_argbuf,Pointer_CTf'''''''''_f'''''''''_Bool) */
  \Pointer_CTf'''''''''_f'''''''''_Bool_t  lizzieLet32_6MQVal_bufchan_d;
  logic lizzieLet32_6MQVal_bufchan_r;
  assign lizzieLet32_6MQVal_r = ((! lizzieLet32_6MQVal_bufchan_d[0]) || lizzieLet32_6MQVal_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet32_6MQVal_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet32_6MQVal_r)
        lizzieLet32_6MQVal_bufchan_d <= lizzieLet32_6MQVal_d;
  \Pointer_CTf'''''''''_f'''''''''_Bool_t  lizzieLet32_6MQVal_bufchan_buf;
  assign lizzieLet32_6MQVal_bufchan_r = (! lizzieLet32_6MQVal_bufchan_buf[0]);
  assign lizzieLet32_6MQVal_1_argbuf_d = (lizzieLet32_6MQVal_bufchan_buf[0] ? lizzieLet32_6MQVal_bufchan_buf :
                                          lizzieLet32_6MQVal_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet32_6MQVal_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet32_6MQVal_1_argbuf_r && lizzieLet32_6MQVal_bufchan_buf[0]))
        lizzieLet32_6MQVal_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet32_6MQVal_1_argbuf_r) && (! lizzieLet32_6MQVal_bufchan_buf[0])))
        lizzieLet32_6MQVal_bufchan_buf <= lizzieLet32_6MQVal_bufchan_d;
  
  /* destruct (Ty CTf,
          Dcon Lcall_f0) : (lizzieLet43_1Lcall_f0,CTf) > [(es_9_destruct,Pointer_QTree_Bool),
                                                          (es_10_1_destruct,Pointer_QTree_Bool),
                                                          (es_11_2_destruct,Pointer_QTree_Bool),
                                                          (sc_0_6_destruct,Pointer_CTf)] */
  logic [3:0] lizzieLet43_1Lcall_f0_emitted;
  logic [3:0] lizzieLet43_1Lcall_f0_done;
  assign es_9_destruct_d = {lizzieLet43_1Lcall_f0_d[19:4],
                            (lizzieLet43_1Lcall_f0_d[0] && (! lizzieLet43_1Lcall_f0_emitted[0]))};
  assign es_10_1_destruct_d = {lizzieLet43_1Lcall_f0_d[35:20],
                               (lizzieLet43_1Lcall_f0_d[0] && (! lizzieLet43_1Lcall_f0_emitted[1]))};
  assign es_11_2_destruct_d = {lizzieLet43_1Lcall_f0_d[51:36],
                               (lizzieLet43_1Lcall_f0_d[0] && (! lizzieLet43_1Lcall_f0_emitted[2]))};
  assign sc_0_6_destruct_d = {lizzieLet43_1Lcall_f0_d[67:52],
                              (lizzieLet43_1Lcall_f0_d[0] && (! lizzieLet43_1Lcall_f0_emitted[3]))};
  assign lizzieLet43_1Lcall_f0_done = (lizzieLet43_1Lcall_f0_emitted | ({sc_0_6_destruct_d[0],
                                                                         es_11_2_destruct_d[0],
                                                                         es_10_1_destruct_d[0],
                                                                         es_9_destruct_d[0]} & {sc_0_6_destruct_r,
                                                                                                es_11_2_destruct_r,
                                                                                                es_10_1_destruct_r,
                                                                                                es_9_destruct_r}));
  assign lizzieLet43_1Lcall_f0_r = (& lizzieLet43_1Lcall_f0_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet43_1Lcall_f0_emitted <= 4'd0;
    else
      lizzieLet43_1Lcall_f0_emitted <= (lizzieLet43_1Lcall_f0_r ? 4'd0 :
                                        lizzieLet43_1Lcall_f0_done);
  
  /* destruct (Ty CTf,
          Dcon Lcall_f1) : (lizzieLet43_1Lcall_f1,CTf) > [(es_10_destruct,Pointer_QTree_Bool),
                                                          (es_11_1_destruct,Pointer_QTree_Bool),
                                                          (sc_0_5_destruct,Pointer_CTf),
                                                          (q1a88_3_destruct,Pointer_MaskQTree),
                                                          (q1'a8n_3_destruct,Pointer_QTree_Bool),
                                                          (t1a8s_3_destruct,Pointer_QTree_Bool)] */
  logic [5:0] lizzieLet43_1Lcall_f1_emitted;
  logic [5:0] lizzieLet43_1Lcall_f1_done;
  assign es_10_destruct_d = {lizzieLet43_1Lcall_f1_d[19:4],
                             (lizzieLet43_1Lcall_f1_d[0] && (! lizzieLet43_1Lcall_f1_emitted[0]))};
  assign es_11_1_destruct_d = {lizzieLet43_1Lcall_f1_d[35:20],
                               (lizzieLet43_1Lcall_f1_d[0] && (! lizzieLet43_1Lcall_f1_emitted[1]))};
  assign sc_0_5_destruct_d = {lizzieLet43_1Lcall_f1_d[51:36],
                              (lizzieLet43_1Lcall_f1_d[0] && (! lizzieLet43_1Lcall_f1_emitted[2]))};
  assign q1a88_3_destruct_d = {lizzieLet43_1Lcall_f1_d[67:52],
                               (lizzieLet43_1Lcall_f1_d[0] && (! lizzieLet43_1Lcall_f1_emitted[3]))};
  assign \q1'a8n_3_destruct_d  = {lizzieLet43_1Lcall_f1_d[83:68],
                                  (lizzieLet43_1Lcall_f1_d[0] && (! lizzieLet43_1Lcall_f1_emitted[4]))};
  assign t1a8s_3_destruct_d = {lizzieLet43_1Lcall_f1_d[99:84],
                               (lizzieLet43_1Lcall_f1_d[0] && (! lizzieLet43_1Lcall_f1_emitted[5]))};
  assign lizzieLet43_1Lcall_f1_done = (lizzieLet43_1Lcall_f1_emitted | ({t1a8s_3_destruct_d[0],
                                                                         \q1'a8n_3_destruct_d [0],
                                                                         q1a88_3_destruct_d[0],
                                                                         sc_0_5_destruct_d[0],
                                                                         es_11_1_destruct_d[0],
                                                                         es_10_destruct_d[0]} & {t1a8s_3_destruct_r,
                                                                                                 \q1'a8n_3_destruct_r ,
                                                                                                 q1a88_3_destruct_r,
                                                                                                 sc_0_5_destruct_r,
                                                                                                 es_11_1_destruct_r,
                                                                                                 es_10_destruct_r}));
  assign lizzieLet43_1Lcall_f1_r = (& lizzieLet43_1Lcall_f1_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet43_1Lcall_f1_emitted <= 6'd0;
    else
      lizzieLet43_1Lcall_f1_emitted <= (lizzieLet43_1Lcall_f1_r ? 6'd0 :
                                        lizzieLet43_1Lcall_f1_done);
  
  /* destruct (Ty CTf,
          Dcon Lcall_f2) : (lizzieLet43_1Lcall_f2,CTf) > [(es_11_destruct,Pointer_QTree_Bool),
                                                          (sc_0_4_destruct,Pointer_CTf),
                                                          (q1a88_2_destruct,Pointer_MaskQTree),
                                                          (q1'a8n_2_destruct,Pointer_QTree_Bool),
                                                          (t1a8s_2_destruct,Pointer_QTree_Bool),
                                                          (q2a89_2_destruct,Pointer_MaskQTree),
                                                          (q2'a8o_2_destruct,Pointer_QTree_Bool),
                                                          (t2a8t_2_destruct,Pointer_QTree_Bool)] */
  logic [7:0] lizzieLet43_1Lcall_f2_emitted;
  logic [7:0] lizzieLet43_1Lcall_f2_done;
  assign es_11_destruct_d = {lizzieLet43_1Lcall_f2_d[19:4],
                             (lizzieLet43_1Lcall_f2_d[0] && (! lizzieLet43_1Lcall_f2_emitted[0]))};
  assign sc_0_4_destruct_d = {lizzieLet43_1Lcall_f2_d[35:20],
                              (lizzieLet43_1Lcall_f2_d[0] && (! lizzieLet43_1Lcall_f2_emitted[1]))};
  assign q1a88_2_destruct_d = {lizzieLet43_1Lcall_f2_d[51:36],
                               (lizzieLet43_1Lcall_f2_d[0] && (! lizzieLet43_1Lcall_f2_emitted[2]))};
  assign \q1'a8n_2_destruct_d  = {lizzieLet43_1Lcall_f2_d[67:52],
                                  (lizzieLet43_1Lcall_f2_d[0] && (! lizzieLet43_1Lcall_f2_emitted[3]))};
  assign t1a8s_2_destruct_d = {lizzieLet43_1Lcall_f2_d[83:68],
                               (lizzieLet43_1Lcall_f2_d[0] && (! lizzieLet43_1Lcall_f2_emitted[4]))};
  assign q2a89_2_destruct_d = {lizzieLet43_1Lcall_f2_d[99:84],
                               (lizzieLet43_1Lcall_f2_d[0] && (! lizzieLet43_1Lcall_f2_emitted[5]))};
  assign \q2'a8o_2_destruct_d  = {lizzieLet43_1Lcall_f2_d[115:100],
                                  (lizzieLet43_1Lcall_f2_d[0] && (! lizzieLet43_1Lcall_f2_emitted[6]))};
  assign t2a8t_2_destruct_d = {lizzieLet43_1Lcall_f2_d[131:116],
                               (lizzieLet43_1Lcall_f2_d[0] && (! lizzieLet43_1Lcall_f2_emitted[7]))};
  assign lizzieLet43_1Lcall_f2_done = (lizzieLet43_1Lcall_f2_emitted | ({t2a8t_2_destruct_d[0],
                                                                         \q2'a8o_2_destruct_d [0],
                                                                         q2a89_2_destruct_d[0],
                                                                         t1a8s_2_destruct_d[0],
                                                                         \q1'a8n_2_destruct_d [0],
                                                                         q1a88_2_destruct_d[0],
                                                                         sc_0_4_destruct_d[0],
                                                                         es_11_destruct_d[0]} & {t2a8t_2_destruct_r,
                                                                                                 \q2'a8o_2_destruct_r ,
                                                                                                 q2a89_2_destruct_r,
                                                                                                 t1a8s_2_destruct_r,
                                                                                                 \q1'a8n_2_destruct_r ,
                                                                                                 q1a88_2_destruct_r,
                                                                                                 sc_0_4_destruct_r,
                                                                                                 es_11_destruct_r}));
  assign lizzieLet43_1Lcall_f2_r = (& lizzieLet43_1Lcall_f2_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet43_1Lcall_f2_emitted <= 8'd0;
    else
      lizzieLet43_1Lcall_f2_emitted <= (lizzieLet43_1Lcall_f2_r ? 8'd0 :
                                        lizzieLet43_1Lcall_f2_done);
  
  /* destruct (Ty CTf,
          Dcon Lcall_f3) : (lizzieLet43_1Lcall_f3,CTf) > [(sc_0_3_destruct,Pointer_CTf),
                                                          (q1a88_1_destruct,Pointer_MaskQTree),
                                                          (q1'a8n_1_destruct,Pointer_QTree_Bool),
                                                          (t1a8s_1_destruct,Pointer_QTree_Bool),
                                                          (q2a89_1_destruct,Pointer_MaskQTree),
                                                          (q2'a8o_1_destruct,Pointer_QTree_Bool),
                                                          (t2a8t_1_destruct,Pointer_QTree_Bool),
                                                          (q3a8a_1_destruct,Pointer_MaskQTree),
                                                          (q3'a8p_1_destruct,Pointer_QTree_Bool),
                                                          (t3a8u_1_destruct,Pointer_QTree_Bool)] */
  logic [9:0] lizzieLet43_1Lcall_f3_emitted;
  logic [9:0] lizzieLet43_1Lcall_f3_done;
  assign sc_0_3_destruct_d = {lizzieLet43_1Lcall_f3_d[19:4],
                              (lizzieLet43_1Lcall_f3_d[0] && (! lizzieLet43_1Lcall_f3_emitted[0]))};
  assign q1a88_1_destruct_d = {lizzieLet43_1Lcall_f3_d[35:20],
                               (lizzieLet43_1Lcall_f3_d[0] && (! lizzieLet43_1Lcall_f3_emitted[1]))};
  assign \q1'a8n_1_destruct_d  = {lizzieLet43_1Lcall_f3_d[51:36],
                                  (lizzieLet43_1Lcall_f3_d[0] && (! lizzieLet43_1Lcall_f3_emitted[2]))};
  assign t1a8s_1_destruct_d = {lizzieLet43_1Lcall_f3_d[67:52],
                               (lizzieLet43_1Lcall_f3_d[0] && (! lizzieLet43_1Lcall_f3_emitted[3]))};
  assign q2a89_1_destruct_d = {lizzieLet43_1Lcall_f3_d[83:68],
                               (lizzieLet43_1Lcall_f3_d[0] && (! lizzieLet43_1Lcall_f3_emitted[4]))};
  assign \q2'a8o_1_destruct_d  = {lizzieLet43_1Lcall_f3_d[99:84],
                                  (lizzieLet43_1Lcall_f3_d[0] && (! lizzieLet43_1Lcall_f3_emitted[5]))};
  assign t2a8t_1_destruct_d = {lizzieLet43_1Lcall_f3_d[115:100],
                               (lizzieLet43_1Lcall_f3_d[0] && (! lizzieLet43_1Lcall_f3_emitted[6]))};
  assign q3a8a_1_destruct_d = {lizzieLet43_1Lcall_f3_d[131:116],
                               (lizzieLet43_1Lcall_f3_d[0] && (! lizzieLet43_1Lcall_f3_emitted[7]))};
  assign \q3'a8p_1_destruct_d  = {lizzieLet43_1Lcall_f3_d[147:132],
                                  (lizzieLet43_1Lcall_f3_d[0] && (! lizzieLet43_1Lcall_f3_emitted[8]))};
  assign t3a8u_1_destruct_d = {lizzieLet43_1Lcall_f3_d[163:148],
                               (lizzieLet43_1Lcall_f3_d[0] && (! lizzieLet43_1Lcall_f3_emitted[9]))};
  assign lizzieLet43_1Lcall_f3_done = (lizzieLet43_1Lcall_f3_emitted | ({t3a8u_1_destruct_d[0],
                                                                         \q3'a8p_1_destruct_d [0],
                                                                         q3a8a_1_destruct_d[0],
                                                                         t2a8t_1_destruct_d[0],
                                                                         \q2'a8o_1_destruct_d [0],
                                                                         q2a89_1_destruct_d[0],
                                                                         t1a8s_1_destruct_d[0],
                                                                         \q1'a8n_1_destruct_d [0],
                                                                         q1a88_1_destruct_d[0],
                                                                         sc_0_3_destruct_d[0]} & {t3a8u_1_destruct_r,
                                                                                                  \q3'a8p_1_destruct_r ,
                                                                                                  q3a8a_1_destruct_r,
                                                                                                  t2a8t_1_destruct_r,
                                                                                                  \q2'a8o_1_destruct_r ,
                                                                                                  q2a89_1_destruct_r,
                                                                                                  t1a8s_1_destruct_r,
                                                                                                  \q1'a8n_1_destruct_r ,
                                                                                                  q1a88_1_destruct_r,
                                                                                                  sc_0_3_destruct_r}));
  assign lizzieLet43_1Lcall_f3_r = (& lizzieLet43_1Lcall_f3_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet43_1Lcall_f3_emitted <= 10'd0;
    else
      lizzieLet43_1Lcall_f3_emitted <= (lizzieLet43_1Lcall_f3_r ? 10'd0 :
                                        lizzieLet43_1Lcall_f3_done);
  
  /* demux (Ty CTf,
       Ty CTf) : (lizzieLet43_2,CTf) (lizzieLet43_1,CTf) > [(_5,CTf),
                                                            (lizzieLet43_1Lcall_f3,CTf),
                                                            (lizzieLet43_1Lcall_f2,CTf),
                                                            (lizzieLet43_1Lcall_f1,CTf),
                                                            (lizzieLet43_1Lcall_f0,CTf)] */
  logic [4:0] lizzieLet43_1_onehotd;
  always_comb
    if ((lizzieLet43_2_d[0] && lizzieLet43_1_d[0]))
      unique case (lizzieLet43_2_d[3:1])
        3'd0: lizzieLet43_1_onehotd = 5'd1;
        3'd1: lizzieLet43_1_onehotd = 5'd2;
        3'd2: lizzieLet43_1_onehotd = 5'd4;
        3'd3: lizzieLet43_1_onehotd = 5'd8;
        3'd4: lizzieLet43_1_onehotd = 5'd16;
        default: lizzieLet43_1_onehotd = 5'd0;
      endcase
    else lizzieLet43_1_onehotd = 5'd0;
  assign _5_d = {lizzieLet43_1_d[163:1], lizzieLet43_1_onehotd[0]};
  assign lizzieLet43_1Lcall_f3_d = {lizzieLet43_1_d[163:1],
                                    lizzieLet43_1_onehotd[1]};
  assign lizzieLet43_1Lcall_f2_d = {lizzieLet43_1_d[163:1],
                                    lizzieLet43_1_onehotd[2]};
  assign lizzieLet43_1Lcall_f1_d = {lizzieLet43_1_d[163:1],
                                    lizzieLet43_1_onehotd[3]};
  assign lizzieLet43_1Lcall_f0_d = {lizzieLet43_1_d[163:1],
                                    lizzieLet43_1_onehotd[4]};
  assign lizzieLet43_1_r = (| (lizzieLet43_1_onehotd & {lizzieLet43_1Lcall_f0_r,
                                                        lizzieLet43_1Lcall_f1_r,
                                                        lizzieLet43_1Lcall_f2_r,
                                                        lizzieLet43_1Lcall_f3_r,
                                                        _5_r}));
  assign lizzieLet43_2_r = lizzieLet43_1_r;
  
  /* demux (Ty CTf,
       Ty Go) : (lizzieLet43_3,CTf) (go_9_goMux_data,Go) > [(_4,Go),
                                                            (lizzieLet43_3Lcall_f3,Go),
                                                            (lizzieLet43_3Lcall_f2,Go),
                                                            (lizzieLet43_3Lcall_f1,Go),
                                                            (lizzieLet43_3Lcall_f0,Go)] */
  logic [4:0] go_9_goMux_data_onehotd;
  always_comb
    if ((lizzieLet43_3_d[0] && go_9_goMux_data_d[0]))
      unique case (lizzieLet43_3_d[3:1])
        3'd0: go_9_goMux_data_onehotd = 5'd1;
        3'd1: go_9_goMux_data_onehotd = 5'd2;
        3'd2: go_9_goMux_data_onehotd = 5'd4;
        3'd3: go_9_goMux_data_onehotd = 5'd8;
        3'd4: go_9_goMux_data_onehotd = 5'd16;
        default: go_9_goMux_data_onehotd = 5'd0;
      endcase
    else go_9_goMux_data_onehotd = 5'd0;
  assign _4_d = go_9_goMux_data_onehotd[0];
  assign lizzieLet43_3Lcall_f3_d = go_9_goMux_data_onehotd[1];
  assign lizzieLet43_3Lcall_f2_d = go_9_goMux_data_onehotd[2];
  assign lizzieLet43_3Lcall_f1_d = go_9_goMux_data_onehotd[3];
  assign lizzieLet43_3Lcall_f0_d = go_9_goMux_data_onehotd[4];
  assign go_9_goMux_data_r = (| (go_9_goMux_data_onehotd & {lizzieLet43_3Lcall_f0_r,
                                                            lizzieLet43_3Lcall_f1_r,
                                                            lizzieLet43_3Lcall_f2_r,
                                                            lizzieLet43_3Lcall_f3_r,
                                                            _4_r}));
  assign lizzieLet43_3_r = go_9_goMux_data_r;
  
  /* buf (Ty Go) : (lizzieLet43_3Lcall_f0,Go) > (lizzieLet43_3Lcall_f0_1_argbuf,Go) */
  Go_t lizzieLet43_3Lcall_f0_bufchan_d;
  logic lizzieLet43_3Lcall_f0_bufchan_r;
  assign lizzieLet43_3Lcall_f0_r = ((! lizzieLet43_3Lcall_f0_bufchan_d[0]) || lizzieLet43_3Lcall_f0_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet43_3Lcall_f0_bufchan_d <= 1'd0;
    else
      if (lizzieLet43_3Lcall_f0_r)
        lizzieLet43_3Lcall_f0_bufchan_d <= lizzieLet43_3Lcall_f0_d;
  Go_t lizzieLet43_3Lcall_f0_bufchan_buf;
  assign lizzieLet43_3Lcall_f0_bufchan_r = (! lizzieLet43_3Lcall_f0_bufchan_buf[0]);
  assign lizzieLet43_3Lcall_f0_1_argbuf_d = (lizzieLet43_3Lcall_f0_bufchan_buf[0] ? lizzieLet43_3Lcall_f0_bufchan_buf :
                                             lizzieLet43_3Lcall_f0_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet43_3Lcall_f0_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet43_3Lcall_f0_1_argbuf_r && lizzieLet43_3Lcall_f0_bufchan_buf[0]))
        lizzieLet43_3Lcall_f0_bufchan_buf <= 1'd0;
      else if (((! lizzieLet43_3Lcall_f0_1_argbuf_r) && (! lizzieLet43_3Lcall_f0_bufchan_buf[0])))
        lizzieLet43_3Lcall_f0_bufchan_buf <= lizzieLet43_3Lcall_f0_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet43_3Lcall_f1,Go) > (lizzieLet43_3Lcall_f1_1_argbuf,Go) */
  Go_t lizzieLet43_3Lcall_f1_bufchan_d;
  logic lizzieLet43_3Lcall_f1_bufchan_r;
  assign lizzieLet43_3Lcall_f1_r = ((! lizzieLet43_3Lcall_f1_bufchan_d[0]) || lizzieLet43_3Lcall_f1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet43_3Lcall_f1_bufchan_d <= 1'd0;
    else
      if (lizzieLet43_3Lcall_f1_r)
        lizzieLet43_3Lcall_f1_bufchan_d <= lizzieLet43_3Lcall_f1_d;
  Go_t lizzieLet43_3Lcall_f1_bufchan_buf;
  assign lizzieLet43_3Lcall_f1_bufchan_r = (! lizzieLet43_3Lcall_f1_bufchan_buf[0]);
  assign lizzieLet43_3Lcall_f1_1_argbuf_d = (lizzieLet43_3Lcall_f1_bufchan_buf[0] ? lizzieLet43_3Lcall_f1_bufchan_buf :
                                             lizzieLet43_3Lcall_f1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet43_3Lcall_f1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet43_3Lcall_f1_1_argbuf_r && lizzieLet43_3Lcall_f1_bufchan_buf[0]))
        lizzieLet43_3Lcall_f1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet43_3Lcall_f1_1_argbuf_r) && (! lizzieLet43_3Lcall_f1_bufchan_buf[0])))
        lizzieLet43_3Lcall_f1_bufchan_buf <= lizzieLet43_3Lcall_f1_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet43_3Lcall_f2,Go) > (lizzieLet43_3Lcall_f2_1_argbuf,Go) */
  Go_t lizzieLet43_3Lcall_f2_bufchan_d;
  logic lizzieLet43_3Lcall_f2_bufchan_r;
  assign lizzieLet43_3Lcall_f2_r = ((! lizzieLet43_3Lcall_f2_bufchan_d[0]) || lizzieLet43_3Lcall_f2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet43_3Lcall_f2_bufchan_d <= 1'd0;
    else
      if (lizzieLet43_3Lcall_f2_r)
        lizzieLet43_3Lcall_f2_bufchan_d <= lizzieLet43_3Lcall_f2_d;
  Go_t lizzieLet43_3Lcall_f2_bufchan_buf;
  assign lizzieLet43_3Lcall_f2_bufchan_r = (! lizzieLet43_3Lcall_f2_bufchan_buf[0]);
  assign lizzieLet43_3Lcall_f2_1_argbuf_d = (lizzieLet43_3Lcall_f2_bufchan_buf[0] ? lizzieLet43_3Lcall_f2_bufchan_buf :
                                             lizzieLet43_3Lcall_f2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet43_3Lcall_f2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet43_3Lcall_f2_1_argbuf_r && lizzieLet43_3Lcall_f2_bufchan_buf[0]))
        lizzieLet43_3Lcall_f2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet43_3Lcall_f2_1_argbuf_r) && (! lizzieLet43_3Lcall_f2_bufchan_buf[0])))
        lizzieLet43_3Lcall_f2_bufchan_buf <= lizzieLet43_3Lcall_f2_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet43_3Lcall_f3,Go) > (lizzieLet43_3Lcall_f3_1_argbuf,Go) */
  Go_t lizzieLet43_3Lcall_f3_bufchan_d;
  logic lizzieLet43_3Lcall_f3_bufchan_r;
  assign lizzieLet43_3Lcall_f3_r = ((! lizzieLet43_3Lcall_f3_bufchan_d[0]) || lizzieLet43_3Lcall_f3_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet43_3Lcall_f3_bufchan_d <= 1'd0;
    else
      if (lizzieLet43_3Lcall_f3_r)
        lizzieLet43_3Lcall_f3_bufchan_d <= lizzieLet43_3Lcall_f3_d;
  Go_t lizzieLet43_3Lcall_f3_bufchan_buf;
  assign lizzieLet43_3Lcall_f3_bufchan_r = (! lizzieLet43_3Lcall_f3_bufchan_buf[0]);
  assign lizzieLet43_3Lcall_f3_1_argbuf_d = (lizzieLet43_3Lcall_f3_bufchan_buf[0] ? lizzieLet43_3Lcall_f3_bufchan_buf :
                                             lizzieLet43_3Lcall_f3_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet43_3Lcall_f3_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet43_3Lcall_f3_1_argbuf_r && lizzieLet43_3Lcall_f3_bufchan_buf[0]))
        lizzieLet43_3Lcall_f3_bufchan_buf <= 1'd0;
      else if (((! lizzieLet43_3Lcall_f3_1_argbuf_r) && (! lizzieLet43_3Lcall_f3_bufchan_buf[0])))
        lizzieLet43_3Lcall_f3_bufchan_buf <= lizzieLet43_3Lcall_f3_bufchan_d;
  
  /* demux (Ty CTf,
       Ty Pointer_QTree_Bool) : (lizzieLet43_4,CTf) (srtarg_0_goMux_mux,Pointer_QTree_Bool) > [(lizzieLet43_4Lfsbos,Pointer_QTree_Bool),
                                                                                               (lizzieLet43_4Lcall_f3,Pointer_QTree_Bool),
                                                                                               (lizzieLet43_4Lcall_f2,Pointer_QTree_Bool),
                                                                                               (lizzieLet43_4Lcall_f1,Pointer_QTree_Bool),
                                                                                               (lizzieLet43_4Lcall_f0,Pointer_QTree_Bool)] */
  logic [4:0] srtarg_0_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet43_4_d[0] && srtarg_0_goMux_mux_d[0]))
      unique case (lizzieLet43_4_d[3:1])
        3'd0: srtarg_0_goMux_mux_onehotd = 5'd1;
        3'd1: srtarg_0_goMux_mux_onehotd = 5'd2;
        3'd2: srtarg_0_goMux_mux_onehotd = 5'd4;
        3'd3: srtarg_0_goMux_mux_onehotd = 5'd8;
        3'd4: srtarg_0_goMux_mux_onehotd = 5'd16;
        default: srtarg_0_goMux_mux_onehotd = 5'd0;
      endcase
    else srtarg_0_goMux_mux_onehotd = 5'd0;
  assign lizzieLet43_4Lfsbos_d = {srtarg_0_goMux_mux_d[16:1],
                                  srtarg_0_goMux_mux_onehotd[0]};
  assign lizzieLet43_4Lcall_f3_d = {srtarg_0_goMux_mux_d[16:1],
                                    srtarg_0_goMux_mux_onehotd[1]};
  assign lizzieLet43_4Lcall_f2_d = {srtarg_0_goMux_mux_d[16:1],
                                    srtarg_0_goMux_mux_onehotd[2]};
  assign lizzieLet43_4Lcall_f1_d = {srtarg_0_goMux_mux_d[16:1],
                                    srtarg_0_goMux_mux_onehotd[3]};
  assign lizzieLet43_4Lcall_f0_d = {srtarg_0_goMux_mux_d[16:1],
                                    srtarg_0_goMux_mux_onehotd[4]};
  assign srtarg_0_goMux_mux_r = (| (srtarg_0_goMux_mux_onehotd & {lizzieLet43_4Lcall_f0_r,
                                                                  lizzieLet43_4Lcall_f1_r,
                                                                  lizzieLet43_4Lcall_f2_r,
                                                                  lizzieLet43_4Lcall_f3_r,
                                                                  lizzieLet43_4Lfsbos_r}));
  assign lizzieLet43_4_r = srtarg_0_goMux_mux_r;
  
  /* dcon (Ty QTree_Bool,
      Dcon QNode_Bool) : [(lizzieLet43_4Lcall_f0,Pointer_QTree_Bool),
                          (es_9_destruct,Pointer_QTree_Bool),
                          (es_10_1_destruct,Pointer_QTree_Bool),
                          (es_11_2_destruct,Pointer_QTree_Bool)] > (lizzieLet43_4Lcall_f0_1es_9_1es_10_1_1es_11_2_1QNode_Bool,QTree_Bool) */
  assign lizzieLet43_4Lcall_f0_1es_9_1es_10_1_1es_11_2_1QNode_Bool_d = QNode_Bool_dc((& {lizzieLet43_4Lcall_f0_d[0],
                                                                                         es_9_destruct_d[0],
                                                                                         es_10_1_destruct_d[0],
                                                                                         es_11_2_destruct_d[0]}), lizzieLet43_4Lcall_f0_d, es_9_destruct_d, es_10_1_destruct_d, es_11_2_destruct_d);
  assign {lizzieLet43_4Lcall_f0_r,
          es_9_destruct_r,
          es_10_1_destruct_r,
          es_11_2_destruct_r} = {4 {(lizzieLet43_4Lcall_f0_1es_9_1es_10_1_1es_11_2_1QNode_Bool_r && lizzieLet43_4Lcall_f0_1es_9_1es_10_1_1es_11_2_1QNode_Bool_d[0])}};
  
  /* buf (Ty QTree_Bool) : (lizzieLet43_4Lcall_f0_1es_9_1es_10_1_1es_11_2_1QNode_Bool,QTree_Bool) > (lizzieLet47_1_argbuf,QTree_Bool) */
  QTree_Bool_t lizzieLet43_4Lcall_f0_1es_9_1es_10_1_1es_11_2_1QNode_Bool_bufchan_d;
  logic lizzieLet43_4Lcall_f0_1es_9_1es_10_1_1es_11_2_1QNode_Bool_bufchan_r;
  assign lizzieLet43_4Lcall_f0_1es_9_1es_10_1_1es_11_2_1QNode_Bool_r = ((! lizzieLet43_4Lcall_f0_1es_9_1es_10_1_1es_11_2_1QNode_Bool_bufchan_d[0]) || lizzieLet43_4Lcall_f0_1es_9_1es_10_1_1es_11_2_1QNode_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet43_4Lcall_f0_1es_9_1es_10_1_1es_11_2_1QNode_Bool_bufchan_d <= {66'd0,
                                                                              1'd0};
    else
      if (lizzieLet43_4Lcall_f0_1es_9_1es_10_1_1es_11_2_1QNode_Bool_r)
        lizzieLet43_4Lcall_f0_1es_9_1es_10_1_1es_11_2_1QNode_Bool_bufchan_d <= lizzieLet43_4Lcall_f0_1es_9_1es_10_1_1es_11_2_1QNode_Bool_d;
  QTree_Bool_t lizzieLet43_4Lcall_f0_1es_9_1es_10_1_1es_11_2_1QNode_Bool_bufchan_buf;
  assign lizzieLet43_4Lcall_f0_1es_9_1es_10_1_1es_11_2_1QNode_Bool_bufchan_r = (! lizzieLet43_4Lcall_f0_1es_9_1es_10_1_1es_11_2_1QNode_Bool_bufchan_buf[0]);
  assign lizzieLet47_1_argbuf_d = (lizzieLet43_4Lcall_f0_1es_9_1es_10_1_1es_11_2_1QNode_Bool_bufchan_buf[0] ? lizzieLet43_4Lcall_f0_1es_9_1es_10_1_1es_11_2_1QNode_Bool_bufchan_buf :
                                   lizzieLet43_4Lcall_f0_1es_9_1es_10_1_1es_11_2_1QNode_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet43_4Lcall_f0_1es_9_1es_10_1_1es_11_2_1QNode_Bool_bufchan_buf <= {66'd0,
                                                                                1'd0};
    else
      if ((lizzieLet47_1_argbuf_r && lizzieLet43_4Lcall_f0_1es_9_1es_10_1_1es_11_2_1QNode_Bool_bufchan_buf[0]))
        lizzieLet43_4Lcall_f0_1es_9_1es_10_1_1es_11_2_1QNode_Bool_bufchan_buf <= {66'd0,
                                                                                  1'd0};
      else if (((! lizzieLet47_1_argbuf_r) && (! lizzieLet43_4Lcall_f0_1es_9_1es_10_1_1es_11_2_1QNode_Bool_bufchan_buf[0])))
        lizzieLet43_4Lcall_f0_1es_9_1es_10_1_1es_11_2_1QNode_Bool_bufchan_buf <= lizzieLet43_4Lcall_f0_1es_9_1es_10_1_1es_11_2_1QNode_Bool_bufchan_d;
  
  /* dcon (Ty CTf,
      Dcon Lcall_f0) : [(lizzieLet43_4Lcall_f1,Pointer_QTree_Bool),
                        (es_10_destruct,Pointer_QTree_Bool),
                        (es_11_1_destruct,Pointer_QTree_Bool),
                        (sc_0_5_destruct,Pointer_CTf)] > (lizzieLet43_4Lcall_f1_1es_10_1es_11_1_1sc_0_5_1Lcall_f0,CTf) */
  assign lizzieLet43_4Lcall_f1_1es_10_1es_11_1_1sc_0_5_1Lcall_f0_d = Lcall_f0_dc((& {lizzieLet43_4Lcall_f1_d[0],
                                                                                     es_10_destruct_d[0],
                                                                                     es_11_1_destruct_d[0],
                                                                                     sc_0_5_destruct_d[0]}), lizzieLet43_4Lcall_f1_d, es_10_destruct_d, es_11_1_destruct_d, sc_0_5_destruct_d);
  assign {lizzieLet43_4Lcall_f1_r,
          es_10_destruct_r,
          es_11_1_destruct_r,
          sc_0_5_destruct_r} = {4 {(lizzieLet43_4Lcall_f1_1es_10_1es_11_1_1sc_0_5_1Lcall_f0_r && lizzieLet43_4Lcall_f1_1es_10_1es_11_1_1sc_0_5_1Lcall_f0_d[0])}};
  
  /* buf (Ty CTf) : (lizzieLet43_4Lcall_f1_1es_10_1es_11_1_1sc_0_5_1Lcall_f0,CTf) > (lizzieLet46_1_argbuf,CTf) */
  CTf_t lizzieLet43_4Lcall_f1_1es_10_1es_11_1_1sc_0_5_1Lcall_f0_bufchan_d;
  logic lizzieLet43_4Lcall_f1_1es_10_1es_11_1_1sc_0_5_1Lcall_f0_bufchan_r;
  assign lizzieLet43_4Lcall_f1_1es_10_1es_11_1_1sc_0_5_1Lcall_f0_r = ((! lizzieLet43_4Lcall_f1_1es_10_1es_11_1_1sc_0_5_1Lcall_f0_bufchan_d[0]) || lizzieLet43_4Lcall_f1_1es_10_1es_11_1_1sc_0_5_1Lcall_f0_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet43_4Lcall_f1_1es_10_1es_11_1_1sc_0_5_1Lcall_f0_bufchan_d <= {163'd0,
                                                                            1'd0};
    else
      if (lizzieLet43_4Lcall_f1_1es_10_1es_11_1_1sc_0_5_1Lcall_f0_r)
        lizzieLet43_4Lcall_f1_1es_10_1es_11_1_1sc_0_5_1Lcall_f0_bufchan_d <= lizzieLet43_4Lcall_f1_1es_10_1es_11_1_1sc_0_5_1Lcall_f0_d;
  CTf_t lizzieLet43_4Lcall_f1_1es_10_1es_11_1_1sc_0_5_1Lcall_f0_bufchan_buf;
  assign lizzieLet43_4Lcall_f1_1es_10_1es_11_1_1sc_0_5_1Lcall_f0_bufchan_r = (! lizzieLet43_4Lcall_f1_1es_10_1es_11_1_1sc_0_5_1Lcall_f0_bufchan_buf[0]);
  assign lizzieLet46_1_argbuf_d = (lizzieLet43_4Lcall_f1_1es_10_1es_11_1_1sc_0_5_1Lcall_f0_bufchan_buf[0] ? lizzieLet43_4Lcall_f1_1es_10_1es_11_1_1sc_0_5_1Lcall_f0_bufchan_buf :
                                   lizzieLet43_4Lcall_f1_1es_10_1es_11_1_1sc_0_5_1Lcall_f0_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet43_4Lcall_f1_1es_10_1es_11_1_1sc_0_5_1Lcall_f0_bufchan_buf <= {163'd0,
                                                                              1'd0};
    else
      if ((lizzieLet46_1_argbuf_r && lizzieLet43_4Lcall_f1_1es_10_1es_11_1_1sc_0_5_1Lcall_f0_bufchan_buf[0]))
        lizzieLet43_4Lcall_f1_1es_10_1es_11_1_1sc_0_5_1Lcall_f0_bufchan_buf <= {163'd0,
                                                                                1'd0};
      else if (((! lizzieLet46_1_argbuf_r) && (! lizzieLet43_4Lcall_f1_1es_10_1es_11_1_1sc_0_5_1Lcall_f0_bufchan_buf[0])))
        lizzieLet43_4Lcall_f1_1es_10_1es_11_1_1sc_0_5_1Lcall_f0_bufchan_buf <= lizzieLet43_4Lcall_f1_1es_10_1es_11_1_1sc_0_5_1Lcall_f0_bufchan_d;
  
  /* dcon (Ty CTf,
      Dcon Lcall_f1) : [(lizzieLet43_4Lcall_f2,Pointer_QTree_Bool),
                        (es_11_destruct,Pointer_QTree_Bool),
                        (sc_0_4_destruct,Pointer_CTf),
                        (q1a88_2_destruct,Pointer_MaskQTree),
                        (q1'a8n_2_destruct,Pointer_QTree_Bool),
                        (t1a8s_2_destruct,Pointer_QTree_Bool)] > (lizzieLet43_4Lcall_f2_1es_11_1sc_0_4_1q1a88_2_1q1'a8n_2_1t1a8s_2_1Lcall_f1,CTf) */
  assign \lizzieLet43_4Lcall_f2_1es_11_1sc_0_4_1q1a88_2_1q1'a8n_2_1t1a8s_2_1Lcall_f1_d  = Lcall_f1_dc((& {lizzieLet43_4Lcall_f2_d[0],
                                                                                                          es_11_destruct_d[0],
                                                                                                          sc_0_4_destruct_d[0],
                                                                                                          q1a88_2_destruct_d[0],
                                                                                                          \q1'a8n_2_destruct_d [0],
                                                                                                          t1a8s_2_destruct_d[0]}), lizzieLet43_4Lcall_f2_d, es_11_destruct_d, sc_0_4_destruct_d, q1a88_2_destruct_d, \q1'a8n_2_destruct_d , t1a8s_2_destruct_d);
  assign {lizzieLet43_4Lcall_f2_r,
          es_11_destruct_r,
          sc_0_4_destruct_r,
          q1a88_2_destruct_r,
          \q1'a8n_2_destruct_r ,
          t1a8s_2_destruct_r} = {6 {(\lizzieLet43_4Lcall_f2_1es_11_1sc_0_4_1q1a88_2_1q1'a8n_2_1t1a8s_2_1Lcall_f1_r  && \lizzieLet43_4Lcall_f2_1es_11_1sc_0_4_1q1a88_2_1q1'a8n_2_1t1a8s_2_1Lcall_f1_d [0])}};
  
  /* buf (Ty CTf) : (lizzieLet43_4Lcall_f2_1es_11_1sc_0_4_1q1a88_2_1q1'a8n_2_1t1a8s_2_1Lcall_f1,CTf) > (lizzieLet45_1_argbuf,CTf) */
  CTf_t \lizzieLet43_4Lcall_f2_1es_11_1sc_0_4_1q1a88_2_1q1'a8n_2_1t1a8s_2_1Lcall_f1_bufchan_d ;
  logic \lizzieLet43_4Lcall_f2_1es_11_1sc_0_4_1q1a88_2_1q1'a8n_2_1t1a8s_2_1Lcall_f1_bufchan_r ;
  assign \lizzieLet43_4Lcall_f2_1es_11_1sc_0_4_1q1a88_2_1q1'a8n_2_1t1a8s_2_1Lcall_f1_r  = ((! \lizzieLet43_4Lcall_f2_1es_11_1sc_0_4_1q1a88_2_1q1'a8n_2_1t1a8s_2_1Lcall_f1_bufchan_d [0]) || \lizzieLet43_4Lcall_f2_1es_11_1sc_0_4_1q1a88_2_1q1'a8n_2_1t1a8s_2_1Lcall_f1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet43_4Lcall_f2_1es_11_1sc_0_4_1q1a88_2_1q1'a8n_2_1t1a8s_2_1Lcall_f1_bufchan_d  <= {163'd0,
                                                                                                 1'd0};
    else
      if (\lizzieLet43_4Lcall_f2_1es_11_1sc_0_4_1q1a88_2_1q1'a8n_2_1t1a8s_2_1Lcall_f1_r )
        \lizzieLet43_4Lcall_f2_1es_11_1sc_0_4_1q1a88_2_1q1'a8n_2_1t1a8s_2_1Lcall_f1_bufchan_d  <= \lizzieLet43_4Lcall_f2_1es_11_1sc_0_4_1q1a88_2_1q1'a8n_2_1t1a8s_2_1Lcall_f1_d ;
  CTf_t \lizzieLet43_4Lcall_f2_1es_11_1sc_0_4_1q1a88_2_1q1'a8n_2_1t1a8s_2_1Lcall_f1_bufchan_buf ;
  assign \lizzieLet43_4Lcall_f2_1es_11_1sc_0_4_1q1a88_2_1q1'a8n_2_1t1a8s_2_1Lcall_f1_bufchan_r  = (! \lizzieLet43_4Lcall_f2_1es_11_1sc_0_4_1q1a88_2_1q1'a8n_2_1t1a8s_2_1Lcall_f1_bufchan_buf [0]);
  assign lizzieLet45_1_argbuf_d = (\lizzieLet43_4Lcall_f2_1es_11_1sc_0_4_1q1a88_2_1q1'a8n_2_1t1a8s_2_1Lcall_f1_bufchan_buf [0] ? \lizzieLet43_4Lcall_f2_1es_11_1sc_0_4_1q1a88_2_1q1'a8n_2_1t1a8s_2_1Lcall_f1_bufchan_buf  :
                                   \lizzieLet43_4Lcall_f2_1es_11_1sc_0_4_1q1a88_2_1q1'a8n_2_1t1a8s_2_1Lcall_f1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet43_4Lcall_f2_1es_11_1sc_0_4_1q1a88_2_1q1'a8n_2_1t1a8s_2_1Lcall_f1_bufchan_buf  <= {163'd0,
                                                                                                   1'd0};
    else
      if ((lizzieLet45_1_argbuf_r && \lizzieLet43_4Lcall_f2_1es_11_1sc_0_4_1q1a88_2_1q1'a8n_2_1t1a8s_2_1Lcall_f1_bufchan_buf [0]))
        \lizzieLet43_4Lcall_f2_1es_11_1sc_0_4_1q1a88_2_1q1'a8n_2_1t1a8s_2_1Lcall_f1_bufchan_buf  <= {163'd0,
                                                                                                     1'd0};
      else if (((! lizzieLet45_1_argbuf_r) && (! \lizzieLet43_4Lcall_f2_1es_11_1sc_0_4_1q1a88_2_1q1'a8n_2_1t1a8s_2_1Lcall_f1_bufchan_buf [0])))
        \lizzieLet43_4Lcall_f2_1es_11_1sc_0_4_1q1a88_2_1q1'a8n_2_1t1a8s_2_1Lcall_f1_bufchan_buf  <= \lizzieLet43_4Lcall_f2_1es_11_1sc_0_4_1q1a88_2_1q1'a8n_2_1t1a8s_2_1Lcall_f1_bufchan_d ;
  
  /* dcon (Ty CTf,
      Dcon Lcall_f2) : [(lizzieLet43_4Lcall_f3,Pointer_QTree_Bool),
                        (sc_0_3_destruct,Pointer_CTf),
                        (q1a88_1_destruct,Pointer_MaskQTree),
                        (q1'a8n_1_destruct,Pointer_QTree_Bool),
                        (t1a8s_1_destruct,Pointer_QTree_Bool),
                        (q2a89_1_destruct,Pointer_MaskQTree),
                        (q2'a8o_1_destruct,Pointer_QTree_Bool),
                        (t2a8t_1_destruct,Pointer_QTree_Bool)] > (lizzieLet43_4Lcall_f3_1sc_0_3_1q1a88_1_1q1'a8n_1_1t1a8s_1_1q2a89_1_1q2'a8o_1_1t2a8t_1_1Lcall_f2,CTf) */
  assign \lizzieLet43_4Lcall_f3_1sc_0_3_1q1a88_1_1q1'a8n_1_1t1a8s_1_1q2a89_1_1q2'a8o_1_1t2a8t_1_1Lcall_f2_d  = Lcall_f2_dc((& {lizzieLet43_4Lcall_f3_d[0],
                                                                                                                               sc_0_3_destruct_d[0],
                                                                                                                               q1a88_1_destruct_d[0],
                                                                                                                               \q1'a8n_1_destruct_d [0],
                                                                                                                               t1a8s_1_destruct_d[0],
                                                                                                                               q2a89_1_destruct_d[0],
                                                                                                                               \q2'a8o_1_destruct_d [0],
                                                                                                                               t2a8t_1_destruct_d[0]}), lizzieLet43_4Lcall_f3_d, sc_0_3_destruct_d, q1a88_1_destruct_d, \q1'a8n_1_destruct_d , t1a8s_1_destruct_d, q2a89_1_destruct_d, \q2'a8o_1_destruct_d , t2a8t_1_destruct_d);
  assign {lizzieLet43_4Lcall_f3_r,
          sc_0_3_destruct_r,
          q1a88_1_destruct_r,
          \q1'a8n_1_destruct_r ,
          t1a8s_1_destruct_r,
          q2a89_1_destruct_r,
          \q2'a8o_1_destruct_r ,
          t2a8t_1_destruct_r} = {8 {(\lizzieLet43_4Lcall_f3_1sc_0_3_1q1a88_1_1q1'a8n_1_1t1a8s_1_1q2a89_1_1q2'a8o_1_1t2a8t_1_1Lcall_f2_r  && \lizzieLet43_4Lcall_f3_1sc_0_3_1q1a88_1_1q1'a8n_1_1t1a8s_1_1q2a89_1_1q2'a8o_1_1t2a8t_1_1Lcall_f2_d [0])}};
  
  /* buf (Ty CTf) : (lizzieLet43_4Lcall_f3_1sc_0_3_1q1a88_1_1q1'a8n_1_1t1a8s_1_1q2a89_1_1q2'a8o_1_1t2a8t_1_1Lcall_f2,CTf) > (lizzieLet44_1_argbuf,CTf) */
  CTf_t \lizzieLet43_4Lcall_f3_1sc_0_3_1q1a88_1_1q1'a8n_1_1t1a8s_1_1q2a89_1_1q2'a8o_1_1t2a8t_1_1Lcall_f2_bufchan_d ;
  logic \lizzieLet43_4Lcall_f3_1sc_0_3_1q1a88_1_1q1'a8n_1_1t1a8s_1_1q2a89_1_1q2'a8o_1_1t2a8t_1_1Lcall_f2_bufchan_r ;
  assign \lizzieLet43_4Lcall_f3_1sc_0_3_1q1a88_1_1q1'a8n_1_1t1a8s_1_1q2a89_1_1q2'a8o_1_1t2a8t_1_1Lcall_f2_r  = ((! \lizzieLet43_4Lcall_f3_1sc_0_3_1q1a88_1_1q1'a8n_1_1t1a8s_1_1q2a89_1_1q2'a8o_1_1t2a8t_1_1Lcall_f2_bufchan_d [0]) || \lizzieLet43_4Lcall_f3_1sc_0_3_1q1a88_1_1q1'a8n_1_1t1a8s_1_1q2a89_1_1q2'a8o_1_1t2a8t_1_1Lcall_f2_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet43_4Lcall_f3_1sc_0_3_1q1a88_1_1q1'a8n_1_1t1a8s_1_1q2a89_1_1q2'a8o_1_1t2a8t_1_1Lcall_f2_bufchan_d  <= {163'd0,
                                                                                                                      1'd0};
    else
      if (\lizzieLet43_4Lcall_f3_1sc_0_3_1q1a88_1_1q1'a8n_1_1t1a8s_1_1q2a89_1_1q2'a8o_1_1t2a8t_1_1Lcall_f2_r )
        \lizzieLet43_4Lcall_f3_1sc_0_3_1q1a88_1_1q1'a8n_1_1t1a8s_1_1q2a89_1_1q2'a8o_1_1t2a8t_1_1Lcall_f2_bufchan_d  <= \lizzieLet43_4Lcall_f3_1sc_0_3_1q1a88_1_1q1'a8n_1_1t1a8s_1_1q2a89_1_1q2'a8o_1_1t2a8t_1_1Lcall_f2_d ;
  CTf_t \lizzieLet43_4Lcall_f3_1sc_0_3_1q1a88_1_1q1'a8n_1_1t1a8s_1_1q2a89_1_1q2'a8o_1_1t2a8t_1_1Lcall_f2_bufchan_buf ;
  assign \lizzieLet43_4Lcall_f3_1sc_0_3_1q1a88_1_1q1'a8n_1_1t1a8s_1_1q2a89_1_1q2'a8o_1_1t2a8t_1_1Lcall_f2_bufchan_r  = (! \lizzieLet43_4Lcall_f3_1sc_0_3_1q1a88_1_1q1'a8n_1_1t1a8s_1_1q2a89_1_1q2'a8o_1_1t2a8t_1_1Lcall_f2_bufchan_buf [0]);
  assign lizzieLet44_1_argbuf_d = (\lizzieLet43_4Lcall_f3_1sc_0_3_1q1a88_1_1q1'a8n_1_1t1a8s_1_1q2a89_1_1q2'a8o_1_1t2a8t_1_1Lcall_f2_bufchan_buf [0] ? \lizzieLet43_4Lcall_f3_1sc_0_3_1q1a88_1_1q1'a8n_1_1t1a8s_1_1q2a89_1_1q2'a8o_1_1t2a8t_1_1Lcall_f2_bufchan_buf  :
                                   \lizzieLet43_4Lcall_f3_1sc_0_3_1q1a88_1_1q1'a8n_1_1t1a8s_1_1q2a89_1_1q2'a8o_1_1t2a8t_1_1Lcall_f2_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet43_4Lcall_f3_1sc_0_3_1q1a88_1_1q1'a8n_1_1t1a8s_1_1q2a89_1_1q2'a8o_1_1t2a8t_1_1Lcall_f2_bufchan_buf  <= {163'd0,
                                                                                                                        1'd0};
    else
      if ((lizzieLet44_1_argbuf_r && \lizzieLet43_4Lcall_f3_1sc_0_3_1q1a88_1_1q1'a8n_1_1t1a8s_1_1q2a89_1_1q2'a8o_1_1t2a8t_1_1Lcall_f2_bufchan_buf [0]))
        \lizzieLet43_4Lcall_f3_1sc_0_3_1q1a88_1_1q1'a8n_1_1t1a8s_1_1q2a89_1_1q2'a8o_1_1t2a8t_1_1Lcall_f2_bufchan_buf  <= {163'd0,
                                                                                                                          1'd0};
      else if (((! lizzieLet44_1_argbuf_r) && (! \lizzieLet43_4Lcall_f3_1sc_0_3_1q1a88_1_1q1'a8n_1_1t1a8s_1_1q2a89_1_1q2'a8o_1_1t2a8t_1_1Lcall_f2_bufchan_buf [0])))
        \lizzieLet43_4Lcall_f3_1sc_0_3_1q1a88_1_1q1'a8n_1_1t1a8s_1_1q2a89_1_1q2'a8o_1_1t2a8t_1_1Lcall_f2_bufchan_buf  <= \lizzieLet43_4Lcall_f3_1sc_0_3_1q1a88_1_1q1'a8n_1_1t1a8s_1_1q2a89_1_1q2'a8o_1_1t2a8t_1_1Lcall_f2_bufchan_d ;
  
  /* fork (Ty Pointer_QTree_Bool) : (lizzieLet43_4Lfsbos,Pointer_QTree_Bool) > [(lizzieLet43_4Lfsbos_1_merge_merge_fork_1,Pointer_QTree_Bool),
                                                                           (lizzieLet43_4Lfsbos_1_merge_merge_fork_2,Pointer_QTree_Bool)] */
  logic [1:0] lizzieLet43_4Lfsbos_emitted;
  logic [1:0] lizzieLet43_4Lfsbos_done;
  assign lizzieLet43_4Lfsbos_1_merge_merge_fork_1_d = {lizzieLet43_4Lfsbos_d[16:1],
                                                       (lizzieLet43_4Lfsbos_d[0] && (! lizzieLet43_4Lfsbos_emitted[0]))};
  assign lizzieLet43_4Lfsbos_1_merge_merge_fork_2_d = {lizzieLet43_4Lfsbos_d[16:1],
                                                       (lizzieLet43_4Lfsbos_d[0] && (! lizzieLet43_4Lfsbos_emitted[1]))};
  assign lizzieLet43_4Lfsbos_done = (lizzieLet43_4Lfsbos_emitted | ({lizzieLet43_4Lfsbos_1_merge_merge_fork_2_d[0],
                                                                     lizzieLet43_4Lfsbos_1_merge_merge_fork_1_d[0]} & {lizzieLet43_4Lfsbos_1_merge_merge_fork_2_r,
                                                                                                                       lizzieLet43_4Lfsbos_1_merge_merge_fork_1_r}));
  assign lizzieLet43_4Lfsbos_r = (& lizzieLet43_4Lfsbos_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet43_4Lfsbos_emitted <= 2'd0;
    else
      lizzieLet43_4Lfsbos_emitted <= (lizzieLet43_4Lfsbos_r ? 2'd0 :
                                      lizzieLet43_4Lfsbos_done);
  
  /* togo (Ty Pointer_QTree_Bool) : (lizzieLet43_4Lfsbos_1_merge_merge_fork_1,Pointer_QTree_Bool) > (call_f_goConst,Go) */
  assign call_f_goConst_d = lizzieLet43_4Lfsbos_1_merge_merge_fork_1_d[0];
  assign lizzieLet43_4Lfsbos_1_merge_merge_fork_1_r = call_f_goConst_r;
  
  /* buf (Ty Pointer_QTree_Bool) : (lizzieLet43_4Lfsbos_1_merge_merge_fork_2,Pointer_QTree_Bool) > (f_resbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t lizzieLet43_4Lfsbos_1_merge_merge_fork_2_bufchan_d;
  logic lizzieLet43_4Lfsbos_1_merge_merge_fork_2_bufchan_r;
  assign lizzieLet43_4Lfsbos_1_merge_merge_fork_2_r = ((! lizzieLet43_4Lfsbos_1_merge_merge_fork_2_bufchan_d[0]) || lizzieLet43_4Lfsbos_1_merge_merge_fork_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet43_4Lfsbos_1_merge_merge_fork_2_bufchan_d <= {16'd0,
                                                             1'd0};
    else
      if (lizzieLet43_4Lfsbos_1_merge_merge_fork_2_r)
        lizzieLet43_4Lfsbos_1_merge_merge_fork_2_bufchan_d <= lizzieLet43_4Lfsbos_1_merge_merge_fork_2_d;
  Pointer_QTree_Bool_t lizzieLet43_4Lfsbos_1_merge_merge_fork_2_bufchan_buf;
  assign lizzieLet43_4Lfsbos_1_merge_merge_fork_2_bufchan_r = (! lizzieLet43_4Lfsbos_1_merge_merge_fork_2_bufchan_buf[0]);
  assign f_resbuf_d = (lizzieLet43_4Lfsbos_1_merge_merge_fork_2_bufchan_buf[0] ? lizzieLet43_4Lfsbos_1_merge_merge_fork_2_bufchan_buf :
                       lizzieLet43_4Lfsbos_1_merge_merge_fork_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet43_4Lfsbos_1_merge_merge_fork_2_bufchan_buf <= {16'd0,
                                                               1'd0};
    else
      if ((f_resbuf_r && lizzieLet43_4Lfsbos_1_merge_merge_fork_2_bufchan_buf[0]))
        lizzieLet43_4Lfsbos_1_merge_merge_fork_2_bufchan_buf <= {16'd0,
                                                                 1'd0};
      else if (((! f_resbuf_r) && (! lizzieLet43_4Lfsbos_1_merge_merge_fork_2_bufchan_buf[0])))
        lizzieLet43_4Lfsbos_1_merge_merge_fork_2_bufchan_buf <= lizzieLet43_4Lfsbos_1_merge_merge_fork_2_bufchan_d;
  
  /* destruct (Ty CTf',
          Dcon Lcall_f'0) : (lizzieLet48_1Lcall_f'0,CTf') > [(es_1_1_destruct,Pointer_QTree_Bool),
                                                             (es_2_2_destruct,Pointer_QTree_Bool),
                                                             (es_3_3_destruct,Pointer_QTree_Bool),
                                                             (sc_0_10_destruct,Pointer_CTf')] */
  logic [3:0] \lizzieLet48_1Lcall_f'0_emitted ;
  logic [3:0] \lizzieLet48_1Lcall_f'0_done ;
  assign es_1_1_destruct_d = {\lizzieLet48_1Lcall_f'0_d [19:4],
                              (\lizzieLet48_1Lcall_f'0_d [0] && (! \lizzieLet48_1Lcall_f'0_emitted [0]))};
  assign es_2_2_destruct_d = {\lizzieLet48_1Lcall_f'0_d [35:20],
                              (\lizzieLet48_1Lcall_f'0_d [0] && (! \lizzieLet48_1Lcall_f'0_emitted [1]))};
  assign es_3_3_destruct_d = {\lizzieLet48_1Lcall_f'0_d [51:36],
                              (\lizzieLet48_1Lcall_f'0_d [0] && (! \lizzieLet48_1Lcall_f'0_emitted [2]))};
  assign sc_0_10_destruct_d = {\lizzieLet48_1Lcall_f'0_d [67:52],
                               (\lizzieLet48_1Lcall_f'0_d [0] && (! \lizzieLet48_1Lcall_f'0_emitted [3]))};
  assign \lizzieLet48_1Lcall_f'0_done  = (\lizzieLet48_1Lcall_f'0_emitted  | ({sc_0_10_destruct_d[0],
                                                                               es_3_3_destruct_d[0],
                                                                               es_2_2_destruct_d[0],
                                                                               es_1_1_destruct_d[0]} & {sc_0_10_destruct_r,
                                                                                                        es_3_3_destruct_r,
                                                                                                        es_2_2_destruct_r,
                                                                                                        es_1_1_destruct_r}));
  assign \lizzieLet48_1Lcall_f'0_r  = (& \lizzieLet48_1Lcall_f'0_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \lizzieLet48_1Lcall_f'0_emitted  <= 4'd0;
    else
      \lizzieLet48_1Lcall_f'0_emitted  <= (\lizzieLet48_1Lcall_f'0_r  ? 4'd0 :
                                           \lizzieLet48_1Lcall_f'0_done );
  
  /* destruct (Ty CTf',
          Dcon Lcall_f'1) : (lizzieLet48_1Lcall_f'1,CTf') > [(es_2_1_destruct,Pointer_QTree_Bool),
                                                             (es_3_2_destruct,Pointer_QTree_Bool),
                                                             (sc_0_9_destruct,Pointer_CTf'),
                                                             (q1a8P_3_destruct,Pointer_QTree_Bool),
                                                             (t1a8U_3_destruct,Pointer_QTree_Bool)] */
  logic [4:0] \lizzieLet48_1Lcall_f'1_emitted ;
  logic [4:0] \lizzieLet48_1Lcall_f'1_done ;
  assign es_2_1_destruct_d = {\lizzieLet48_1Lcall_f'1_d [19:4],
                              (\lizzieLet48_1Lcall_f'1_d [0] && (! \lizzieLet48_1Lcall_f'1_emitted [0]))};
  assign es_3_2_destruct_d = {\lizzieLet48_1Lcall_f'1_d [35:20],
                              (\lizzieLet48_1Lcall_f'1_d [0] && (! \lizzieLet48_1Lcall_f'1_emitted [1]))};
  assign sc_0_9_destruct_d = {\lizzieLet48_1Lcall_f'1_d [51:36],
                              (\lizzieLet48_1Lcall_f'1_d [0] && (! \lizzieLet48_1Lcall_f'1_emitted [2]))};
  assign q1a8P_3_destruct_d = {\lizzieLet48_1Lcall_f'1_d [67:52],
                               (\lizzieLet48_1Lcall_f'1_d [0] && (! \lizzieLet48_1Lcall_f'1_emitted [3]))};
  assign t1a8U_3_destruct_d = {\lizzieLet48_1Lcall_f'1_d [83:68],
                               (\lizzieLet48_1Lcall_f'1_d [0] && (! \lizzieLet48_1Lcall_f'1_emitted [4]))};
  assign \lizzieLet48_1Lcall_f'1_done  = (\lizzieLet48_1Lcall_f'1_emitted  | ({t1a8U_3_destruct_d[0],
                                                                               q1a8P_3_destruct_d[0],
                                                                               sc_0_9_destruct_d[0],
                                                                               es_3_2_destruct_d[0],
                                                                               es_2_1_destruct_d[0]} & {t1a8U_3_destruct_r,
                                                                                                        q1a8P_3_destruct_r,
                                                                                                        sc_0_9_destruct_r,
                                                                                                        es_3_2_destruct_r,
                                                                                                        es_2_1_destruct_r}));
  assign \lizzieLet48_1Lcall_f'1_r  = (& \lizzieLet48_1Lcall_f'1_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \lizzieLet48_1Lcall_f'1_emitted  <= 5'd0;
    else
      \lizzieLet48_1Lcall_f'1_emitted  <= (\lizzieLet48_1Lcall_f'1_r  ? 5'd0 :
                                           \lizzieLet48_1Lcall_f'1_done );
  
  /* destruct (Ty CTf',
          Dcon Lcall_f'2) : (lizzieLet48_1Lcall_f'2,CTf') > [(es_3_1_destruct,Pointer_QTree_Bool),
                                                             (sc_0_8_destruct,Pointer_CTf'),
                                                             (q1a8P_2_destruct,Pointer_QTree_Bool),
                                                             (t1a8U_2_destruct,Pointer_QTree_Bool),
                                                             (q2a8Q_2_destruct,Pointer_QTree_Bool),
                                                             (t2a8V_2_destruct,Pointer_QTree_Bool)] */
  logic [5:0] \lizzieLet48_1Lcall_f'2_emitted ;
  logic [5:0] \lizzieLet48_1Lcall_f'2_done ;
  assign es_3_1_destruct_d = {\lizzieLet48_1Lcall_f'2_d [19:4],
                              (\lizzieLet48_1Lcall_f'2_d [0] && (! \lizzieLet48_1Lcall_f'2_emitted [0]))};
  assign sc_0_8_destruct_d = {\lizzieLet48_1Lcall_f'2_d [35:20],
                              (\lizzieLet48_1Lcall_f'2_d [0] && (! \lizzieLet48_1Lcall_f'2_emitted [1]))};
  assign q1a8P_2_destruct_d = {\lizzieLet48_1Lcall_f'2_d [51:36],
                               (\lizzieLet48_1Lcall_f'2_d [0] && (! \lizzieLet48_1Lcall_f'2_emitted [2]))};
  assign t1a8U_2_destruct_d = {\lizzieLet48_1Lcall_f'2_d [67:52],
                               (\lizzieLet48_1Lcall_f'2_d [0] && (! \lizzieLet48_1Lcall_f'2_emitted [3]))};
  assign q2a8Q_2_destruct_d = {\lizzieLet48_1Lcall_f'2_d [83:68],
                               (\lizzieLet48_1Lcall_f'2_d [0] && (! \lizzieLet48_1Lcall_f'2_emitted [4]))};
  assign t2a8V_2_destruct_d = {\lizzieLet48_1Lcall_f'2_d [99:84],
                               (\lizzieLet48_1Lcall_f'2_d [0] && (! \lizzieLet48_1Lcall_f'2_emitted [5]))};
  assign \lizzieLet48_1Lcall_f'2_done  = (\lizzieLet48_1Lcall_f'2_emitted  | ({t2a8V_2_destruct_d[0],
                                                                               q2a8Q_2_destruct_d[0],
                                                                               t1a8U_2_destruct_d[0],
                                                                               q1a8P_2_destruct_d[0],
                                                                               sc_0_8_destruct_d[0],
                                                                               es_3_1_destruct_d[0]} & {t2a8V_2_destruct_r,
                                                                                                        q2a8Q_2_destruct_r,
                                                                                                        t1a8U_2_destruct_r,
                                                                                                        q1a8P_2_destruct_r,
                                                                                                        sc_0_8_destruct_r,
                                                                                                        es_3_1_destruct_r}));
  assign \lizzieLet48_1Lcall_f'2_r  = (& \lizzieLet48_1Lcall_f'2_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \lizzieLet48_1Lcall_f'2_emitted  <= 6'd0;
    else
      \lizzieLet48_1Lcall_f'2_emitted  <= (\lizzieLet48_1Lcall_f'2_r  ? 6'd0 :
                                           \lizzieLet48_1Lcall_f'2_done );
  
  /* destruct (Ty CTf',
          Dcon Lcall_f'3) : (lizzieLet48_1Lcall_f'3,CTf') > [(sc_0_7_destruct,Pointer_CTf'),
                                                             (q1a8P_1_destruct,Pointer_QTree_Bool),
                                                             (t1a8U_1_destruct,Pointer_QTree_Bool),
                                                             (q2a8Q_1_destruct,Pointer_QTree_Bool),
                                                             (t2a8V_1_destruct,Pointer_QTree_Bool),
                                                             (q3a8R_1_destruct,Pointer_QTree_Bool),
                                                             (t3a8W_1_destruct,Pointer_QTree_Bool)] */
  logic [6:0] \lizzieLet48_1Lcall_f'3_emitted ;
  logic [6:0] \lizzieLet48_1Lcall_f'3_done ;
  assign sc_0_7_destruct_d = {\lizzieLet48_1Lcall_f'3_d [19:4],
                              (\lizzieLet48_1Lcall_f'3_d [0] && (! \lizzieLet48_1Lcall_f'3_emitted [0]))};
  assign q1a8P_1_destruct_d = {\lizzieLet48_1Lcall_f'3_d [35:20],
                               (\lizzieLet48_1Lcall_f'3_d [0] && (! \lizzieLet48_1Lcall_f'3_emitted [1]))};
  assign t1a8U_1_destruct_d = {\lizzieLet48_1Lcall_f'3_d [51:36],
                               (\lizzieLet48_1Lcall_f'3_d [0] && (! \lizzieLet48_1Lcall_f'3_emitted [2]))};
  assign q2a8Q_1_destruct_d = {\lizzieLet48_1Lcall_f'3_d [67:52],
                               (\lizzieLet48_1Lcall_f'3_d [0] && (! \lizzieLet48_1Lcall_f'3_emitted [3]))};
  assign t2a8V_1_destruct_d = {\lizzieLet48_1Lcall_f'3_d [83:68],
                               (\lizzieLet48_1Lcall_f'3_d [0] && (! \lizzieLet48_1Lcall_f'3_emitted [4]))};
  assign q3a8R_1_destruct_d = {\lizzieLet48_1Lcall_f'3_d [99:84],
                               (\lizzieLet48_1Lcall_f'3_d [0] && (! \lizzieLet48_1Lcall_f'3_emitted [5]))};
  assign t3a8W_1_destruct_d = {\lizzieLet48_1Lcall_f'3_d [115:100],
                               (\lizzieLet48_1Lcall_f'3_d [0] && (! \lizzieLet48_1Lcall_f'3_emitted [6]))};
  assign \lizzieLet48_1Lcall_f'3_done  = (\lizzieLet48_1Lcall_f'3_emitted  | ({t3a8W_1_destruct_d[0],
                                                                               q3a8R_1_destruct_d[0],
                                                                               t2a8V_1_destruct_d[0],
                                                                               q2a8Q_1_destruct_d[0],
                                                                               t1a8U_1_destruct_d[0],
                                                                               q1a8P_1_destruct_d[0],
                                                                               sc_0_7_destruct_d[0]} & {t3a8W_1_destruct_r,
                                                                                                        q3a8R_1_destruct_r,
                                                                                                        t2a8V_1_destruct_r,
                                                                                                        q2a8Q_1_destruct_r,
                                                                                                        t1a8U_1_destruct_r,
                                                                                                        q1a8P_1_destruct_r,
                                                                                                        sc_0_7_destruct_r}));
  assign \lizzieLet48_1Lcall_f'3_r  = (& \lizzieLet48_1Lcall_f'3_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \lizzieLet48_1Lcall_f'3_emitted  <= 7'd0;
    else
      \lizzieLet48_1Lcall_f'3_emitted  <= (\lizzieLet48_1Lcall_f'3_r  ? 7'd0 :
                                           \lizzieLet48_1Lcall_f'3_done );
  
  /* demux (Ty CTf',
       Ty CTf') : (lizzieLet48_2,CTf') (lizzieLet48_1,CTf') > [(_3,CTf'),
                                                               (lizzieLet48_1Lcall_f'3,CTf'),
                                                               (lizzieLet48_1Lcall_f'2,CTf'),
                                                               (lizzieLet48_1Lcall_f'1,CTf'),
                                                               (lizzieLet48_1Lcall_f'0,CTf')] */
  logic [4:0] lizzieLet48_1_onehotd;
  always_comb
    if ((lizzieLet48_2_d[0] && lizzieLet48_1_d[0]))
      unique case (lizzieLet48_2_d[3:1])
        3'd0: lizzieLet48_1_onehotd = 5'd1;
        3'd1: lizzieLet48_1_onehotd = 5'd2;
        3'd2: lizzieLet48_1_onehotd = 5'd4;
        3'd3: lizzieLet48_1_onehotd = 5'd8;
        3'd4: lizzieLet48_1_onehotd = 5'd16;
        default: lizzieLet48_1_onehotd = 5'd0;
      endcase
    else lizzieLet48_1_onehotd = 5'd0;
  assign _3_d = {lizzieLet48_1_d[115:1], lizzieLet48_1_onehotd[0]};
  assign \lizzieLet48_1Lcall_f'3_d  = {lizzieLet48_1_d[115:1],
                                       lizzieLet48_1_onehotd[1]};
  assign \lizzieLet48_1Lcall_f'2_d  = {lizzieLet48_1_d[115:1],
                                       lizzieLet48_1_onehotd[2]};
  assign \lizzieLet48_1Lcall_f'1_d  = {lizzieLet48_1_d[115:1],
                                       lizzieLet48_1_onehotd[3]};
  assign \lizzieLet48_1Lcall_f'0_d  = {lizzieLet48_1_d[115:1],
                                       lizzieLet48_1_onehotd[4]};
  assign lizzieLet48_1_r = (| (lizzieLet48_1_onehotd & {\lizzieLet48_1Lcall_f'0_r ,
                                                        \lizzieLet48_1Lcall_f'1_r ,
                                                        \lizzieLet48_1Lcall_f'2_r ,
                                                        \lizzieLet48_1Lcall_f'3_r ,
                                                        _3_r}));
  assign lizzieLet48_2_r = lizzieLet48_1_r;
  
  /* demux (Ty CTf',
       Ty Go) : (lizzieLet48_3,CTf') (go_10_goMux_data,Go) > [(_2,Go),
                                                              (lizzieLet48_3Lcall_f'3,Go),
                                                              (lizzieLet48_3Lcall_f'2,Go),
                                                              (lizzieLet48_3Lcall_f'1,Go),
                                                              (lizzieLet48_3Lcall_f'0,Go)] */
  logic [4:0] go_10_goMux_data_onehotd;
  always_comb
    if ((lizzieLet48_3_d[0] && go_10_goMux_data_d[0]))
      unique case (lizzieLet48_3_d[3:1])
        3'd0: go_10_goMux_data_onehotd = 5'd1;
        3'd1: go_10_goMux_data_onehotd = 5'd2;
        3'd2: go_10_goMux_data_onehotd = 5'd4;
        3'd3: go_10_goMux_data_onehotd = 5'd8;
        3'd4: go_10_goMux_data_onehotd = 5'd16;
        default: go_10_goMux_data_onehotd = 5'd0;
      endcase
    else go_10_goMux_data_onehotd = 5'd0;
  assign _2_d = go_10_goMux_data_onehotd[0];
  assign \lizzieLet48_3Lcall_f'3_d  = go_10_goMux_data_onehotd[1];
  assign \lizzieLet48_3Lcall_f'2_d  = go_10_goMux_data_onehotd[2];
  assign \lizzieLet48_3Lcall_f'1_d  = go_10_goMux_data_onehotd[3];
  assign \lizzieLet48_3Lcall_f'0_d  = go_10_goMux_data_onehotd[4];
  assign go_10_goMux_data_r = (| (go_10_goMux_data_onehotd & {\lizzieLet48_3Lcall_f'0_r ,
                                                              \lizzieLet48_3Lcall_f'1_r ,
                                                              \lizzieLet48_3Lcall_f'2_r ,
                                                              \lizzieLet48_3Lcall_f'3_r ,
                                                              _2_r}));
  assign lizzieLet48_3_r = go_10_goMux_data_r;
  
  /* buf (Ty Go) : (lizzieLet48_3Lcall_f'0,Go) > (lizzieLet48_3Lcall_f'0_1_argbuf,Go) */
  Go_t \lizzieLet48_3Lcall_f'0_bufchan_d ;
  logic \lizzieLet48_3Lcall_f'0_bufchan_r ;
  assign \lizzieLet48_3Lcall_f'0_r  = ((! \lizzieLet48_3Lcall_f'0_bufchan_d [0]) || \lizzieLet48_3Lcall_f'0_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \lizzieLet48_3Lcall_f'0_bufchan_d  <= 1'd0;
    else
      if (\lizzieLet48_3Lcall_f'0_r )
        \lizzieLet48_3Lcall_f'0_bufchan_d  <= \lizzieLet48_3Lcall_f'0_d ;
  Go_t \lizzieLet48_3Lcall_f'0_bufchan_buf ;
  assign \lizzieLet48_3Lcall_f'0_bufchan_r  = (! \lizzieLet48_3Lcall_f'0_bufchan_buf [0]);
  assign \lizzieLet48_3Lcall_f'0_1_argbuf_d  = (\lizzieLet48_3Lcall_f'0_bufchan_buf [0] ? \lizzieLet48_3Lcall_f'0_bufchan_buf  :
                                                \lizzieLet48_3Lcall_f'0_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \lizzieLet48_3Lcall_f'0_bufchan_buf  <= 1'd0;
    else
      if ((\lizzieLet48_3Lcall_f'0_1_argbuf_r  && \lizzieLet48_3Lcall_f'0_bufchan_buf [0]))
        \lizzieLet48_3Lcall_f'0_bufchan_buf  <= 1'd0;
      else if (((! \lizzieLet48_3Lcall_f'0_1_argbuf_r ) && (! \lizzieLet48_3Lcall_f'0_bufchan_buf [0])))
        \lizzieLet48_3Lcall_f'0_bufchan_buf  <= \lizzieLet48_3Lcall_f'0_bufchan_d ;
  
  /* buf (Ty Go) : (lizzieLet48_3Lcall_f'1,Go) > (lizzieLet48_3Lcall_f'1_1_argbuf,Go) */
  Go_t \lizzieLet48_3Lcall_f'1_bufchan_d ;
  logic \lizzieLet48_3Lcall_f'1_bufchan_r ;
  assign \lizzieLet48_3Lcall_f'1_r  = ((! \lizzieLet48_3Lcall_f'1_bufchan_d [0]) || \lizzieLet48_3Lcall_f'1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \lizzieLet48_3Lcall_f'1_bufchan_d  <= 1'd0;
    else
      if (\lizzieLet48_3Lcall_f'1_r )
        \lizzieLet48_3Lcall_f'1_bufchan_d  <= \lizzieLet48_3Lcall_f'1_d ;
  Go_t \lizzieLet48_3Lcall_f'1_bufchan_buf ;
  assign \lizzieLet48_3Lcall_f'1_bufchan_r  = (! \lizzieLet48_3Lcall_f'1_bufchan_buf [0]);
  assign \lizzieLet48_3Lcall_f'1_1_argbuf_d  = (\lizzieLet48_3Lcall_f'1_bufchan_buf [0] ? \lizzieLet48_3Lcall_f'1_bufchan_buf  :
                                                \lizzieLet48_3Lcall_f'1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \lizzieLet48_3Lcall_f'1_bufchan_buf  <= 1'd0;
    else
      if ((\lizzieLet48_3Lcall_f'1_1_argbuf_r  && \lizzieLet48_3Lcall_f'1_bufchan_buf [0]))
        \lizzieLet48_3Lcall_f'1_bufchan_buf  <= 1'd0;
      else if (((! \lizzieLet48_3Lcall_f'1_1_argbuf_r ) && (! \lizzieLet48_3Lcall_f'1_bufchan_buf [0])))
        \lizzieLet48_3Lcall_f'1_bufchan_buf  <= \lizzieLet48_3Lcall_f'1_bufchan_d ;
  
  /* buf (Ty Go) : (lizzieLet48_3Lcall_f'2,Go) > (lizzieLet48_3Lcall_f'2_1_argbuf,Go) */
  Go_t \lizzieLet48_3Lcall_f'2_bufchan_d ;
  logic \lizzieLet48_3Lcall_f'2_bufchan_r ;
  assign \lizzieLet48_3Lcall_f'2_r  = ((! \lizzieLet48_3Lcall_f'2_bufchan_d [0]) || \lizzieLet48_3Lcall_f'2_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \lizzieLet48_3Lcall_f'2_bufchan_d  <= 1'd0;
    else
      if (\lizzieLet48_3Lcall_f'2_r )
        \lizzieLet48_3Lcall_f'2_bufchan_d  <= \lizzieLet48_3Lcall_f'2_d ;
  Go_t \lizzieLet48_3Lcall_f'2_bufchan_buf ;
  assign \lizzieLet48_3Lcall_f'2_bufchan_r  = (! \lizzieLet48_3Lcall_f'2_bufchan_buf [0]);
  assign \lizzieLet48_3Lcall_f'2_1_argbuf_d  = (\lizzieLet48_3Lcall_f'2_bufchan_buf [0] ? \lizzieLet48_3Lcall_f'2_bufchan_buf  :
                                                \lizzieLet48_3Lcall_f'2_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \lizzieLet48_3Lcall_f'2_bufchan_buf  <= 1'd0;
    else
      if ((\lizzieLet48_3Lcall_f'2_1_argbuf_r  && \lizzieLet48_3Lcall_f'2_bufchan_buf [0]))
        \lizzieLet48_3Lcall_f'2_bufchan_buf  <= 1'd0;
      else if (((! \lizzieLet48_3Lcall_f'2_1_argbuf_r ) && (! \lizzieLet48_3Lcall_f'2_bufchan_buf [0])))
        \lizzieLet48_3Lcall_f'2_bufchan_buf  <= \lizzieLet48_3Lcall_f'2_bufchan_d ;
  
  /* buf (Ty Go) : (lizzieLet48_3Lcall_f'3,Go) > (lizzieLet48_3Lcall_f'3_1_argbuf,Go) */
  Go_t \lizzieLet48_3Lcall_f'3_bufchan_d ;
  logic \lizzieLet48_3Lcall_f'3_bufchan_r ;
  assign \lizzieLet48_3Lcall_f'3_r  = ((! \lizzieLet48_3Lcall_f'3_bufchan_d [0]) || \lizzieLet48_3Lcall_f'3_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \lizzieLet48_3Lcall_f'3_bufchan_d  <= 1'd0;
    else
      if (\lizzieLet48_3Lcall_f'3_r )
        \lizzieLet48_3Lcall_f'3_bufchan_d  <= \lizzieLet48_3Lcall_f'3_d ;
  Go_t \lizzieLet48_3Lcall_f'3_bufchan_buf ;
  assign \lizzieLet48_3Lcall_f'3_bufchan_r  = (! \lizzieLet48_3Lcall_f'3_bufchan_buf [0]);
  assign \lizzieLet48_3Lcall_f'3_1_argbuf_d  = (\lizzieLet48_3Lcall_f'3_bufchan_buf [0] ? \lizzieLet48_3Lcall_f'3_bufchan_buf  :
                                                \lizzieLet48_3Lcall_f'3_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \lizzieLet48_3Lcall_f'3_bufchan_buf  <= 1'd0;
    else
      if ((\lizzieLet48_3Lcall_f'3_1_argbuf_r  && \lizzieLet48_3Lcall_f'3_bufchan_buf [0]))
        \lizzieLet48_3Lcall_f'3_bufchan_buf  <= 1'd0;
      else if (((! \lizzieLet48_3Lcall_f'3_1_argbuf_r ) && (! \lizzieLet48_3Lcall_f'3_bufchan_buf [0])))
        \lizzieLet48_3Lcall_f'3_bufchan_buf  <= \lizzieLet48_3Lcall_f'3_bufchan_d ;
  
  /* demux (Ty CTf',
       Ty Pointer_QTree_Bool) : (lizzieLet48_4,CTf') (srtarg_0_1_goMux_mux,Pointer_QTree_Bool) > [(lizzieLet48_4Lf'sbos,Pointer_QTree_Bool),
                                                                                                  (lizzieLet48_4Lcall_f'3,Pointer_QTree_Bool),
                                                                                                  (lizzieLet48_4Lcall_f'2,Pointer_QTree_Bool),
                                                                                                  (lizzieLet48_4Lcall_f'1,Pointer_QTree_Bool),
                                                                                                  (lizzieLet48_4Lcall_f'0,Pointer_QTree_Bool)] */
  logic [4:0] srtarg_0_1_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet48_4_d[0] && srtarg_0_1_goMux_mux_d[0]))
      unique case (lizzieLet48_4_d[3:1])
        3'd0: srtarg_0_1_goMux_mux_onehotd = 5'd1;
        3'd1: srtarg_0_1_goMux_mux_onehotd = 5'd2;
        3'd2: srtarg_0_1_goMux_mux_onehotd = 5'd4;
        3'd3: srtarg_0_1_goMux_mux_onehotd = 5'd8;
        3'd4: srtarg_0_1_goMux_mux_onehotd = 5'd16;
        default: srtarg_0_1_goMux_mux_onehotd = 5'd0;
      endcase
    else srtarg_0_1_goMux_mux_onehotd = 5'd0;
  assign \lizzieLet48_4Lf'sbos_d  = {srtarg_0_1_goMux_mux_d[16:1],
                                     srtarg_0_1_goMux_mux_onehotd[0]};
  assign \lizzieLet48_4Lcall_f'3_d  = {srtarg_0_1_goMux_mux_d[16:1],
                                       srtarg_0_1_goMux_mux_onehotd[1]};
  assign \lizzieLet48_4Lcall_f'2_d  = {srtarg_0_1_goMux_mux_d[16:1],
                                       srtarg_0_1_goMux_mux_onehotd[2]};
  assign \lizzieLet48_4Lcall_f'1_d  = {srtarg_0_1_goMux_mux_d[16:1],
                                       srtarg_0_1_goMux_mux_onehotd[3]};
  assign \lizzieLet48_4Lcall_f'0_d  = {srtarg_0_1_goMux_mux_d[16:1],
                                       srtarg_0_1_goMux_mux_onehotd[4]};
  assign srtarg_0_1_goMux_mux_r = (| (srtarg_0_1_goMux_mux_onehotd & {\lizzieLet48_4Lcall_f'0_r ,
                                                                      \lizzieLet48_4Lcall_f'1_r ,
                                                                      \lizzieLet48_4Lcall_f'2_r ,
                                                                      \lizzieLet48_4Lcall_f'3_r ,
                                                                      \lizzieLet48_4Lf'sbos_r }));
  assign lizzieLet48_4_r = srtarg_0_1_goMux_mux_r;
  
  /* dcon (Ty QTree_Bool,
      Dcon QNode_Bool) : [(lizzieLet48_4Lcall_f'0,Pointer_QTree_Bool),
                          (es_1_1_destruct,Pointer_QTree_Bool),
                          (es_2_2_destruct,Pointer_QTree_Bool),
                          (es_3_3_destruct,Pointer_QTree_Bool)] > (lizzieLet48_4Lcall_f'0_1es_1_1_1es_2_2_1es_3_3_1QNode_Bool,QTree_Bool) */
  assign \lizzieLet48_4Lcall_f'0_1es_1_1_1es_2_2_1es_3_3_1QNode_Bool_d  = QNode_Bool_dc((& {\lizzieLet48_4Lcall_f'0_d [0],
                                                                                            es_1_1_destruct_d[0],
                                                                                            es_2_2_destruct_d[0],
                                                                                            es_3_3_destruct_d[0]}), \lizzieLet48_4Lcall_f'0_d , es_1_1_destruct_d, es_2_2_destruct_d, es_3_3_destruct_d);
  assign {\lizzieLet48_4Lcall_f'0_r ,
          es_1_1_destruct_r,
          es_2_2_destruct_r,
          es_3_3_destruct_r} = {4 {(\lizzieLet48_4Lcall_f'0_1es_1_1_1es_2_2_1es_3_3_1QNode_Bool_r  && \lizzieLet48_4Lcall_f'0_1es_1_1_1es_2_2_1es_3_3_1QNode_Bool_d [0])}};
  
  /* buf (Ty QTree_Bool) : (lizzieLet48_4Lcall_f'0_1es_1_1_1es_2_2_1es_3_3_1QNode_Bool,QTree_Bool) > (lizzieLet52_1_argbuf,QTree_Bool) */
  QTree_Bool_t \lizzieLet48_4Lcall_f'0_1es_1_1_1es_2_2_1es_3_3_1QNode_Bool_bufchan_d ;
  logic \lizzieLet48_4Lcall_f'0_1es_1_1_1es_2_2_1es_3_3_1QNode_Bool_bufchan_r ;
  assign \lizzieLet48_4Lcall_f'0_1es_1_1_1es_2_2_1es_3_3_1QNode_Bool_r  = ((! \lizzieLet48_4Lcall_f'0_1es_1_1_1es_2_2_1es_3_3_1QNode_Bool_bufchan_d [0]) || \lizzieLet48_4Lcall_f'0_1es_1_1_1es_2_2_1es_3_3_1QNode_Bool_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet48_4Lcall_f'0_1es_1_1_1es_2_2_1es_3_3_1QNode_Bool_bufchan_d  <= {66'd0,
                                                                                 1'd0};
    else
      if (\lizzieLet48_4Lcall_f'0_1es_1_1_1es_2_2_1es_3_3_1QNode_Bool_r )
        \lizzieLet48_4Lcall_f'0_1es_1_1_1es_2_2_1es_3_3_1QNode_Bool_bufchan_d  <= \lizzieLet48_4Lcall_f'0_1es_1_1_1es_2_2_1es_3_3_1QNode_Bool_d ;
  QTree_Bool_t \lizzieLet48_4Lcall_f'0_1es_1_1_1es_2_2_1es_3_3_1QNode_Bool_bufchan_buf ;
  assign \lizzieLet48_4Lcall_f'0_1es_1_1_1es_2_2_1es_3_3_1QNode_Bool_bufchan_r  = (! \lizzieLet48_4Lcall_f'0_1es_1_1_1es_2_2_1es_3_3_1QNode_Bool_bufchan_buf [0]);
  assign lizzieLet52_1_argbuf_d = (\lizzieLet48_4Lcall_f'0_1es_1_1_1es_2_2_1es_3_3_1QNode_Bool_bufchan_buf [0] ? \lizzieLet48_4Lcall_f'0_1es_1_1_1es_2_2_1es_3_3_1QNode_Bool_bufchan_buf  :
                                   \lizzieLet48_4Lcall_f'0_1es_1_1_1es_2_2_1es_3_3_1QNode_Bool_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet48_4Lcall_f'0_1es_1_1_1es_2_2_1es_3_3_1QNode_Bool_bufchan_buf  <= {66'd0,
                                                                                   1'd0};
    else
      if ((lizzieLet52_1_argbuf_r && \lizzieLet48_4Lcall_f'0_1es_1_1_1es_2_2_1es_3_3_1QNode_Bool_bufchan_buf [0]))
        \lizzieLet48_4Lcall_f'0_1es_1_1_1es_2_2_1es_3_3_1QNode_Bool_bufchan_buf  <= {66'd0,
                                                                                     1'd0};
      else if (((! lizzieLet52_1_argbuf_r) && (! \lizzieLet48_4Lcall_f'0_1es_1_1_1es_2_2_1es_3_3_1QNode_Bool_bufchan_buf [0])))
        \lizzieLet48_4Lcall_f'0_1es_1_1_1es_2_2_1es_3_3_1QNode_Bool_bufchan_buf  <= \lizzieLet48_4Lcall_f'0_1es_1_1_1es_2_2_1es_3_3_1QNode_Bool_bufchan_d ;
  
  /* dcon (Ty CTf',
      Dcon Lcall_f'0) : [(lizzieLet48_4Lcall_f'1,Pointer_QTree_Bool),
                         (es_2_1_destruct,Pointer_QTree_Bool),
                         (es_3_2_destruct,Pointer_QTree_Bool),
                         (sc_0_9_destruct,Pointer_CTf')] > (lizzieLet48_4Lcall_f'1_1es_2_1_1es_3_2_1sc_0_9_1Lcall_f'0,CTf') */
  assign \lizzieLet48_4Lcall_f'1_1es_2_1_1es_3_2_1sc_0_9_1Lcall_f'0_d  = \Lcall_f'0_dc ((& {\lizzieLet48_4Lcall_f'1_d [0],
                                                                                            es_2_1_destruct_d[0],
                                                                                            es_3_2_destruct_d[0],
                                                                                            sc_0_9_destruct_d[0]}), \lizzieLet48_4Lcall_f'1_d , es_2_1_destruct_d, es_3_2_destruct_d, sc_0_9_destruct_d);
  assign {\lizzieLet48_4Lcall_f'1_r ,
          es_2_1_destruct_r,
          es_3_2_destruct_r,
          sc_0_9_destruct_r} = {4 {(\lizzieLet48_4Lcall_f'1_1es_2_1_1es_3_2_1sc_0_9_1Lcall_f'0_r  && \lizzieLet48_4Lcall_f'1_1es_2_1_1es_3_2_1sc_0_9_1Lcall_f'0_d [0])}};
  
  /* buf (Ty CTf') : (lizzieLet48_4Lcall_f'1_1es_2_1_1es_3_2_1sc_0_9_1Lcall_f'0,CTf') > (lizzieLet51_1_argbuf,CTf') */
  \CTf'_t  \lizzieLet48_4Lcall_f'1_1es_2_1_1es_3_2_1sc_0_9_1Lcall_f'0_bufchan_d ;
  logic \lizzieLet48_4Lcall_f'1_1es_2_1_1es_3_2_1sc_0_9_1Lcall_f'0_bufchan_r ;
  assign \lizzieLet48_4Lcall_f'1_1es_2_1_1es_3_2_1sc_0_9_1Lcall_f'0_r  = ((! \lizzieLet48_4Lcall_f'1_1es_2_1_1es_3_2_1sc_0_9_1Lcall_f'0_bufchan_d [0]) || \lizzieLet48_4Lcall_f'1_1es_2_1_1es_3_2_1sc_0_9_1Lcall_f'0_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet48_4Lcall_f'1_1es_2_1_1es_3_2_1sc_0_9_1Lcall_f'0_bufchan_d  <= {115'd0,
                                                                                1'd0};
    else
      if (\lizzieLet48_4Lcall_f'1_1es_2_1_1es_3_2_1sc_0_9_1Lcall_f'0_r )
        \lizzieLet48_4Lcall_f'1_1es_2_1_1es_3_2_1sc_0_9_1Lcall_f'0_bufchan_d  <= \lizzieLet48_4Lcall_f'1_1es_2_1_1es_3_2_1sc_0_9_1Lcall_f'0_d ;
  \CTf'_t  \lizzieLet48_4Lcall_f'1_1es_2_1_1es_3_2_1sc_0_9_1Lcall_f'0_bufchan_buf ;
  assign \lizzieLet48_4Lcall_f'1_1es_2_1_1es_3_2_1sc_0_9_1Lcall_f'0_bufchan_r  = (! \lizzieLet48_4Lcall_f'1_1es_2_1_1es_3_2_1sc_0_9_1Lcall_f'0_bufchan_buf [0]);
  assign lizzieLet51_1_argbuf_d = (\lizzieLet48_4Lcall_f'1_1es_2_1_1es_3_2_1sc_0_9_1Lcall_f'0_bufchan_buf [0] ? \lizzieLet48_4Lcall_f'1_1es_2_1_1es_3_2_1sc_0_9_1Lcall_f'0_bufchan_buf  :
                                   \lizzieLet48_4Lcall_f'1_1es_2_1_1es_3_2_1sc_0_9_1Lcall_f'0_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet48_4Lcall_f'1_1es_2_1_1es_3_2_1sc_0_9_1Lcall_f'0_bufchan_buf  <= {115'd0,
                                                                                  1'd0};
    else
      if ((lizzieLet51_1_argbuf_r && \lizzieLet48_4Lcall_f'1_1es_2_1_1es_3_2_1sc_0_9_1Lcall_f'0_bufchan_buf [0]))
        \lizzieLet48_4Lcall_f'1_1es_2_1_1es_3_2_1sc_0_9_1Lcall_f'0_bufchan_buf  <= {115'd0,
                                                                                    1'd0};
      else if (((! lizzieLet51_1_argbuf_r) && (! \lizzieLet48_4Lcall_f'1_1es_2_1_1es_3_2_1sc_0_9_1Lcall_f'0_bufchan_buf [0])))
        \lizzieLet48_4Lcall_f'1_1es_2_1_1es_3_2_1sc_0_9_1Lcall_f'0_bufchan_buf  <= \lizzieLet48_4Lcall_f'1_1es_2_1_1es_3_2_1sc_0_9_1Lcall_f'0_bufchan_d ;
  
  /* dcon (Ty CTf',
      Dcon Lcall_f'1) : [(lizzieLet48_4Lcall_f'2,Pointer_QTree_Bool),
                         (es_3_1_destruct,Pointer_QTree_Bool),
                         (sc_0_8_destruct,Pointer_CTf'),
                         (q1a8P_2_destruct,Pointer_QTree_Bool),
                         (t1a8U_2_destruct,Pointer_QTree_Bool)] > (lizzieLet48_4Lcall_f'2_1es_3_1_1sc_0_8_1q1a8P_2_1t1a8U_2_1Lcall_f'1,CTf') */
  assign \lizzieLet48_4Lcall_f'2_1es_3_1_1sc_0_8_1q1a8P_2_1t1a8U_2_1Lcall_f'1_d  = \Lcall_f'1_dc ((& {\lizzieLet48_4Lcall_f'2_d [0],
                                                                                                      es_3_1_destruct_d[0],
                                                                                                      sc_0_8_destruct_d[0],
                                                                                                      q1a8P_2_destruct_d[0],
                                                                                                      t1a8U_2_destruct_d[0]}), \lizzieLet48_4Lcall_f'2_d , es_3_1_destruct_d, sc_0_8_destruct_d, q1a8P_2_destruct_d, t1a8U_2_destruct_d);
  assign {\lizzieLet48_4Lcall_f'2_r ,
          es_3_1_destruct_r,
          sc_0_8_destruct_r,
          q1a8P_2_destruct_r,
          t1a8U_2_destruct_r} = {5 {(\lizzieLet48_4Lcall_f'2_1es_3_1_1sc_0_8_1q1a8P_2_1t1a8U_2_1Lcall_f'1_r  && \lizzieLet48_4Lcall_f'2_1es_3_1_1sc_0_8_1q1a8P_2_1t1a8U_2_1Lcall_f'1_d [0])}};
  
  /* buf (Ty CTf') : (lizzieLet48_4Lcall_f'2_1es_3_1_1sc_0_8_1q1a8P_2_1t1a8U_2_1Lcall_f'1,CTf') > (lizzieLet50_1_argbuf,CTf') */
  \CTf'_t  \lizzieLet48_4Lcall_f'2_1es_3_1_1sc_0_8_1q1a8P_2_1t1a8U_2_1Lcall_f'1_bufchan_d ;
  logic \lizzieLet48_4Lcall_f'2_1es_3_1_1sc_0_8_1q1a8P_2_1t1a8U_2_1Lcall_f'1_bufchan_r ;
  assign \lizzieLet48_4Lcall_f'2_1es_3_1_1sc_0_8_1q1a8P_2_1t1a8U_2_1Lcall_f'1_r  = ((! \lizzieLet48_4Lcall_f'2_1es_3_1_1sc_0_8_1q1a8P_2_1t1a8U_2_1Lcall_f'1_bufchan_d [0]) || \lizzieLet48_4Lcall_f'2_1es_3_1_1sc_0_8_1q1a8P_2_1t1a8U_2_1Lcall_f'1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet48_4Lcall_f'2_1es_3_1_1sc_0_8_1q1a8P_2_1t1a8U_2_1Lcall_f'1_bufchan_d  <= {115'd0,
                                                                                          1'd0};
    else
      if (\lizzieLet48_4Lcall_f'2_1es_3_1_1sc_0_8_1q1a8P_2_1t1a8U_2_1Lcall_f'1_r )
        \lizzieLet48_4Lcall_f'2_1es_3_1_1sc_0_8_1q1a8P_2_1t1a8U_2_1Lcall_f'1_bufchan_d  <= \lizzieLet48_4Lcall_f'2_1es_3_1_1sc_0_8_1q1a8P_2_1t1a8U_2_1Lcall_f'1_d ;
  \CTf'_t  \lizzieLet48_4Lcall_f'2_1es_3_1_1sc_0_8_1q1a8P_2_1t1a8U_2_1Lcall_f'1_bufchan_buf ;
  assign \lizzieLet48_4Lcall_f'2_1es_3_1_1sc_0_8_1q1a8P_2_1t1a8U_2_1Lcall_f'1_bufchan_r  = (! \lizzieLet48_4Lcall_f'2_1es_3_1_1sc_0_8_1q1a8P_2_1t1a8U_2_1Lcall_f'1_bufchan_buf [0]);
  assign lizzieLet50_1_argbuf_d = (\lizzieLet48_4Lcall_f'2_1es_3_1_1sc_0_8_1q1a8P_2_1t1a8U_2_1Lcall_f'1_bufchan_buf [0] ? \lizzieLet48_4Lcall_f'2_1es_3_1_1sc_0_8_1q1a8P_2_1t1a8U_2_1Lcall_f'1_bufchan_buf  :
                                   \lizzieLet48_4Lcall_f'2_1es_3_1_1sc_0_8_1q1a8P_2_1t1a8U_2_1Lcall_f'1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet48_4Lcall_f'2_1es_3_1_1sc_0_8_1q1a8P_2_1t1a8U_2_1Lcall_f'1_bufchan_buf  <= {115'd0,
                                                                                            1'd0};
    else
      if ((lizzieLet50_1_argbuf_r && \lizzieLet48_4Lcall_f'2_1es_3_1_1sc_0_8_1q1a8P_2_1t1a8U_2_1Lcall_f'1_bufchan_buf [0]))
        \lizzieLet48_4Lcall_f'2_1es_3_1_1sc_0_8_1q1a8P_2_1t1a8U_2_1Lcall_f'1_bufchan_buf  <= {115'd0,
                                                                                              1'd0};
      else if (((! lizzieLet50_1_argbuf_r) && (! \lizzieLet48_4Lcall_f'2_1es_3_1_1sc_0_8_1q1a8P_2_1t1a8U_2_1Lcall_f'1_bufchan_buf [0])))
        \lizzieLet48_4Lcall_f'2_1es_3_1_1sc_0_8_1q1a8P_2_1t1a8U_2_1Lcall_f'1_bufchan_buf  <= \lizzieLet48_4Lcall_f'2_1es_3_1_1sc_0_8_1q1a8P_2_1t1a8U_2_1Lcall_f'1_bufchan_d ;
  
  /* dcon (Ty CTf',
      Dcon Lcall_f'2) : [(lizzieLet48_4Lcall_f'3,Pointer_QTree_Bool),
                         (sc_0_7_destruct,Pointer_CTf'),
                         (q1a8P_1_destruct,Pointer_QTree_Bool),
                         (t1a8U_1_destruct,Pointer_QTree_Bool),
                         (q2a8Q_1_destruct,Pointer_QTree_Bool),
                         (t2a8V_1_destruct,Pointer_QTree_Bool)] > (lizzieLet48_4Lcall_f'3_1sc_0_7_1q1a8P_1_1t1a8U_1_1q2a8Q_1_1t2a8V_1_1Lcall_f'2,CTf') */
  assign \lizzieLet48_4Lcall_f'3_1sc_0_7_1q1a8P_1_1t1a8U_1_1q2a8Q_1_1t2a8V_1_1Lcall_f'2_d  = \Lcall_f'2_dc ((& {\lizzieLet48_4Lcall_f'3_d [0],
                                                                                                                sc_0_7_destruct_d[0],
                                                                                                                q1a8P_1_destruct_d[0],
                                                                                                                t1a8U_1_destruct_d[0],
                                                                                                                q2a8Q_1_destruct_d[0],
                                                                                                                t2a8V_1_destruct_d[0]}), \lizzieLet48_4Lcall_f'3_d , sc_0_7_destruct_d, q1a8P_1_destruct_d, t1a8U_1_destruct_d, q2a8Q_1_destruct_d, t2a8V_1_destruct_d);
  assign {\lizzieLet48_4Lcall_f'3_r ,
          sc_0_7_destruct_r,
          q1a8P_1_destruct_r,
          t1a8U_1_destruct_r,
          q2a8Q_1_destruct_r,
          t2a8V_1_destruct_r} = {6 {(\lizzieLet48_4Lcall_f'3_1sc_0_7_1q1a8P_1_1t1a8U_1_1q2a8Q_1_1t2a8V_1_1Lcall_f'2_r  && \lizzieLet48_4Lcall_f'3_1sc_0_7_1q1a8P_1_1t1a8U_1_1q2a8Q_1_1t2a8V_1_1Lcall_f'2_d [0])}};
  
  /* buf (Ty CTf') : (lizzieLet48_4Lcall_f'3_1sc_0_7_1q1a8P_1_1t1a8U_1_1q2a8Q_1_1t2a8V_1_1Lcall_f'2,CTf') > (lizzieLet49_1_argbuf,CTf') */
  \CTf'_t  \lizzieLet48_4Lcall_f'3_1sc_0_7_1q1a8P_1_1t1a8U_1_1q2a8Q_1_1t2a8V_1_1Lcall_f'2_bufchan_d ;
  logic \lizzieLet48_4Lcall_f'3_1sc_0_7_1q1a8P_1_1t1a8U_1_1q2a8Q_1_1t2a8V_1_1Lcall_f'2_bufchan_r ;
  assign \lizzieLet48_4Lcall_f'3_1sc_0_7_1q1a8P_1_1t1a8U_1_1q2a8Q_1_1t2a8V_1_1Lcall_f'2_r  = ((! \lizzieLet48_4Lcall_f'3_1sc_0_7_1q1a8P_1_1t1a8U_1_1q2a8Q_1_1t2a8V_1_1Lcall_f'2_bufchan_d [0]) || \lizzieLet48_4Lcall_f'3_1sc_0_7_1q1a8P_1_1t1a8U_1_1q2a8Q_1_1t2a8V_1_1Lcall_f'2_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet48_4Lcall_f'3_1sc_0_7_1q1a8P_1_1t1a8U_1_1q2a8Q_1_1t2a8V_1_1Lcall_f'2_bufchan_d  <= {115'd0,
                                                                                                    1'd0};
    else
      if (\lizzieLet48_4Lcall_f'3_1sc_0_7_1q1a8P_1_1t1a8U_1_1q2a8Q_1_1t2a8V_1_1Lcall_f'2_r )
        \lizzieLet48_4Lcall_f'3_1sc_0_7_1q1a8P_1_1t1a8U_1_1q2a8Q_1_1t2a8V_1_1Lcall_f'2_bufchan_d  <= \lizzieLet48_4Lcall_f'3_1sc_0_7_1q1a8P_1_1t1a8U_1_1q2a8Q_1_1t2a8V_1_1Lcall_f'2_d ;
  \CTf'_t  \lizzieLet48_4Lcall_f'3_1sc_0_7_1q1a8P_1_1t1a8U_1_1q2a8Q_1_1t2a8V_1_1Lcall_f'2_bufchan_buf ;
  assign \lizzieLet48_4Lcall_f'3_1sc_0_7_1q1a8P_1_1t1a8U_1_1q2a8Q_1_1t2a8V_1_1Lcall_f'2_bufchan_r  = (! \lizzieLet48_4Lcall_f'3_1sc_0_7_1q1a8P_1_1t1a8U_1_1q2a8Q_1_1t2a8V_1_1Lcall_f'2_bufchan_buf [0]);
  assign lizzieLet49_1_argbuf_d = (\lizzieLet48_4Lcall_f'3_1sc_0_7_1q1a8P_1_1t1a8U_1_1q2a8Q_1_1t2a8V_1_1Lcall_f'2_bufchan_buf [0] ? \lizzieLet48_4Lcall_f'3_1sc_0_7_1q1a8P_1_1t1a8U_1_1q2a8Q_1_1t2a8V_1_1Lcall_f'2_bufchan_buf  :
                                   \lizzieLet48_4Lcall_f'3_1sc_0_7_1q1a8P_1_1t1a8U_1_1q2a8Q_1_1t2a8V_1_1Lcall_f'2_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet48_4Lcall_f'3_1sc_0_7_1q1a8P_1_1t1a8U_1_1q2a8Q_1_1t2a8V_1_1Lcall_f'2_bufchan_buf  <= {115'd0,
                                                                                                      1'd0};
    else
      if ((lizzieLet49_1_argbuf_r && \lizzieLet48_4Lcall_f'3_1sc_0_7_1q1a8P_1_1t1a8U_1_1q2a8Q_1_1t2a8V_1_1Lcall_f'2_bufchan_buf [0]))
        \lizzieLet48_4Lcall_f'3_1sc_0_7_1q1a8P_1_1t1a8U_1_1q2a8Q_1_1t2a8V_1_1Lcall_f'2_bufchan_buf  <= {115'd0,
                                                                                                        1'd0};
      else if (((! lizzieLet49_1_argbuf_r) && (! \lizzieLet48_4Lcall_f'3_1sc_0_7_1q1a8P_1_1t1a8U_1_1q2a8Q_1_1t2a8V_1_1Lcall_f'2_bufchan_buf [0])))
        \lizzieLet48_4Lcall_f'3_1sc_0_7_1q1a8P_1_1t1a8U_1_1q2a8Q_1_1t2a8V_1_1Lcall_f'2_bufchan_buf  <= \lizzieLet48_4Lcall_f'3_1sc_0_7_1q1a8P_1_1t1a8U_1_1q2a8Q_1_1t2a8V_1_1Lcall_f'2_bufchan_d ;
  
  /* fork (Ty Pointer_QTree_Bool) : (lizzieLet48_4Lf'sbos,Pointer_QTree_Bool) > [(lizzieLet48_4Lf'sbos_1_merge_merge_fork_1,Pointer_QTree_Bool),
                                                                            (lizzieLet48_4Lf'sbos_1_merge_merge_fork_2,Pointer_QTree_Bool)] */
  logic [1:0] \lizzieLet48_4Lf'sbos_emitted ;
  logic [1:0] \lizzieLet48_4Lf'sbos_done ;
  assign \lizzieLet48_4Lf'sbos_1_merge_merge_fork_1_d  = {\lizzieLet48_4Lf'sbos_d [16:1],
                                                          (\lizzieLet48_4Lf'sbos_d [0] && (! \lizzieLet48_4Lf'sbos_emitted [0]))};
  assign \lizzieLet48_4Lf'sbos_1_merge_merge_fork_2_d  = {\lizzieLet48_4Lf'sbos_d [16:1],
                                                          (\lizzieLet48_4Lf'sbos_d [0] && (! \lizzieLet48_4Lf'sbos_emitted [1]))};
  assign \lizzieLet48_4Lf'sbos_done  = (\lizzieLet48_4Lf'sbos_emitted  | ({\lizzieLet48_4Lf'sbos_1_merge_merge_fork_2_d [0],
                                                                           \lizzieLet48_4Lf'sbos_1_merge_merge_fork_1_d [0]} & {\lizzieLet48_4Lf'sbos_1_merge_merge_fork_2_r ,
                                                                                                                                \lizzieLet48_4Lf'sbos_1_merge_merge_fork_1_r }));
  assign \lizzieLet48_4Lf'sbos_r  = (& \lizzieLet48_4Lf'sbos_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \lizzieLet48_4Lf'sbos_emitted  <= 2'd0;
    else
      \lizzieLet48_4Lf'sbos_emitted  <= (\lizzieLet48_4Lf'sbos_r  ? 2'd0 :
                                         \lizzieLet48_4Lf'sbos_done );
  
  /* togo (Ty Pointer_QTree_Bool) : (lizzieLet48_4Lf'sbos_1_merge_merge_fork_1,Pointer_QTree_Bool) > (call_f'_goConst,Go) */
  assign \call_f'_goConst_d  = \lizzieLet48_4Lf'sbos_1_merge_merge_fork_1_d [0];
  assign \lizzieLet48_4Lf'sbos_1_merge_merge_fork_1_r  = \call_f'_goConst_r ;
  
  /* buf (Ty Pointer_QTree_Bool) : (lizzieLet48_4Lf'sbos_1_merge_merge_fork_2,Pointer_QTree_Bool) > (f'_resbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t \lizzieLet48_4Lf'sbos_1_merge_merge_fork_2_bufchan_d ;
  logic \lizzieLet48_4Lf'sbos_1_merge_merge_fork_2_bufchan_r ;
  assign \lizzieLet48_4Lf'sbos_1_merge_merge_fork_2_r  = ((! \lizzieLet48_4Lf'sbos_1_merge_merge_fork_2_bufchan_d [0]) || \lizzieLet48_4Lf'sbos_1_merge_merge_fork_2_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet48_4Lf'sbos_1_merge_merge_fork_2_bufchan_d  <= {16'd0,
                                                                1'd0};
    else
      if (\lizzieLet48_4Lf'sbos_1_merge_merge_fork_2_r )
        \lizzieLet48_4Lf'sbos_1_merge_merge_fork_2_bufchan_d  <= \lizzieLet48_4Lf'sbos_1_merge_merge_fork_2_d ;
  Pointer_QTree_Bool_t \lizzieLet48_4Lf'sbos_1_merge_merge_fork_2_bufchan_buf ;
  assign \lizzieLet48_4Lf'sbos_1_merge_merge_fork_2_bufchan_r  = (! \lizzieLet48_4Lf'sbos_1_merge_merge_fork_2_bufchan_buf [0]);
  assign \f'_resbuf_d  = (\lizzieLet48_4Lf'sbos_1_merge_merge_fork_2_bufchan_buf [0] ? \lizzieLet48_4Lf'sbos_1_merge_merge_fork_2_bufchan_buf  :
                          \lizzieLet48_4Lf'sbos_1_merge_merge_fork_2_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet48_4Lf'sbos_1_merge_merge_fork_2_bufchan_buf  <= {16'd0,
                                                                  1'd0};
    else
      if ((\f'_resbuf_r  && \lizzieLet48_4Lf'sbos_1_merge_merge_fork_2_bufchan_buf [0]))
        \lizzieLet48_4Lf'sbos_1_merge_merge_fork_2_bufchan_buf  <= {16'd0,
                                                                    1'd0};
      else if (((! \f'_resbuf_r ) && (! \lizzieLet48_4Lf'sbos_1_merge_merge_fork_2_bufchan_buf [0])))
        \lizzieLet48_4Lf'sbos_1_merge_merge_fork_2_bufchan_buf  <= \lizzieLet48_4Lf'sbos_1_merge_merge_fork_2_bufchan_d ;
  
  /* destruct (Ty CTf'''''''''_f'''''''''_Bool,
          Dcon Lcall_f'''''''''_f'''''''''_Bool0) : (lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool0,CTf'''''''''_f'''''''''_Bool) > [(es_1_2_destruct,Pointer_QTree_Bool),
                                                                                                                                     (es_2_4_destruct,Pointer_QTree_Bool),
                                                                                                                                     (es_3_6_destruct,Pointer_QTree_Bool),
                                                                                                                                     (sc_0_14_destruct,Pointer_CTf'''''''''_f'''''''''_Bool)] */
  logic [3:0] \lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool0_emitted ;
  logic [3:0] \lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool0_done ;
  assign es_1_2_destruct_d = {\lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool0_d [19:4],
                              (\lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool0_d [0] && (! \lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool0_emitted [0]))};
  assign es_2_4_destruct_d = {\lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool0_d [35:20],
                              (\lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool0_d [0] && (! \lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool0_emitted [1]))};
  assign es_3_6_destruct_d = {\lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool0_d [51:36],
                              (\lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool0_d [0] && (! \lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool0_emitted [2]))};
  assign sc_0_14_destruct_d = {\lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool0_d [67:52],
                               (\lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool0_d [0] && (! \lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool0_emitted [3]))};
  assign \lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool0_done  = (\lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool0_emitted  | ({sc_0_14_destruct_d[0],
                                                                                                                               es_3_6_destruct_d[0],
                                                                                                                               es_2_4_destruct_d[0],
                                                                                                                               es_1_2_destruct_d[0]} & {sc_0_14_destruct_r,
                                                                                                                                                        es_3_6_destruct_r,
                                                                                                                                                        es_2_4_destruct_r,
                                                                                                                                                        es_1_2_destruct_r}));
  assign \lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool0_r  = (& \lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool0_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool0_emitted  <= 4'd0;
    else
      \lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool0_emitted  <= (\lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool0_r  ? 4'd0 :
                                                                   \lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool0_done );
  
  /* destruct (Ty CTf'''''''''_f'''''''''_Bool,
          Dcon Lcall_f'''''''''_f'''''''''_Bool1) : (lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool1,CTf'''''''''_f'''''''''_Bool) > [(es_2_3_destruct,Pointer_QTree_Bool),
                                                                                                                                     (es_3_5_destruct,Pointer_QTree_Bool),
                                                                                                                                     (sc_0_13_destruct,Pointer_CTf'''''''''_f'''''''''_Bool),
                                                                                                                                     (q1a8y_3_destruct,Pointer_MaskQTree),
                                                                                                                                     (t1a8D_3_destruct,Pointer_QTree_Bool)] */
  logic [4:0] \lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool1_emitted ;
  logic [4:0] \lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool1_done ;
  assign es_2_3_destruct_d = {\lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool1_d [19:4],
                              (\lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool1_d [0] && (! \lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool1_emitted [0]))};
  assign es_3_5_destruct_d = {\lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool1_d [35:20],
                              (\lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool1_d [0] && (! \lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool1_emitted [1]))};
  assign sc_0_13_destruct_d = {\lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool1_d [51:36],
                               (\lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool1_d [0] && (! \lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool1_emitted [2]))};
  assign q1a8y_3_destruct_d = {\lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool1_d [67:52],
                               (\lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool1_d [0] && (! \lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool1_emitted [3]))};
  assign t1a8D_3_destruct_d = {\lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool1_d [83:68],
                               (\lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool1_d [0] && (! \lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool1_emitted [4]))};
  assign \lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool1_done  = (\lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool1_emitted  | ({t1a8D_3_destruct_d[0],
                                                                                                                               q1a8y_3_destruct_d[0],
                                                                                                                               sc_0_13_destruct_d[0],
                                                                                                                               es_3_5_destruct_d[0],
                                                                                                                               es_2_3_destruct_d[0]} & {t1a8D_3_destruct_r,
                                                                                                                                                        q1a8y_3_destruct_r,
                                                                                                                                                        sc_0_13_destruct_r,
                                                                                                                                                        es_3_5_destruct_r,
                                                                                                                                                        es_2_3_destruct_r}));
  assign \lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool1_r  = (& \lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool1_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool1_emitted  <= 5'd0;
    else
      \lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool1_emitted  <= (\lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool1_r  ? 5'd0 :
                                                                   \lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool1_done );
  
  /* destruct (Ty CTf'''''''''_f'''''''''_Bool,
          Dcon Lcall_f'''''''''_f'''''''''_Bool2) : (lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool2,CTf'''''''''_f'''''''''_Bool) > [(es_3_4_destruct,Pointer_QTree_Bool),
                                                                                                                                     (sc_0_12_destruct,Pointer_CTf'''''''''_f'''''''''_Bool),
                                                                                                                                     (q1a8y_2_destruct,Pointer_MaskQTree),
                                                                                                                                     (t1a8D_2_destruct,Pointer_QTree_Bool),
                                                                                                                                     (q2a8z_2_destruct,Pointer_MaskQTree),
                                                                                                                                     (t2a8E_2_destruct,Pointer_QTree_Bool)] */
  logic [5:0] \lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool2_emitted ;
  logic [5:0] \lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool2_done ;
  assign es_3_4_destruct_d = {\lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool2_d [19:4],
                              (\lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool2_d [0] && (! \lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool2_emitted [0]))};
  assign sc_0_12_destruct_d = {\lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool2_d [35:20],
                               (\lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool2_d [0] && (! \lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool2_emitted [1]))};
  assign q1a8y_2_destruct_d = {\lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool2_d [51:36],
                               (\lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool2_d [0] && (! \lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool2_emitted [2]))};
  assign t1a8D_2_destruct_d = {\lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool2_d [67:52],
                               (\lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool2_d [0] && (! \lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool2_emitted [3]))};
  assign q2a8z_2_destruct_d = {\lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool2_d [83:68],
                               (\lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool2_d [0] && (! \lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool2_emitted [4]))};
  assign t2a8E_2_destruct_d = {\lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool2_d [99:84],
                               (\lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool2_d [0] && (! \lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool2_emitted [5]))};
  assign \lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool2_done  = (\lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool2_emitted  | ({t2a8E_2_destruct_d[0],
                                                                                                                               q2a8z_2_destruct_d[0],
                                                                                                                               t1a8D_2_destruct_d[0],
                                                                                                                               q1a8y_2_destruct_d[0],
                                                                                                                               sc_0_12_destruct_d[0],
                                                                                                                               es_3_4_destruct_d[0]} & {t2a8E_2_destruct_r,
                                                                                                                                                        q2a8z_2_destruct_r,
                                                                                                                                                        t1a8D_2_destruct_r,
                                                                                                                                                        q1a8y_2_destruct_r,
                                                                                                                                                        sc_0_12_destruct_r,
                                                                                                                                                        es_3_4_destruct_r}));
  assign \lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool2_r  = (& \lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool2_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool2_emitted  <= 6'd0;
    else
      \lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool2_emitted  <= (\lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool2_r  ? 6'd0 :
                                                                   \lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool2_done );
  
  /* destruct (Ty CTf'''''''''_f'''''''''_Bool,
          Dcon Lcall_f'''''''''_f'''''''''_Bool3) : (lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool3,CTf'''''''''_f'''''''''_Bool) > [(sc_0_11_destruct,Pointer_CTf'''''''''_f'''''''''_Bool),
                                                                                                                                     (q1a8y_1_destruct,Pointer_MaskQTree),
                                                                                                                                     (t1a8D_1_destruct,Pointer_QTree_Bool),
                                                                                                                                     (q2a8z_1_destruct,Pointer_MaskQTree),
                                                                                                                                     (t2a8E_1_destruct,Pointer_QTree_Bool),
                                                                                                                                     (q3a8A_1_destruct,Pointer_MaskQTree),
                                                                                                                                     (t3a8F_1_destruct,Pointer_QTree_Bool)] */
  logic [6:0] \lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool3_emitted ;
  logic [6:0] \lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool3_done ;
  assign sc_0_11_destruct_d = {\lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool3_d [19:4],
                               (\lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool3_d [0] && (! \lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool3_emitted [0]))};
  assign q1a8y_1_destruct_d = {\lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool3_d [35:20],
                               (\lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool3_d [0] && (! \lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool3_emitted [1]))};
  assign t1a8D_1_destruct_d = {\lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool3_d [51:36],
                               (\lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool3_d [0] && (! \lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool3_emitted [2]))};
  assign q2a8z_1_destruct_d = {\lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool3_d [67:52],
                               (\lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool3_d [0] && (! \lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool3_emitted [3]))};
  assign t2a8E_1_destruct_d = {\lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool3_d [83:68],
                               (\lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool3_d [0] && (! \lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool3_emitted [4]))};
  assign q3a8A_1_destruct_d = {\lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool3_d [99:84],
                               (\lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool3_d [0] && (! \lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool3_emitted [5]))};
  assign t3a8F_1_destruct_d = {\lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool3_d [115:100],
                               (\lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool3_d [0] && (! \lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool3_emitted [6]))};
  assign \lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool3_done  = (\lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool3_emitted  | ({t3a8F_1_destruct_d[0],
                                                                                                                               q3a8A_1_destruct_d[0],
                                                                                                                               t2a8E_1_destruct_d[0],
                                                                                                                               q2a8z_1_destruct_d[0],
                                                                                                                               t1a8D_1_destruct_d[0],
                                                                                                                               q1a8y_1_destruct_d[0],
                                                                                                                               sc_0_11_destruct_d[0]} & {t3a8F_1_destruct_r,
                                                                                                                                                         q3a8A_1_destruct_r,
                                                                                                                                                         t2a8E_1_destruct_r,
                                                                                                                                                         q2a8z_1_destruct_r,
                                                                                                                                                         t1a8D_1_destruct_r,
                                                                                                                                                         q1a8y_1_destruct_r,
                                                                                                                                                         sc_0_11_destruct_r}));
  assign \lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool3_r  = (& \lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool3_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool3_emitted  <= 7'd0;
    else
      \lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool3_emitted  <= (\lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool3_r  ? 7'd0 :
                                                                   \lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool3_done );
  
  /* demux (Ty CTf'''''''''_f'''''''''_Bool,
       Ty CTf'''''''''_f'''''''''_Bool) : (lizzieLet53_2,CTf'''''''''_f'''''''''_Bool) (lizzieLet53_1,CTf'''''''''_f'''''''''_Bool) > [(_1,CTf'''''''''_f'''''''''_Bool),
                                                                                                                                       (lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool3,CTf'''''''''_f'''''''''_Bool),
                                                                                                                                       (lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool2,CTf'''''''''_f'''''''''_Bool),
                                                                                                                                       (lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool1,CTf'''''''''_f'''''''''_Bool),
                                                                                                                                       (lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool0,CTf'''''''''_f'''''''''_Bool)] */
  logic [4:0] lizzieLet53_1_onehotd;
  always_comb
    if ((lizzieLet53_2_d[0] && lizzieLet53_1_d[0]))
      unique case (lizzieLet53_2_d[3:1])
        3'd0: lizzieLet53_1_onehotd = 5'd1;
        3'd1: lizzieLet53_1_onehotd = 5'd2;
        3'd2: lizzieLet53_1_onehotd = 5'd4;
        3'd3: lizzieLet53_1_onehotd = 5'd8;
        3'd4: lizzieLet53_1_onehotd = 5'd16;
        default: lizzieLet53_1_onehotd = 5'd0;
      endcase
    else lizzieLet53_1_onehotd = 5'd0;
  assign _1_d = {lizzieLet53_1_d[115:1], lizzieLet53_1_onehotd[0]};
  assign \lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool3_d  = {lizzieLet53_1_d[115:1],
                                                               lizzieLet53_1_onehotd[1]};
  assign \lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool2_d  = {lizzieLet53_1_d[115:1],
                                                               lizzieLet53_1_onehotd[2]};
  assign \lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool1_d  = {lizzieLet53_1_d[115:1],
                                                               lizzieLet53_1_onehotd[3]};
  assign \lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool0_d  = {lizzieLet53_1_d[115:1],
                                                               lizzieLet53_1_onehotd[4]};
  assign lizzieLet53_1_r = (| (lizzieLet53_1_onehotd & {\lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool0_r ,
                                                        \lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool1_r ,
                                                        \lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool2_r ,
                                                        \lizzieLet53_1Lcall_f'''''''''_f'''''''''_Bool3_r ,
                                                        _1_r}));
  assign lizzieLet53_2_r = lizzieLet53_1_r;
  
  /* demux (Ty CTf'''''''''_f'''''''''_Bool,
       Ty Go) : (lizzieLet53_3,CTf'''''''''_f'''''''''_Bool) (go_11_goMux_data,Go) > [(_0,Go),
                                                                                      (lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool3,Go),
                                                                                      (lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool2,Go),
                                                                                      (lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool1,Go),
                                                                                      (lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool0,Go)] */
  logic [4:0] go_11_goMux_data_onehotd;
  always_comb
    if ((lizzieLet53_3_d[0] && go_11_goMux_data_d[0]))
      unique case (lizzieLet53_3_d[3:1])
        3'd0: go_11_goMux_data_onehotd = 5'd1;
        3'd1: go_11_goMux_data_onehotd = 5'd2;
        3'd2: go_11_goMux_data_onehotd = 5'd4;
        3'd3: go_11_goMux_data_onehotd = 5'd8;
        3'd4: go_11_goMux_data_onehotd = 5'd16;
        default: go_11_goMux_data_onehotd = 5'd0;
      endcase
    else go_11_goMux_data_onehotd = 5'd0;
  assign _0_d = go_11_goMux_data_onehotd[0];
  assign \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool3_d  = go_11_goMux_data_onehotd[1];
  assign \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool2_d  = go_11_goMux_data_onehotd[2];
  assign \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool1_d  = go_11_goMux_data_onehotd[3];
  assign \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool0_d  = go_11_goMux_data_onehotd[4];
  assign go_11_goMux_data_r = (| (go_11_goMux_data_onehotd & {\lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool0_r ,
                                                              \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool1_r ,
                                                              \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool2_r ,
                                                              \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool3_r ,
                                                              _0_r}));
  assign lizzieLet53_3_r = go_11_goMux_data_r;
  
  /* buf (Ty Go) : (lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool0,Go) > (lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool0_1_argbuf,Go) */
  Go_t \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool0_bufchan_d ;
  logic \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool0_bufchan_r ;
  assign \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool0_r  = ((! \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool0_bufchan_d [0]) || \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool0_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool0_bufchan_d  <= 1'd0;
    else
      if (\lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool0_r )
        \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool0_bufchan_d  <= \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool0_d ;
  Go_t \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool0_bufchan_buf ;
  assign \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool0_bufchan_r  = (! \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool0_bufchan_buf [0]);
  assign \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool0_1_argbuf_d  = (\lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool0_bufchan_buf [0] ? \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool0_bufchan_buf  :
                                                                        \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool0_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool0_bufchan_buf  <= 1'd0;
    else
      if ((\lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool0_1_argbuf_r  && \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool0_bufchan_buf [0]))
        \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool0_bufchan_buf  <= 1'd0;
      else if (((! \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool0_1_argbuf_r ) && (! \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool0_bufchan_buf [0])))
        \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool0_bufchan_buf  <= \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool0_bufchan_d ;
  
  /* buf (Ty Go) : (lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool1,Go) > (lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool1_1_argbuf,Go) */
  Go_t \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool1_bufchan_d ;
  logic \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool1_bufchan_r ;
  assign \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool1_r  = ((! \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool1_bufchan_d [0]) || \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool1_bufchan_d  <= 1'd0;
    else
      if (\lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool1_r )
        \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool1_bufchan_d  <= \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool1_d ;
  Go_t \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool1_bufchan_buf ;
  assign \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool1_bufchan_r  = (! \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool1_bufchan_buf [0]);
  assign \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool1_1_argbuf_d  = (\lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool1_bufchan_buf [0] ? \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool1_bufchan_buf  :
                                                                        \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool1_bufchan_buf  <= 1'd0;
    else
      if ((\lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool1_1_argbuf_r  && \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool1_bufchan_buf [0]))
        \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool1_bufchan_buf  <= 1'd0;
      else if (((! \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool1_1_argbuf_r ) && (! \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool1_bufchan_buf [0])))
        \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool1_bufchan_buf  <= \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool1_bufchan_d ;
  
  /* buf (Ty Go) : (lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool2,Go) > (lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool2_1_argbuf,Go) */
  Go_t \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool2_bufchan_d ;
  logic \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool2_bufchan_r ;
  assign \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool2_r  = ((! \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool2_bufchan_d [0]) || \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool2_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool2_bufchan_d  <= 1'd0;
    else
      if (\lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool2_r )
        \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool2_bufchan_d  <= \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool2_d ;
  Go_t \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool2_bufchan_buf ;
  assign \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool2_bufchan_r  = (! \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool2_bufchan_buf [0]);
  assign \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool2_1_argbuf_d  = (\lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool2_bufchan_buf [0] ? \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool2_bufchan_buf  :
                                                                        \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool2_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool2_bufchan_buf  <= 1'd0;
    else
      if ((\lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool2_1_argbuf_r  && \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool2_bufchan_buf [0]))
        \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool2_bufchan_buf  <= 1'd0;
      else if (((! \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool2_1_argbuf_r ) && (! \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool2_bufchan_buf [0])))
        \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool2_bufchan_buf  <= \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool2_bufchan_d ;
  
  /* buf (Ty Go) : (lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool3,Go) > (lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool3_1_argbuf,Go) */
  Go_t \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool3_bufchan_d ;
  logic \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool3_bufchan_r ;
  assign \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool3_r  = ((! \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool3_bufchan_d [0]) || \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool3_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool3_bufchan_d  <= 1'd0;
    else
      if (\lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool3_r )
        \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool3_bufchan_d  <= \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool3_d ;
  Go_t \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool3_bufchan_buf ;
  assign \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool3_bufchan_r  = (! \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool3_bufchan_buf [0]);
  assign \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool3_1_argbuf_d  = (\lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool3_bufchan_buf [0] ? \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool3_bufchan_buf  :
                                                                        \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool3_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool3_bufchan_buf  <= 1'd0;
    else
      if ((\lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool3_1_argbuf_r  && \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool3_bufchan_buf [0]))
        \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool3_bufchan_buf  <= 1'd0;
      else if (((! \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool3_1_argbuf_r ) && (! \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool3_bufchan_buf [0])))
        \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool3_bufchan_buf  <= \lizzieLet53_3Lcall_f'''''''''_f'''''''''_Bool3_bufchan_d ;
  
  /* demux (Ty CTf'''''''''_f'''''''''_Bool,
       Ty Pointer_QTree_Bool) : (lizzieLet53_4,CTf'''''''''_f'''''''''_Bool) (srtarg_0_2_goMux_mux,Pointer_QTree_Bool) > [(lizzieLet53_4Lf'''''''''_f'''''''''_Boolsbos,Pointer_QTree_Bool),
                                                                                                                          (lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool3,Pointer_QTree_Bool),
                                                                                                                          (lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool2,Pointer_QTree_Bool),
                                                                                                                          (lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool1,Pointer_QTree_Bool),
                                                                                                                          (lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool0,Pointer_QTree_Bool)] */
  logic [4:0] srtarg_0_2_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet53_4_d[0] && srtarg_0_2_goMux_mux_d[0]))
      unique case (lizzieLet53_4_d[3:1])
        3'd0: srtarg_0_2_goMux_mux_onehotd = 5'd1;
        3'd1: srtarg_0_2_goMux_mux_onehotd = 5'd2;
        3'd2: srtarg_0_2_goMux_mux_onehotd = 5'd4;
        3'd3: srtarg_0_2_goMux_mux_onehotd = 5'd8;
        3'd4: srtarg_0_2_goMux_mux_onehotd = 5'd16;
        default: srtarg_0_2_goMux_mux_onehotd = 5'd0;
      endcase
    else srtarg_0_2_goMux_mux_onehotd = 5'd0;
  assign \lizzieLet53_4Lf'''''''''_f'''''''''_Boolsbos_d  = {srtarg_0_2_goMux_mux_d[16:1],
                                                             srtarg_0_2_goMux_mux_onehotd[0]};
  assign \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool3_d  = {srtarg_0_2_goMux_mux_d[16:1],
                                                               srtarg_0_2_goMux_mux_onehotd[1]};
  assign \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool2_d  = {srtarg_0_2_goMux_mux_d[16:1],
                                                               srtarg_0_2_goMux_mux_onehotd[2]};
  assign \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool1_d  = {srtarg_0_2_goMux_mux_d[16:1],
                                                               srtarg_0_2_goMux_mux_onehotd[3]};
  assign \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool0_d  = {srtarg_0_2_goMux_mux_d[16:1],
                                                               srtarg_0_2_goMux_mux_onehotd[4]};
  assign srtarg_0_2_goMux_mux_r = (| (srtarg_0_2_goMux_mux_onehotd & {\lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool0_r ,
                                                                      \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool1_r ,
                                                                      \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool2_r ,
                                                                      \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool3_r ,
                                                                      \lizzieLet53_4Lf'''''''''_f'''''''''_Boolsbos_r }));
  assign lizzieLet53_4_r = srtarg_0_2_goMux_mux_r;
  
  /* dcon (Ty QTree_Bool,
      Dcon QNode_Bool) : [(lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool0,Pointer_QTree_Bool),
                          (es_1_2_destruct,Pointer_QTree_Bool),
                          (es_2_4_destruct,Pointer_QTree_Bool),
                          (es_3_6_destruct,Pointer_QTree_Bool)] > (lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool0_1es_1_2_1es_2_4_1es_3_6_1QNode_Bool,QTree_Bool) */
  assign \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool0_1es_1_2_1es_2_4_1es_3_6_1QNode_Bool_d  = QNode_Bool_dc((& {\lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool0_d [0],
                                                                                                                    es_1_2_destruct_d[0],
                                                                                                                    es_2_4_destruct_d[0],
                                                                                                                    es_3_6_destruct_d[0]}), \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool0_d , es_1_2_destruct_d, es_2_4_destruct_d, es_3_6_destruct_d);
  assign {\lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool0_r ,
          es_1_2_destruct_r,
          es_2_4_destruct_r,
          es_3_6_destruct_r} = {4 {(\lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool0_1es_1_2_1es_2_4_1es_3_6_1QNode_Bool_r  && \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool0_1es_1_2_1es_2_4_1es_3_6_1QNode_Bool_d [0])}};
  
  /* buf (Ty QTree_Bool) : (lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool0_1es_1_2_1es_2_4_1es_3_6_1QNode_Bool,QTree_Bool) > (lizzieLet57_1_argbuf,QTree_Bool) */
  QTree_Bool_t \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool0_1es_1_2_1es_2_4_1es_3_6_1QNode_Bool_bufchan_d ;
  logic \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool0_1es_1_2_1es_2_4_1es_3_6_1QNode_Bool_bufchan_r ;
  assign \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool0_1es_1_2_1es_2_4_1es_3_6_1QNode_Bool_r  = ((! \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool0_1es_1_2_1es_2_4_1es_3_6_1QNode_Bool_bufchan_d [0]) || \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool0_1es_1_2_1es_2_4_1es_3_6_1QNode_Bool_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool0_1es_1_2_1es_2_4_1es_3_6_1QNode_Bool_bufchan_d  <= {66'd0,
                                                                                                         1'd0};
    else
      if (\lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool0_1es_1_2_1es_2_4_1es_3_6_1QNode_Bool_r )
        \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool0_1es_1_2_1es_2_4_1es_3_6_1QNode_Bool_bufchan_d  <= \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool0_1es_1_2_1es_2_4_1es_3_6_1QNode_Bool_d ;
  QTree_Bool_t \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool0_1es_1_2_1es_2_4_1es_3_6_1QNode_Bool_bufchan_buf ;
  assign \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool0_1es_1_2_1es_2_4_1es_3_6_1QNode_Bool_bufchan_r  = (! \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool0_1es_1_2_1es_2_4_1es_3_6_1QNode_Bool_bufchan_buf [0]);
  assign lizzieLet57_1_argbuf_d = (\lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool0_1es_1_2_1es_2_4_1es_3_6_1QNode_Bool_bufchan_buf [0] ? \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool0_1es_1_2_1es_2_4_1es_3_6_1QNode_Bool_bufchan_buf  :
                                   \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool0_1es_1_2_1es_2_4_1es_3_6_1QNode_Bool_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool0_1es_1_2_1es_2_4_1es_3_6_1QNode_Bool_bufchan_buf  <= {66'd0,
                                                                                                           1'd0};
    else
      if ((lizzieLet57_1_argbuf_r && \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool0_1es_1_2_1es_2_4_1es_3_6_1QNode_Bool_bufchan_buf [0]))
        \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool0_1es_1_2_1es_2_4_1es_3_6_1QNode_Bool_bufchan_buf  <= {66'd0,
                                                                                                             1'd0};
      else if (((! lizzieLet57_1_argbuf_r) && (! \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool0_1es_1_2_1es_2_4_1es_3_6_1QNode_Bool_bufchan_buf [0])))
        \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool0_1es_1_2_1es_2_4_1es_3_6_1QNode_Bool_bufchan_buf  <= \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool0_1es_1_2_1es_2_4_1es_3_6_1QNode_Bool_bufchan_d ;
  
  /* dcon (Ty CTf'''''''''_f'''''''''_Bool,
      Dcon Lcall_f'''''''''_f'''''''''_Bool0) : [(lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool1,Pointer_QTree_Bool),
                                                 (es_2_3_destruct,Pointer_QTree_Bool),
                                                 (es_3_5_destruct,Pointer_QTree_Bool),
                                                 (sc_0_13_destruct,Pointer_CTf'''''''''_f'''''''''_Bool)] > (lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool1_1es_2_3_1es_3_5_1sc_0_13_1Lcall_f'''''''''_f'''''''''_Bool0,CTf'''''''''_f'''''''''_Bool) */
  assign \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool1_1es_2_3_1es_3_5_1sc_0_13_1Lcall_f'''''''''_f'''''''''_Bool0_d  = \Lcall_f'''''''''_f'''''''''_Bool0_dc ((& {\lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool1_d [0],
                                                                                                                                                                     es_2_3_destruct_d[0],
                                                                                                                                                                     es_3_5_destruct_d[0],
                                                                                                                                                                     sc_0_13_destruct_d[0]}), \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool1_d , es_2_3_destruct_d, es_3_5_destruct_d, sc_0_13_destruct_d);
  assign {\lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool1_r ,
          es_2_3_destruct_r,
          es_3_5_destruct_r,
          sc_0_13_destruct_r} = {4 {(\lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool1_1es_2_3_1es_3_5_1sc_0_13_1Lcall_f'''''''''_f'''''''''_Bool0_r  && \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool1_1es_2_3_1es_3_5_1sc_0_13_1Lcall_f'''''''''_f'''''''''_Bool0_d [0])}};
  
  /* buf (Ty CTf'''''''''_f'''''''''_Bool) : (lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool1_1es_2_3_1es_3_5_1sc_0_13_1Lcall_f'''''''''_f'''''''''_Bool0,CTf'''''''''_f'''''''''_Bool) > (lizzieLet56_1_argbuf,CTf'''''''''_f'''''''''_Bool) */
  \CTf'''''''''_f'''''''''_Bool_t  \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool1_1es_2_3_1es_3_5_1sc_0_13_1Lcall_f'''''''''_f'''''''''_Bool0_bufchan_d ;
  logic \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool1_1es_2_3_1es_3_5_1sc_0_13_1Lcall_f'''''''''_f'''''''''_Bool0_bufchan_r ;
  assign \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool1_1es_2_3_1es_3_5_1sc_0_13_1Lcall_f'''''''''_f'''''''''_Bool0_r  = ((! \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool1_1es_2_3_1es_3_5_1sc_0_13_1Lcall_f'''''''''_f'''''''''_Bool0_bufchan_d [0]) || \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool1_1es_2_3_1es_3_5_1sc_0_13_1Lcall_f'''''''''_f'''''''''_Bool0_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool1_1es_2_3_1es_3_5_1sc_0_13_1Lcall_f'''''''''_f'''''''''_Bool0_bufchan_d  <= {115'd0,
                                                                                                                                 1'd0};
    else
      if (\lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool1_1es_2_3_1es_3_5_1sc_0_13_1Lcall_f'''''''''_f'''''''''_Bool0_r )
        \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool1_1es_2_3_1es_3_5_1sc_0_13_1Lcall_f'''''''''_f'''''''''_Bool0_bufchan_d  <= \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool1_1es_2_3_1es_3_5_1sc_0_13_1Lcall_f'''''''''_f'''''''''_Bool0_d ;
  \CTf'''''''''_f'''''''''_Bool_t  \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool1_1es_2_3_1es_3_5_1sc_0_13_1Lcall_f'''''''''_f'''''''''_Bool0_bufchan_buf ;
  assign \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool1_1es_2_3_1es_3_5_1sc_0_13_1Lcall_f'''''''''_f'''''''''_Bool0_bufchan_r  = (! \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool1_1es_2_3_1es_3_5_1sc_0_13_1Lcall_f'''''''''_f'''''''''_Bool0_bufchan_buf [0]);
  assign lizzieLet56_1_argbuf_d = (\lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool1_1es_2_3_1es_3_5_1sc_0_13_1Lcall_f'''''''''_f'''''''''_Bool0_bufchan_buf [0] ? \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool1_1es_2_3_1es_3_5_1sc_0_13_1Lcall_f'''''''''_f'''''''''_Bool0_bufchan_buf  :
                                   \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool1_1es_2_3_1es_3_5_1sc_0_13_1Lcall_f'''''''''_f'''''''''_Bool0_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool1_1es_2_3_1es_3_5_1sc_0_13_1Lcall_f'''''''''_f'''''''''_Bool0_bufchan_buf  <= {115'd0,
                                                                                                                                   1'd0};
    else
      if ((lizzieLet56_1_argbuf_r && \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool1_1es_2_3_1es_3_5_1sc_0_13_1Lcall_f'''''''''_f'''''''''_Bool0_bufchan_buf [0]))
        \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool1_1es_2_3_1es_3_5_1sc_0_13_1Lcall_f'''''''''_f'''''''''_Bool0_bufchan_buf  <= {115'd0,
                                                                                                                                     1'd0};
      else if (((! lizzieLet56_1_argbuf_r) && (! \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool1_1es_2_3_1es_3_5_1sc_0_13_1Lcall_f'''''''''_f'''''''''_Bool0_bufchan_buf [0])))
        \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool1_1es_2_3_1es_3_5_1sc_0_13_1Lcall_f'''''''''_f'''''''''_Bool0_bufchan_buf  <= \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool1_1es_2_3_1es_3_5_1sc_0_13_1Lcall_f'''''''''_f'''''''''_Bool0_bufchan_d ;
  
  /* dcon (Ty CTf'''''''''_f'''''''''_Bool,
      Dcon Lcall_f'''''''''_f'''''''''_Bool1) : [(lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool2,Pointer_QTree_Bool),
                                                 (es_3_4_destruct,Pointer_QTree_Bool),
                                                 (sc_0_12_destruct,Pointer_CTf'''''''''_f'''''''''_Bool),
                                                 (q1a8y_2_destruct,Pointer_MaskQTree),
                                                 (t1a8D_2_destruct,Pointer_QTree_Bool)] > (lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool2_1es_3_4_1sc_0_12_1q1a8y_2_1t1a8D_2_1Lcall_f'''''''''_f'''''''''_Bool1,CTf'''''''''_f'''''''''_Bool) */
  assign \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool2_1es_3_4_1sc_0_12_1q1a8y_2_1t1a8D_2_1Lcall_f'''''''''_f'''''''''_Bool1_d  = \Lcall_f'''''''''_f'''''''''_Bool1_dc ((& {\lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool2_d [0],
                                                                                                                                                                               es_3_4_destruct_d[0],
                                                                                                                                                                               sc_0_12_destruct_d[0],
                                                                                                                                                                               q1a8y_2_destruct_d[0],
                                                                                                                                                                               t1a8D_2_destruct_d[0]}), \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool2_d , es_3_4_destruct_d, sc_0_12_destruct_d, q1a8y_2_destruct_d, t1a8D_2_destruct_d);
  assign {\lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool2_r ,
          es_3_4_destruct_r,
          sc_0_12_destruct_r,
          q1a8y_2_destruct_r,
          t1a8D_2_destruct_r} = {5 {(\lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool2_1es_3_4_1sc_0_12_1q1a8y_2_1t1a8D_2_1Lcall_f'''''''''_f'''''''''_Bool1_r  && \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool2_1es_3_4_1sc_0_12_1q1a8y_2_1t1a8D_2_1Lcall_f'''''''''_f'''''''''_Bool1_d [0])}};
  
  /* buf (Ty CTf'''''''''_f'''''''''_Bool) : (lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool2_1es_3_4_1sc_0_12_1q1a8y_2_1t1a8D_2_1Lcall_f'''''''''_f'''''''''_Bool1,CTf'''''''''_f'''''''''_Bool) > (lizzieLet55_1_argbuf,CTf'''''''''_f'''''''''_Bool) */
  \CTf'''''''''_f'''''''''_Bool_t  \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool2_1es_3_4_1sc_0_12_1q1a8y_2_1t1a8D_2_1Lcall_f'''''''''_f'''''''''_Bool1_bufchan_d ;
  logic \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool2_1es_3_4_1sc_0_12_1q1a8y_2_1t1a8D_2_1Lcall_f'''''''''_f'''''''''_Bool1_bufchan_r ;
  assign \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool2_1es_3_4_1sc_0_12_1q1a8y_2_1t1a8D_2_1Lcall_f'''''''''_f'''''''''_Bool1_r  = ((! \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool2_1es_3_4_1sc_0_12_1q1a8y_2_1t1a8D_2_1Lcall_f'''''''''_f'''''''''_Bool1_bufchan_d [0]) || \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool2_1es_3_4_1sc_0_12_1q1a8y_2_1t1a8D_2_1Lcall_f'''''''''_f'''''''''_Bool1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool2_1es_3_4_1sc_0_12_1q1a8y_2_1t1a8D_2_1Lcall_f'''''''''_f'''''''''_Bool1_bufchan_d  <= {115'd0,
                                                                                                                                           1'd0};
    else
      if (\lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool2_1es_3_4_1sc_0_12_1q1a8y_2_1t1a8D_2_1Lcall_f'''''''''_f'''''''''_Bool1_r )
        \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool2_1es_3_4_1sc_0_12_1q1a8y_2_1t1a8D_2_1Lcall_f'''''''''_f'''''''''_Bool1_bufchan_d  <= \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool2_1es_3_4_1sc_0_12_1q1a8y_2_1t1a8D_2_1Lcall_f'''''''''_f'''''''''_Bool1_d ;
  \CTf'''''''''_f'''''''''_Bool_t  \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool2_1es_3_4_1sc_0_12_1q1a8y_2_1t1a8D_2_1Lcall_f'''''''''_f'''''''''_Bool1_bufchan_buf ;
  assign \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool2_1es_3_4_1sc_0_12_1q1a8y_2_1t1a8D_2_1Lcall_f'''''''''_f'''''''''_Bool1_bufchan_r  = (! \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool2_1es_3_4_1sc_0_12_1q1a8y_2_1t1a8D_2_1Lcall_f'''''''''_f'''''''''_Bool1_bufchan_buf [0]);
  assign lizzieLet55_1_argbuf_d = (\lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool2_1es_3_4_1sc_0_12_1q1a8y_2_1t1a8D_2_1Lcall_f'''''''''_f'''''''''_Bool1_bufchan_buf [0] ? \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool2_1es_3_4_1sc_0_12_1q1a8y_2_1t1a8D_2_1Lcall_f'''''''''_f'''''''''_Bool1_bufchan_buf  :
                                   \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool2_1es_3_4_1sc_0_12_1q1a8y_2_1t1a8D_2_1Lcall_f'''''''''_f'''''''''_Bool1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool2_1es_3_4_1sc_0_12_1q1a8y_2_1t1a8D_2_1Lcall_f'''''''''_f'''''''''_Bool1_bufchan_buf  <= {115'd0,
                                                                                                                                             1'd0};
    else
      if ((lizzieLet55_1_argbuf_r && \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool2_1es_3_4_1sc_0_12_1q1a8y_2_1t1a8D_2_1Lcall_f'''''''''_f'''''''''_Bool1_bufchan_buf [0]))
        \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool2_1es_3_4_1sc_0_12_1q1a8y_2_1t1a8D_2_1Lcall_f'''''''''_f'''''''''_Bool1_bufchan_buf  <= {115'd0,
                                                                                                                                               1'd0};
      else if (((! lizzieLet55_1_argbuf_r) && (! \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool2_1es_3_4_1sc_0_12_1q1a8y_2_1t1a8D_2_1Lcall_f'''''''''_f'''''''''_Bool1_bufchan_buf [0])))
        \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool2_1es_3_4_1sc_0_12_1q1a8y_2_1t1a8D_2_1Lcall_f'''''''''_f'''''''''_Bool1_bufchan_buf  <= \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool2_1es_3_4_1sc_0_12_1q1a8y_2_1t1a8D_2_1Lcall_f'''''''''_f'''''''''_Bool1_bufchan_d ;
  
  /* dcon (Ty CTf'''''''''_f'''''''''_Bool,
      Dcon Lcall_f'''''''''_f'''''''''_Bool2) : [(lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool3,Pointer_QTree_Bool),
                                                 (sc_0_11_destruct,Pointer_CTf'''''''''_f'''''''''_Bool),
                                                 (q1a8y_1_destruct,Pointer_MaskQTree),
                                                 (t1a8D_1_destruct,Pointer_QTree_Bool),
                                                 (q2a8z_1_destruct,Pointer_MaskQTree),
                                                 (t2a8E_1_destruct,Pointer_QTree_Bool)] > (lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool3_1sc_0_11_1q1a8y_1_1t1a8D_1_1q2a8z_1_1t2a8E_1_1Lcall_f'''''''''_f'''''''''_Bool2,CTf'''''''''_f'''''''''_Bool) */
  assign \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool3_1sc_0_11_1q1a8y_1_1t1a8D_1_1q2a8z_1_1t2a8E_1_1Lcall_f'''''''''_f'''''''''_Bool2_d  = \Lcall_f'''''''''_f'''''''''_Bool2_dc ((& {\lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool3_d [0],
                                                                                                                                                                                         sc_0_11_destruct_d[0],
                                                                                                                                                                                         q1a8y_1_destruct_d[0],
                                                                                                                                                                                         t1a8D_1_destruct_d[0],
                                                                                                                                                                                         q2a8z_1_destruct_d[0],
                                                                                                                                                                                         t2a8E_1_destruct_d[0]}), \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool3_d , sc_0_11_destruct_d, q1a8y_1_destruct_d, t1a8D_1_destruct_d, q2a8z_1_destruct_d, t2a8E_1_destruct_d);
  assign {\lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool3_r ,
          sc_0_11_destruct_r,
          q1a8y_1_destruct_r,
          t1a8D_1_destruct_r,
          q2a8z_1_destruct_r,
          t2a8E_1_destruct_r} = {6 {(\lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool3_1sc_0_11_1q1a8y_1_1t1a8D_1_1q2a8z_1_1t2a8E_1_1Lcall_f'''''''''_f'''''''''_Bool2_r  && \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool3_1sc_0_11_1q1a8y_1_1t1a8D_1_1q2a8z_1_1t2a8E_1_1Lcall_f'''''''''_f'''''''''_Bool2_d [0])}};
  
  /* buf (Ty CTf'''''''''_f'''''''''_Bool) : (lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool3_1sc_0_11_1q1a8y_1_1t1a8D_1_1q2a8z_1_1t2a8E_1_1Lcall_f'''''''''_f'''''''''_Bool2,CTf'''''''''_f'''''''''_Bool) > (lizzieLet54_1_argbuf,CTf'''''''''_f'''''''''_Bool) */
  \CTf'''''''''_f'''''''''_Bool_t  \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool3_1sc_0_11_1q1a8y_1_1t1a8D_1_1q2a8z_1_1t2a8E_1_1Lcall_f'''''''''_f'''''''''_Bool2_bufchan_d ;
  logic \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool3_1sc_0_11_1q1a8y_1_1t1a8D_1_1q2a8z_1_1t2a8E_1_1Lcall_f'''''''''_f'''''''''_Bool2_bufchan_r ;
  assign \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool3_1sc_0_11_1q1a8y_1_1t1a8D_1_1q2a8z_1_1t2a8E_1_1Lcall_f'''''''''_f'''''''''_Bool2_r  = ((! \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool3_1sc_0_11_1q1a8y_1_1t1a8D_1_1q2a8z_1_1t2a8E_1_1Lcall_f'''''''''_f'''''''''_Bool2_bufchan_d [0]) || \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool3_1sc_0_11_1q1a8y_1_1t1a8D_1_1q2a8z_1_1t2a8E_1_1Lcall_f'''''''''_f'''''''''_Bool2_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool3_1sc_0_11_1q1a8y_1_1t1a8D_1_1q2a8z_1_1t2a8E_1_1Lcall_f'''''''''_f'''''''''_Bool2_bufchan_d  <= {115'd0,
                                                                                                                                                     1'd0};
    else
      if (\lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool3_1sc_0_11_1q1a8y_1_1t1a8D_1_1q2a8z_1_1t2a8E_1_1Lcall_f'''''''''_f'''''''''_Bool2_r )
        \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool3_1sc_0_11_1q1a8y_1_1t1a8D_1_1q2a8z_1_1t2a8E_1_1Lcall_f'''''''''_f'''''''''_Bool2_bufchan_d  <= \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool3_1sc_0_11_1q1a8y_1_1t1a8D_1_1q2a8z_1_1t2a8E_1_1Lcall_f'''''''''_f'''''''''_Bool2_d ;
  \CTf'''''''''_f'''''''''_Bool_t  \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool3_1sc_0_11_1q1a8y_1_1t1a8D_1_1q2a8z_1_1t2a8E_1_1Lcall_f'''''''''_f'''''''''_Bool2_bufchan_buf ;
  assign \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool3_1sc_0_11_1q1a8y_1_1t1a8D_1_1q2a8z_1_1t2a8E_1_1Lcall_f'''''''''_f'''''''''_Bool2_bufchan_r  = (! \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool3_1sc_0_11_1q1a8y_1_1t1a8D_1_1q2a8z_1_1t2a8E_1_1Lcall_f'''''''''_f'''''''''_Bool2_bufchan_buf [0]);
  assign lizzieLet54_1_argbuf_d = (\lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool3_1sc_0_11_1q1a8y_1_1t1a8D_1_1q2a8z_1_1t2a8E_1_1Lcall_f'''''''''_f'''''''''_Bool2_bufchan_buf [0] ? \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool3_1sc_0_11_1q1a8y_1_1t1a8D_1_1q2a8z_1_1t2a8E_1_1Lcall_f'''''''''_f'''''''''_Bool2_bufchan_buf  :
                                   \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool3_1sc_0_11_1q1a8y_1_1t1a8D_1_1q2a8z_1_1t2a8E_1_1Lcall_f'''''''''_f'''''''''_Bool2_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool3_1sc_0_11_1q1a8y_1_1t1a8D_1_1q2a8z_1_1t2a8E_1_1Lcall_f'''''''''_f'''''''''_Bool2_bufchan_buf  <= {115'd0,
                                                                                                                                                       1'd0};
    else
      if ((lizzieLet54_1_argbuf_r && \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool3_1sc_0_11_1q1a8y_1_1t1a8D_1_1q2a8z_1_1t2a8E_1_1Lcall_f'''''''''_f'''''''''_Bool2_bufchan_buf [0]))
        \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool3_1sc_0_11_1q1a8y_1_1t1a8D_1_1q2a8z_1_1t2a8E_1_1Lcall_f'''''''''_f'''''''''_Bool2_bufchan_buf  <= {115'd0,
                                                                                                                                                         1'd0};
      else if (((! lizzieLet54_1_argbuf_r) && (! \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool3_1sc_0_11_1q1a8y_1_1t1a8D_1_1q2a8z_1_1t2a8E_1_1Lcall_f'''''''''_f'''''''''_Bool2_bufchan_buf [0])))
        \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool3_1sc_0_11_1q1a8y_1_1t1a8D_1_1q2a8z_1_1t2a8E_1_1Lcall_f'''''''''_f'''''''''_Bool2_bufchan_buf  <= \lizzieLet53_4Lcall_f'''''''''_f'''''''''_Bool3_1sc_0_11_1q1a8y_1_1t1a8D_1_1q2a8z_1_1t2a8E_1_1Lcall_f'''''''''_f'''''''''_Bool2_bufchan_d ;
  
  /* fork (Ty Pointer_QTree_Bool) : (lizzieLet53_4Lf'''''''''_f'''''''''_Boolsbos,Pointer_QTree_Bool) > [(lizzieLet53_4Lf'''''''''_f'''''''''_Boolsbos_1_merge_merge_fork_1,Pointer_QTree_Bool),
                                                                                                    (lizzieLet53_4Lf'''''''''_f'''''''''_Boolsbos_1_merge_merge_fork_2,Pointer_QTree_Bool)] */
  logic [1:0] \lizzieLet53_4Lf'''''''''_f'''''''''_Boolsbos_emitted ;
  logic [1:0] \lizzieLet53_4Lf'''''''''_f'''''''''_Boolsbos_done ;
  assign \lizzieLet53_4Lf'''''''''_f'''''''''_Boolsbos_1_merge_merge_fork_1_d  = {\lizzieLet53_4Lf'''''''''_f'''''''''_Boolsbos_d [16:1],
                                                                                  (\lizzieLet53_4Lf'''''''''_f'''''''''_Boolsbos_d [0] && (! \lizzieLet53_4Lf'''''''''_f'''''''''_Boolsbos_emitted [0]))};
  assign \lizzieLet53_4Lf'''''''''_f'''''''''_Boolsbos_1_merge_merge_fork_2_d  = {\lizzieLet53_4Lf'''''''''_f'''''''''_Boolsbos_d [16:1],
                                                                                  (\lizzieLet53_4Lf'''''''''_f'''''''''_Boolsbos_d [0] && (! \lizzieLet53_4Lf'''''''''_f'''''''''_Boolsbos_emitted [1]))};
  assign \lizzieLet53_4Lf'''''''''_f'''''''''_Boolsbos_done  = (\lizzieLet53_4Lf'''''''''_f'''''''''_Boolsbos_emitted  | ({\lizzieLet53_4Lf'''''''''_f'''''''''_Boolsbos_1_merge_merge_fork_2_d [0],
                                                                                                                           \lizzieLet53_4Lf'''''''''_f'''''''''_Boolsbos_1_merge_merge_fork_1_d [0]} & {\lizzieLet53_4Lf'''''''''_f'''''''''_Boolsbos_1_merge_merge_fork_2_r ,
                                                                                                                                                                                                        \lizzieLet53_4Lf'''''''''_f'''''''''_Boolsbos_1_merge_merge_fork_1_r }));
  assign \lizzieLet53_4Lf'''''''''_f'''''''''_Boolsbos_r  = (& \lizzieLet53_4Lf'''''''''_f'''''''''_Boolsbos_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet53_4Lf'''''''''_f'''''''''_Boolsbos_emitted  <= 2'd0;
    else
      \lizzieLet53_4Lf'''''''''_f'''''''''_Boolsbos_emitted  <= (\lizzieLet53_4Lf'''''''''_f'''''''''_Boolsbos_r  ? 2'd0 :
                                                                 \lizzieLet53_4Lf'''''''''_f'''''''''_Boolsbos_done );
  
  /* togo (Ty Pointer_QTree_Bool) : (lizzieLet53_4Lf'''''''''_f'''''''''_Boolsbos_1_merge_merge_fork_1,Pointer_QTree_Bool) > (call_f'''''''''_f'''''''''_Bool_goConst,Go) */
  assign \call_f'''''''''_f'''''''''_Bool_goConst_d  = \lizzieLet53_4Lf'''''''''_f'''''''''_Boolsbos_1_merge_merge_fork_1_d [0];
  assign \lizzieLet53_4Lf'''''''''_f'''''''''_Boolsbos_1_merge_merge_fork_1_r  = \call_f'''''''''_f'''''''''_Bool_goConst_r ;
  
  /* mergectrl (Ty C2,Ty TupGo) : [(lvlrcX-0TupGo_1,TupGo),
                              (lvlrcX-0TupGo2,TupGo)] > (lvlrcX-0_choice,C2) (lvlrcX-0_data,TupGo) */
  logic [1:0] \lvlrcX-0TupGo_1_select_d ;
  assign \lvlrcX-0TupGo_1_select_d  = ((| \lvlrcX-0TupGo_1_select_q ) ? \lvlrcX-0TupGo_1_select_q  :
                                       (\lvlrcX-0TupGo_1_d [0] ? 2'd1 :
                                        (\lvlrcX-0TupGo2_d [0] ? 2'd2 :
                                         2'd0)));
  logic [1:0] \lvlrcX-0TupGo_1_select_q ;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \lvlrcX-0TupGo_1_select_q  <= 2'd0;
    else
      \lvlrcX-0TupGo_1_select_q  <= (\lvlrcX-0TupGo_1_done  ? 2'd0 :
                                     \lvlrcX-0TupGo_1_select_d );
  logic [1:0] \lvlrcX-0TupGo_1_emit_q ;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \lvlrcX-0TupGo_1_emit_q  <= 2'd0;
    else
      \lvlrcX-0TupGo_1_emit_q  <= (\lvlrcX-0TupGo_1_done  ? 2'd0 :
                                   \lvlrcX-0TupGo_1_emit_d );
  logic [1:0] \lvlrcX-0TupGo_1_emit_d ;
  assign \lvlrcX-0TupGo_1_emit_d  = (\lvlrcX-0TupGo_1_emit_q  | ({\lvlrcX-0_choice_d [0],
                                                                  \lvlrcX-0_data_d [0]} & {\lvlrcX-0_choice_r ,
                                                                                           \lvlrcX-0_data_r }));
  logic \lvlrcX-0TupGo_1_done ;
  assign \lvlrcX-0TupGo_1_done  = (& \lvlrcX-0TupGo_1_emit_d );
  assign {\lvlrcX-0TupGo2_r ,
          \lvlrcX-0TupGo_1_r } = (\lvlrcX-0TupGo_1_done  ? \lvlrcX-0TupGo_1_select_d  :
                                  2'd0);
  assign \lvlrcX-0_data_d  = ((\lvlrcX-0TupGo_1_select_d [0] && (! \lvlrcX-0TupGo_1_emit_q [0])) ? \lvlrcX-0TupGo_1_d  :
                              ((\lvlrcX-0TupGo_1_select_d [1] && (! \lvlrcX-0TupGo_1_emit_q [0])) ? \lvlrcX-0TupGo2_d  :
                               1'd0));
  assign \lvlrcX-0_choice_d  = ((\lvlrcX-0TupGo_1_select_d [0] && (! \lvlrcX-0TupGo_1_emit_q [1])) ? C1_2_dc(1'd1) :
                                ((\lvlrcX-0TupGo_1_select_d [1] && (! \lvlrcX-0TupGo_1_emit_q [1])) ? C2_2_dc(1'd1) :
                                 {1'd0, 1'd0}));
  
  /* dcon (Ty MyBool,
      Dcon MyTrue) : [(lvlrcX-0TupGogo_8,Go)] > (go_8_1MyTrue,MyBool) */
  assign go_8_1MyTrue_d = MyTrue_dc((& {\lvlrcX-0TupGogo_8_d [0]}), \lvlrcX-0TupGogo_8_d );
  assign {\lvlrcX-0TupGogo_8_r } = {1 {(go_8_1MyTrue_r && go_8_1MyTrue_d[0])}};
  
  /* buf (Ty Pointer_QTree_Bool) : (lvlrcX-0_1,Pointer_QTree_Bool) > (lvlrcX-0_resbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t \lvlrcX-0_1_bufchan_d ;
  logic \lvlrcX-0_1_bufchan_r ;
  assign \lvlrcX-0_1_r  = ((! \lvlrcX-0_1_bufchan_d [0]) || \lvlrcX-0_1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \lvlrcX-0_1_bufchan_d  <= {16'd0, 1'd0};
    else if (\lvlrcX-0_1_r ) \lvlrcX-0_1_bufchan_d  <= \lvlrcX-0_1_d ;
  Pointer_QTree_Bool_t \lvlrcX-0_1_bufchan_buf ;
  assign \lvlrcX-0_1_bufchan_r  = (! \lvlrcX-0_1_bufchan_buf [0]);
  assign \lvlrcX-0_resbuf_d  = (\lvlrcX-0_1_bufchan_buf [0] ? \lvlrcX-0_1_bufchan_buf  :
                                \lvlrcX-0_1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \lvlrcX-0_1_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((\lvlrcX-0_resbuf_r  && \lvlrcX-0_1_bufchan_buf [0]))
        \lvlrcX-0_1_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! \lvlrcX-0_resbuf_r ) && (! \lvlrcX-0_1_bufchan_buf [0])))
        \lvlrcX-0_1_bufchan_buf  <= \lvlrcX-0_1_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Bool) : (lvlrcX-0_2,Pointer_QTree_Bool) > (lvlrcX-0_2_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t \lvlrcX-0_2_bufchan_d ;
  logic \lvlrcX-0_2_bufchan_r ;
  assign \lvlrcX-0_2_r  = ((! \lvlrcX-0_2_bufchan_d [0]) || \lvlrcX-0_2_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \lvlrcX-0_2_bufchan_d  <= {16'd0, 1'd0};
    else if (\lvlrcX-0_2_r ) \lvlrcX-0_2_bufchan_d  <= \lvlrcX-0_2_d ;
  Pointer_QTree_Bool_t \lvlrcX-0_2_bufchan_buf ;
  assign \lvlrcX-0_2_bufchan_r  = (! \lvlrcX-0_2_bufchan_buf [0]);
  assign \lvlrcX-0_2_argbuf_d  = (\lvlrcX-0_2_bufchan_buf [0] ? \lvlrcX-0_2_bufchan_buf  :
                                  \lvlrcX-0_2_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \lvlrcX-0_2_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((\lvlrcX-0_2_argbuf_r  && \lvlrcX-0_2_bufchan_buf [0]))
        \lvlrcX-0_2_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! \lvlrcX-0_2_argbuf_r ) && (! \lvlrcX-0_2_bufchan_buf [0])))
        \lvlrcX-0_2_bufchan_buf  <= \lvlrcX-0_2_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Bool) : (lvlrcX-0_2_argbuf,Pointer_QTree_Bool) > (lizzieLet24_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t \lvlrcX-0_2_argbuf_bufchan_d ;
  logic \lvlrcX-0_2_argbuf_bufchan_r ;
  assign \lvlrcX-0_2_argbuf_r  = ((! \lvlrcX-0_2_argbuf_bufchan_d [0]) || \lvlrcX-0_2_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lvlrcX-0_2_argbuf_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\lvlrcX-0_2_argbuf_r )
        \lvlrcX-0_2_argbuf_bufchan_d  <= \lvlrcX-0_2_argbuf_d ;
  Pointer_QTree_Bool_t \lvlrcX-0_2_argbuf_bufchan_buf ;
  assign \lvlrcX-0_2_argbuf_bufchan_r  = (! \lvlrcX-0_2_argbuf_bufchan_buf [0]);
  assign lizzieLet24_1_1_argbuf_d = (\lvlrcX-0_2_argbuf_bufchan_buf [0] ? \lvlrcX-0_2_argbuf_bufchan_buf  :
                                     \lvlrcX-0_2_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lvlrcX-0_2_argbuf_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((lizzieLet24_1_1_argbuf_r && \lvlrcX-0_2_argbuf_bufchan_buf [0]))
        \lvlrcX-0_2_argbuf_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! lizzieLet24_1_1_argbuf_r) && (! \lvlrcX-0_2_argbuf_bufchan_buf [0])))
        \lvlrcX-0_2_argbuf_bufchan_buf  <= \lvlrcX-0_2_argbuf_bufchan_d ;
  
  /* demux (Ty C2,
       Ty Pointer_QTree_Bool) : (lvlrcX-0_choice,C2) (writeQTree_BoollizzieLet42_1_argbuf_rwb,Pointer_QTree_Bool) > [(lvlrcX-0_1,Pointer_QTree_Bool),
                                                                                                                     (lvlrcX-0_2,Pointer_QTree_Bool)] */
  logic [1:0] writeQTree_BoollizzieLet42_1_argbuf_rwb_onehotd;
  always_comb
    if ((\lvlrcX-0_choice_d [0] && writeQTree_BoollizzieLet42_1_argbuf_rwb_d[0]))
      unique case (\lvlrcX-0_choice_d [1:1])
        1'd0: writeQTree_BoollizzieLet42_1_argbuf_rwb_onehotd = 2'd1;
        1'd1: writeQTree_BoollizzieLet42_1_argbuf_rwb_onehotd = 2'd2;
        default: writeQTree_BoollizzieLet42_1_argbuf_rwb_onehotd = 2'd0;
      endcase
    else writeQTree_BoollizzieLet42_1_argbuf_rwb_onehotd = 2'd0;
  assign \lvlrcX-0_1_d  = {writeQTree_BoollizzieLet42_1_argbuf_rwb_d[16:1],
                           writeQTree_BoollizzieLet42_1_argbuf_rwb_onehotd[0]};
  assign \lvlrcX-0_2_d  = {writeQTree_BoollizzieLet42_1_argbuf_rwb_d[16:1],
                           writeQTree_BoollizzieLet42_1_argbuf_rwb_onehotd[1]};
  assign writeQTree_BoollizzieLet42_1_argbuf_rwb_r = (| (writeQTree_BoollizzieLet42_1_argbuf_rwb_onehotd & {\lvlrcX-0_2_r ,
                                                                                                            \lvlrcX-0_1_r }));
  assign \lvlrcX-0_choice_r  = writeQTree_BoollizzieLet42_1_argbuf_rwb_r;
  
  /* destruct (Ty TupGo,
          Dcon TupGo) : (lvlrcX-0_data,TupGo) > [(lvlrcX-0TupGogo_8,Go)] */
  assign \lvlrcX-0TupGogo_8_d  = \lvlrcX-0_data_d [0];
  assign \lvlrcX-0_data_r  = \lvlrcX-0TupGogo_8_r ;
  
  /* buf (Ty Pointer_QTree_Bool) : (lvlrcX-0_resbuf,Pointer_QTree_Bool) > (lizzieLet23_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t \lvlrcX-0_resbuf_bufchan_d ;
  logic \lvlrcX-0_resbuf_bufchan_r ;
  assign \lvlrcX-0_resbuf_r  = ((! \lvlrcX-0_resbuf_bufchan_d [0]) || \lvlrcX-0_resbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \lvlrcX-0_resbuf_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\lvlrcX-0_resbuf_r )
        \lvlrcX-0_resbuf_bufchan_d  <= \lvlrcX-0_resbuf_d ;
  Pointer_QTree_Bool_t \lvlrcX-0_resbuf_bufchan_buf ;
  assign \lvlrcX-0_resbuf_bufchan_r  = (! \lvlrcX-0_resbuf_bufchan_buf [0]);
  assign lizzieLet23_1_1_argbuf_d = (\lvlrcX-0_resbuf_bufchan_buf [0] ? \lvlrcX-0_resbuf_bufchan_buf  :
                                     \lvlrcX-0_resbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lvlrcX-0_resbuf_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((lizzieLet23_1_1_argbuf_r && \lvlrcX-0_resbuf_bufchan_buf [0]))
        \lvlrcX-0_resbuf_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! lizzieLet23_1_1_argbuf_r) && (! \lvlrcX-0_resbuf_bufchan_buf [0])))
        \lvlrcX-0_resbuf_bufchan_buf  <= \lvlrcX-0_resbuf_bufchan_d ;
  
  /* buf (Ty Pointer_MaskQTree) : (m1a85_goMux_mux,Pointer_MaskQTree) > (m1a85_1_argbuf,Pointer_MaskQTree) */
  Pointer_MaskQTree_t m1a85_goMux_mux_bufchan_d;
  logic m1a85_goMux_mux_bufchan_r;
  assign m1a85_goMux_mux_r = ((! m1a85_goMux_mux_bufchan_d[0]) || m1a85_goMux_mux_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m1a85_goMux_mux_bufchan_d <= {16'd0, 1'd0};
    else
      if (m1a85_goMux_mux_r)
        m1a85_goMux_mux_bufchan_d <= m1a85_goMux_mux_d;
  Pointer_MaskQTree_t m1a85_goMux_mux_bufchan_buf;
  assign m1a85_goMux_mux_bufchan_r = (! m1a85_goMux_mux_bufchan_buf[0]);
  assign m1a85_1_argbuf_d = (m1a85_goMux_mux_bufchan_buf[0] ? m1a85_goMux_mux_bufchan_buf :
                             m1a85_goMux_mux_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m1a85_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((m1a85_1_argbuf_r && m1a85_goMux_mux_bufchan_buf[0]))
        m1a85_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
      else if (((! m1a85_1_argbuf_r) && (! m1a85_goMux_mux_bufchan_buf[0])))
        m1a85_goMux_mux_bufchan_buf <= m1a85_goMux_mux_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (m2a86_1,Pointer_QTree_Bool) > (m2a86_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t m2a86_1_bufchan_d;
  logic m2a86_1_bufchan_r;
  assign m2a86_1_r = ((! m2a86_1_bufchan_d[0]) || m2a86_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m2a86_1_bufchan_d <= {16'd0, 1'd0};
    else if (m2a86_1_r) m2a86_1_bufchan_d <= m2a86_1_d;
  Pointer_QTree_Bool_t m2a86_1_bufchan_buf;
  assign m2a86_1_bufchan_r = (! m2a86_1_bufchan_buf[0]);
  assign m2a86_1_argbuf_d = (m2a86_1_bufchan_buf[0] ? m2a86_1_bufchan_buf :
                             m2a86_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m2a86_1_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((m2a86_1_argbuf_r && m2a86_1_bufchan_buf[0]))
        m2a86_1_bufchan_buf <= {16'd0, 1'd0};
      else if (((! m2a86_1_argbuf_r) && (! m2a86_1_bufchan_buf[0])))
        m2a86_1_bufchan_buf <= m2a86_1_bufchan_d;
  
  /* fork (Ty Pointer_QTree_Bool) : (m2a86_goMux_mux,Pointer_QTree_Bool) > [(m2a86_1,Pointer_QTree_Bool),
                                                                       (m2a86_2,Pointer_QTree_Bool)] */
  logic [1:0] m2a86_goMux_mux_emitted;
  logic [1:0] m2a86_goMux_mux_done;
  assign m2a86_1_d = {m2a86_goMux_mux_d[16:1],
                      (m2a86_goMux_mux_d[0] && (! m2a86_goMux_mux_emitted[0]))};
  assign m2a86_2_d = {m2a86_goMux_mux_d[16:1],
                      (m2a86_goMux_mux_d[0] && (! m2a86_goMux_mux_emitted[1]))};
  assign m2a86_goMux_mux_done = (m2a86_goMux_mux_emitted | ({m2a86_2_d[0],
                                                             m2a86_1_d[0]} & {m2a86_2_r,
                                                                              m2a86_1_r}));
  assign m2a86_goMux_mux_r = (& m2a86_goMux_mux_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m2a86_goMux_mux_emitted <= 2'd0;
    else
      m2a86_goMux_mux_emitted <= (m2a86_goMux_mux_r ? 2'd0 :
                                  m2a86_goMux_mux_done);
  
  /* buf (Ty Pointer_QTree_Bool) : (m2a8H_1,Pointer_QTree_Bool) > (m2a8H_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t m2a8H_1_bufchan_d;
  logic m2a8H_1_bufchan_r;
  assign m2a8H_1_r = ((! m2a8H_1_bufchan_d[0]) || m2a8H_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m2a8H_1_bufchan_d <= {16'd0, 1'd0};
    else if (m2a8H_1_r) m2a8H_1_bufchan_d <= m2a8H_1_d;
  Pointer_QTree_Bool_t m2a8H_1_bufchan_buf;
  assign m2a8H_1_bufchan_r = (! m2a8H_1_bufchan_buf[0]);
  assign m2a8H_1_argbuf_d = (m2a8H_1_bufchan_buf[0] ? m2a8H_1_bufchan_buf :
                             m2a8H_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m2a8H_1_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((m2a8H_1_argbuf_r && m2a8H_1_bufchan_buf[0]))
        m2a8H_1_bufchan_buf <= {16'd0, 1'd0};
      else if (((! m2a8H_1_argbuf_r) && (! m2a8H_1_bufchan_buf[0])))
        m2a8H_1_bufchan_buf <= m2a8H_1_bufchan_d;
  
  /* fork (Ty Pointer_QTree_Bool) : (m2a8H_goMux_mux,Pointer_QTree_Bool) > [(m2a8H_1,Pointer_QTree_Bool),
                                                                       (m2a8H_2,Pointer_QTree_Bool)] */
  logic [1:0] m2a8H_goMux_mux_emitted;
  logic [1:0] m2a8H_goMux_mux_done;
  assign m2a8H_1_d = {m2a8H_goMux_mux_d[16:1],
                      (m2a8H_goMux_mux_d[0] && (! m2a8H_goMux_mux_emitted[0]))};
  assign m2a8H_2_d = {m2a8H_goMux_mux_d[16:1],
                      (m2a8H_goMux_mux_d[0] && (! m2a8H_goMux_mux_emitted[1]))};
  assign m2a8H_goMux_mux_done = (m2a8H_goMux_mux_emitted | ({m2a8H_2_d[0],
                                                             m2a8H_1_d[0]} & {m2a8H_2_r,
                                                                              m2a8H_1_r}));
  assign m2a8H_goMux_mux_r = (& m2a8H_goMux_mux_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m2a8H_goMux_mux_emitted <= 2'd0;
    else
      m2a8H_goMux_mux_emitted <= (m2a8H_goMux_mux_r ? 2'd0 :
                                  m2a8H_goMux_mux_done);
  
  /* buf (Ty Pointer_QTree_Bool) : (m3a87_1,Pointer_QTree_Bool) > (m3a87_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t m3a87_1_bufchan_d;
  logic m3a87_1_bufchan_r;
  assign m3a87_1_r = ((! m3a87_1_bufchan_d[0]) || m3a87_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m3a87_1_bufchan_d <= {16'd0, 1'd0};
    else if (m3a87_1_r) m3a87_1_bufchan_d <= m3a87_1_d;
  Pointer_QTree_Bool_t m3a87_1_bufchan_buf;
  assign m3a87_1_bufchan_r = (! m3a87_1_bufchan_buf[0]);
  assign m3a87_1_argbuf_d = (m3a87_1_bufchan_buf[0] ? m3a87_1_bufchan_buf :
                             m3a87_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m3a87_1_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((m3a87_1_argbuf_r && m3a87_1_bufchan_buf[0]))
        m3a87_1_bufchan_buf <= {16'd0, 1'd0};
      else if (((! m3a87_1_argbuf_r) && (! m3a87_1_bufchan_buf[0])))
        m3a87_1_bufchan_buf <= m3a87_1_bufchan_d;
  
  /* fork (Ty Pointer_QTree_Bool) : (m3a87_goMux_mux,Pointer_QTree_Bool) > [(m3a87_1,Pointer_QTree_Bool),
                                                                       (m3a87_2,Pointer_QTree_Bool)] */
  logic [1:0] m3a87_goMux_mux_emitted;
  logic [1:0] m3a87_goMux_mux_done;
  assign m3a87_1_d = {m3a87_goMux_mux_d[16:1],
                      (m3a87_goMux_mux_d[0] && (! m3a87_goMux_mux_emitted[0]))};
  assign m3a87_2_d = {m3a87_goMux_mux_d[16:1],
                      (m3a87_goMux_mux_d[0] && (! m3a87_goMux_mux_emitted[1]))};
  assign m3a87_goMux_mux_done = (m3a87_goMux_mux_emitted | ({m3a87_2_d[0],
                                                             m3a87_1_d[0]} & {m3a87_2_r,
                                                                              m3a87_1_r}));
  assign m3a87_goMux_mux_r = (& m3a87_goMux_mux_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m3a87_goMux_mux_emitted <= 2'd0;
    else
      m3a87_goMux_mux_emitted <= (m3a87_goMux_mux_r ? 2'd0 :
                                  m3a87_goMux_mux_done);
  
  /* buf (Ty Pointer_QTree_Bool) : (m3a8I_1,Pointer_QTree_Bool) > (m3a8I_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t m3a8I_1_bufchan_d;
  logic m3a8I_1_bufchan_r;
  assign m3a8I_1_r = ((! m3a8I_1_bufchan_d[0]) || m3a8I_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m3a8I_1_bufchan_d <= {16'd0, 1'd0};
    else if (m3a8I_1_r) m3a8I_1_bufchan_d <= m3a8I_1_d;
  Pointer_QTree_Bool_t m3a8I_1_bufchan_buf;
  assign m3a8I_1_bufchan_r = (! m3a8I_1_bufchan_buf[0]);
  assign m3a8I_1_argbuf_d = (m3a8I_1_bufchan_buf[0] ? m3a8I_1_bufchan_buf :
                             m3a8I_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m3a8I_1_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((m3a8I_1_argbuf_r && m3a8I_1_bufchan_buf[0]))
        m3a8I_1_bufchan_buf <= {16'd0, 1'd0};
      else if (((! m3a8I_1_argbuf_r) && (! m3a8I_1_bufchan_buf[0])))
        m3a8I_1_bufchan_buf <= m3a8I_1_bufchan_d;
  
  /* fork (Ty Pointer_QTree_Bool) : (m3a8I_goMux_mux,Pointer_QTree_Bool) > [(m3a8I_1,Pointer_QTree_Bool),
                                                                       (m3a8I_2,Pointer_QTree_Bool)] */
  logic [1:0] m3a8I_goMux_mux_emitted;
  logic [1:0] m3a8I_goMux_mux_done;
  assign m3a8I_1_d = {m3a8I_goMux_mux_d[16:1],
                      (m3a8I_goMux_mux_d[0] && (! m3a8I_goMux_mux_emitted[0]))};
  assign m3a8I_2_d = {m3a8I_goMux_mux_d[16:1],
                      (m3a8I_goMux_mux_d[0] && (! m3a8I_goMux_mux_emitted[1]))};
  assign m3a8I_goMux_mux_done = (m3a8I_goMux_mux_emitted | ({m3a8I_2_d[0],
                                                             m3a8I_1_d[0]} & {m3a8I_2_r,
                                                                              m3a8I_1_r}));
  assign m3a8I_goMux_mux_r = (& m3a8I_goMux_mux_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m3a8I_goMux_mux_emitted <= 2'd0;
    else
      m3a8I_goMux_mux_emitted <= (m3a8I_goMux_mux_r ? 2'd0 :
                                  m3a8I_goMux_mux_done);
  
  /* buf (Ty Pointer_QTree_Bool) : (q1'a8n_3_destruct,Pointer_QTree_Bool) > (q1'a8n_3_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t \q1'a8n_3_destruct_bufchan_d ;
  logic \q1'a8n_3_destruct_bufchan_r ;
  assign \q1'a8n_3_destruct_r  = ((! \q1'a8n_3_destruct_bufchan_d [0]) || \q1'a8n_3_destruct_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \q1'a8n_3_destruct_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\q1'a8n_3_destruct_r )
        \q1'a8n_3_destruct_bufchan_d  <= \q1'a8n_3_destruct_d ;
  Pointer_QTree_Bool_t \q1'a8n_3_destruct_bufchan_buf ;
  assign \q1'a8n_3_destruct_bufchan_r  = (! \q1'a8n_3_destruct_bufchan_buf [0]);
  assign \q1'a8n_3_1_argbuf_d  = (\q1'a8n_3_destruct_bufchan_buf [0] ? \q1'a8n_3_destruct_bufchan_buf  :
                                  \q1'a8n_3_destruct_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \q1'a8n_3_destruct_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((\q1'a8n_3_1_argbuf_r  && \q1'a8n_3_destruct_bufchan_buf [0]))
        \q1'a8n_3_destruct_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! \q1'a8n_3_1_argbuf_r ) && (! \q1'a8n_3_destruct_bufchan_buf [0])))
        \q1'a8n_3_destruct_bufchan_buf  <= \q1'a8n_3_destruct_bufchan_d ;
  
  /* buf (Ty Pointer_MaskQTree) : (q1a88_3_destruct,Pointer_MaskQTree) > (q1a88_3_1_argbuf,Pointer_MaskQTree) */
  Pointer_MaskQTree_t q1a88_3_destruct_bufchan_d;
  logic q1a88_3_destruct_bufchan_r;
  assign q1a88_3_destruct_r = ((! q1a88_3_destruct_bufchan_d[0]) || q1a88_3_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q1a88_3_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q1a88_3_destruct_r)
        q1a88_3_destruct_bufchan_d <= q1a88_3_destruct_d;
  Pointer_MaskQTree_t q1a88_3_destruct_bufchan_buf;
  assign q1a88_3_destruct_bufchan_r = (! q1a88_3_destruct_bufchan_buf[0]);
  assign q1a88_3_1_argbuf_d = (q1a88_3_destruct_bufchan_buf[0] ? q1a88_3_destruct_bufchan_buf :
                               q1a88_3_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q1a88_3_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q1a88_3_1_argbuf_r && q1a88_3_destruct_bufchan_buf[0]))
        q1a88_3_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q1a88_3_1_argbuf_r) && (! q1a88_3_destruct_bufchan_buf[0])))
        q1a88_3_destruct_bufchan_buf <= q1a88_3_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (q1a8P_3_destruct,Pointer_QTree_Bool) > (q1a8P_3_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t q1a8P_3_destruct_bufchan_d;
  logic q1a8P_3_destruct_bufchan_r;
  assign q1a8P_3_destruct_r = ((! q1a8P_3_destruct_bufchan_d[0]) || q1a8P_3_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q1a8P_3_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q1a8P_3_destruct_r)
        q1a8P_3_destruct_bufchan_d <= q1a8P_3_destruct_d;
  Pointer_QTree_Bool_t q1a8P_3_destruct_bufchan_buf;
  assign q1a8P_3_destruct_bufchan_r = (! q1a8P_3_destruct_bufchan_buf[0]);
  assign q1a8P_3_1_argbuf_d = (q1a8P_3_destruct_bufchan_buf[0] ? q1a8P_3_destruct_bufchan_buf :
                               q1a8P_3_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q1a8P_3_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q1a8P_3_1_argbuf_r && q1a8P_3_destruct_bufchan_buf[0]))
        q1a8P_3_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q1a8P_3_1_argbuf_r) && (! q1a8P_3_destruct_bufchan_buf[0])))
        q1a8P_3_destruct_bufchan_buf <= q1a8P_3_destruct_bufchan_d;
  
  /* buf (Ty Pointer_MaskQTree) : (q1a8y_3_destruct,Pointer_MaskQTree) > (q1a8y_3_1_argbuf,Pointer_MaskQTree) */
  Pointer_MaskQTree_t q1a8y_3_destruct_bufchan_d;
  logic q1a8y_3_destruct_bufchan_r;
  assign q1a8y_3_destruct_r = ((! q1a8y_3_destruct_bufchan_d[0]) || q1a8y_3_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q1a8y_3_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q1a8y_3_destruct_r)
        q1a8y_3_destruct_bufchan_d <= q1a8y_3_destruct_d;
  Pointer_MaskQTree_t q1a8y_3_destruct_bufchan_buf;
  assign q1a8y_3_destruct_bufchan_r = (! q1a8y_3_destruct_bufchan_buf[0]);
  assign q1a8y_3_1_argbuf_d = (q1a8y_3_destruct_bufchan_buf[0] ? q1a8y_3_destruct_bufchan_buf :
                               q1a8y_3_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q1a8y_3_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q1a8y_3_1_argbuf_r && q1a8y_3_destruct_bufchan_buf[0]))
        q1a8y_3_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q1a8y_3_1_argbuf_r) && (! q1a8y_3_destruct_bufchan_buf[0])))
        q1a8y_3_destruct_bufchan_buf <= q1a8y_3_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (q2'a8o_2_destruct,Pointer_QTree_Bool) > (q2'a8o_2_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t \q2'a8o_2_destruct_bufchan_d ;
  logic \q2'a8o_2_destruct_bufchan_r ;
  assign \q2'a8o_2_destruct_r  = ((! \q2'a8o_2_destruct_bufchan_d [0]) || \q2'a8o_2_destruct_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \q2'a8o_2_destruct_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\q2'a8o_2_destruct_r )
        \q2'a8o_2_destruct_bufchan_d  <= \q2'a8o_2_destruct_d ;
  Pointer_QTree_Bool_t \q2'a8o_2_destruct_bufchan_buf ;
  assign \q2'a8o_2_destruct_bufchan_r  = (! \q2'a8o_2_destruct_bufchan_buf [0]);
  assign \q2'a8o_2_1_argbuf_d  = (\q2'a8o_2_destruct_bufchan_buf [0] ? \q2'a8o_2_destruct_bufchan_buf  :
                                  \q2'a8o_2_destruct_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \q2'a8o_2_destruct_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((\q2'a8o_2_1_argbuf_r  && \q2'a8o_2_destruct_bufchan_buf [0]))
        \q2'a8o_2_destruct_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! \q2'a8o_2_1_argbuf_r ) && (! \q2'a8o_2_destruct_bufchan_buf [0])))
        \q2'a8o_2_destruct_bufchan_buf  <= \q2'a8o_2_destruct_bufchan_d ;
  
  /* buf (Ty Pointer_MaskQTree) : (q2a89_2_destruct,Pointer_MaskQTree) > (q2a89_2_1_argbuf,Pointer_MaskQTree) */
  Pointer_MaskQTree_t q2a89_2_destruct_bufchan_d;
  logic q2a89_2_destruct_bufchan_r;
  assign q2a89_2_destruct_r = ((! q2a89_2_destruct_bufchan_d[0]) || q2a89_2_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q2a89_2_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q2a89_2_destruct_r)
        q2a89_2_destruct_bufchan_d <= q2a89_2_destruct_d;
  Pointer_MaskQTree_t q2a89_2_destruct_bufchan_buf;
  assign q2a89_2_destruct_bufchan_r = (! q2a89_2_destruct_bufchan_buf[0]);
  assign q2a89_2_1_argbuf_d = (q2a89_2_destruct_bufchan_buf[0] ? q2a89_2_destruct_bufchan_buf :
                               q2a89_2_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q2a89_2_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q2a89_2_1_argbuf_r && q2a89_2_destruct_bufchan_buf[0]))
        q2a89_2_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q2a89_2_1_argbuf_r) && (! q2a89_2_destruct_bufchan_buf[0])))
        q2a89_2_destruct_bufchan_buf <= q2a89_2_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (q2a8Q_2_destruct,Pointer_QTree_Bool) > (q2a8Q_2_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t q2a8Q_2_destruct_bufchan_d;
  logic q2a8Q_2_destruct_bufchan_r;
  assign q2a8Q_2_destruct_r = ((! q2a8Q_2_destruct_bufchan_d[0]) || q2a8Q_2_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q2a8Q_2_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q2a8Q_2_destruct_r)
        q2a8Q_2_destruct_bufchan_d <= q2a8Q_2_destruct_d;
  Pointer_QTree_Bool_t q2a8Q_2_destruct_bufchan_buf;
  assign q2a8Q_2_destruct_bufchan_r = (! q2a8Q_2_destruct_bufchan_buf[0]);
  assign q2a8Q_2_1_argbuf_d = (q2a8Q_2_destruct_bufchan_buf[0] ? q2a8Q_2_destruct_bufchan_buf :
                               q2a8Q_2_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q2a8Q_2_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q2a8Q_2_1_argbuf_r && q2a8Q_2_destruct_bufchan_buf[0]))
        q2a8Q_2_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q2a8Q_2_1_argbuf_r) && (! q2a8Q_2_destruct_bufchan_buf[0])))
        q2a8Q_2_destruct_bufchan_buf <= q2a8Q_2_destruct_bufchan_d;
  
  /* buf (Ty Pointer_MaskQTree) : (q2a8z_2_destruct,Pointer_MaskQTree) > (q2a8z_2_1_argbuf,Pointer_MaskQTree) */
  Pointer_MaskQTree_t q2a8z_2_destruct_bufchan_d;
  logic q2a8z_2_destruct_bufchan_r;
  assign q2a8z_2_destruct_r = ((! q2a8z_2_destruct_bufchan_d[0]) || q2a8z_2_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q2a8z_2_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q2a8z_2_destruct_r)
        q2a8z_2_destruct_bufchan_d <= q2a8z_2_destruct_d;
  Pointer_MaskQTree_t q2a8z_2_destruct_bufchan_buf;
  assign q2a8z_2_destruct_bufchan_r = (! q2a8z_2_destruct_bufchan_buf[0]);
  assign q2a8z_2_1_argbuf_d = (q2a8z_2_destruct_bufchan_buf[0] ? q2a8z_2_destruct_bufchan_buf :
                               q2a8z_2_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q2a8z_2_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q2a8z_2_1_argbuf_r && q2a8z_2_destruct_bufchan_buf[0]))
        q2a8z_2_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q2a8z_2_1_argbuf_r) && (! q2a8z_2_destruct_bufchan_buf[0])))
        q2a8z_2_destruct_bufchan_buf <= q2a8z_2_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (q3'a8p_1_destruct,Pointer_QTree_Bool) > (q3'a8p_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t \q3'a8p_1_destruct_bufchan_d ;
  logic \q3'a8p_1_destruct_bufchan_r ;
  assign \q3'a8p_1_destruct_r  = ((! \q3'a8p_1_destruct_bufchan_d [0]) || \q3'a8p_1_destruct_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \q3'a8p_1_destruct_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\q3'a8p_1_destruct_r )
        \q3'a8p_1_destruct_bufchan_d  <= \q3'a8p_1_destruct_d ;
  Pointer_QTree_Bool_t \q3'a8p_1_destruct_bufchan_buf ;
  assign \q3'a8p_1_destruct_bufchan_r  = (! \q3'a8p_1_destruct_bufchan_buf [0]);
  assign \q3'a8p_1_1_argbuf_d  = (\q3'a8p_1_destruct_bufchan_buf [0] ? \q3'a8p_1_destruct_bufchan_buf  :
                                  \q3'a8p_1_destruct_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \q3'a8p_1_destruct_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((\q3'a8p_1_1_argbuf_r  && \q3'a8p_1_destruct_bufchan_buf [0]))
        \q3'a8p_1_destruct_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! \q3'a8p_1_1_argbuf_r ) && (! \q3'a8p_1_destruct_bufchan_buf [0])))
        \q3'a8p_1_destruct_bufchan_buf  <= \q3'a8p_1_destruct_bufchan_d ;
  
  /* buf (Ty Pointer_MaskQTree) : (q3a8A_1_destruct,Pointer_MaskQTree) > (q3a8A_1_1_argbuf,Pointer_MaskQTree) */
  Pointer_MaskQTree_t q3a8A_1_destruct_bufchan_d;
  logic q3a8A_1_destruct_bufchan_r;
  assign q3a8A_1_destruct_r = ((! q3a8A_1_destruct_bufchan_d[0]) || q3a8A_1_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q3a8A_1_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q3a8A_1_destruct_r)
        q3a8A_1_destruct_bufchan_d <= q3a8A_1_destruct_d;
  Pointer_MaskQTree_t q3a8A_1_destruct_bufchan_buf;
  assign q3a8A_1_destruct_bufchan_r = (! q3a8A_1_destruct_bufchan_buf[0]);
  assign q3a8A_1_1_argbuf_d = (q3a8A_1_destruct_bufchan_buf[0] ? q3a8A_1_destruct_bufchan_buf :
                               q3a8A_1_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q3a8A_1_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q3a8A_1_1_argbuf_r && q3a8A_1_destruct_bufchan_buf[0]))
        q3a8A_1_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q3a8A_1_1_argbuf_r) && (! q3a8A_1_destruct_bufchan_buf[0])))
        q3a8A_1_destruct_bufchan_buf <= q3a8A_1_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (q3a8R_1_destruct,Pointer_QTree_Bool) > (q3a8R_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t q3a8R_1_destruct_bufchan_d;
  logic q3a8R_1_destruct_bufchan_r;
  assign q3a8R_1_destruct_r = ((! q3a8R_1_destruct_bufchan_d[0]) || q3a8R_1_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q3a8R_1_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q3a8R_1_destruct_r)
        q3a8R_1_destruct_bufchan_d <= q3a8R_1_destruct_d;
  Pointer_QTree_Bool_t q3a8R_1_destruct_bufchan_buf;
  assign q3a8R_1_destruct_bufchan_r = (! q3a8R_1_destruct_bufchan_buf[0]);
  assign q3a8R_1_1_argbuf_d = (q3a8R_1_destruct_bufchan_buf[0] ? q3a8R_1_destruct_bufchan_buf :
                               q3a8R_1_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q3a8R_1_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q3a8R_1_1_argbuf_r && q3a8R_1_destruct_bufchan_buf[0]))
        q3a8R_1_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q3a8R_1_1_argbuf_r) && (! q3a8R_1_destruct_bufchan_buf[0])))
        q3a8R_1_destruct_bufchan_buf <= q3a8R_1_destruct_bufchan_d;
  
  /* buf (Ty Pointer_MaskQTree) : (q3a8a_1_destruct,Pointer_MaskQTree) > (q3a8a_1_1_argbuf,Pointer_MaskQTree) */
  Pointer_MaskQTree_t q3a8a_1_destruct_bufchan_d;
  logic q3a8a_1_destruct_bufchan_r;
  assign q3a8a_1_destruct_r = ((! q3a8a_1_destruct_bufchan_d[0]) || q3a8a_1_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q3a8a_1_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q3a8a_1_destruct_r)
        q3a8a_1_destruct_bufchan_d <= q3a8a_1_destruct_d;
  Pointer_MaskQTree_t q3a8a_1_destruct_bufchan_buf;
  assign q3a8a_1_destruct_bufchan_r = (! q3a8a_1_destruct_bufchan_buf[0]);
  assign q3a8a_1_1_argbuf_d = (q3a8a_1_destruct_bufchan_buf[0] ? q3a8a_1_destruct_bufchan_buf :
                               q3a8a_1_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q3a8a_1_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q3a8a_1_1_argbuf_r && q3a8a_1_destruct_bufchan_buf[0]))
        q3a8a_1_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q3a8a_1_1_argbuf_r) && (! q3a8a_1_destruct_bufchan_buf[0])))
        q3a8a_1_destruct_bufchan_buf <= q3a8a_1_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (q4'a8x_1,Pointer_QTree_Bool) > (q4'a8x_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t \q4'a8x_1_bufchan_d ;
  logic \q4'a8x_1_bufchan_r ;
  assign \q4'a8x_1_r  = ((! \q4'a8x_1_bufchan_d [0]) || \q4'a8x_1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \q4'a8x_1_bufchan_d  <= {16'd0, 1'd0};
    else if (\q4'a8x_1_r ) \q4'a8x_1_bufchan_d  <= \q4'a8x_1_d ;
  Pointer_QTree_Bool_t \q4'a8x_1_bufchan_buf ;
  assign \q4'a8x_1_bufchan_r  = (! \q4'a8x_1_bufchan_buf [0]);
  assign \q4'a8x_1_argbuf_d  = (\q4'a8x_1_bufchan_buf [0] ? \q4'a8x_1_bufchan_buf  :
                                \q4'a8x_1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \q4'a8x_1_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((\q4'a8x_1_argbuf_r  && \q4'a8x_1_bufchan_buf [0]))
        \q4'a8x_1_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! \q4'a8x_1_argbuf_r ) && (! \q4'a8x_1_bufchan_buf [0])))
        \q4'a8x_1_bufchan_buf  <= \q4'a8x_1_bufchan_d ;
  
  /* fork (Ty Pointer_QTree_Bool) : (q4'a8x_goMux_mux,Pointer_QTree_Bool) > [(q4'a8x_1,Pointer_QTree_Bool),
                                                                        (q4'a8x_2,Pointer_QTree_Bool)] */
  logic [1:0] \q4'a8x_goMux_mux_emitted ;
  logic [1:0] \q4'a8x_goMux_mux_done ;
  assign \q4'a8x_1_d  = {\q4'a8x_goMux_mux_d [16:1],
                         (\q4'a8x_goMux_mux_d [0] && (! \q4'a8x_goMux_mux_emitted [0]))};
  assign \q4'a8x_2_d  = {\q4'a8x_goMux_mux_d [16:1],
                         (\q4'a8x_goMux_mux_d [0] && (! \q4'a8x_goMux_mux_emitted [1]))};
  assign \q4'a8x_goMux_mux_done  = (\q4'a8x_goMux_mux_emitted  | ({\q4'a8x_2_d [0],
                                                                   \q4'a8x_1_d [0]} & {\q4'a8x_2_r ,
                                                                                       \q4'a8x_1_r }));
  assign \q4'a8x_goMux_mux_r  = (& \q4'a8x_goMux_mux_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \q4'a8x_goMux_mux_emitted  <= 2'd0;
    else
      \q4'a8x_goMux_mux_emitted  <= (\q4'a8x_goMux_mux_r  ? 2'd0 :
                                     \q4'a8x_goMux_mux_done );
  
  /* buf (Ty Pointer_MaskQTree) : (q4a8w_goMux_mux,Pointer_MaskQTree) > (q4a8w_1_argbuf,Pointer_MaskQTree) */
  Pointer_MaskQTree_t q4a8w_goMux_mux_bufchan_d;
  logic q4a8w_goMux_mux_bufchan_r;
  assign q4a8w_goMux_mux_r = ((! q4a8w_goMux_mux_bufchan_d[0]) || q4a8w_goMux_mux_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q4a8w_goMux_mux_bufchan_d <= {16'd0, 1'd0};
    else
      if (q4a8w_goMux_mux_r)
        q4a8w_goMux_mux_bufchan_d <= q4a8w_goMux_mux_d;
  Pointer_MaskQTree_t q4a8w_goMux_mux_bufchan_buf;
  assign q4a8w_goMux_mux_bufchan_r = (! q4a8w_goMux_mux_bufchan_buf[0]);
  assign q4a8w_1_argbuf_d = (q4a8w_goMux_mux_bufchan_buf[0] ? q4a8w_goMux_mux_bufchan_buf :
                             q4a8w_goMux_mux_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q4a8w_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q4a8w_1_argbuf_r && q4a8w_goMux_mux_bufchan_buf[0]))
        q4a8w_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q4a8w_1_argbuf_r) && (! q4a8w_goMux_mux_bufchan_buf[0])))
        q4a8w_goMux_mux_bufchan_buf <= q4a8w_goMux_mux_bufchan_d;
  
  /* buf (Ty CTf'''''''''_f'''''''''_Bool) : (readPointer_CTf'''''''''_f'''''''''_Boolscfarg_0_2_1_argbuf,CTf'''''''''_f'''''''''_Bool) > (readPointer_CTf'''''''''_f'''''''''_Boolscfarg_0_2_1_argbuf_rwb,CTf'''''''''_f'''''''''_Bool) */
  \CTf'''''''''_f'''''''''_Bool_t  \readPointer_CTf'''''''''_f'''''''''_Boolscfarg_0_2_1_argbuf_bufchan_d ;
  logic \readPointer_CTf'''''''''_f'''''''''_Boolscfarg_0_2_1_argbuf_bufchan_r ;
  assign \readPointer_CTf'''''''''_f'''''''''_Boolscfarg_0_2_1_argbuf_r  = ((! \readPointer_CTf'''''''''_f'''''''''_Boolscfarg_0_2_1_argbuf_bufchan_d [0]) || \readPointer_CTf'''''''''_f'''''''''_Boolscfarg_0_2_1_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \readPointer_CTf'''''''''_f'''''''''_Boolscfarg_0_2_1_argbuf_bufchan_d  <= {115'd0,
                                                                                  1'd0};
    else
      if (\readPointer_CTf'''''''''_f'''''''''_Boolscfarg_0_2_1_argbuf_r )
        \readPointer_CTf'''''''''_f'''''''''_Boolscfarg_0_2_1_argbuf_bufchan_d  <= \readPointer_CTf'''''''''_f'''''''''_Boolscfarg_0_2_1_argbuf_d ;
  \CTf'''''''''_f'''''''''_Bool_t  \readPointer_CTf'''''''''_f'''''''''_Boolscfarg_0_2_1_argbuf_bufchan_buf ;
  assign \readPointer_CTf'''''''''_f'''''''''_Boolscfarg_0_2_1_argbuf_bufchan_r  = (! \readPointer_CTf'''''''''_f'''''''''_Boolscfarg_0_2_1_argbuf_bufchan_buf [0]);
  assign \readPointer_CTf'''''''''_f'''''''''_Boolscfarg_0_2_1_argbuf_rwb_d  = (\readPointer_CTf'''''''''_f'''''''''_Boolscfarg_0_2_1_argbuf_bufchan_buf [0] ? \readPointer_CTf'''''''''_f'''''''''_Boolscfarg_0_2_1_argbuf_bufchan_buf  :
                                                                                \readPointer_CTf'''''''''_f'''''''''_Boolscfarg_0_2_1_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \readPointer_CTf'''''''''_f'''''''''_Boolscfarg_0_2_1_argbuf_bufchan_buf  <= {115'd0,
                                                                                    1'd0};
    else
      if ((\readPointer_CTf'''''''''_f'''''''''_Boolscfarg_0_2_1_argbuf_rwb_r  && \readPointer_CTf'''''''''_f'''''''''_Boolscfarg_0_2_1_argbuf_bufchan_buf [0]))
        \readPointer_CTf'''''''''_f'''''''''_Boolscfarg_0_2_1_argbuf_bufchan_buf  <= {115'd0,
                                                                                      1'd0};
      else if (((! \readPointer_CTf'''''''''_f'''''''''_Boolscfarg_0_2_1_argbuf_rwb_r ) && (! \readPointer_CTf'''''''''_f'''''''''_Boolscfarg_0_2_1_argbuf_bufchan_buf [0])))
        \readPointer_CTf'''''''''_f'''''''''_Boolscfarg_0_2_1_argbuf_bufchan_buf  <= \readPointer_CTf'''''''''_f'''''''''_Boolscfarg_0_2_1_argbuf_bufchan_d ;
  
  /* fork (Ty CTf'''''''''_f'''''''''_Bool) : (readPointer_CTf'''''''''_f'''''''''_Boolscfarg_0_2_1_argbuf_rwb,CTf'''''''''_f'''''''''_Bool) > [(lizzieLet53_1,CTf'''''''''_f'''''''''_Bool),
                                                                                                                                           (lizzieLet53_2,CTf'''''''''_f'''''''''_Bool),
                                                                                                                                           (lizzieLet53_3,CTf'''''''''_f'''''''''_Bool),
                                                                                                                                           (lizzieLet53_4,CTf'''''''''_f'''''''''_Bool)] */
  logic [3:0] \readPointer_CTf'''''''''_f'''''''''_Boolscfarg_0_2_1_argbuf_rwb_emitted ;
  logic [3:0] \readPointer_CTf'''''''''_f'''''''''_Boolscfarg_0_2_1_argbuf_rwb_done ;
  assign lizzieLet53_1_d = {\readPointer_CTf'''''''''_f'''''''''_Boolscfarg_0_2_1_argbuf_rwb_d [115:1],
                            (\readPointer_CTf'''''''''_f'''''''''_Boolscfarg_0_2_1_argbuf_rwb_d [0] && (! \readPointer_CTf'''''''''_f'''''''''_Boolscfarg_0_2_1_argbuf_rwb_emitted [0]))};
  assign lizzieLet53_2_d = {\readPointer_CTf'''''''''_f'''''''''_Boolscfarg_0_2_1_argbuf_rwb_d [115:1],
                            (\readPointer_CTf'''''''''_f'''''''''_Boolscfarg_0_2_1_argbuf_rwb_d [0] && (! \readPointer_CTf'''''''''_f'''''''''_Boolscfarg_0_2_1_argbuf_rwb_emitted [1]))};
  assign lizzieLet53_3_d = {\readPointer_CTf'''''''''_f'''''''''_Boolscfarg_0_2_1_argbuf_rwb_d [115:1],
                            (\readPointer_CTf'''''''''_f'''''''''_Boolscfarg_0_2_1_argbuf_rwb_d [0] && (! \readPointer_CTf'''''''''_f'''''''''_Boolscfarg_0_2_1_argbuf_rwb_emitted [2]))};
  assign lizzieLet53_4_d = {\readPointer_CTf'''''''''_f'''''''''_Boolscfarg_0_2_1_argbuf_rwb_d [115:1],
                            (\readPointer_CTf'''''''''_f'''''''''_Boolscfarg_0_2_1_argbuf_rwb_d [0] && (! \readPointer_CTf'''''''''_f'''''''''_Boolscfarg_0_2_1_argbuf_rwb_emitted [3]))};
  assign \readPointer_CTf'''''''''_f'''''''''_Boolscfarg_0_2_1_argbuf_rwb_done  = (\readPointer_CTf'''''''''_f'''''''''_Boolscfarg_0_2_1_argbuf_rwb_emitted  | ({lizzieLet53_4_d[0],
                                                                                                                                                                 lizzieLet53_3_d[0],
                                                                                                                                                                 lizzieLet53_2_d[0],
                                                                                                                                                                 lizzieLet53_1_d[0]} & {lizzieLet53_4_r,
                                                                                                                                                                                        lizzieLet53_3_r,
                                                                                                                                                                                        lizzieLet53_2_r,
                                                                                                                                                                                        lizzieLet53_1_r}));
  assign \readPointer_CTf'''''''''_f'''''''''_Boolscfarg_0_2_1_argbuf_rwb_r  = (& \readPointer_CTf'''''''''_f'''''''''_Boolscfarg_0_2_1_argbuf_rwb_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \readPointer_CTf'''''''''_f'''''''''_Boolscfarg_0_2_1_argbuf_rwb_emitted  <= 4'd0;
    else
      \readPointer_CTf'''''''''_f'''''''''_Boolscfarg_0_2_1_argbuf_rwb_emitted  <= (\readPointer_CTf'''''''''_f'''''''''_Boolscfarg_0_2_1_argbuf_rwb_r  ? 4'd0 :
                                                                                    \readPointer_CTf'''''''''_f'''''''''_Boolscfarg_0_2_1_argbuf_rwb_done );
  
  /* buf (Ty CTf') : (readPointer_CTf'scfarg_0_1_1_argbuf,CTf') > (readPointer_CTf'scfarg_0_1_1_argbuf_rwb,CTf') */
  \CTf'_t  \readPointer_CTf'scfarg_0_1_1_argbuf_bufchan_d ;
  logic \readPointer_CTf'scfarg_0_1_1_argbuf_bufchan_r ;
  assign \readPointer_CTf'scfarg_0_1_1_argbuf_r  = ((! \readPointer_CTf'scfarg_0_1_1_argbuf_bufchan_d [0]) || \readPointer_CTf'scfarg_0_1_1_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \readPointer_CTf'scfarg_0_1_1_argbuf_bufchan_d  <= {115'd0, 1'd0};
    else
      if (\readPointer_CTf'scfarg_0_1_1_argbuf_r )
        \readPointer_CTf'scfarg_0_1_1_argbuf_bufchan_d  <= \readPointer_CTf'scfarg_0_1_1_argbuf_d ;
  \CTf'_t  \readPointer_CTf'scfarg_0_1_1_argbuf_bufchan_buf ;
  assign \readPointer_CTf'scfarg_0_1_1_argbuf_bufchan_r  = (! \readPointer_CTf'scfarg_0_1_1_argbuf_bufchan_buf [0]);
  assign \readPointer_CTf'scfarg_0_1_1_argbuf_rwb_d  = (\readPointer_CTf'scfarg_0_1_1_argbuf_bufchan_buf [0] ? \readPointer_CTf'scfarg_0_1_1_argbuf_bufchan_buf  :
                                                        \readPointer_CTf'scfarg_0_1_1_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \readPointer_CTf'scfarg_0_1_1_argbuf_bufchan_buf  <= {115'd0,
                                                            1'd0};
    else
      if ((\readPointer_CTf'scfarg_0_1_1_argbuf_rwb_r  && \readPointer_CTf'scfarg_0_1_1_argbuf_bufchan_buf [0]))
        \readPointer_CTf'scfarg_0_1_1_argbuf_bufchan_buf  <= {115'd0,
                                                              1'd0};
      else if (((! \readPointer_CTf'scfarg_0_1_1_argbuf_rwb_r ) && (! \readPointer_CTf'scfarg_0_1_1_argbuf_bufchan_buf [0])))
        \readPointer_CTf'scfarg_0_1_1_argbuf_bufchan_buf  <= \readPointer_CTf'scfarg_0_1_1_argbuf_bufchan_d ;
  
  /* fork (Ty CTf') : (readPointer_CTf'scfarg_0_1_1_argbuf_rwb,CTf') > [(lizzieLet48_1,CTf'),
                                                                   (lizzieLet48_2,CTf'),
                                                                   (lizzieLet48_3,CTf'),
                                                                   (lizzieLet48_4,CTf')] */
  logic [3:0] \readPointer_CTf'scfarg_0_1_1_argbuf_rwb_emitted ;
  logic [3:0] \readPointer_CTf'scfarg_0_1_1_argbuf_rwb_done ;
  assign lizzieLet48_1_d = {\readPointer_CTf'scfarg_0_1_1_argbuf_rwb_d [115:1],
                            (\readPointer_CTf'scfarg_0_1_1_argbuf_rwb_d [0] && (! \readPointer_CTf'scfarg_0_1_1_argbuf_rwb_emitted [0]))};
  assign lizzieLet48_2_d = {\readPointer_CTf'scfarg_0_1_1_argbuf_rwb_d [115:1],
                            (\readPointer_CTf'scfarg_0_1_1_argbuf_rwb_d [0] && (! \readPointer_CTf'scfarg_0_1_1_argbuf_rwb_emitted [1]))};
  assign lizzieLet48_3_d = {\readPointer_CTf'scfarg_0_1_1_argbuf_rwb_d [115:1],
                            (\readPointer_CTf'scfarg_0_1_1_argbuf_rwb_d [0] && (! \readPointer_CTf'scfarg_0_1_1_argbuf_rwb_emitted [2]))};
  assign lizzieLet48_4_d = {\readPointer_CTf'scfarg_0_1_1_argbuf_rwb_d [115:1],
                            (\readPointer_CTf'scfarg_0_1_1_argbuf_rwb_d [0] && (! \readPointer_CTf'scfarg_0_1_1_argbuf_rwb_emitted [3]))};
  assign \readPointer_CTf'scfarg_0_1_1_argbuf_rwb_done  = (\readPointer_CTf'scfarg_0_1_1_argbuf_rwb_emitted  | ({lizzieLet48_4_d[0],
                                                                                                                 lizzieLet48_3_d[0],
                                                                                                                 lizzieLet48_2_d[0],
                                                                                                                 lizzieLet48_1_d[0]} & {lizzieLet48_4_r,
                                                                                                                                        lizzieLet48_3_r,
                                                                                                                                        lizzieLet48_2_r,
                                                                                                                                        lizzieLet48_1_r}));
  assign \readPointer_CTf'scfarg_0_1_1_argbuf_rwb_r  = (& \readPointer_CTf'scfarg_0_1_1_argbuf_rwb_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \readPointer_CTf'scfarg_0_1_1_argbuf_rwb_emitted  <= 4'd0;
    else
      \readPointer_CTf'scfarg_0_1_1_argbuf_rwb_emitted  <= (\readPointer_CTf'scfarg_0_1_1_argbuf_rwb_r  ? 4'd0 :
                                                            \readPointer_CTf'scfarg_0_1_1_argbuf_rwb_done );
  
  /* buf (Ty CTf) : (readPointer_CTfscfarg_0_1_argbuf,CTf) > (readPointer_CTfscfarg_0_1_argbuf_rwb,CTf) */
  CTf_t readPointer_CTfscfarg_0_1_argbuf_bufchan_d;
  logic readPointer_CTfscfarg_0_1_argbuf_bufchan_r;
  assign readPointer_CTfscfarg_0_1_argbuf_r = ((! readPointer_CTfscfarg_0_1_argbuf_bufchan_d[0]) || readPointer_CTfscfarg_0_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_CTfscfarg_0_1_argbuf_bufchan_d <= {163'd0, 1'd0};
    else
      if (readPointer_CTfscfarg_0_1_argbuf_r)
        readPointer_CTfscfarg_0_1_argbuf_bufchan_d <= readPointer_CTfscfarg_0_1_argbuf_d;
  CTf_t readPointer_CTfscfarg_0_1_argbuf_bufchan_buf;
  assign readPointer_CTfscfarg_0_1_argbuf_bufchan_r = (! readPointer_CTfscfarg_0_1_argbuf_bufchan_buf[0]);
  assign readPointer_CTfscfarg_0_1_argbuf_rwb_d = (readPointer_CTfscfarg_0_1_argbuf_bufchan_buf[0] ? readPointer_CTfscfarg_0_1_argbuf_bufchan_buf :
                                                   readPointer_CTfscfarg_0_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_CTfscfarg_0_1_argbuf_bufchan_buf <= {163'd0, 1'd0};
    else
      if ((readPointer_CTfscfarg_0_1_argbuf_rwb_r && readPointer_CTfscfarg_0_1_argbuf_bufchan_buf[0]))
        readPointer_CTfscfarg_0_1_argbuf_bufchan_buf <= {163'd0, 1'd0};
      else if (((! readPointer_CTfscfarg_0_1_argbuf_rwb_r) && (! readPointer_CTfscfarg_0_1_argbuf_bufchan_buf[0])))
        readPointer_CTfscfarg_0_1_argbuf_bufchan_buf <= readPointer_CTfscfarg_0_1_argbuf_bufchan_d;
  
  /* fork (Ty CTf) : (readPointer_CTfscfarg_0_1_argbuf_rwb,CTf) > [(lizzieLet43_1,CTf),
                                                              (lizzieLet43_2,CTf),
                                                              (lizzieLet43_3,CTf),
                                                              (lizzieLet43_4,CTf)] */
  logic [3:0] readPointer_CTfscfarg_0_1_argbuf_rwb_emitted;
  logic [3:0] readPointer_CTfscfarg_0_1_argbuf_rwb_done;
  assign lizzieLet43_1_d = {readPointer_CTfscfarg_0_1_argbuf_rwb_d[163:1],
                            (readPointer_CTfscfarg_0_1_argbuf_rwb_d[0] && (! readPointer_CTfscfarg_0_1_argbuf_rwb_emitted[0]))};
  assign lizzieLet43_2_d = {readPointer_CTfscfarg_0_1_argbuf_rwb_d[163:1],
                            (readPointer_CTfscfarg_0_1_argbuf_rwb_d[0] && (! readPointer_CTfscfarg_0_1_argbuf_rwb_emitted[1]))};
  assign lizzieLet43_3_d = {readPointer_CTfscfarg_0_1_argbuf_rwb_d[163:1],
                            (readPointer_CTfscfarg_0_1_argbuf_rwb_d[0] && (! readPointer_CTfscfarg_0_1_argbuf_rwb_emitted[2]))};
  assign lizzieLet43_4_d = {readPointer_CTfscfarg_0_1_argbuf_rwb_d[163:1],
                            (readPointer_CTfscfarg_0_1_argbuf_rwb_d[0] && (! readPointer_CTfscfarg_0_1_argbuf_rwb_emitted[3]))};
  assign readPointer_CTfscfarg_0_1_argbuf_rwb_done = (readPointer_CTfscfarg_0_1_argbuf_rwb_emitted | ({lizzieLet43_4_d[0],
                                                                                                       lizzieLet43_3_d[0],
                                                                                                       lizzieLet43_2_d[0],
                                                                                                       lizzieLet43_1_d[0]} & {lizzieLet43_4_r,
                                                                                                                              lizzieLet43_3_r,
                                                                                                                              lizzieLet43_2_r,
                                                                                                                              lizzieLet43_1_r}));
  assign readPointer_CTfscfarg_0_1_argbuf_rwb_r = (& readPointer_CTfscfarg_0_1_argbuf_rwb_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_CTfscfarg_0_1_argbuf_rwb_emitted <= 4'd0;
    else
      readPointer_CTfscfarg_0_1_argbuf_rwb_emitted <= (readPointer_CTfscfarg_0_1_argbuf_rwb_r ? 4'd0 :
                                                       readPointer_CTfscfarg_0_1_argbuf_rwb_done);
  
  /* buf (Ty MaskQTree) : (readPointer_MaskQTreem1a85_1_argbuf,MaskQTree) > (readPointer_MaskQTreem1a85_1_argbuf_rwb,MaskQTree) */
  MaskQTree_t readPointer_MaskQTreem1a85_1_argbuf_bufchan_d;
  logic readPointer_MaskQTreem1a85_1_argbuf_bufchan_r;
  assign readPointer_MaskQTreem1a85_1_argbuf_r = ((! readPointer_MaskQTreem1a85_1_argbuf_bufchan_d[0]) || readPointer_MaskQTreem1a85_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_MaskQTreem1a85_1_argbuf_bufchan_d <= {66'd0, 1'd0};
    else
      if (readPointer_MaskQTreem1a85_1_argbuf_r)
        readPointer_MaskQTreem1a85_1_argbuf_bufchan_d <= readPointer_MaskQTreem1a85_1_argbuf_d;
  MaskQTree_t readPointer_MaskQTreem1a85_1_argbuf_bufchan_buf;
  assign readPointer_MaskQTreem1a85_1_argbuf_bufchan_r = (! readPointer_MaskQTreem1a85_1_argbuf_bufchan_buf[0]);
  assign readPointer_MaskQTreem1a85_1_argbuf_rwb_d = (readPointer_MaskQTreem1a85_1_argbuf_bufchan_buf[0] ? readPointer_MaskQTreem1a85_1_argbuf_bufchan_buf :
                                                      readPointer_MaskQTreem1a85_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_MaskQTreem1a85_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((readPointer_MaskQTreem1a85_1_argbuf_rwb_r && readPointer_MaskQTreem1a85_1_argbuf_bufchan_buf[0]))
        readPointer_MaskQTreem1a85_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
      else if (((! readPointer_MaskQTreem1a85_1_argbuf_rwb_r) && (! readPointer_MaskQTreem1a85_1_argbuf_bufchan_buf[0])))
        readPointer_MaskQTreem1a85_1_argbuf_bufchan_buf <= readPointer_MaskQTreem1a85_1_argbuf_bufchan_d;
  
  /* fork (Ty MaskQTree) : (readPointer_MaskQTreem1a85_1_argbuf_rwb,MaskQTree) > [(lizzieLet0_1,MaskQTree),
                                                                             (lizzieLet0_2,MaskQTree),
                                                                             (lizzieLet0_3,MaskQTree),
                                                                             (lizzieLet0_4,MaskQTree),
                                                                             (lizzieLet0_5,MaskQTree),
                                                                             (lizzieLet0_6,MaskQTree),
                                                                             (lizzieLet0_7,MaskQTree),
                                                                             (lizzieLet0_8,MaskQTree)] */
  logic [7:0] readPointer_MaskQTreem1a85_1_argbuf_rwb_emitted;
  logic [7:0] readPointer_MaskQTreem1a85_1_argbuf_rwb_done;
  assign lizzieLet0_1_d = {readPointer_MaskQTreem1a85_1_argbuf_rwb_d[66:1],
                           (readPointer_MaskQTreem1a85_1_argbuf_rwb_d[0] && (! readPointer_MaskQTreem1a85_1_argbuf_rwb_emitted[0]))};
  assign lizzieLet0_2_d = {readPointer_MaskQTreem1a85_1_argbuf_rwb_d[66:1],
                           (readPointer_MaskQTreem1a85_1_argbuf_rwb_d[0] && (! readPointer_MaskQTreem1a85_1_argbuf_rwb_emitted[1]))};
  assign lizzieLet0_3_d = {readPointer_MaskQTreem1a85_1_argbuf_rwb_d[66:1],
                           (readPointer_MaskQTreem1a85_1_argbuf_rwb_d[0] && (! readPointer_MaskQTreem1a85_1_argbuf_rwb_emitted[2]))};
  assign lizzieLet0_4_d = {readPointer_MaskQTreem1a85_1_argbuf_rwb_d[66:1],
                           (readPointer_MaskQTreem1a85_1_argbuf_rwb_d[0] && (! readPointer_MaskQTreem1a85_1_argbuf_rwb_emitted[3]))};
  assign lizzieLet0_5_d = {readPointer_MaskQTreem1a85_1_argbuf_rwb_d[66:1],
                           (readPointer_MaskQTreem1a85_1_argbuf_rwb_d[0] && (! readPointer_MaskQTreem1a85_1_argbuf_rwb_emitted[4]))};
  assign lizzieLet0_6_d = {readPointer_MaskQTreem1a85_1_argbuf_rwb_d[66:1],
                           (readPointer_MaskQTreem1a85_1_argbuf_rwb_d[0] && (! readPointer_MaskQTreem1a85_1_argbuf_rwb_emitted[5]))};
  assign lizzieLet0_7_d = {readPointer_MaskQTreem1a85_1_argbuf_rwb_d[66:1],
                           (readPointer_MaskQTreem1a85_1_argbuf_rwb_d[0] && (! readPointer_MaskQTreem1a85_1_argbuf_rwb_emitted[6]))};
  assign lizzieLet0_8_d = {readPointer_MaskQTreem1a85_1_argbuf_rwb_d[66:1],
                           (readPointer_MaskQTreem1a85_1_argbuf_rwb_d[0] && (! readPointer_MaskQTreem1a85_1_argbuf_rwb_emitted[7]))};
  assign readPointer_MaskQTreem1a85_1_argbuf_rwb_done = (readPointer_MaskQTreem1a85_1_argbuf_rwb_emitted | ({lizzieLet0_8_d[0],
                                                                                                             lizzieLet0_7_d[0],
                                                                                                             lizzieLet0_6_d[0],
                                                                                                             lizzieLet0_5_d[0],
                                                                                                             lizzieLet0_4_d[0],
                                                                                                             lizzieLet0_3_d[0],
                                                                                                             lizzieLet0_2_d[0],
                                                                                                             lizzieLet0_1_d[0]} & {lizzieLet0_8_r,
                                                                                                                                   lizzieLet0_7_r,
                                                                                                                                   lizzieLet0_6_r,
                                                                                                                                   lizzieLet0_5_r,
                                                                                                                                   lizzieLet0_4_r,
                                                                                                                                   lizzieLet0_3_r,
                                                                                                                                   lizzieLet0_2_r,
                                                                                                                                   lizzieLet0_1_r}));
  assign readPointer_MaskQTreem1a85_1_argbuf_rwb_r = (& readPointer_MaskQTreem1a85_1_argbuf_rwb_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_MaskQTreem1a85_1_argbuf_rwb_emitted <= 8'd0;
    else
      readPointer_MaskQTreem1a85_1_argbuf_rwb_emitted <= (readPointer_MaskQTreem1a85_1_argbuf_rwb_r ? 8'd0 :
                                                          readPointer_MaskQTreem1a85_1_argbuf_rwb_done);
  
  /* buf (Ty MaskQTree) : (readPointer_MaskQTreeq4a8w_1_argbuf,MaskQTree) > (readPointer_MaskQTreeq4a8w_1_argbuf_rwb,MaskQTree) */
  MaskQTree_t readPointer_MaskQTreeq4a8w_1_argbuf_bufchan_d;
  logic readPointer_MaskQTreeq4a8w_1_argbuf_bufchan_r;
  assign readPointer_MaskQTreeq4a8w_1_argbuf_r = ((! readPointer_MaskQTreeq4a8w_1_argbuf_bufchan_d[0]) || readPointer_MaskQTreeq4a8w_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_MaskQTreeq4a8w_1_argbuf_bufchan_d <= {66'd0, 1'd0};
    else
      if (readPointer_MaskQTreeq4a8w_1_argbuf_r)
        readPointer_MaskQTreeq4a8w_1_argbuf_bufchan_d <= readPointer_MaskQTreeq4a8w_1_argbuf_d;
  MaskQTree_t readPointer_MaskQTreeq4a8w_1_argbuf_bufchan_buf;
  assign readPointer_MaskQTreeq4a8w_1_argbuf_bufchan_r = (! readPointer_MaskQTreeq4a8w_1_argbuf_bufchan_buf[0]);
  assign readPointer_MaskQTreeq4a8w_1_argbuf_rwb_d = (readPointer_MaskQTreeq4a8w_1_argbuf_bufchan_buf[0] ? readPointer_MaskQTreeq4a8w_1_argbuf_bufchan_buf :
                                                      readPointer_MaskQTreeq4a8w_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_MaskQTreeq4a8w_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((readPointer_MaskQTreeq4a8w_1_argbuf_rwb_r && readPointer_MaskQTreeq4a8w_1_argbuf_bufchan_buf[0]))
        readPointer_MaskQTreeq4a8w_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
      else if (((! readPointer_MaskQTreeq4a8w_1_argbuf_rwb_r) && (! readPointer_MaskQTreeq4a8w_1_argbuf_bufchan_buf[0])))
        readPointer_MaskQTreeq4a8w_1_argbuf_bufchan_buf <= readPointer_MaskQTreeq4a8w_1_argbuf_bufchan_d;
  
  /* fork (Ty MaskQTree) : (readPointer_MaskQTreeq4a8w_1_argbuf_rwb,MaskQTree) > [(lizzieLet32_1,MaskQTree),
                                                                             (lizzieLet32_2,MaskQTree),
                                                                             (lizzieLet32_3,MaskQTree),
                                                                             (lizzieLet32_4,MaskQTree),
                                                                             (lizzieLet32_5,MaskQTree),
                                                                             (lizzieLet32_6,MaskQTree)] */
  logic [5:0] readPointer_MaskQTreeq4a8w_1_argbuf_rwb_emitted;
  logic [5:0] readPointer_MaskQTreeq4a8w_1_argbuf_rwb_done;
  assign lizzieLet32_1_d = {readPointer_MaskQTreeq4a8w_1_argbuf_rwb_d[66:1],
                            (readPointer_MaskQTreeq4a8w_1_argbuf_rwb_d[0] && (! readPointer_MaskQTreeq4a8w_1_argbuf_rwb_emitted[0]))};
  assign lizzieLet32_2_d = {readPointer_MaskQTreeq4a8w_1_argbuf_rwb_d[66:1],
                            (readPointer_MaskQTreeq4a8w_1_argbuf_rwb_d[0] && (! readPointer_MaskQTreeq4a8w_1_argbuf_rwb_emitted[1]))};
  assign lizzieLet32_3_d = {readPointer_MaskQTreeq4a8w_1_argbuf_rwb_d[66:1],
                            (readPointer_MaskQTreeq4a8w_1_argbuf_rwb_d[0] && (! readPointer_MaskQTreeq4a8w_1_argbuf_rwb_emitted[2]))};
  assign lizzieLet32_4_d = {readPointer_MaskQTreeq4a8w_1_argbuf_rwb_d[66:1],
                            (readPointer_MaskQTreeq4a8w_1_argbuf_rwb_d[0] && (! readPointer_MaskQTreeq4a8w_1_argbuf_rwb_emitted[3]))};
  assign lizzieLet32_5_d = {readPointer_MaskQTreeq4a8w_1_argbuf_rwb_d[66:1],
                            (readPointer_MaskQTreeq4a8w_1_argbuf_rwb_d[0] && (! readPointer_MaskQTreeq4a8w_1_argbuf_rwb_emitted[4]))};
  assign lizzieLet32_6_d = {readPointer_MaskQTreeq4a8w_1_argbuf_rwb_d[66:1],
                            (readPointer_MaskQTreeq4a8w_1_argbuf_rwb_d[0] && (! readPointer_MaskQTreeq4a8w_1_argbuf_rwb_emitted[5]))};
  assign readPointer_MaskQTreeq4a8w_1_argbuf_rwb_done = (readPointer_MaskQTreeq4a8w_1_argbuf_rwb_emitted | ({lizzieLet32_6_d[0],
                                                                                                             lizzieLet32_5_d[0],
                                                                                                             lizzieLet32_4_d[0],
                                                                                                             lizzieLet32_3_d[0],
                                                                                                             lizzieLet32_2_d[0],
                                                                                                             lizzieLet32_1_d[0]} & {lizzieLet32_6_r,
                                                                                                                                    lizzieLet32_5_r,
                                                                                                                                    lizzieLet32_4_r,
                                                                                                                                    lizzieLet32_3_r,
                                                                                                                                    lizzieLet32_2_r,
                                                                                                                                    lizzieLet32_1_r}));
  assign readPointer_MaskQTreeq4a8w_1_argbuf_rwb_r = (& readPointer_MaskQTreeq4a8w_1_argbuf_rwb_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_MaskQTreeq4a8w_1_argbuf_rwb_emitted <= 6'd0;
    else
      readPointer_MaskQTreeq4a8w_1_argbuf_rwb_emitted <= (readPointer_MaskQTreeq4a8w_1_argbuf_rwb_r ? 6'd0 :
                                                          readPointer_MaskQTreeq4a8w_1_argbuf_rwb_done);
  
  /* buf (Ty QTree_Bool) : (readPointer_QTree_Boolm2a86_1_argbuf,QTree_Bool) > (readPointer_QTree_Boolm2a86_1_argbuf_rwb,QTree_Bool) */
  QTree_Bool_t readPointer_QTree_Boolm2a86_1_argbuf_bufchan_d;
  logic readPointer_QTree_Boolm2a86_1_argbuf_bufchan_r;
  assign readPointer_QTree_Boolm2a86_1_argbuf_r = ((! readPointer_QTree_Boolm2a86_1_argbuf_bufchan_d[0]) || readPointer_QTree_Boolm2a86_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Boolm2a86_1_argbuf_bufchan_d <= {66'd0, 1'd0};
    else
      if (readPointer_QTree_Boolm2a86_1_argbuf_r)
        readPointer_QTree_Boolm2a86_1_argbuf_bufchan_d <= readPointer_QTree_Boolm2a86_1_argbuf_d;
  QTree_Bool_t readPointer_QTree_Boolm2a86_1_argbuf_bufchan_buf;
  assign readPointer_QTree_Boolm2a86_1_argbuf_bufchan_r = (! readPointer_QTree_Boolm2a86_1_argbuf_bufchan_buf[0]);
  assign readPointer_QTree_Boolm2a86_1_argbuf_rwb_d = (readPointer_QTree_Boolm2a86_1_argbuf_bufchan_buf[0] ? readPointer_QTree_Boolm2a86_1_argbuf_bufchan_buf :
                                                       readPointer_QTree_Boolm2a86_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Boolm2a86_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((readPointer_QTree_Boolm2a86_1_argbuf_rwb_r && readPointer_QTree_Boolm2a86_1_argbuf_bufchan_buf[0]))
        readPointer_QTree_Boolm2a86_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
      else if (((! readPointer_QTree_Boolm2a86_1_argbuf_rwb_r) && (! readPointer_QTree_Boolm2a86_1_argbuf_bufchan_buf[0])))
        readPointer_QTree_Boolm2a86_1_argbuf_bufchan_buf <= readPointer_QTree_Boolm2a86_1_argbuf_bufchan_d;
  
  /* buf (Ty QTree_Bool) : (readPointer_QTree_Boolm2a8H_1_argbuf,QTree_Bool) > (readPointer_QTree_Boolm2a8H_1_argbuf_rwb,QTree_Bool) */
  QTree_Bool_t readPointer_QTree_Boolm2a8H_1_argbuf_bufchan_d;
  logic readPointer_QTree_Boolm2a8H_1_argbuf_bufchan_r;
  assign readPointer_QTree_Boolm2a8H_1_argbuf_r = ((! readPointer_QTree_Boolm2a8H_1_argbuf_bufchan_d[0]) || readPointer_QTree_Boolm2a8H_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Boolm2a8H_1_argbuf_bufchan_d <= {66'd0, 1'd0};
    else
      if (readPointer_QTree_Boolm2a8H_1_argbuf_r)
        readPointer_QTree_Boolm2a8H_1_argbuf_bufchan_d <= readPointer_QTree_Boolm2a8H_1_argbuf_d;
  QTree_Bool_t readPointer_QTree_Boolm2a8H_1_argbuf_bufchan_buf;
  assign readPointer_QTree_Boolm2a8H_1_argbuf_bufchan_r = (! readPointer_QTree_Boolm2a8H_1_argbuf_bufchan_buf[0]);
  assign readPointer_QTree_Boolm2a8H_1_argbuf_rwb_d = (readPointer_QTree_Boolm2a8H_1_argbuf_bufchan_buf[0] ? readPointer_QTree_Boolm2a8H_1_argbuf_bufchan_buf :
                                                       readPointer_QTree_Boolm2a8H_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Boolm2a8H_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((readPointer_QTree_Boolm2a8H_1_argbuf_rwb_r && readPointer_QTree_Boolm2a8H_1_argbuf_bufchan_buf[0]))
        readPointer_QTree_Boolm2a8H_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
      else if (((! readPointer_QTree_Boolm2a8H_1_argbuf_rwb_r) && (! readPointer_QTree_Boolm2a8H_1_argbuf_bufchan_buf[0])))
        readPointer_QTree_Boolm2a8H_1_argbuf_bufchan_buf <= readPointer_QTree_Boolm2a8H_1_argbuf_bufchan_d;
  
  /* fork (Ty QTree_Bool) : (readPointer_QTree_Boolm2a8H_1_argbuf_rwb,QTree_Bool) > [(lizzieLet20_1_1,QTree_Bool),
                                                                                (lizzieLet20_1_2,QTree_Bool),
                                                                                (lizzieLet20_1_3,QTree_Bool),
                                                                                (lizzieLet20_1_4,QTree_Bool),
                                                                                (lizzieLet20_1_5,QTree_Bool),
                                                                                (lizzieLet20_1_6,QTree_Bool),
                                                                                (lizzieLet20_1_7,QTree_Bool)] */
  logic [6:0] readPointer_QTree_Boolm2a8H_1_argbuf_rwb_emitted;
  logic [6:0] readPointer_QTree_Boolm2a8H_1_argbuf_rwb_done;
  assign lizzieLet20_1_1_d = {readPointer_QTree_Boolm2a8H_1_argbuf_rwb_d[66:1],
                              (readPointer_QTree_Boolm2a8H_1_argbuf_rwb_d[0] && (! readPointer_QTree_Boolm2a8H_1_argbuf_rwb_emitted[0]))};
  assign lizzieLet20_1_2_d = {readPointer_QTree_Boolm2a8H_1_argbuf_rwb_d[66:1],
                              (readPointer_QTree_Boolm2a8H_1_argbuf_rwb_d[0] && (! readPointer_QTree_Boolm2a8H_1_argbuf_rwb_emitted[1]))};
  assign lizzieLet20_1_3_d = {readPointer_QTree_Boolm2a8H_1_argbuf_rwb_d[66:1],
                              (readPointer_QTree_Boolm2a8H_1_argbuf_rwb_d[0] && (! readPointer_QTree_Boolm2a8H_1_argbuf_rwb_emitted[2]))};
  assign lizzieLet20_1_4_d = {readPointer_QTree_Boolm2a8H_1_argbuf_rwb_d[66:1],
                              (readPointer_QTree_Boolm2a8H_1_argbuf_rwb_d[0] && (! readPointer_QTree_Boolm2a8H_1_argbuf_rwb_emitted[3]))};
  assign lizzieLet20_1_5_d = {readPointer_QTree_Boolm2a8H_1_argbuf_rwb_d[66:1],
                              (readPointer_QTree_Boolm2a8H_1_argbuf_rwb_d[0] && (! readPointer_QTree_Boolm2a8H_1_argbuf_rwb_emitted[4]))};
  assign lizzieLet20_1_6_d = {readPointer_QTree_Boolm2a8H_1_argbuf_rwb_d[66:1],
                              (readPointer_QTree_Boolm2a8H_1_argbuf_rwb_d[0] && (! readPointer_QTree_Boolm2a8H_1_argbuf_rwb_emitted[5]))};
  assign lizzieLet20_1_7_d = {readPointer_QTree_Boolm2a8H_1_argbuf_rwb_d[66:1],
                              (readPointer_QTree_Boolm2a8H_1_argbuf_rwb_d[0] && (! readPointer_QTree_Boolm2a8H_1_argbuf_rwb_emitted[6]))};
  assign readPointer_QTree_Boolm2a8H_1_argbuf_rwb_done = (readPointer_QTree_Boolm2a8H_1_argbuf_rwb_emitted | ({lizzieLet20_1_7_d[0],
                                                                                                               lizzieLet20_1_6_d[0],
                                                                                                               lizzieLet20_1_5_d[0],
                                                                                                               lizzieLet20_1_4_d[0],
                                                                                                               lizzieLet20_1_3_d[0],
                                                                                                               lizzieLet20_1_2_d[0],
                                                                                                               lizzieLet20_1_1_d[0]} & {lizzieLet20_1_7_r,
                                                                                                                                        lizzieLet20_1_6_r,
                                                                                                                                        lizzieLet20_1_5_r,
                                                                                                                                        lizzieLet20_1_4_r,
                                                                                                                                        lizzieLet20_1_3_r,
                                                                                                                                        lizzieLet20_1_2_r,
                                                                                                                                        lizzieLet20_1_1_r}));
  assign readPointer_QTree_Boolm2a8H_1_argbuf_rwb_r = (& readPointer_QTree_Boolm2a8H_1_argbuf_rwb_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Boolm2a8H_1_argbuf_rwb_emitted <= 7'd0;
    else
      readPointer_QTree_Boolm2a8H_1_argbuf_rwb_emitted <= (readPointer_QTree_Boolm2a8H_1_argbuf_rwb_r ? 7'd0 :
                                                           readPointer_QTree_Boolm2a8H_1_argbuf_rwb_done);
  
  /* buf (Ty QTree_Bool) : (readPointer_QTree_Boolm3a87_1_argbuf,QTree_Bool) > (readPointer_QTree_Boolm3a87_1_argbuf_rwb,QTree_Bool) */
  QTree_Bool_t readPointer_QTree_Boolm3a87_1_argbuf_bufchan_d;
  logic readPointer_QTree_Boolm3a87_1_argbuf_bufchan_r;
  assign readPointer_QTree_Boolm3a87_1_argbuf_r = ((! readPointer_QTree_Boolm3a87_1_argbuf_bufchan_d[0]) || readPointer_QTree_Boolm3a87_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Boolm3a87_1_argbuf_bufchan_d <= {66'd0, 1'd0};
    else
      if (readPointer_QTree_Boolm3a87_1_argbuf_r)
        readPointer_QTree_Boolm3a87_1_argbuf_bufchan_d <= readPointer_QTree_Boolm3a87_1_argbuf_d;
  QTree_Bool_t readPointer_QTree_Boolm3a87_1_argbuf_bufchan_buf;
  assign readPointer_QTree_Boolm3a87_1_argbuf_bufchan_r = (! readPointer_QTree_Boolm3a87_1_argbuf_bufchan_buf[0]);
  assign readPointer_QTree_Boolm3a87_1_argbuf_rwb_d = (readPointer_QTree_Boolm3a87_1_argbuf_bufchan_buf[0] ? readPointer_QTree_Boolm3a87_1_argbuf_bufchan_buf :
                                                       readPointer_QTree_Boolm3a87_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Boolm3a87_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((readPointer_QTree_Boolm3a87_1_argbuf_rwb_r && readPointer_QTree_Boolm3a87_1_argbuf_bufchan_buf[0]))
        readPointer_QTree_Boolm3a87_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
      else if (((! readPointer_QTree_Boolm3a87_1_argbuf_rwb_r) && (! readPointer_QTree_Boolm3a87_1_argbuf_bufchan_buf[0])))
        readPointer_QTree_Boolm3a87_1_argbuf_bufchan_buf <= readPointer_QTree_Boolm3a87_1_argbuf_bufchan_d;
  
  /* buf (Ty QTree_Bool) : (readPointer_QTree_Boolm3a8I_1_argbuf,QTree_Bool) > (readPointer_QTree_Boolm3a8I_1_argbuf_rwb,QTree_Bool) */
  QTree_Bool_t readPointer_QTree_Boolm3a8I_1_argbuf_bufchan_d;
  logic readPointer_QTree_Boolm3a8I_1_argbuf_bufchan_r;
  assign readPointer_QTree_Boolm3a8I_1_argbuf_r = ((! readPointer_QTree_Boolm3a8I_1_argbuf_bufchan_d[0]) || readPointer_QTree_Boolm3a8I_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Boolm3a8I_1_argbuf_bufchan_d <= {66'd0, 1'd0};
    else
      if (readPointer_QTree_Boolm3a8I_1_argbuf_r)
        readPointer_QTree_Boolm3a8I_1_argbuf_bufchan_d <= readPointer_QTree_Boolm3a8I_1_argbuf_d;
  QTree_Bool_t readPointer_QTree_Boolm3a8I_1_argbuf_bufchan_buf;
  assign readPointer_QTree_Boolm3a8I_1_argbuf_bufchan_r = (! readPointer_QTree_Boolm3a8I_1_argbuf_bufchan_buf[0]);
  assign readPointer_QTree_Boolm3a8I_1_argbuf_rwb_d = (readPointer_QTree_Boolm3a8I_1_argbuf_bufchan_buf[0] ? readPointer_QTree_Boolm3a8I_1_argbuf_bufchan_buf :
                                                       readPointer_QTree_Boolm3a8I_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Boolm3a8I_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((readPointer_QTree_Boolm3a8I_1_argbuf_rwb_r && readPointer_QTree_Boolm3a8I_1_argbuf_bufchan_buf[0]))
        readPointer_QTree_Boolm3a8I_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
      else if (((! readPointer_QTree_Boolm3a8I_1_argbuf_rwb_r) && (! readPointer_QTree_Boolm3a8I_1_argbuf_bufchan_buf[0])))
        readPointer_QTree_Boolm3a8I_1_argbuf_bufchan_buf <= readPointer_QTree_Boolm3a8I_1_argbuf_bufchan_d;
  
  /* buf (Ty QTree_Bool) : (readPointer_QTree_Boolq4'a8x_1_argbuf,QTree_Bool) > (readPointer_QTree_Boolq4'a8x_1_argbuf_rwb,QTree_Bool) */
  QTree_Bool_t \readPointer_QTree_Boolq4'a8x_1_argbuf_bufchan_d ;
  logic \readPointer_QTree_Boolq4'a8x_1_argbuf_bufchan_r ;
  assign \readPointer_QTree_Boolq4'a8x_1_argbuf_r  = ((! \readPointer_QTree_Boolq4'a8x_1_argbuf_bufchan_d [0]) || \readPointer_QTree_Boolq4'a8x_1_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \readPointer_QTree_Boolq4'a8x_1_argbuf_bufchan_d  <= {66'd0, 1'd0};
    else
      if (\readPointer_QTree_Boolq4'a8x_1_argbuf_r )
        \readPointer_QTree_Boolq4'a8x_1_argbuf_bufchan_d  <= \readPointer_QTree_Boolq4'a8x_1_argbuf_d ;
  QTree_Bool_t \readPointer_QTree_Boolq4'a8x_1_argbuf_bufchan_buf ;
  assign \readPointer_QTree_Boolq4'a8x_1_argbuf_bufchan_r  = (! \readPointer_QTree_Boolq4'a8x_1_argbuf_bufchan_buf [0]);
  assign \readPointer_QTree_Boolq4'a8x_1_argbuf_rwb_d  = (\readPointer_QTree_Boolq4'a8x_1_argbuf_bufchan_buf [0] ? \readPointer_QTree_Boolq4'a8x_1_argbuf_bufchan_buf  :
                                                          \readPointer_QTree_Boolq4'a8x_1_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \readPointer_QTree_Boolq4'a8x_1_argbuf_bufchan_buf  <= {66'd0,
                                                              1'd0};
    else
      if ((\readPointer_QTree_Boolq4'a8x_1_argbuf_rwb_r  && \readPointer_QTree_Boolq4'a8x_1_argbuf_bufchan_buf [0]))
        \readPointer_QTree_Boolq4'a8x_1_argbuf_bufchan_buf  <= {66'd0,
                                                                1'd0};
      else if (((! \readPointer_QTree_Boolq4'a8x_1_argbuf_rwb_r ) && (! \readPointer_QTree_Boolq4'a8x_1_argbuf_bufchan_buf [0])))
        \readPointer_QTree_Boolq4'a8x_1_argbuf_bufchan_buf  <= \readPointer_QTree_Boolq4'a8x_1_argbuf_bufchan_d ;
  
  /* buf (Ty Pointer_CTf') : (sc_0_10_destruct,Pointer_CTf') > (sc_0_10_1_argbuf,Pointer_CTf') */
  \Pointer_CTf'_t  sc_0_10_destruct_bufchan_d;
  logic sc_0_10_destruct_bufchan_r;
  assign sc_0_10_destruct_r = ((! sc_0_10_destruct_bufchan_d[0]) || sc_0_10_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) sc_0_10_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (sc_0_10_destruct_r)
        sc_0_10_destruct_bufchan_d <= sc_0_10_destruct_d;
  \Pointer_CTf'_t  sc_0_10_destruct_bufchan_buf;
  assign sc_0_10_destruct_bufchan_r = (! sc_0_10_destruct_bufchan_buf[0]);
  assign sc_0_10_1_argbuf_d = (sc_0_10_destruct_bufchan_buf[0] ? sc_0_10_destruct_bufchan_buf :
                               sc_0_10_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) sc_0_10_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((sc_0_10_1_argbuf_r && sc_0_10_destruct_bufchan_buf[0]))
        sc_0_10_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! sc_0_10_1_argbuf_r) && (! sc_0_10_destruct_bufchan_buf[0])))
        sc_0_10_destruct_bufchan_buf <= sc_0_10_destruct_bufchan_d;
  
  /* buf (Ty Pointer_CTf'''''''''_f'''''''''_Bool) : (sc_0_14_destruct,Pointer_CTf'''''''''_f'''''''''_Bool) > (sc_0_14_1_argbuf,Pointer_CTf'''''''''_f'''''''''_Bool) */
  \Pointer_CTf'''''''''_f'''''''''_Bool_t  sc_0_14_destruct_bufchan_d;
  logic sc_0_14_destruct_bufchan_r;
  assign sc_0_14_destruct_r = ((! sc_0_14_destruct_bufchan_d[0]) || sc_0_14_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) sc_0_14_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (sc_0_14_destruct_r)
        sc_0_14_destruct_bufchan_d <= sc_0_14_destruct_d;
  \Pointer_CTf'''''''''_f'''''''''_Bool_t  sc_0_14_destruct_bufchan_buf;
  assign sc_0_14_destruct_bufchan_r = (! sc_0_14_destruct_bufchan_buf[0]);
  assign sc_0_14_1_argbuf_d = (sc_0_14_destruct_bufchan_buf[0] ? sc_0_14_destruct_bufchan_buf :
                               sc_0_14_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) sc_0_14_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((sc_0_14_1_argbuf_r && sc_0_14_destruct_bufchan_buf[0]))
        sc_0_14_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! sc_0_14_1_argbuf_r) && (! sc_0_14_destruct_bufchan_buf[0])))
        sc_0_14_destruct_bufchan_buf <= sc_0_14_destruct_bufchan_d;
  
  /* buf (Ty Pointer_CTf) : (sc_0_6_destruct,Pointer_CTf) > (sc_0_6_1_argbuf,Pointer_CTf) */
  Pointer_CTf_t sc_0_6_destruct_bufchan_d;
  logic sc_0_6_destruct_bufchan_r;
  assign sc_0_6_destruct_r = ((! sc_0_6_destruct_bufchan_d[0]) || sc_0_6_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) sc_0_6_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (sc_0_6_destruct_r)
        sc_0_6_destruct_bufchan_d <= sc_0_6_destruct_d;
  Pointer_CTf_t sc_0_6_destruct_bufchan_buf;
  assign sc_0_6_destruct_bufchan_r = (! sc_0_6_destruct_bufchan_buf[0]);
  assign sc_0_6_1_argbuf_d = (sc_0_6_destruct_bufchan_buf[0] ? sc_0_6_destruct_bufchan_buf :
                              sc_0_6_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) sc_0_6_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((sc_0_6_1_argbuf_r && sc_0_6_destruct_bufchan_buf[0]))
        sc_0_6_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! sc_0_6_1_argbuf_r) && (! sc_0_6_destruct_bufchan_buf[0])))
        sc_0_6_destruct_bufchan_buf <= sc_0_6_destruct_bufchan_d;
  
  /* buf (Ty Pointer_CTf') : (scfarg_0_1_goMux_mux,Pointer_CTf') > (scfarg_0_1_1_argbuf,Pointer_CTf') */
  \Pointer_CTf'_t  scfarg_0_1_goMux_mux_bufchan_d;
  logic scfarg_0_1_goMux_mux_bufchan_r;
  assign scfarg_0_1_goMux_mux_r = ((! scfarg_0_1_goMux_mux_bufchan_d[0]) || scfarg_0_1_goMux_mux_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      scfarg_0_1_goMux_mux_bufchan_d <= {16'd0, 1'd0};
    else
      if (scfarg_0_1_goMux_mux_r)
        scfarg_0_1_goMux_mux_bufchan_d <= scfarg_0_1_goMux_mux_d;
  \Pointer_CTf'_t  scfarg_0_1_goMux_mux_bufchan_buf;
  assign scfarg_0_1_goMux_mux_bufchan_r = (! scfarg_0_1_goMux_mux_bufchan_buf[0]);
  assign scfarg_0_1_1_argbuf_d = (scfarg_0_1_goMux_mux_bufchan_buf[0] ? scfarg_0_1_goMux_mux_bufchan_buf :
                                  scfarg_0_1_goMux_mux_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      scfarg_0_1_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((scfarg_0_1_1_argbuf_r && scfarg_0_1_goMux_mux_bufchan_buf[0]))
        scfarg_0_1_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
      else if (((! scfarg_0_1_1_argbuf_r) && (! scfarg_0_1_goMux_mux_bufchan_buf[0])))
        scfarg_0_1_goMux_mux_bufchan_buf <= scfarg_0_1_goMux_mux_bufchan_d;
  
  /* buf (Ty Pointer_CTf'''''''''_f'''''''''_Bool) : (scfarg_0_2_goMux_mux,Pointer_CTf'''''''''_f'''''''''_Bool) > (scfarg_0_2_1_argbuf,Pointer_CTf'''''''''_f'''''''''_Bool) */
  \Pointer_CTf'''''''''_f'''''''''_Bool_t  scfarg_0_2_goMux_mux_bufchan_d;
  logic scfarg_0_2_goMux_mux_bufchan_r;
  assign scfarg_0_2_goMux_mux_r = ((! scfarg_0_2_goMux_mux_bufchan_d[0]) || scfarg_0_2_goMux_mux_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      scfarg_0_2_goMux_mux_bufchan_d <= {16'd0, 1'd0};
    else
      if (scfarg_0_2_goMux_mux_r)
        scfarg_0_2_goMux_mux_bufchan_d <= scfarg_0_2_goMux_mux_d;
  \Pointer_CTf'''''''''_f'''''''''_Bool_t  scfarg_0_2_goMux_mux_bufchan_buf;
  assign scfarg_0_2_goMux_mux_bufchan_r = (! scfarg_0_2_goMux_mux_bufchan_buf[0]);
  assign scfarg_0_2_1_argbuf_d = (scfarg_0_2_goMux_mux_bufchan_buf[0] ? scfarg_0_2_goMux_mux_bufchan_buf :
                                  scfarg_0_2_goMux_mux_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      scfarg_0_2_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((scfarg_0_2_1_argbuf_r && scfarg_0_2_goMux_mux_bufchan_buf[0]))
        scfarg_0_2_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
      else if (((! scfarg_0_2_1_argbuf_r) && (! scfarg_0_2_goMux_mux_bufchan_buf[0])))
        scfarg_0_2_goMux_mux_bufchan_buf <= scfarg_0_2_goMux_mux_bufchan_d;
  
  /* buf (Ty Pointer_CTf) : (scfarg_0_goMux_mux,Pointer_CTf) > (scfarg_0_1_argbuf,Pointer_CTf) */
  Pointer_CTf_t scfarg_0_goMux_mux_bufchan_d;
  logic scfarg_0_goMux_mux_bufchan_r;
  assign scfarg_0_goMux_mux_r = ((! scfarg_0_goMux_mux_bufchan_d[0]) || scfarg_0_goMux_mux_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) scfarg_0_goMux_mux_bufchan_d <= {16'd0, 1'd0};
    else
      if (scfarg_0_goMux_mux_r)
        scfarg_0_goMux_mux_bufchan_d <= scfarg_0_goMux_mux_d;
  Pointer_CTf_t scfarg_0_goMux_mux_bufchan_buf;
  assign scfarg_0_goMux_mux_bufchan_r = (! scfarg_0_goMux_mux_bufchan_buf[0]);
  assign scfarg_0_1_argbuf_d = (scfarg_0_goMux_mux_bufchan_buf[0] ? scfarg_0_goMux_mux_bufchan_buf :
                                scfarg_0_goMux_mux_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      scfarg_0_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((scfarg_0_1_argbuf_r && scfarg_0_goMux_mux_bufchan_buf[0]))
        scfarg_0_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
      else if (((! scfarg_0_1_argbuf_r) && (! scfarg_0_goMux_mux_bufchan_buf[0])))
        scfarg_0_goMux_mux_bufchan_buf <= scfarg_0_goMux_mux_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (t1a8D_3_destruct,Pointer_QTree_Bool) > (t1a8D_3_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t t1a8D_3_destruct_bufchan_d;
  logic t1a8D_3_destruct_bufchan_r;
  assign t1a8D_3_destruct_r = ((! t1a8D_3_destruct_bufchan_d[0]) || t1a8D_3_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t1a8D_3_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (t1a8D_3_destruct_r)
        t1a8D_3_destruct_bufchan_d <= t1a8D_3_destruct_d;
  Pointer_QTree_Bool_t t1a8D_3_destruct_bufchan_buf;
  assign t1a8D_3_destruct_bufchan_r = (! t1a8D_3_destruct_bufchan_buf[0]);
  assign t1a8D_3_1_argbuf_d = (t1a8D_3_destruct_bufchan_buf[0] ? t1a8D_3_destruct_bufchan_buf :
                               t1a8D_3_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t1a8D_3_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((t1a8D_3_1_argbuf_r && t1a8D_3_destruct_bufchan_buf[0]))
        t1a8D_3_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! t1a8D_3_1_argbuf_r) && (! t1a8D_3_destruct_bufchan_buf[0])))
        t1a8D_3_destruct_bufchan_buf <= t1a8D_3_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (t1a8U_3_destruct,Pointer_QTree_Bool) > (t1a8U_3_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t t1a8U_3_destruct_bufchan_d;
  logic t1a8U_3_destruct_bufchan_r;
  assign t1a8U_3_destruct_r = ((! t1a8U_3_destruct_bufchan_d[0]) || t1a8U_3_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t1a8U_3_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (t1a8U_3_destruct_r)
        t1a8U_3_destruct_bufchan_d <= t1a8U_3_destruct_d;
  Pointer_QTree_Bool_t t1a8U_3_destruct_bufchan_buf;
  assign t1a8U_3_destruct_bufchan_r = (! t1a8U_3_destruct_bufchan_buf[0]);
  assign t1a8U_3_1_argbuf_d = (t1a8U_3_destruct_bufchan_buf[0] ? t1a8U_3_destruct_bufchan_buf :
                               t1a8U_3_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t1a8U_3_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((t1a8U_3_1_argbuf_r && t1a8U_3_destruct_bufchan_buf[0]))
        t1a8U_3_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! t1a8U_3_1_argbuf_r) && (! t1a8U_3_destruct_bufchan_buf[0])))
        t1a8U_3_destruct_bufchan_buf <= t1a8U_3_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (t1a8d_destruct,Pointer_QTree_Bool) > (t1a8d_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t t1a8d_destruct_bufchan_d;
  logic t1a8d_destruct_bufchan_r;
  assign t1a8d_destruct_r = ((! t1a8d_destruct_bufchan_d[0]) || t1a8d_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t1a8d_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (t1a8d_destruct_r) t1a8d_destruct_bufchan_d <= t1a8d_destruct_d;
  Pointer_QTree_Bool_t t1a8d_destruct_bufchan_buf;
  assign t1a8d_destruct_bufchan_r = (! t1a8d_destruct_bufchan_buf[0]);
  assign t1a8d_1_argbuf_d = (t1a8d_destruct_bufchan_buf[0] ? t1a8d_destruct_bufchan_buf :
                             t1a8d_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t1a8d_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((t1a8d_1_argbuf_r && t1a8d_destruct_bufchan_buf[0]))
        t1a8d_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! t1a8d_1_argbuf_r) && (! t1a8d_destruct_bufchan_buf[0])))
        t1a8d_destruct_bufchan_buf <= t1a8d_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (t1a8s_3_destruct,Pointer_QTree_Bool) > (t1a8s_3_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t t1a8s_3_destruct_bufchan_d;
  logic t1a8s_3_destruct_bufchan_r;
  assign t1a8s_3_destruct_r = ((! t1a8s_3_destruct_bufchan_d[0]) || t1a8s_3_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t1a8s_3_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (t1a8s_3_destruct_r)
        t1a8s_3_destruct_bufchan_d <= t1a8s_3_destruct_d;
  Pointer_QTree_Bool_t t1a8s_3_destruct_bufchan_buf;
  assign t1a8s_3_destruct_bufchan_r = (! t1a8s_3_destruct_bufchan_buf[0]);
  assign t1a8s_3_1_argbuf_d = (t1a8s_3_destruct_bufchan_buf[0] ? t1a8s_3_destruct_bufchan_buf :
                               t1a8s_3_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t1a8s_3_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((t1a8s_3_1_argbuf_r && t1a8s_3_destruct_bufchan_buf[0]))
        t1a8s_3_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! t1a8s_3_1_argbuf_r) && (! t1a8s_3_destruct_bufchan_buf[0])))
        t1a8s_3_destruct_bufchan_buf <= t1a8s_3_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (t2a8E_2_destruct,Pointer_QTree_Bool) > (t2a8E_2_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t t2a8E_2_destruct_bufchan_d;
  logic t2a8E_2_destruct_bufchan_r;
  assign t2a8E_2_destruct_r = ((! t2a8E_2_destruct_bufchan_d[0]) || t2a8E_2_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t2a8E_2_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (t2a8E_2_destruct_r)
        t2a8E_2_destruct_bufchan_d <= t2a8E_2_destruct_d;
  Pointer_QTree_Bool_t t2a8E_2_destruct_bufchan_buf;
  assign t2a8E_2_destruct_bufchan_r = (! t2a8E_2_destruct_bufchan_buf[0]);
  assign t2a8E_2_1_argbuf_d = (t2a8E_2_destruct_bufchan_buf[0] ? t2a8E_2_destruct_bufchan_buf :
                               t2a8E_2_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t2a8E_2_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((t2a8E_2_1_argbuf_r && t2a8E_2_destruct_bufchan_buf[0]))
        t2a8E_2_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! t2a8E_2_1_argbuf_r) && (! t2a8E_2_destruct_bufchan_buf[0])))
        t2a8E_2_destruct_bufchan_buf <= t2a8E_2_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (t2a8V_2_destruct,Pointer_QTree_Bool) > (t2a8V_2_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t t2a8V_2_destruct_bufchan_d;
  logic t2a8V_2_destruct_bufchan_r;
  assign t2a8V_2_destruct_r = ((! t2a8V_2_destruct_bufchan_d[0]) || t2a8V_2_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t2a8V_2_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (t2a8V_2_destruct_r)
        t2a8V_2_destruct_bufchan_d <= t2a8V_2_destruct_d;
  Pointer_QTree_Bool_t t2a8V_2_destruct_bufchan_buf;
  assign t2a8V_2_destruct_bufchan_r = (! t2a8V_2_destruct_bufchan_buf[0]);
  assign t2a8V_2_1_argbuf_d = (t2a8V_2_destruct_bufchan_buf[0] ? t2a8V_2_destruct_bufchan_buf :
                               t2a8V_2_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t2a8V_2_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((t2a8V_2_1_argbuf_r && t2a8V_2_destruct_bufchan_buf[0]))
        t2a8V_2_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! t2a8V_2_1_argbuf_r) && (! t2a8V_2_destruct_bufchan_buf[0])))
        t2a8V_2_destruct_bufchan_buf <= t2a8V_2_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (t2a8e_destruct,Pointer_QTree_Bool) > (t2a8e_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t t2a8e_destruct_bufchan_d;
  logic t2a8e_destruct_bufchan_r;
  assign t2a8e_destruct_r = ((! t2a8e_destruct_bufchan_d[0]) || t2a8e_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t2a8e_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (t2a8e_destruct_r) t2a8e_destruct_bufchan_d <= t2a8e_destruct_d;
  Pointer_QTree_Bool_t t2a8e_destruct_bufchan_buf;
  assign t2a8e_destruct_bufchan_r = (! t2a8e_destruct_bufchan_buf[0]);
  assign t2a8e_1_argbuf_d = (t2a8e_destruct_bufchan_buf[0] ? t2a8e_destruct_bufchan_buf :
                             t2a8e_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t2a8e_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((t2a8e_1_argbuf_r && t2a8e_destruct_bufchan_buf[0]))
        t2a8e_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! t2a8e_1_argbuf_r) && (! t2a8e_destruct_bufchan_buf[0])))
        t2a8e_destruct_bufchan_buf <= t2a8e_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (t2a8t_2_destruct,Pointer_QTree_Bool) > (t2a8t_2_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t t2a8t_2_destruct_bufchan_d;
  logic t2a8t_2_destruct_bufchan_r;
  assign t2a8t_2_destruct_r = ((! t2a8t_2_destruct_bufchan_d[0]) || t2a8t_2_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t2a8t_2_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (t2a8t_2_destruct_r)
        t2a8t_2_destruct_bufchan_d <= t2a8t_2_destruct_d;
  Pointer_QTree_Bool_t t2a8t_2_destruct_bufchan_buf;
  assign t2a8t_2_destruct_bufchan_r = (! t2a8t_2_destruct_bufchan_buf[0]);
  assign t2a8t_2_1_argbuf_d = (t2a8t_2_destruct_bufchan_buf[0] ? t2a8t_2_destruct_bufchan_buf :
                               t2a8t_2_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t2a8t_2_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((t2a8t_2_1_argbuf_r && t2a8t_2_destruct_bufchan_buf[0]))
        t2a8t_2_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! t2a8t_2_1_argbuf_r) && (! t2a8t_2_destruct_bufchan_buf[0])))
        t2a8t_2_destruct_bufchan_buf <= t2a8t_2_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (t3a8F_1_destruct,Pointer_QTree_Bool) > (t3a8F_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t t3a8F_1_destruct_bufchan_d;
  logic t3a8F_1_destruct_bufchan_r;
  assign t3a8F_1_destruct_r = ((! t3a8F_1_destruct_bufchan_d[0]) || t3a8F_1_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t3a8F_1_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (t3a8F_1_destruct_r)
        t3a8F_1_destruct_bufchan_d <= t3a8F_1_destruct_d;
  Pointer_QTree_Bool_t t3a8F_1_destruct_bufchan_buf;
  assign t3a8F_1_destruct_bufchan_r = (! t3a8F_1_destruct_bufchan_buf[0]);
  assign t3a8F_1_1_argbuf_d = (t3a8F_1_destruct_bufchan_buf[0] ? t3a8F_1_destruct_bufchan_buf :
                               t3a8F_1_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t3a8F_1_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((t3a8F_1_1_argbuf_r && t3a8F_1_destruct_bufchan_buf[0]))
        t3a8F_1_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! t3a8F_1_1_argbuf_r) && (! t3a8F_1_destruct_bufchan_buf[0])))
        t3a8F_1_destruct_bufchan_buf <= t3a8F_1_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (t3a8W_1_destruct,Pointer_QTree_Bool) > (t3a8W_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t t3a8W_1_destruct_bufchan_d;
  logic t3a8W_1_destruct_bufchan_r;
  assign t3a8W_1_destruct_r = ((! t3a8W_1_destruct_bufchan_d[0]) || t3a8W_1_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t3a8W_1_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (t3a8W_1_destruct_r)
        t3a8W_1_destruct_bufchan_d <= t3a8W_1_destruct_d;
  Pointer_QTree_Bool_t t3a8W_1_destruct_bufchan_buf;
  assign t3a8W_1_destruct_bufchan_r = (! t3a8W_1_destruct_bufchan_buf[0]);
  assign t3a8W_1_1_argbuf_d = (t3a8W_1_destruct_bufchan_buf[0] ? t3a8W_1_destruct_bufchan_buf :
                               t3a8W_1_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t3a8W_1_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((t3a8W_1_1_argbuf_r && t3a8W_1_destruct_bufchan_buf[0]))
        t3a8W_1_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! t3a8W_1_1_argbuf_r) && (! t3a8W_1_destruct_bufchan_buf[0])))
        t3a8W_1_destruct_bufchan_buf <= t3a8W_1_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (t3a8f_destruct,Pointer_QTree_Bool) > (t3a8f_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t t3a8f_destruct_bufchan_d;
  logic t3a8f_destruct_bufchan_r;
  assign t3a8f_destruct_r = ((! t3a8f_destruct_bufchan_d[0]) || t3a8f_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t3a8f_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (t3a8f_destruct_r) t3a8f_destruct_bufchan_d <= t3a8f_destruct_d;
  Pointer_QTree_Bool_t t3a8f_destruct_bufchan_buf;
  assign t3a8f_destruct_bufchan_r = (! t3a8f_destruct_bufchan_buf[0]);
  assign t3a8f_1_argbuf_d = (t3a8f_destruct_bufchan_buf[0] ? t3a8f_destruct_bufchan_buf :
                             t3a8f_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t3a8f_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((t3a8f_1_argbuf_r && t3a8f_destruct_bufchan_buf[0]))
        t3a8f_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! t3a8f_1_argbuf_r) && (! t3a8f_destruct_bufchan_buf[0])))
        t3a8f_destruct_bufchan_buf <= t3a8f_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (t3a8u_1_destruct,Pointer_QTree_Bool) > (t3a8u_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t t3a8u_1_destruct_bufchan_d;
  logic t3a8u_1_destruct_bufchan_r;
  assign t3a8u_1_destruct_r = ((! t3a8u_1_destruct_bufchan_d[0]) || t3a8u_1_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t3a8u_1_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (t3a8u_1_destruct_r)
        t3a8u_1_destruct_bufchan_d <= t3a8u_1_destruct_d;
  Pointer_QTree_Bool_t t3a8u_1_destruct_bufchan_buf;
  assign t3a8u_1_destruct_bufchan_r = (! t3a8u_1_destruct_bufchan_buf[0]);
  assign t3a8u_1_1_argbuf_d = (t3a8u_1_destruct_bufchan_buf[0] ? t3a8u_1_destruct_bufchan_buf :
                               t3a8u_1_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t3a8u_1_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((t3a8u_1_1_argbuf_r && t3a8u_1_destruct_bufchan_buf[0]))
        t3a8u_1_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! t3a8u_1_1_argbuf_r) && (! t3a8u_1_destruct_bufchan_buf[0])))
        t3a8u_1_destruct_bufchan_buf <= t3a8u_1_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (t4a8G_destruct,Pointer_QTree_Bool) > (t4a8G_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t t4a8G_destruct_bufchan_d;
  logic t4a8G_destruct_bufchan_r;
  assign t4a8G_destruct_r = ((! t4a8G_destruct_bufchan_d[0]) || t4a8G_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t4a8G_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (t4a8G_destruct_r) t4a8G_destruct_bufchan_d <= t4a8G_destruct_d;
  Pointer_QTree_Bool_t t4a8G_destruct_bufchan_buf;
  assign t4a8G_destruct_bufchan_r = (! t4a8G_destruct_bufchan_buf[0]);
  assign t4a8G_1_argbuf_d = (t4a8G_destruct_bufchan_buf[0] ? t4a8G_destruct_bufchan_buf :
                             t4a8G_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t4a8G_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((t4a8G_1_argbuf_r && t4a8G_destruct_bufchan_buf[0]))
        t4a8G_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! t4a8G_1_argbuf_r) && (! t4a8G_destruct_bufchan_buf[0])))
        t4a8G_destruct_bufchan_buf <= t4a8G_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (t4a8X_destruct,Pointer_QTree_Bool) > (t4a8X_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t t4a8X_destruct_bufchan_d;
  logic t4a8X_destruct_bufchan_r;
  assign t4a8X_destruct_r = ((! t4a8X_destruct_bufchan_d[0]) || t4a8X_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t4a8X_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (t4a8X_destruct_r) t4a8X_destruct_bufchan_d <= t4a8X_destruct_d;
  Pointer_QTree_Bool_t t4a8X_destruct_bufchan_buf;
  assign t4a8X_destruct_bufchan_r = (! t4a8X_destruct_bufchan_buf[0]);
  assign t4a8X_1_argbuf_d = (t4a8X_destruct_bufchan_buf[0] ? t4a8X_destruct_bufchan_buf :
                             t4a8X_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t4a8X_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((t4a8X_1_argbuf_r && t4a8X_destruct_bufchan_buf[0]))
        t4a8X_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! t4a8X_1_argbuf_r) && (! t4a8X_destruct_bufchan_buf[0])))
        t4a8X_destruct_bufchan_buf <= t4a8X_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (t4a8g_destruct,Pointer_QTree_Bool) > (t4a8g_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t t4a8g_destruct_bufchan_d;
  logic t4a8g_destruct_bufchan_r;
  assign t4a8g_destruct_r = ((! t4a8g_destruct_bufchan_d[0]) || t4a8g_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t4a8g_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (t4a8g_destruct_r) t4a8g_destruct_bufchan_d <= t4a8g_destruct_d;
  Pointer_QTree_Bool_t t4a8g_destruct_bufchan_buf;
  assign t4a8g_destruct_bufchan_r = (! t4a8g_destruct_bufchan_buf[0]);
  assign t4a8g_1_argbuf_d = (t4a8g_destruct_bufchan_buf[0] ? t4a8g_destruct_bufchan_buf :
                             t4a8g_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t4a8g_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((t4a8g_1_argbuf_r && t4a8g_destruct_bufchan_buf[0]))
        t4a8g_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! t4a8g_1_argbuf_r) && (! t4a8g_destruct_bufchan_buf[0])))
        t4a8g_destruct_bufchan_buf <= t4a8g_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (t4a8v_destruct,Pointer_QTree_Bool) > (t4a8v_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t t4a8v_destruct_bufchan_d;
  logic t4a8v_destruct_bufchan_r;
  assign t4a8v_destruct_r = ((! t4a8v_destruct_bufchan_d[0]) || t4a8v_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t4a8v_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (t4a8v_destruct_r) t4a8v_destruct_bufchan_d <= t4a8v_destruct_d;
  Pointer_QTree_Bool_t t4a8v_destruct_bufchan_buf;
  assign t4a8v_destruct_bufchan_r = (! t4a8v_destruct_bufchan_buf[0]);
  assign t4a8v_1_argbuf_d = (t4a8v_destruct_bufchan_buf[0] ? t4a8v_destruct_bufchan_buf :
                             t4a8v_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t4a8v_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((t4a8v_1_argbuf_r && t4a8v_destruct_bufchan_buf[0]))
        t4a8v_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! t4a8v_1_argbuf_r) && (! t4a8v_destruct_bufchan_buf[0])))
        t4a8v_destruct_bufchan_buf <= t4a8v_destruct_bufchan_d;
  
  /* buf (Ty Pointer_CTf'''''''''_f'''''''''_Bool) : (writeCTf'''''''''_f'''''''''_BoollizzieLet37_1_argbuf,Pointer_CTf'''''''''_f'''''''''_Bool) > (writeCTf'''''''''_f'''''''''_BoollizzieLet37_1_argbuf_rwb,Pointer_CTf'''''''''_f'''''''''_Bool) */
  \Pointer_CTf'''''''''_f'''''''''_Bool_t  \writeCTf'''''''''_f'''''''''_BoollizzieLet37_1_argbuf_bufchan_d ;
  logic \writeCTf'''''''''_f'''''''''_BoollizzieLet37_1_argbuf_bufchan_r ;
  assign \writeCTf'''''''''_f'''''''''_BoollizzieLet37_1_argbuf_r  = ((! \writeCTf'''''''''_f'''''''''_BoollizzieLet37_1_argbuf_bufchan_d [0]) || \writeCTf'''''''''_f'''''''''_BoollizzieLet37_1_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf'''''''''_f'''''''''_BoollizzieLet37_1_argbuf_bufchan_d  <= {16'd0,
                                                                            1'd0};
    else
      if (\writeCTf'''''''''_f'''''''''_BoollizzieLet37_1_argbuf_r )
        \writeCTf'''''''''_f'''''''''_BoollizzieLet37_1_argbuf_bufchan_d  <= \writeCTf'''''''''_f'''''''''_BoollizzieLet37_1_argbuf_d ;
  \Pointer_CTf'''''''''_f'''''''''_Bool_t  \writeCTf'''''''''_f'''''''''_BoollizzieLet37_1_argbuf_bufchan_buf ;
  assign \writeCTf'''''''''_f'''''''''_BoollizzieLet37_1_argbuf_bufchan_r  = (! \writeCTf'''''''''_f'''''''''_BoollizzieLet37_1_argbuf_bufchan_buf [0]);
  assign \writeCTf'''''''''_f'''''''''_BoollizzieLet37_1_argbuf_rwb_d  = (\writeCTf'''''''''_f'''''''''_BoollizzieLet37_1_argbuf_bufchan_buf [0] ? \writeCTf'''''''''_f'''''''''_BoollizzieLet37_1_argbuf_bufchan_buf  :
                                                                          \writeCTf'''''''''_f'''''''''_BoollizzieLet37_1_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf'''''''''_f'''''''''_BoollizzieLet37_1_argbuf_bufchan_buf  <= {16'd0,
                                                                              1'd0};
    else
      if ((\writeCTf'''''''''_f'''''''''_BoollizzieLet37_1_argbuf_rwb_r  && \writeCTf'''''''''_f'''''''''_BoollizzieLet37_1_argbuf_bufchan_buf [0]))
        \writeCTf'''''''''_f'''''''''_BoollizzieLet37_1_argbuf_bufchan_buf  <= {16'd0,
                                                                                1'd0};
      else if (((! \writeCTf'''''''''_f'''''''''_BoollizzieLet37_1_argbuf_rwb_r ) && (! \writeCTf'''''''''_f'''''''''_BoollizzieLet37_1_argbuf_bufchan_buf [0])))
        \writeCTf'''''''''_f'''''''''_BoollizzieLet37_1_argbuf_bufchan_buf  <= \writeCTf'''''''''_f'''''''''_BoollizzieLet37_1_argbuf_bufchan_d ;
  
  /* buf (Ty Pointer_CTf'''''''''_f'''''''''_Bool) : (writeCTf'''''''''_f'''''''''_BoollizzieLet37_1_argbuf_rwb,Pointer_CTf'''''''''_f'''''''''_Bool) > (sca3_2_1_argbuf,Pointer_CTf'''''''''_f'''''''''_Bool) */
  \Pointer_CTf'''''''''_f'''''''''_Bool_t  \writeCTf'''''''''_f'''''''''_BoollizzieLet37_1_argbuf_rwb_bufchan_d ;
  logic \writeCTf'''''''''_f'''''''''_BoollizzieLet37_1_argbuf_rwb_bufchan_r ;
  assign \writeCTf'''''''''_f'''''''''_BoollizzieLet37_1_argbuf_rwb_r  = ((! \writeCTf'''''''''_f'''''''''_BoollizzieLet37_1_argbuf_rwb_bufchan_d [0]) || \writeCTf'''''''''_f'''''''''_BoollizzieLet37_1_argbuf_rwb_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf'''''''''_f'''''''''_BoollizzieLet37_1_argbuf_rwb_bufchan_d  <= {16'd0,
                                                                                1'd0};
    else
      if (\writeCTf'''''''''_f'''''''''_BoollizzieLet37_1_argbuf_rwb_r )
        \writeCTf'''''''''_f'''''''''_BoollizzieLet37_1_argbuf_rwb_bufchan_d  <= \writeCTf'''''''''_f'''''''''_BoollizzieLet37_1_argbuf_rwb_d ;
  \Pointer_CTf'''''''''_f'''''''''_Bool_t  \writeCTf'''''''''_f'''''''''_BoollizzieLet37_1_argbuf_rwb_bufchan_buf ;
  assign \writeCTf'''''''''_f'''''''''_BoollizzieLet37_1_argbuf_rwb_bufchan_r  = (! \writeCTf'''''''''_f'''''''''_BoollizzieLet37_1_argbuf_rwb_bufchan_buf [0]);
  assign sca3_2_1_argbuf_d = (\writeCTf'''''''''_f'''''''''_BoollizzieLet37_1_argbuf_rwb_bufchan_buf [0] ? \writeCTf'''''''''_f'''''''''_BoollizzieLet37_1_argbuf_rwb_bufchan_buf  :
                              \writeCTf'''''''''_f'''''''''_BoollizzieLet37_1_argbuf_rwb_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf'''''''''_f'''''''''_BoollizzieLet37_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                                  1'd0};
    else
      if ((sca3_2_1_argbuf_r && \writeCTf'''''''''_f'''''''''_BoollizzieLet37_1_argbuf_rwb_bufchan_buf [0]))
        \writeCTf'''''''''_f'''''''''_BoollizzieLet37_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                                    1'd0};
      else if (((! sca3_2_1_argbuf_r) && (! \writeCTf'''''''''_f'''''''''_BoollizzieLet37_1_argbuf_rwb_bufchan_buf [0])))
        \writeCTf'''''''''_f'''''''''_BoollizzieLet37_1_argbuf_rwb_bufchan_buf  <= \writeCTf'''''''''_f'''''''''_BoollizzieLet37_1_argbuf_rwb_bufchan_d ;
  
  /* buf (Ty Pointer_CTf'''''''''_f'''''''''_Bool) : (writeCTf'''''''''_f'''''''''_BoollizzieLet41_1_argbuf,Pointer_CTf'''''''''_f'''''''''_Bool) > (writeCTf'''''''''_f'''''''''_BoollizzieLet41_1_argbuf_rwb,Pointer_CTf'''''''''_f'''''''''_Bool) */
  \Pointer_CTf'''''''''_f'''''''''_Bool_t  \writeCTf'''''''''_f'''''''''_BoollizzieLet41_1_argbuf_bufchan_d ;
  logic \writeCTf'''''''''_f'''''''''_BoollizzieLet41_1_argbuf_bufchan_r ;
  assign \writeCTf'''''''''_f'''''''''_BoollizzieLet41_1_argbuf_r  = ((! \writeCTf'''''''''_f'''''''''_BoollizzieLet41_1_argbuf_bufchan_d [0]) || \writeCTf'''''''''_f'''''''''_BoollizzieLet41_1_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf'''''''''_f'''''''''_BoollizzieLet41_1_argbuf_bufchan_d  <= {16'd0,
                                                                            1'd0};
    else
      if (\writeCTf'''''''''_f'''''''''_BoollizzieLet41_1_argbuf_r )
        \writeCTf'''''''''_f'''''''''_BoollizzieLet41_1_argbuf_bufchan_d  <= \writeCTf'''''''''_f'''''''''_BoollizzieLet41_1_argbuf_d ;
  \Pointer_CTf'''''''''_f'''''''''_Bool_t  \writeCTf'''''''''_f'''''''''_BoollizzieLet41_1_argbuf_bufchan_buf ;
  assign \writeCTf'''''''''_f'''''''''_BoollizzieLet41_1_argbuf_bufchan_r  = (! \writeCTf'''''''''_f'''''''''_BoollizzieLet41_1_argbuf_bufchan_buf [0]);
  assign \writeCTf'''''''''_f'''''''''_BoollizzieLet41_1_argbuf_rwb_d  = (\writeCTf'''''''''_f'''''''''_BoollizzieLet41_1_argbuf_bufchan_buf [0] ? \writeCTf'''''''''_f'''''''''_BoollizzieLet41_1_argbuf_bufchan_buf  :
                                                                          \writeCTf'''''''''_f'''''''''_BoollizzieLet41_1_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf'''''''''_f'''''''''_BoollizzieLet41_1_argbuf_bufchan_buf  <= {16'd0,
                                                                              1'd0};
    else
      if ((\writeCTf'''''''''_f'''''''''_BoollizzieLet41_1_argbuf_rwb_r  && \writeCTf'''''''''_f'''''''''_BoollizzieLet41_1_argbuf_bufchan_buf [0]))
        \writeCTf'''''''''_f'''''''''_BoollizzieLet41_1_argbuf_bufchan_buf  <= {16'd0,
                                                                                1'd0};
      else if (((! \writeCTf'''''''''_f'''''''''_BoollizzieLet41_1_argbuf_rwb_r ) && (! \writeCTf'''''''''_f'''''''''_BoollizzieLet41_1_argbuf_bufchan_buf [0])))
        \writeCTf'''''''''_f'''''''''_BoollizzieLet41_1_argbuf_bufchan_buf  <= \writeCTf'''''''''_f'''''''''_BoollizzieLet41_1_argbuf_bufchan_d ;
  
  /* buf (Ty Pointer_CTf'''''''''_f'''''''''_Bool) : (writeCTf'''''''''_f'''''''''_BoollizzieLet41_1_argbuf_rwb,Pointer_CTf'''''''''_f'''''''''_Bool) > (lizzieLet5_1_1_argbuf,Pointer_CTf'''''''''_f'''''''''_Bool) */
  \Pointer_CTf'''''''''_f'''''''''_Bool_t  \writeCTf'''''''''_f'''''''''_BoollizzieLet41_1_argbuf_rwb_bufchan_d ;
  logic \writeCTf'''''''''_f'''''''''_BoollizzieLet41_1_argbuf_rwb_bufchan_r ;
  assign \writeCTf'''''''''_f'''''''''_BoollizzieLet41_1_argbuf_rwb_r  = ((! \writeCTf'''''''''_f'''''''''_BoollizzieLet41_1_argbuf_rwb_bufchan_d [0]) || \writeCTf'''''''''_f'''''''''_BoollizzieLet41_1_argbuf_rwb_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf'''''''''_f'''''''''_BoollizzieLet41_1_argbuf_rwb_bufchan_d  <= {16'd0,
                                                                                1'd0};
    else
      if (\writeCTf'''''''''_f'''''''''_BoollizzieLet41_1_argbuf_rwb_r )
        \writeCTf'''''''''_f'''''''''_BoollizzieLet41_1_argbuf_rwb_bufchan_d  <= \writeCTf'''''''''_f'''''''''_BoollizzieLet41_1_argbuf_rwb_d ;
  \Pointer_CTf'''''''''_f'''''''''_Bool_t  \writeCTf'''''''''_f'''''''''_BoollizzieLet41_1_argbuf_rwb_bufchan_buf ;
  assign \writeCTf'''''''''_f'''''''''_BoollizzieLet41_1_argbuf_rwb_bufchan_r  = (! \writeCTf'''''''''_f'''''''''_BoollizzieLet41_1_argbuf_rwb_bufchan_buf [0]);
  assign lizzieLet5_1_1_argbuf_d = (\writeCTf'''''''''_f'''''''''_BoollizzieLet41_1_argbuf_rwb_bufchan_buf [0] ? \writeCTf'''''''''_f'''''''''_BoollizzieLet41_1_argbuf_rwb_bufchan_buf  :
                                    \writeCTf'''''''''_f'''''''''_BoollizzieLet41_1_argbuf_rwb_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf'''''''''_f'''''''''_BoollizzieLet41_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                                  1'd0};
    else
      if ((lizzieLet5_1_1_argbuf_r && \writeCTf'''''''''_f'''''''''_BoollizzieLet41_1_argbuf_rwb_bufchan_buf [0]))
        \writeCTf'''''''''_f'''''''''_BoollizzieLet41_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                                    1'd0};
      else if (((! lizzieLet5_1_1_argbuf_r) && (! \writeCTf'''''''''_f'''''''''_BoollizzieLet41_1_argbuf_rwb_bufchan_buf [0])))
        \writeCTf'''''''''_f'''''''''_BoollizzieLet41_1_argbuf_rwb_bufchan_buf  <= \writeCTf'''''''''_f'''''''''_BoollizzieLet41_1_argbuf_rwb_bufchan_d ;
  
  /* buf (Ty Pointer_CTf'''''''''_f'''''''''_Bool) : (writeCTf'''''''''_f'''''''''_BoollizzieLet54_1_argbuf,Pointer_CTf'''''''''_f'''''''''_Bool) > (writeCTf'''''''''_f'''''''''_BoollizzieLet54_1_argbuf_rwb,Pointer_CTf'''''''''_f'''''''''_Bool) */
  \Pointer_CTf'''''''''_f'''''''''_Bool_t  \writeCTf'''''''''_f'''''''''_BoollizzieLet54_1_argbuf_bufchan_d ;
  logic \writeCTf'''''''''_f'''''''''_BoollizzieLet54_1_argbuf_bufchan_r ;
  assign \writeCTf'''''''''_f'''''''''_BoollizzieLet54_1_argbuf_r  = ((! \writeCTf'''''''''_f'''''''''_BoollizzieLet54_1_argbuf_bufchan_d [0]) || \writeCTf'''''''''_f'''''''''_BoollizzieLet54_1_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf'''''''''_f'''''''''_BoollizzieLet54_1_argbuf_bufchan_d  <= {16'd0,
                                                                            1'd0};
    else
      if (\writeCTf'''''''''_f'''''''''_BoollizzieLet54_1_argbuf_r )
        \writeCTf'''''''''_f'''''''''_BoollizzieLet54_1_argbuf_bufchan_d  <= \writeCTf'''''''''_f'''''''''_BoollizzieLet54_1_argbuf_d ;
  \Pointer_CTf'''''''''_f'''''''''_Bool_t  \writeCTf'''''''''_f'''''''''_BoollizzieLet54_1_argbuf_bufchan_buf ;
  assign \writeCTf'''''''''_f'''''''''_BoollizzieLet54_1_argbuf_bufchan_r  = (! \writeCTf'''''''''_f'''''''''_BoollizzieLet54_1_argbuf_bufchan_buf [0]);
  assign \writeCTf'''''''''_f'''''''''_BoollizzieLet54_1_argbuf_rwb_d  = (\writeCTf'''''''''_f'''''''''_BoollizzieLet54_1_argbuf_bufchan_buf [0] ? \writeCTf'''''''''_f'''''''''_BoollizzieLet54_1_argbuf_bufchan_buf  :
                                                                          \writeCTf'''''''''_f'''''''''_BoollizzieLet54_1_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf'''''''''_f'''''''''_BoollizzieLet54_1_argbuf_bufchan_buf  <= {16'd0,
                                                                              1'd0};
    else
      if ((\writeCTf'''''''''_f'''''''''_BoollizzieLet54_1_argbuf_rwb_r  && \writeCTf'''''''''_f'''''''''_BoollizzieLet54_1_argbuf_bufchan_buf [0]))
        \writeCTf'''''''''_f'''''''''_BoollizzieLet54_1_argbuf_bufchan_buf  <= {16'd0,
                                                                                1'd0};
      else if (((! \writeCTf'''''''''_f'''''''''_BoollizzieLet54_1_argbuf_rwb_r ) && (! \writeCTf'''''''''_f'''''''''_BoollizzieLet54_1_argbuf_bufchan_buf [0])))
        \writeCTf'''''''''_f'''''''''_BoollizzieLet54_1_argbuf_bufchan_buf  <= \writeCTf'''''''''_f'''''''''_BoollizzieLet54_1_argbuf_bufchan_d ;
  
  /* buf (Ty Pointer_CTf'''''''''_f'''''''''_Bool) : (writeCTf'''''''''_f'''''''''_BoollizzieLet54_1_argbuf_rwb,Pointer_CTf'''''''''_f'''''''''_Bool) > (sca2_2_1_argbuf,Pointer_CTf'''''''''_f'''''''''_Bool) */
  \Pointer_CTf'''''''''_f'''''''''_Bool_t  \writeCTf'''''''''_f'''''''''_BoollizzieLet54_1_argbuf_rwb_bufchan_d ;
  logic \writeCTf'''''''''_f'''''''''_BoollizzieLet54_1_argbuf_rwb_bufchan_r ;
  assign \writeCTf'''''''''_f'''''''''_BoollizzieLet54_1_argbuf_rwb_r  = ((! \writeCTf'''''''''_f'''''''''_BoollizzieLet54_1_argbuf_rwb_bufchan_d [0]) || \writeCTf'''''''''_f'''''''''_BoollizzieLet54_1_argbuf_rwb_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf'''''''''_f'''''''''_BoollizzieLet54_1_argbuf_rwb_bufchan_d  <= {16'd0,
                                                                                1'd0};
    else
      if (\writeCTf'''''''''_f'''''''''_BoollizzieLet54_1_argbuf_rwb_r )
        \writeCTf'''''''''_f'''''''''_BoollizzieLet54_1_argbuf_rwb_bufchan_d  <= \writeCTf'''''''''_f'''''''''_BoollizzieLet54_1_argbuf_rwb_d ;
  \Pointer_CTf'''''''''_f'''''''''_Bool_t  \writeCTf'''''''''_f'''''''''_BoollizzieLet54_1_argbuf_rwb_bufchan_buf ;
  assign \writeCTf'''''''''_f'''''''''_BoollizzieLet54_1_argbuf_rwb_bufchan_r  = (! \writeCTf'''''''''_f'''''''''_BoollizzieLet54_1_argbuf_rwb_bufchan_buf [0]);
  assign sca2_2_1_argbuf_d = (\writeCTf'''''''''_f'''''''''_BoollizzieLet54_1_argbuf_rwb_bufchan_buf [0] ? \writeCTf'''''''''_f'''''''''_BoollizzieLet54_1_argbuf_rwb_bufchan_buf  :
                              \writeCTf'''''''''_f'''''''''_BoollizzieLet54_1_argbuf_rwb_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf'''''''''_f'''''''''_BoollizzieLet54_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                                  1'd0};
    else
      if ((sca2_2_1_argbuf_r && \writeCTf'''''''''_f'''''''''_BoollizzieLet54_1_argbuf_rwb_bufchan_buf [0]))
        \writeCTf'''''''''_f'''''''''_BoollizzieLet54_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                                    1'd0};
      else if (((! sca2_2_1_argbuf_r) && (! \writeCTf'''''''''_f'''''''''_BoollizzieLet54_1_argbuf_rwb_bufchan_buf [0])))
        \writeCTf'''''''''_f'''''''''_BoollizzieLet54_1_argbuf_rwb_bufchan_buf  <= \writeCTf'''''''''_f'''''''''_BoollizzieLet54_1_argbuf_rwb_bufchan_d ;
  
  /* buf (Ty Pointer_CTf'''''''''_f'''''''''_Bool) : (writeCTf'''''''''_f'''''''''_BoollizzieLet55_1_argbuf,Pointer_CTf'''''''''_f'''''''''_Bool) > (writeCTf'''''''''_f'''''''''_BoollizzieLet55_1_argbuf_rwb,Pointer_CTf'''''''''_f'''''''''_Bool) */
  \Pointer_CTf'''''''''_f'''''''''_Bool_t  \writeCTf'''''''''_f'''''''''_BoollizzieLet55_1_argbuf_bufchan_d ;
  logic \writeCTf'''''''''_f'''''''''_BoollizzieLet55_1_argbuf_bufchan_r ;
  assign \writeCTf'''''''''_f'''''''''_BoollizzieLet55_1_argbuf_r  = ((! \writeCTf'''''''''_f'''''''''_BoollizzieLet55_1_argbuf_bufchan_d [0]) || \writeCTf'''''''''_f'''''''''_BoollizzieLet55_1_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf'''''''''_f'''''''''_BoollizzieLet55_1_argbuf_bufchan_d  <= {16'd0,
                                                                            1'd0};
    else
      if (\writeCTf'''''''''_f'''''''''_BoollizzieLet55_1_argbuf_r )
        \writeCTf'''''''''_f'''''''''_BoollizzieLet55_1_argbuf_bufchan_d  <= \writeCTf'''''''''_f'''''''''_BoollizzieLet55_1_argbuf_d ;
  \Pointer_CTf'''''''''_f'''''''''_Bool_t  \writeCTf'''''''''_f'''''''''_BoollizzieLet55_1_argbuf_bufchan_buf ;
  assign \writeCTf'''''''''_f'''''''''_BoollizzieLet55_1_argbuf_bufchan_r  = (! \writeCTf'''''''''_f'''''''''_BoollizzieLet55_1_argbuf_bufchan_buf [0]);
  assign \writeCTf'''''''''_f'''''''''_BoollizzieLet55_1_argbuf_rwb_d  = (\writeCTf'''''''''_f'''''''''_BoollizzieLet55_1_argbuf_bufchan_buf [0] ? \writeCTf'''''''''_f'''''''''_BoollizzieLet55_1_argbuf_bufchan_buf  :
                                                                          \writeCTf'''''''''_f'''''''''_BoollizzieLet55_1_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf'''''''''_f'''''''''_BoollizzieLet55_1_argbuf_bufchan_buf  <= {16'd0,
                                                                              1'd0};
    else
      if ((\writeCTf'''''''''_f'''''''''_BoollizzieLet55_1_argbuf_rwb_r  && \writeCTf'''''''''_f'''''''''_BoollizzieLet55_1_argbuf_bufchan_buf [0]))
        \writeCTf'''''''''_f'''''''''_BoollizzieLet55_1_argbuf_bufchan_buf  <= {16'd0,
                                                                                1'd0};
      else if (((! \writeCTf'''''''''_f'''''''''_BoollizzieLet55_1_argbuf_rwb_r ) && (! \writeCTf'''''''''_f'''''''''_BoollizzieLet55_1_argbuf_bufchan_buf [0])))
        \writeCTf'''''''''_f'''''''''_BoollizzieLet55_1_argbuf_bufchan_buf  <= \writeCTf'''''''''_f'''''''''_BoollizzieLet55_1_argbuf_bufchan_d ;
  
  /* buf (Ty Pointer_CTf'''''''''_f'''''''''_Bool) : (writeCTf'''''''''_f'''''''''_BoollizzieLet55_1_argbuf_rwb,Pointer_CTf'''''''''_f'''''''''_Bool) > (sca1_2_1_argbuf,Pointer_CTf'''''''''_f'''''''''_Bool) */
  \Pointer_CTf'''''''''_f'''''''''_Bool_t  \writeCTf'''''''''_f'''''''''_BoollizzieLet55_1_argbuf_rwb_bufchan_d ;
  logic \writeCTf'''''''''_f'''''''''_BoollizzieLet55_1_argbuf_rwb_bufchan_r ;
  assign \writeCTf'''''''''_f'''''''''_BoollizzieLet55_1_argbuf_rwb_r  = ((! \writeCTf'''''''''_f'''''''''_BoollizzieLet55_1_argbuf_rwb_bufchan_d [0]) || \writeCTf'''''''''_f'''''''''_BoollizzieLet55_1_argbuf_rwb_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf'''''''''_f'''''''''_BoollizzieLet55_1_argbuf_rwb_bufchan_d  <= {16'd0,
                                                                                1'd0};
    else
      if (\writeCTf'''''''''_f'''''''''_BoollizzieLet55_1_argbuf_rwb_r )
        \writeCTf'''''''''_f'''''''''_BoollizzieLet55_1_argbuf_rwb_bufchan_d  <= \writeCTf'''''''''_f'''''''''_BoollizzieLet55_1_argbuf_rwb_d ;
  \Pointer_CTf'''''''''_f'''''''''_Bool_t  \writeCTf'''''''''_f'''''''''_BoollizzieLet55_1_argbuf_rwb_bufchan_buf ;
  assign \writeCTf'''''''''_f'''''''''_BoollizzieLet55_1_argbuf_rwb_bufchan_r  = (! \writeCTf'''''''''_f'''''''''_BoollizzieLet55_1_argbuf_rwb_bufchan_buf [0]);
  assign sca1_2_1_argbuf_d = (\writeCTf'''''''''_f'''''''''_BoollizzieLet55_1_argbuf_rwb_bufchan_buf [0] ? \writeCTf'''''''''_f'''''''''_BoollizzieLet55_1_argbuf_rwb_bufchan_buf  :
                              \writeCTf'''''''''_f'''''''''_BoollizzieLet55_1_argbuf_rwb_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf'''''''''_f'''''''''_BoollizzieLet55_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                                  1'd0};
    else
      if ((sca1_2_1_argbuf_r && \writeCTf'''''''''_f'''''''''_BoollizzieLet55_1_argbuf_rwb_bufchan_buf [0]))
        \writeCTf'''''''''_f'''''''''_BoollizzieLet55_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                                    1'd0};
      else if (((! sca1_2_1_argbuf_r) && (! \writeCTf'''''''''_f'''''''''_BoollizzieLet55_1_argbuf_rwb_bufchan_buf [0])))
        \writeCTf'''''''''_f'''''''''_BoollizzieLet55_1_argbuf_rwb_bufchan_buf  <= \writeCTf'''''''''_f'''''''''_BoollizzieLet55_1_argbuf_rwb_bufchan_d ;
  
  /* buf (Ty Pointer_CTf'''''''''_f'''''''''_Bool) : (writeCTf'''''''''_f'''''''''_BoollizzieLet56_1_argbuf,Pointer_CTf'''''''''_f'''''''''_Bool) > (writeCTf'''''''''_f'''''''''_BoollizzieLet56_1_argbuf_rwb,Pointer_CTf'''''''''_f'''''''''_Bool) */
  \Pointer_CTf'''''''''_f'''''''''_Bool_t  \writeCTf'''''''''_f'''''''''_BoollizzieLet56_1_argbuf_bufchan_d ;
  logic \writeCTf'''''''''_f'''''''''_BoollizzieLet56_1_argbuf_bufchan_r ;
  assign \writeCTf'''''''''_f'''''''''_BoollizzieLet56_1_argbuf_r  = ((! \writeCTf'''''''''_f'''''''''_BoollizzieLet56_1_argbuf_bufchan_d [0]) || \writeCTf'''''''''_f'''''''''_BoollizzieLet56_1_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf'''''''''_f'''''''''_BoollizzieLet56_1_argbuf_bufchan_d  <= {16'd0,
                                                                            1'd0};
    else
      if (\writeCTf'''''''''_f'''''''''_BoollizzieLet56_1_argbuf_r )
        \writeCTf'''''''''_f'''''''''_BoollizzieLet56_1_argbuf_bufchan_d  <= \writeCTf'''''''''_f'''''''''_BoollizzieLet56_1_argbuf_d ;
  \Pointer_CTf'''''''''_f'''''''''_Bool_t  \writeCTf'''''''''_f'''''''''_BoollizzieLet56_1_argbuf_bufchan_buf ;
  assign \writeCTf'''''''''_f'''''''''_BoollizzieLet56_1_argbuf_bufchan_r  = (! \writeCTf'''''''''_f'''''''''_BoollizzieLet56_1_argbuf_bufchan_buf [0]);
  assign \writeCTf'''''''''_f'''''''''_BoollizzieLet56_1_argbuf_rwb_d  = (\writeCTf'''''''''_f'''''''''_BoollizzieLet56_1_argbuf_bufchan_buf [0] ? \writeCTf'''''''''_f'''''''''_BoollizzieLet56_1_argbuf_bufchan_buf  :
                                                                          \writeCTf'''''''''_f'''''''''_BoollizzieLet56_1_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf'''''''''_f'''''''''_BoollizzieLet56_1_argbuf_bufchan_buf  <= {16'd0,
                                                                              1'd0};
    else
      if ((\writeCTf'''''''''_f'''''''''_BoollizzieLet56_1_argbuf_rwb_r  && \writeCTf'''''''''_f'''''''''_BoollizzieLet56_1_argbuf_bufchan_buf [0]))
        \writeCTf'''''''''_f'''''''''_BoollizzieLet56_1_argbuf_bufchan_buf  <= {16'd0,
                                                                                1'd0};
      else if (((! \writeCTf'''''''''_f'''''''''_BoollizzieLet56_1_argbuf_rwb_r ) && (! \writeCTf'''''''''_f'''''''''_BoollizzieLet56_1_argbuf_bufchan_buf [0])))
        \writeCTf'''''''''_f'''''''''_BoollizzieLet56_1_argbuf_bufchan_buf  <= \writeCTf'''''''''_f'''''''''_BoollizzieLet56_1_argbuf_bufchan_d ;
  
  /* buf (Ty Pointer_CTf'''''''''_f'''''''''_Bool) : (writeCTf'''''''''_f'''''''''_BoollizzieLet56_1_argbuf_rwb,Pointer_CTf'''''''''_f'''''''''_Bool) > (sca0_2_1_argbuf,Pointer_CTf'''''''''_f'''''''''_Bool) */
  \Pointer_CTf'''''''''_f'''''''''_Bool_t  \writeCTf'''''''''_f'''''''''_BoollizzieLet56_1_argbuf_rwb_bufchan_d ;
  logic \writeCTf'''''''''_f'''''''''_BoollizzieLet56_1_argbuf_rwb_bufchan_r ;
  assign \writeCTf'''''''''_f'''''''''_BoollizzieLet56_1_argbuf_rwb_r  = ((! \writeCTf'''''''''_f'''''''''_BoollizzieLet56_1_argbuf_rwb_bufchan_d [0]) || \writeCTf'''''''''_f'''''''''_BoollizzieLet56_1_argbuf_rwb_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf'''''''''_f'''''''''_BoollizzieLet56_1_argbuf_rwb_bufchan_d  <= {16'd0,
                                                                                1'd0};
    else
      if (\writeCTf'''''''''_f'''''''''_BoollizzieLet56_1_argbuf_rwb_r )
        \writeCTf'''''''''_f'''''''''_BoollizzieLet56_1_argbuf_rwb_bufchan_d  <= \writeCTf'''''''''_f'''''''''_BoollizzieLet56_1_argbuf_rwb_d ;
  \Pointer_CTf'''''''''_f'''''''''_Bool_t  \writeCTf'''''''''_f'''''''''_BoollizzieLet56_1_argbuf_rwb_bufchan_buf ;
  assign \writeCTf'''''''''_f'''''''''_BoollizzieLet56_1_argbuf_rwb_bufchan_r  = (! \writeCTf'''''''''_f'''''''''_BoollizzieLet56_1_argbuf_rwb_bufchan_buf [0]);
  assign sca0_2_1_argbuf_d = (\writeCTf'''''''''_f'''''''''_BoollizzieLet56_1_argbuf_rwb_bufchan_buf [0] ? \writeCTf'''''''''_f'''''''''_BoollizzieLet56_1_argbuf_rwb_bufchan_buf  :
                              \writeCTf'''''''''_f'''''''''_BoollizzieLet56_1_argbuf_rwb_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf'''''''''_f'''''''''_BoollizzieLet56_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                                  1'd0};
    else
      if ((sca0_2_1_argbuf_r && \writeCTf'''''''''_f'''''''''_BoollizzieLet56_1_argbuf_rwb_bufchan_buf [0]))
        \writeCTf'''''''''_f'''''''''_BoollizzieLet56_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                                    1'd0};
      else if (((! sca0_2_1_argbuf_r) && (! \writeCTf'''''''''_f'''''''''_BoollizzieLet56_1_argbuf_rwb_bufchan_buf [0])))
        \writeCTf'''''''''_f'''''''''_BoollizzieLet56_1_argbuf_rwb_bufchan_buf  <= \writeCTf'''''''''_f'''''''''_BoollizzieLet56_1_argbuf_rwb_bufchan_d ;
  
  /* buf (Ty Pointer_CTf') : (writeCTf'lizzieLet29_1_argbuf,Pointer_CTf') > (writeCTf'lizzieLet29_1_argbuf_rwb,Pointer_CTf') */
  \Pointer_CTf'_t  \writeCTf'lizzieLet29_1_argbuf_bufchan_d ;
  logic \writeCTf'lizzieLet29_1_argbuf_bufchan_r ;
  assign \writeCTf'lizzieLet29_1_argbuf_r  = ((! \writeCTf'lizzieLet29_1_argbuf_bufchan_d [0]) || \writeCTf'lizzieLet29_1_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf'lizzieLet29_1_argbuf_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\writeCTf'lizzieLet29_1_argbuf_r )
        \writeCTf'lizzieLet29_1_argbuf_bufchan_d  <= \writeCTf'lizzieLet29_1_argbuf_d ;
  \Pointer_CTf'_t  \writeCTf'lizzieLet29_1_argbuf_bufchan_buf ;
  assign \writeCTf'lizzieLet29_1_argbuf_bufchan_r  = (! \writeCTf'lizzieLet29_1_argbuf_bufchan_buf [0]);
  assign \writeCTf'lizzieLet29_1_argbuf_rwb_d  = (\writeCTf'lizzieLet29_1_argbuf_bufchan_buf [0] ? \writeCTf'lizzieLet29_1_argbuf_bufchan_buf  :
                                                  \writeCTf'lizzieLet29_1_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf'lizzieLet29_1_argbuf_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((\writeCTf'lizzieLet29_1_argbuf_rwb_r  && \writeCTf'lizzieLet29_1_argbuf_bufchan_buf [0]))
        \writeCTf'lizzieLet29_1_argbuf_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! \writeCTf'lizzieLet29_1_argbuf_rwb_r ) && (! \writeCTf'lizzieLet29_1_argbuf_bufchan_buf [0])))
        \writeCTf'lizzieLet29_1_argbuf_bufchan_buf  <= \writeCTf'lizzieLet29_1_argbuf_bufchan_d ;
  
  /* buf (Ty Pointer_CTf') : (writeCTf'lizzieLet29_1_argbuf_rwb,Pointer_CTf') > (sca3_1_1_argbuf,Pointer_CTf') */
  \Pointer_CTf'_t  \writeCTf'lizzieLet29_1_argbuf_rwb_bufchan_d ;
  logic \writeCTf'lizzieLet29_1_argbuf_rwb_bufchan_r ;
  assign \writeCTf'lizzieLet29_1_argbuf_rwb_r  = ((! \writeCTf'lizzieLet29_1_argbuf_rwb_bufchan_d [0]) || \writeCTf'lizzieLet29_1_argbuf_rwb_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf'lizzieLet29_1_argbuf_rwb_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\writeCTf'lizzieLet29_1_argbuf_rwb_r )
        \writeCTf'lizzieLet29_1_argbuf_rwb_bufchan_d  <= \writeCTf'lizzieLet29_1_argbuf_rwb_d ;
  \Pointer_CTf'_t  \writeCTf'lizzieLet29_1_argbuf_rwb_bufchan_buf ;
  assign \writeCTf'lizzieLet29_1_argbuf_rwb_bufchan_r  = (! \writeCTf'lizzieLet29_1_argbuf_rwb_bufchan_buf [0]);
  assign sca3_1_1_argbuf_d = (\writeCTf'lizzieLet29_1_argbuf_rwb_bufchan_buf [0] ? \writeCTf'lizzieLet29_1_argbuf_rwb_bufchan_buf  :
                              \writeCTf'lizzieLet29_1_argbuf_rwb_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf'lizzieLet29_1_argbuf_rwb_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((sca3_1_1_argbuf_r && \writeCTf'lizzieLet29_1_argbuf_rwb_bufchan_buf [0]))
        \writeCTf'lizzieLet29_1_argbuf_rwb_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! sca3_1_1_argbuf_r) && (! \writeCTf'lizzieLet29_1_argbuf_rwb_bufchan_buf [0])))
        \writeCTf'lizzieLet29_1_argbuf_rwb_bufchan_buf  <= \writeCTf'lizzieLet29_1_argbuf_rwb_bufchan_d ;
  
  /* buf (Ty Pointer_CTf') : (writeCTf'lizzieLet40_1_argbuf,Pointer_CTf') > (writeCTf'lizzieLet40_1_argbuf_rwb,Pointer_CTf') */
  \Pointer_CTf'_t  \writeCTf'lizzieLet40_1_argbuf_bufchan_d ;
  logic \writeCTf'lizzieLet40_1_argbuf_bufchan_r ;
  assign \writeCTf'lizzieLet40_1_argbuf_r  = ((! \writeCTf'lizzieLet40_1_argbuf_bufchan_d [0]) || \writeCTf'lizzieLet40_1_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf'lizzieLet40_1_argbuf_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\writeCTf'lizzieLet40_1_argbuf_r )
        \writeCTf'lizzieLet40_1_argbuf_bufchan_d  <= \writeCTf'lizzieLet40_1_argbuf_d ;
  \Pointer_CTf'_t  \writeCTf'lizzieLet40_1_argbuf_bufchan_buf ;
  assign \writeCTf'lizzieLet40_1_argbuf_bufchan_r  = (! \writeCTf'lizzieLet40_1_argbuf_bufchan_buf [0]);
  assign \writeCTf'lizzieLet40_1_argbuf_rwb_d  = (\writeCTf'lizzieLet40_1_argbuf_bufchan_buf [0] ? \writeCTf'lizzieLet40_1_argbuf_bufchan_buf  :
                                                  \writeCTf'lizzieLet40_1_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf'lizzieLet40_1_argbuf_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((\writeCTf'lizzieLet40_1_argbuf_rwb_r  && \writeCTf'lizzieLet40_1_argbuf_bufchan_buf [0]))
        \writeCTf'lizzieLet40_1_argbuf_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! \writeCTf'lizzieLet40_1_argbuf_rwb_r ) && (! \writeCTf'lizzieLet40_1_argbuf_bufchan_buf [0])))
        \writeCTf'lizzieLet40_1_argbuf_bufchan_buf  <= \writeCTf'lizzieLet40_1_argbuf_bufchan_d ;
  
  /* buf (Ty Pointer_CTf') : (writeCTf'lizzieLet40_1_argbuf_rwb,Pointer_CTf') > (lizzieLet12_1_1_argbuf,Pointer_CTf') */
  \Pointer_CTf'_t  \writeCTf'lizzieLet40_1_argbuf_rwb_bufchan_d ;
  logic \writeCTf'lizzieLet40_1_argbuf_rwb_bufchan_r ;
  assign \writeCTf'lizzieLet40_1_argbuf_rwb_r  = ((! \writeCTf'lizzieLet40_1_argbuf_rwb_bufchan_d [0]) || \writeCTf'lizzieLet40_1_argbuf_rwb_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf'lizzieLet40_1_argbuf_rwb_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\writeCTf'lizzieLet40_1_argbuf_rwb_r )
        \writeCTf'lizzieLet40_1_argbuf_rwb_bufchan_d  <= \writeCTf'lizzieLet40_1_argbuf_rwb_d ;
  \Pointer_CTf'_t  \writeCTf'lizzieLet40_1_argbuf_rwb_bufchan_buf ;
  assign \writeCTf'lizzieLet40_1_argbuf_rwb_bufchan_r  = (! \writeCTf'lizzieLet40_1_argbuf_rwb_bufchan_buf [0]);
  assign lizzieLet12_1_1_argbuf_d = (\writeCTf'lizzieLet40_1_argbuf_rwb_bufchan_buf [0] ? \writeCTf'lizzieLet40_1_argbuf_rwb_bufchan_buf  :
                                     \writeCTf'lizzieLet40_1_argbuf_rwb_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf'lizzieLet40_1_argbuf_rwb_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((lizzieLet12_1_1_argbuf_r && \writeCTf'lizzieLet40_1_argbuf_rwb_bufchan_buf [0]))
        \writeCTf'lizzieLet40_1_argbuf_rwb_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! lizzieLet12_1_1_argbuf_r) && (! \writeCTf'lizzieLet40_1_argbuf_rwb_bufchan_buf [0])))
        \writeCTf'lizzieLet40_1_argbuf_rwb_bufchan_buf  <= \writeCTf'lizzieLet40_1_argbuf_rwb_bufchan_d ;
  
  /* buf (Ty Pointer_CTf') : (writeCTf'lizzieLet49_1_argbuf,Pointer_CTf') > (writeCTf'lizzieLet49_1_argbuf_rwb,Pointer_CTf') */
  \Pointer_CTf'_t  \writeCTf'lizzieLet49_1_argbuf_bufchan_d ;
  logic \writeCTf'lizzieLet49_1_argbuf_bufchan_r ;
  assign \writeCTf'lizzieLet49_1_argbuf_r  = ((! \writeCTf'lizzieLet49_1_argbuf_bufchan_d [0]) || \writeCTf'lizzieLet49_1_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf'lizzieLet49_1_argbuf_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\writeCTf'lizzieLet49_1_argbuf_r )
        \writeCTf'lizzieLet49_1_argbuf_bufchan_d  <= \writeCTf'lizzieLet49_1_argbuf_d ;
  \Pointer_CTf'_t  \writeCTf'lizzieLet49_1_argbuf_bufchan_buf ;
  assign \writeCTf'lizzieLet49_1_argbuf_bufchan_r  = (! \writeCTf'lizzieLet49_1_argbuf_bufchan_buf [0]);
  assign \writeCTf'lizzieLet49_1_argbuf_rwb_d  = (\writeCTf'lizzieLet49_1_argbuf_bufchan_buf [0] ? \writeCTf'lizzieLet49_1_argbuf_bufchan_buf  :
                                                  \writeCTf'lizzieLet49_1_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf'lizzieLet49_1_argbuf_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((\writeCTf'lizzieLet49_1_argbuf_rwb_r  && \writeCTf'lizzieLet49_1_argbuf_bufchan_buf [0]))
        \writeCTf'lizzieLet49_1_argbuf_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! \writeCTf'lizzieLet49_1_argbuf_rwb_r ) && (! \writeCTf'lizzieLet49_1_argbuf_bufchan_buf [0])))
        \writeCTf'lizzieLet49_1_argbuf_bufchan_buf  <= \writeCTf'lizzieLet49_1_argbuf_bufchan_d ;
  
  /* buf (Ty Pointer_CTf') : (writeCTf'lizzieLet49_1_argbuf_rwb,Pointer_CTf') > (sca2_1_1_argbuf,Pointer_CTf') */
  \Pointer_CTf'_t  \writeCTf'lizzieLet49_1_argbuf_rwb_bufchan_d ;
  logic \writeCTf'lizzieLet49_1_argbuf_rwb_bufchan_r ;
  assign \writeCTf'lizzieLet49_1_argbuf_rwb_r  = ((! \writeCTf'lizzieLet49_1_argbuf_rwb_bufchan_d [0]) || \writeCTf'lizzieLet49_1_argbuf_rwb_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf'lizzieLet49_1_argbuf_rwb_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\writeCTf'lizzieLet49_1_argbuf_rwb_r )
        \writeCTf'lizzieLet49_1_argbuf_rwb_bufchan_d  <= \writeCTf'lizzieLet49_1_argbuf_rwb_d ;
  \Pointer_CTf'_t  \writeCTf'lizzieLet49_1_argbuf_rwb_bufchan_buf ;
  assign \writeCTf'lizzieLet49_1_argbuf_rwb_bufchan_r  = (! \writeCTf'lizzieLet49_1_argbuf_rwb_bufchan_buf [0]);
  assign sca2_1_1_argbuf_d = (\writeCTf'lizzieLet49_1_argbuf_rwb_bufchan_buf [0] ? \writeCTf'lizzieLet49_1_argbuf_rwb_bufchan_buf  :
                              \writeCTf'lizzieLet49_1_argbuf_rwb_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf'lizzieLet49_1_argbuf_rwb_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((sca2_1_1_argbuf_r && \writeCTf'lizzieLet49_1_argbuf_rwb_bufchan_buf [0]))
        \writeCTf'lizzieLet49_1_argbuf_rwb_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! sca2_1_1_argbuf_r) && (! \writeCTf'lizzieLet49_1_argbuf_rwb_bufchan_buf [0])))
        \writeCTf'lizzieLet49_1_argbuf_rwb_bufchan_buf  <= \writeCTf'lizzieLet49_1_argbuf_rwb_bufchan_d ;
  
  /* buf (Ty Pointer_CTf') : (writeCTf'lizzieLet50_1_argbuf,Pointer_CTf') > (writeCTf'lizzieLet50_1_argbuf_rwb,Pointer_CTf') */
  \Pointer_CTf'_t  \writeCTf'lizzieLet50_1_argbuf_bufchan_d ;
  logic \writeCTf'lizzieLet50_1_argbuf_bufchan_r ;
  assign \writeCTf'lizzieLet50_1_argbuf_r  = ((! \writeCTf'lizzieLet50_1_argbuf_bufchan_d [0]) || \writeCTf'lizzieLet50_1_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf'lizzieLet50_1_argbuf_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\writeCTf'lizzieLet50_1_argbuf_r )
        \writeCTf'lizzieLet50_1_argbuf_bufchan_d  <= \writeCTf'lizzieLet50_1_argbuf_d ;
  \Pointer_CTf'_t  \writeCTf'lizzieLet50_1_argbuf_bufchan_buf ;
  assign \writeCTf'lizzieLet50_1_argbuf_bufchan_r  = (! \writeCTf'lizzieLet50_1_argbuf_bufchan_buf [0]);
  assign \writeCTf'lizzieLet50_1_argbuf_rwb_d  = (\writeCTf'lizzieLet50_1_argbuf_bufchan_buf [0] ? \writeCTf'lizzieLet50_1_argbuf_bufchan_buf  :
                                                  \writeCTf'lizzieLet50_1_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf'lizzieLet50_1_argbuf_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((\writeCTf'lizzieLet50_1_argbuf_rwb_r  && \writeCTf'lizzieLet50_1_argbuf_bufchan_buf [0]))
        \writeCTf'lizzieLet50_1_argbuf_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! \writeCTf'lizzieLet50_1_argbuf_rwb_r ) && (! \writeCTf'lizzieLet50_1_argbuf_bufchan_buf [0])))
        \writeCTf'lizzieLet50_1_argbuf_bufchan_buf  <= \writeCTf'lizzieLet50_1_argbuf_bufchan_d ;
  
  /* buf (Ty Pointer_CTf') : (writeCTf'lizzieLet50_1_argbuf_rwb,Pointer_CTf') > (sca1_1_1_argbuf,Pointer_CTf') */
  \Pointer_CTf'_t  \writeCTf'lizzieLet50_1_argbuf_rwb_bufchan_d ;
  logic \writeCTf'lizzieLet50_1_argbuf_rwb_bufchan_r ;
  assign \writeCTf'lizzieLet50_1_argbuf_rwb_r  = ((! \writeCTf'lizzieLet50_1_argbuf_rwb_bufchan_d [0]) || \writeCTf'lizzieLet50_1_argbuf_rwb_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf'lizzieLet50_1_argbuf_rwb_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\writeCTf'lizzieLet50_1_argbuf_rwb_r )
        \writeCTf'lizzieLet50_1_argbuf_rwb_bufchan_d  <= \writeCTf'lizzieLet50_1_argbuf_rwb_d ;
  \Pointer_CTf'_t  \writeCTf'lizzieLet50_1_argbuf_rwb_bufchan_buf ;
  assign \writeCTf'lizzieLet50_1_argbuf_rwb_bufchan_r  = (! \writeCTf'lizzieLet50_1_argbuf_rwb_bufchan_buf [0]);
  assign sca1_1_1_argbuf_d = (\writeCTf'lizzieLet50_1_argbuf_rwb_bufchan_buf [0] ? \writeCTf'lizzieLet50_1_argbuf_rwb_bufchan_buf  :
                              \writeCTf'lizzieLet50_1_argbuf_rwb_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf'lizzieLet50_1_argbuf_rwb_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((sca1_1_1_argbuf_r && \writeCTf'lizzieLet50_1_argbuf_rwb_bufchan_buf [0]))
        \writeCTf'lizzieLet50_1_argbuf_rwb_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! sca1_1_1_argbuf_r) && (! \writeCTf'lizzieLet50_1_argbuf_rwb_bufchan_buf [0])))
        \writeCTf'lizzieLet50_1_argbuf_rwb_bufchan_buf  <= \writeCTf'lizzieLet50_1_argbuf_rwb_bufchan_d ;
  
  /* buf (Ty Pointer_CTf') : (writeCTf'lizzieLet51_1_argbuf,Pointer_CTf') > (writeCTf'lizzieLet51_1_argbuf_rwb,Pointer_CTf') */
  \Pointer_CTf'_t  \writeCTf'lizzieLet51_1_argbuf_bufchan_d ;
  logic \writeCTf'lizzieLet51_1_argbuf_bufchan_r ;
  assign \writeCTf'lizzieLet51_1_argbuf_r  = ((! \writeCTf'lizzieLet51_1_argbuf_bufchan_d [0]) || \writeCTf'lizzieLet51_1_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf'lizzieLet51_1_argbuf_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\writeCTf'lizzieLet51_1_argbuf_r )
        \writeCTf'lizzieLet51_1_argbuf_bufchan_d  <= \writeCTf'lizzieLet51_1_argbuf_d ;
  \Pointer_CTf'_t  \writeCTf'lizzieLet51_1_argbuf_bufchan_buf ;
  assign \writeCTf'lizzieLet51_1_argbuf_bufchan_r  = (! \writeCTf'lizzieLet51_1_argbuf_bufchan_buf [0]);
  assign \writeCTf'lizzieLet51_1_argbuf_rwb_d  = (\writeCTf'lizzieLet51_1_argbuf_bufchan_buf [0] ? \writeCTf'lizzieLet51_1_argbuf_bufchan_buf  :
                                                  \writeCTf'lizzieLet51_1_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf'lizzieLet51_1_argbuf_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((\writeCTf'lizzieLet51_1_argbuf_rwb_r  && \writeCTf'lizzieLet51_1_argbuf_bufchan_buf [0]))
        \writeCTf'lizzieLet51_1_argbuf_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! \writeCTf'lizzieLet51_1_argbuf_rwb_r ) && (! \writeCTf'lizzieLet51_1_argbuf_bufchan_buf [0])))
        \writeCTf'lizzieLet51_1_argbuf_bufchan_buf  <= \writeCTf'lizzieLet51_1_argbuf_bufchan_d ;
  
  /* buf (Ty Pointer_CTf') : (writeCTf'lizzieLet51_1_argbuf_rwb,Pointer_CTf') > (sca0_1_1_argbuf,Pointer_CTf') */
  \Pointer_CTf'_t  \writeCTf'lizzieLet51_1_argbuf_rwb_bufchan_d ;
  logic \writeCTf'lizzieLet51_1_argbuf_rwb_bufchan_r ;
  assign \writeCTf'lizzieLet51_1_argbuf_rwb_r  = ((! \writeCTf'lizzieLet51_1_argbuf_rwb_bufchan_d [0]) || \writeCTf'lizzieLet51_1_argbuf_rwb_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf'lizzieLet51_1_argbuf_rwb_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\writeCTf'lizzieLet51_1_argbuf_rwb_r )
        \writeCTf'lizzieLet51_1_argbuf_rwb_bufchan_d  <= \writeCTf'lizzieLet51_1_argbuf_rwb_d ;
  \Pointer_CTf'_t  \writeCTf'lizzieLet51_1_argbuf_rwb_bufchan_buf ;
  assign \writeCTf'lizzieLet51_1_argbuf_rwb_bufchan_r  = (! \writeCTf'lizzieLet51_1_argbuf_rwb_bufchan_buf [0]);
  assign sca0_1_1_argbuf_d = (\writeCTf'lizzieLet51_1_argbuf_rwb_bufchan_buf [0] ? \writeCTf'lizzieLet51_1_argbuf_rwb_bufchan_buf  :
                              \writeCTf'lizzieLet51_1_argbuf_rwb_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf'lizzieLet51_1_argbuf_rwb_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((sca0_1_1_argbuf_r && \writeCTf'lizzieLet51_1_argbuf_rwb_bufchan_buf [0]))
        \writeCTf'lizzieLet51_1_argbuf_rwb_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! sca0_1_1_argbuf_r) && (! \writeCTf'lizzieLet51_1_argbuf_rwb_bufchan_buf [0])))
        \writeCTf'lizzieLet51_1_argbuf_rwb_bufchan_buf  <= \writeCTf'lizzieLet51_1_argbuf_rwb_bufchan_d ;
  
  /* buf (Ty Pointer_CTf) : (writeCTflizzieLet17_1_1_argbuf,Pointer_CTf) > (writeCTflizzieLet17_1_1_argbuf_rwb,Pointer_CTf) */
  Pointer_CTf_t writeCTflizzieLet17_1_1_argbuf_bufchan_d;
  logic writeCTflizzieLet17_1_1_argbuf_bufchan_r;
  assign writeCTflizzieLet17_1_1_argbuf_r = ((! writeCTflizzieLet17_1_1_argbuf_bufchan_d[0]) || writeCTflizzieLet17_1_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTflizzieLet17_1_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCTflizzieLet17_1_1_argbuf_r)
        writeCTflizzieLet17_1_1_argbuf_bufchan_d <= writeCTflizzieLet17_1_1_argbuf_d;
  Pointer_CTf_t writeCTflizzieLet17_1_1_argbuf_bufchan_buf;
  assign writeCTflizzieLet17_1_1_argbuf_bufchan_r = (! writeCTflizzieLet17_1_1_argbuf_bufchan_buf[0]);
  assign writeCTflizzieLet17_1_1_argbuf_rwb_d = (writeCTflizzieLet17_1_1_argbuf_bufchan_buf[0] ? writeCTflizzieLet17_1_1_argbuf_bufchan_buf :
                                                 writeCTflizzieLet17_1_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTflizzieLet17_1_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeCTflizzieLet17_1_1_argbuf_rwb_r && writeCTflizzieLet17_1_1_argbuf_bufchan_buf[0]))
        writeCTflizzieLet17_1_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeCTflizzieLet17_1_1_argbuf_rwb_r) && (! writeCTflizzieLet17_1_1_argbuf_bufchan_buf[0])))
        writeCTflizzieLet17_1_1_argbuf_bufchan_buf <= writeCTflizzieLet17_1_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CTf) : (writeCTflizzieLet17_1_1_argbuf_rwb,Pointer_CTf) > (sca3_1_argbuf,Pointer_CTf) */
  Pointer_CTf_t writeCTflizzieLet17_1_1_argbuf_rwb_bufchan_d;
  logic writeCTflizzieLet17_1_1_argbuf_rwb_bufchan_r;
  assign writeCTflizzieLet17_1_1_argbuf_rwb_r = ((! writeCTflizzieLet17_1_1_argbuf_rwb_bufchan_d[0]) || writeCTflizzieLet17_1_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTflizzieLet17_1_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCTflizzieLet17_1_1_argbuf_rwb_r)
        writeCTflizzieLet17_1_1_argbuf_rwb_bufchan_d <= writeCTflizzieLet17_1_1_argbuf_rwb_d;
  Pointer_CTf_t writeCTflizzieLet17_1_1_argbuf_rwb_bufchan_buf;
  assign writeCTflizzieLet17_1_1_argbuf_rwb_bufchan_r = (! writeCTflizzieLet17_1_1_argbuf_rwb_bufchan_buf[0]);
  assign sca3_1_argbuf_d = (writeCTflizzieLet17_1_1_argbuf_rwb_bufchan_buf[0] ? writeCTflizzieLet17_1_1_argbuf_rwb_bufchan_buf :
                            writeCTflizzieLet17_1_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTflizzieLet17_1_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((sca3_1_argbuf_r && writeCTflizzieLet17_1_1_argbuf_rwb_bufchan_buf[0]))
        writeCTflizzieLet17_1_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
      else if (((! sca3_1_argbuf_r) && (! writeCTflizzieLet17_1_1_argbuf_rwb_bufchan_buf[0])))
        writeCTflizzieLet17_1_1_argbuf_rwb_bufchan_buf <= writeCTflizzieLet17_1_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CTf) : (writeCTflizzieLet39_1_argbuf,Pointer_CTf) > (writeCTflizzieLet39_1_argbuf_rwb,Pointer_CTf) */
  Pointer_CTf_t writeCTflizzieLet39_1_argbuf_bufchan_d;
  logic writeCTflizzieLet39_1_argbuf_bufchan_r;
  assign writeCTflizzieLet39_1_argbuf_r = ((! writeCTflizzieLet39_1_argbuf_bufchan_d[0]) || writeCTflizzieLet39_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTflizzieLet39_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCTflizzieLet39_1_argbuf_r)
        writeCTflizzieLet39_1_argbuf_bufchan_d <= writeCTflizzieLet39_1_argbuf_d;
  Pointer_CTf_t writeCTflizzieLet39_1_argbuf_bufchan_buf;
  assign writeCTflizzieLet39_1_argbuf_bufchan_r = (! writeCTflizzieLet39_1_argbuf_bufchan_buf[0]);
  assign writeCTflizzieLet39_1_argbuf_rwb_d = (writeCTflizzieLet39_1_argbuf_bufchan_buf[0] ? writeCTflizzieLet39_1_argbuf_bufchan_buf :
                                               writeCTflizzieLet39_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTflizzieLet39_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeCTflizzieLet39_1_argbuf_rwb_r && writeCTflizzieLet39_1_argbuf_bufchan_buf[0]))
        writeCTflizzieLet39_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeCTflizzieLet39_1_argbuf_rwb_r) && (! writeCTflizzieLet39_1_argbuf_bufchan_buf[0])))
        writeCTflizzieLet39_1_argbuf_bufchan_buf <= writeCTflizzieLet39_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CTf) : (writeCTflizzieLet39_1_argbuf_rwb,Pointer_CTf) > (lizzieLet28_1_1_argbuf,Pointer_CTf) */
  Pointer_CTf_t writeCTflizzieLet39_1_argbuf_rwb_bufchan_d;
  logic writeCTflizzieLet39_1_argbuf_rwb_bufchan_r;
  assign writeCTflizzieLet39_1_argbuf_rwb_r = ((! writeCTflizzieLet39_1_argbuf_rwb_bufchan_d[0]) || writeCTflizzieLet39_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTflizzieLet39_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCTflizzieLet39_1_argbuf_rwb_r)
        writeCTflizzieLet39_1_argbuf_rwb_bufchan_d <= writeCTflizzieLet39_1_argbuf_rwb_d;
  Pointer_CTf_t writeCTflizzieLet39_1_argbuf_rwb_bufchan_buf;
  assign writeCTflizzieLet39_1_argbuf_rwb_bufchan_r = (! writeCTflizzieLet39_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet28_1_1_argbuf_d = (writeCTflizzieLet39_1_argbuf_rwb_bufchan_buf[0] ? writeCTflizzieLet39_1_argbuf_rwb_bufchan_buf :
                                     writeCTflizzieLet39_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTflizzieLet39_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet28_1_1_argbuf_r && writeCTflizzieLet39_1_argbuf_rwb_bufchan_buf[0]))
        writeCTflizzieLet39_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet28_1_1_argbuf_r) && (! writeCTflizzieLet39_1_argbuf_rwb_bufchan_buf[0])))
        writeCTflizzieLet39_1_argbuf_rwb_bufchan_buf <= writeCTflizzieLet39_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CTf) : (writeCTflizzieLet44_1_argbuf,Pointer_CTf) > (writeCTflizzieLet44_1_argbuf_rwb,Pointer_CTf) */
  Pointer_CTf_t writeCTflizzieLet44_1_argbuf_bufchan_d;
  logic writeCTflizzieLet44_1_argbuf_bufchan_r;
  assign writeCTflizzieLet44_1_argbuf_r = ((! writeCTflizzieLet44_1_argbuf_bufchan_d[0]) || writeCTflizzieLet44_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTflizzieLet44_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCTflizzieLet44_1_argbuf_r)
        writeCTflizzieLet44_1_argbuf_bufchan_d <= writeCTflizzieLet44_1_argbuf_d;
  Pointer_CTf_t writeCTflizzieLet44_1_argbuf_bufchan_buf;
  assign writeCTflizzieLet44_1_argbuf_bufchan_r = (! writeCTflizzieLet44_1_argbuf_bufchan_buf[0]);
  assign writeCTflizzieLet44_1_argbuf_rwb_d = (writeCTflizzieLet44_1_argbuf_bufchan_buf[0] ? writeCTflizzieLet44_1_argbuf_bufchan_buf :
                                               writeCTflizzieLet44_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTflizzieLet44_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeCTflizzieLet44_1_argbuf_rwb_r && writeCTflizzieLet44_1_argbuf_bufchan_buf[0]))
        writeCTflizzieLet44_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeCTflizzieLet44_1_argbuf_rwb_r) && (! writeCTflizzieLet44_1_argbuf_bufchan_buf[0])))
        writeCTflizzieLet44_1_argbuf_bufchan_buf <= writeCTflizzieLet44_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CTf) : (writeCTflizzieLet44_1_argbuf_rwb,Pointer_CTf) > (sca2_1_argbuf,Pointer_CTf) */
  Pointer_CTf_t writeCTflizzieLet44_1_argbuf_rwb_bufchan_d;
  logic writeCTflizzieLet44_1_argbuf_rwb_bufchan_r;
  assign writeCTflizzieLet44_1_argbuf_rwb_r = ((! writeCTflizzieLet44_1_argbuf_rwb_bufchan_d[0]) || writeCTflizzieLet44_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTflizzieLet44_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCTflizzieLet44_1_argbuf_rwb_r)
        writeCTflizzieLet44_1_argbuf_rwb_bufchan_d <= writeCTflizzieLet44_1_argbuf_rwb_d;
  Pointer_CTf_t writeCTflizzieLet44_1_argbuf_rwb_bufchan_buf;
  assign writeCTflizzieLet44_1_argbuf_rwb_bufchan_r = (! writeCTflizzieLet44_1_argbuf_rwb_bufchan_buf[0]);
  assign sca2_1_argbuf_d = (writeCTflizzieLet44_1_argbuf_rwb_bufchan_buf[0] ? writeCTflizzieLet44_1_argbuf_rwb_bufchan_buf :
                            writeCTflizzieLet44_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTflizzieLet44_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((sca2_1_argbuf_r && writeCTflizzieLet44_1_argbuf_rwb_bufchan_buf[0]))
        writeCTflizzieLet44_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
      else if (((! sca2_1_argbuf_r) && (! writeCTflizzieLet44_1_argbuf_rwb_bufchan_buf[0])))
        writeCTflizzieLet44_1_argbuf_rwb_bufchan_buf <= writeCTflizzieLet44_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CTf) : (writeCTflizzieLet45_1_argbuf,Pointer_CTf) > (writeCTflizzieLet45_1_argbuf_rwb,Pointer_CTf) */
  Pointer_CTf_t writeCTflizzieLet45_1_argbuf_bufchan_d;
  logic writeCTflizzieLet45_1_argbuf_bufchan_r;
  assign writeCTflizzieLet45_1_argbuf_r = ((! writeCTflizzieLet45_1_argbuf_bufchan_d[0]) || writeCTflizzieLet45_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTflizzieLet45_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCTflizzieLet45_1_argbuf_r)
        writeCTflizzieLet45_1_argbuf_bufchan_d <= writeCTflizzieLet45_1_argbuf_d;
  Pointer_CTf_t writeCTflizzieLet45_1_argbuf_bufchan_buf;
  assign writeCTflizzieLet45_1_argbuf_bufchan_r = (! writeCTflizzieLet45_1_argbuf_bufchan_buf[0]);
  assign writeCTflizzieLet45_1_argbuf_rwb_d = (writeCTflizzieLet45_1_argbuf_bufchan_buf[0] ? writeCTflizzieLet45_1_argbuf_bufchan_buf :
                                               writeCTflizzieLet45_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTflizzieLet45_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeCTflizzieLet45_1_argbuf_rwb_r && writeCTflizzieLet45_1_argbuf_bufchan_buf[0]))
        writeCTflizzieLet45_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeCTflizzieLet45_1_argbuf_rwb_r) && (! writeCTflizzieLet45_1_argbuf_bufchan_buf[0])))
        writeCTflizzieLet45_1_argbuf_bufchan_buf <= writeCTflizzieLet45_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CTf) : (writeCTflizzieLet45_1_argbuf_rwb,Pointer_CTf) > (sca1_1_argbuf,Pointer_CTf) */
  Pointer_CTf_t writeCTflizzieLet45_1_argbuf_rwb_bufchan_d;
  logic writeCTflizzieLet45_1_argbuf_rwb_bufchan_r;
  assign writeCTflizzieLet45_1_argbuf_rwb_r = ((! writeCTflizzieLet45_1_argbuf_rwb_bufchan_d[0]) || writeCTflizzieLet45_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTflizzieLet45_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCTflizzieLet45_1_argbuf_rwb_r)
        writeCTflizzieLet45_1_argbuf_rwb_bufchan_d <= writeCTflizzieLet45_1_argbuf_rwb_d;
  Pointer_CTf_t writeCTflizzieLet45_1_argbuf_rwb_bufchan_buf;
  assign writeCTflizzieLet45_1_argbuf_rwb_bufchan_r = (! writeCTflizzieLet45_1_argbuf_rwb_bufchan_buf[0]);
  assign sca1_1_argbuf_d = (writeCTflizzieLet45_1_argbuf_rwb_bufchan_buf[0] ? writeCTflizzieLet45_1_argbuf_rwb_bufchan_buf :
                            writeCTflizzieLet45_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTflizzieLet45_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((sca1_1_argbuf_r && writeCTflizzieLet45_1_argbuf_rwb_bufchan_buf[0]))
        writeCTflizzieLet45_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
      else if (((! sca1_1_argbuf_r) && (! writeCTflizzieLet45_1_argbuf_rwb_bufchan_buf[0])))
        writeCTflizzieLet45_1_argbuf_rwb_bufchan_buf <= writeCTflizzieLet45_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CTf) : (writeCTflizzieLet46_1_argbuf,Pointer_CTf) > (writeCTflizzieLet46_1_argbuf_rwb,Pointer_CTf) */
  Pointer_CTf_t writeCTflizzieLet46_1_argbuf_bufchan_d;
  logic writeCTflizzieLet46_1_argbuf_bufchan_r;
  assign writeCTflizzieLet46_1_argbuf_r = ((! writeCTflizzieLet46_1_argbuf_bufchan_d[0]) || writeCTflizzieLet46_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTflizzieLet46_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCTflizzieLet46_1_argbuf_r)
        writeCTflizzieLet46_1_argbuf_bufchan_d <= writeCTflizzieLet46_1_argbuf_d;
  Pointer_CTf_t writeCTflizzieLet46_1_argbuf_bufchan_buf;
  assign writeCTflizzieLet46_1_argbuf_bufchan_r = (! writeCTflizzieLet46_1_argbuf_bufchan_buf[0]);
  assign writeCTflizzieLet46_1_argbuf_rwb_d = (writeCTflizzieLet46_1_argbuf_bufchan_buf[0] ? writeCTflizzieLet46_1_argbuf_bufchan_buf :
                                               writeCTflizzieLet46_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTflizzieLet46_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeCTflizzieLet46_1_argbuf_rwb_r && writeCTflizzieLet46_1_argbuf_bufchan_buf[0]))
        writeCTflizzieLet46_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeCTflizzieLet46_1_argbuf_rwb_r) && (! writeCTflizzieLet46_1_argbuf_bufchan_buf[0])))
        writeCTflizzieLet46_1_argbuf_bufchan_buf <= writeCTflizzieLet46_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CTf) : (writeCTflizzieLet46_1_argbuf_rwb,Pointer_CTf) > (sca0_1_argbuf,Pointer_CTf) */
  Pointer_CTf_t writeCTflizzieLet46_1_argbuf_rwb_bufchan_d;
  logic writeCTflizzieLet46_1_argbuf_rwb_bufchan_r;
  assign writeCTflizzieLet46_1_argbuf_rwb_r = ((! writeCTflizzieLet46_1_argbuf_rwb_bufchan_d[0]) || writeCTflizzieLet46_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTflizzieLet46_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCTflizzieLet46_1_argbuf_rwb_r)
        writeCTflizzieLet46_1_argbuf_rwb_bufchan_d <= writeCTflizzieLet46_1_argbuf_rwb_d;
  Pointer_CTf_t writeCTflizzieLet46_1_argbuf_rwb_bufchan_buf;
  assign writeCTflizzieLet46_1_argbuf_rwb_bufchan_r = (! writeCTflizzieLet46_1_argbuf_rwb_bufchan_buf[0]);
  assign sca0_1_argbuf_d = (writeCTflizzieLet46_1_argbuf_rwb_bufchan_buf[0] ? writeCTflizzieLet46_1_argbuf_rwb_bufchan_buf :
                            writeCTflizzieLet46_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTflizzieLet46_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((sca0_1_argbuf_r && writeCTflizzieLet46_1_argbuf_rwb_bufchan_buf[0]))
        writeCTflizzieLet46_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
      else if (((! sca0_1_argbuf_r) && (! writeCTflizzieLet46_1_argbuf_rwb_bufchan_buf[0])))
        writeCTflizzieLet46_1_argbuf_rwb_bufchan_buf <= writeCTflizzieLet46_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet10_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet10_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet10_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet10_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet10_1_argbuf_r = ((! writeQTree_BoollizzieLet10_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet10_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet10_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet10_1_argbuf_r)
        writeQTree_BoollizzieLet10_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet10_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet10_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet10_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet10_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet10_1_argbuf_rwb_d = (writeQTree_BoollizzieLet10_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet10_1_argbuf_bufchan_buf :
                                                      writeQTree_BoollizzieLet10_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet10_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet10_1_argbuf_rwb_r && writeQTree_BoollizzieLet10_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet10_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet10_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet10_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet10_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet10_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet10_1_argbuf_rwb,Pointer_QTree_Bool) > (lizzieLet20_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet10_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet10_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet10_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet10_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet10_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet10_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet10_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet10_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet10_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet10_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet10_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet10_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet20_1_argbuf_d = (writeQTree_BoollizzieLet10_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet10_1_argbuf_rwb_bufchan_buf :
                                   writeQTree_BoollizzieLet10_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet10_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                              1'd0};
    else
      if ((lizzieLet20_1_argbuf_r && writeQTree_BoollizzieLet10_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet10_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
      else if (((! lizzieLet20_1_argbuf_r) && (! writeQTree_BoollizzieLet10_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet10_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet10_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet11_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet11_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet11_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet11_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet11_1_argbuf_r = ((! writeQTree_BoollizzieLet11_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet11_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet11_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet11_1_argbuf_r)
        writeQTree_BoollizzieLet11_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet11_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet11_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet11_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet11_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet11_1_argbuf_rwb_d = (writeQTree_BoollizzieLet11_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet11_1_argbuf_bufchan_buf :
                                                      writeQTree_BoollizzieLet11_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet11_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet11_1_argbuf_rwb_r && writeQTree_BoollizzieLet11_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet11_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet11_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet11_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet11_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet11_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet11_1_argbuf_rwb,Pointer_QTree_Bool) > (lizzieLet21_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet11_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet11_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet11_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet11_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet11_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet11_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet11_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet11_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet11_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet11_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet11_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet11_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet21_1_argbuf_d = (writeQTree_BoollizzieLet11_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet11_1_argbuf_rwb_bufchan_buf :
                                   writeQTree_BoollizzieLet11_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet11_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                              1'd0};
    else
      if ((lizzieLet21_1_argbuf_r && writeQTree_BoollizzieLet11_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet11_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
      else if (((! lizzieLet21_1_argbuf_r) && (! writeQTree_BoollizzieLet11_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet11_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet11_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet12_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet12_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet12_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet12_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet12_1_argbuf_r = ((! writeQTree_BoollizzieLet12_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet12_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet12_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet12_1_argbuf_r)
        writeQTree_BoollizzieLet12_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet12_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet12_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet12_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet12_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet12_1_argbuf_rwb_d = (writeQTree_BoollizzieLet12_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet12_1_argbuf_bufchan_buf :
                                                      writeQTree_BoollizzieLet12_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet12_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet12_1_argbuf_rwb_r && writeQTree_BoollizzieLet12_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet12_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet12_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet12_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet12_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet12_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet12_1_argbuf_rwb,Pointer_QTree_Bool) > (lizzieLet22_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet12_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet12_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet12_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet12_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet12_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet12_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet12_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet12_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet12_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet12_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet12_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet12_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet22_1_argbuf_d = (writeQTree_BoollizzieLet12_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet12_1_argbuf_rwb_bufchan_buf :
                                   writeQTree_BoollizzieLet12_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet12_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                              1'd0};
    else
      if ((lizzieLet22_1_argbuf_r && writeQTree_BoollizzieLet12_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet12_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
      else if (((! lizzieLet22_1_argbuf_r) && (! writeQTree_BoollizzieLet12_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet12_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet12_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet13_1_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet13_1_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet13_1_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet13_1_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet13_1_1_argbuf_r = ((! writeQTree_BoollizzieLet13_1_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet13_1_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet13_1_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet13_1_1_argbuf_r)
        writeQTree_BoollizzieLet13_1_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet13_1_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet13_1_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet13_1_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet13_1_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet13_1_1_argbuf_rwb_d = (writeQTree_BoollizzieLet13_1_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet13_1_1_argbuf_bufchan_buf :
                                                        writeQTree_BoollizzieLet13_1_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet13_1_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet13_1_1_argbuf_rwb_r && writeQTree_BoollizzieLet13_1_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet13_1_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet13_1_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet13_1_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet13_1_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet13_1_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet13_1_1_argbuf_rwb,Pointer_QTree_Bool) > (lizzieLet23_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet13_1_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet13_1_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet13_1_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet13_1_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet13_1_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet13_1_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                              1'd0};
    else
      if (writeQTree_BoollizzieLet13_1_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet13_1_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet13_1_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet13_1_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet13_1_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet13_1_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet23_1_argbuf_d = (writeQTree_BoollizzieLet13_1_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet13_1_1_argbuf_rwb_bufchan_buf :
                                   writeQTree_BoollizzieLet13_1_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet13_1_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
    else
      if ((lizzieLet23_1_argbuf_r && writeQTree_BoollizzieLet13_1_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet13_1_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                  1'd0};
      else if (((! lizzieLet23_1_argbuf_r) && (! writeQTree_BoollizzieLet13_1_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet13_1_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet13_1_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet15_1_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet15_1_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet15_1_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet15_1_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet15_1_1_argbuf_r = ((! writeQTree_BoollizzieLet15_1_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet15_1_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet15_1_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet15_1_1_argbuf_r)
        writeQTree_BoollizzieLet15_1_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet15_1_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet15_1_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet15_1_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet15_1_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet15_1_1_argbuf_rwb_d = (writeQTree_BoollizzieLet15_1_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet15_1_1_argbuf_bufchan_buf :
                                                        writeQTree_BoollizzieLet15_1_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet15_1_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet15_1_1_argbuf_rwb_r && writeQTree_BoollizzieLet15_1_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet15_1_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet15_1_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet15_1_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet15_1_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet15_1_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet15_1_1_argbuf_rwb,Pointer_QTree_Bool) > (lizzieLet24_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet15_1_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet15_1_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet15_1_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet15_1_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet15_1_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet15_1_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                              1'd0};
    else
      if (writeQTree_BoollizzieLet15_1_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet15_1_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet15_1_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet15_1_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet15_1_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet15_1_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet24_1_argbuf_d = (writeQTree_BoollizzieLet15_1_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet15_1_1_argbuf_rwb_bufchan_buf :
                                   writeQTree_BoollizzieLet15_1_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet15_1_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
    else
      if ((lizzieLet24_1_argbuf_r && writeQTree_BoollizzieLet15_1_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet15_1_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                  1'd0};
      else if (((! lizzieLet24_1_argbuf_r) && (! writeQTree_BoollizzieLet15_1_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet15_1_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet15_1_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet16_1_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet16_1_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet16_1_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet16_1_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet16_1_1_argbuf_r = ((! writeQTree_BoollizzieLet16_1_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet16_1_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet16_1_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet16_1_1_argbuf_r)
        writeQTree_BoollizzieLet16_1_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet16_1_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet16_1_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet16_1_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet16_1_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet16_1_1_argbuf_rwb_d = (writeQTree_BoollizzieLet16_1_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet16_1_1_argbuf_bufchan_buf :
                                                        writeQTree_BoollizzieLet16_1_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet16_1_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet16_1_1_argbuf_rwb_r && writeQTree_BoollizzieLet16_1_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet16_1_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet16_1_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet16_1_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet16_1_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet16_1_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet16_1_1_argbuf_rwb,Pointer_QTree_Bool) > (lizzieLet25_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet16_1_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet16_1_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet16_1_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet16_1_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet16_1_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet16_1_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                              1'd0};
    else
      if (writeQTree_BoollizzieLet16_1_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet16_1_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet16_1_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet16_1_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet16_1_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet16_1_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet25_1_argbuf_d = (writeQTree_BoollizzieLet16_1_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet16_1_1_argbuf_rwb_bufchan_buf :
                                   writeQTree_BoollizzieLet16_1_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet16_1_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
    else
      if ((lizzieLet25_1_argbuf_r && writeQTree_BoollizzieLet16_1_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet16_1_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                  1'd0};
      else if (((! lizzieLet25_1_argbuf_r) && (! writeQTree_BoollizzieLet16_1_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet16_1_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet16_1_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet18_1_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet18_1_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet18_1_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet18_1_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet18_1_1_argbuf_r = ((! writeQTree_BoollizzieLet18_1_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet18_1_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet18_1_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet18_1_1_argbuf_r)
        writeQTree_BoollizzieLet18_1_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet18_1_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet18_1_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet18_1_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet18_1_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet18_1_1_argbuf_rwb_d = (writeQTree_BoollizzieLet18_1_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet18_1_1_argbuf_bufchan_buf :
                                                        writeQTree_BoollizzieLet18_1_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet18_1_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet18_1_1_argbuf_rwb_r && writeQTree_BoollizzieLet18_1_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet18_1_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet18_1_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet18_1_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet18_1_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet18_1_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet18_1_1_argbuf_rwb,Pointer_QTree_Bool) > (lizzieLet26_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet18_1_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet18_1_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet18_1_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet18_1_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet18_1_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet18_1_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                              1'd0};
    else
      if (writeQTree_BoollizzieLet18_1_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet18_1_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet18_1_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet18_1_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet18_1_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet18_1_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet26_1_argbuf_d = (writeQTree_BoollizzieLet18_1_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet18_1_1_argbuf_rwb_bufchan_buf :
                                   writeQTree_BoollizzieLet18_1_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet18_1_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
    else
      if ((lizzieLet26_1_argbuf_r && writeQTree_BoollizzieLet18_1_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet18_1_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                  1'd0};
      else if (((! lizzieLet26_1_argbuf_r) && (! writeQTree_BoollizzieLet18_1_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet18_1_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet18_1_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet19_2_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet19_2_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet19_2_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet19_2_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet19_2_1_argbuf_r = ((! writeQTree_BoollizzieLet19_2_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet19_2_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet19_2_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet19_2_1_argbuf_r)
        writeQTree_BoollizzieLet19_2_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet19_2_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet19_2_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet19_2_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet19_2_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet19_2_1_argbuf_rwb_d = (writeQTree_BoollizzieLet19_2_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet19_2_1_argbuf_bufchan_buf :
                                                        writeQTree_BoollizzieLet19_2_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet19_2_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet19_2_1_argbuf_rwb_r && writeQTree_BoollizzieLet19_2_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet19_2_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet19_2_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet19_2_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet19_2_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet19_2_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet19_2_1_argbuf_rwb,Pointer_QTree_Bool) > (lizzieLet27_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet19_2_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet19_2_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet19_2_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet19_2_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet19_2_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet19_2_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                              1'd0};
    else
      if (writeQTree_BoollizzieLet19_2_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet19_2_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet19_2_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet19_2_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet19_2_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet19_2_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet27_1_argbuf_d = (writeQTree_BoollizzieLet19_2_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet19_2_1_argbuf_rwb_bufchan_buf :
                                   writeQTree_BoollizzieLet19_2_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet19_2_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
    else
      if ((lizzieLet27_1_argbuf_r && writeQTree_BoollizzieLet19_2_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet19_2_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                  1'd0};
      else if (((! lizzieLet27_1_argbuf_r) && (! writeQTree_BoollizzieLet19_2_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet19_2_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet19_2_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet1_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet1_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet1_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet1_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet1_1_argbuf_r = ((! writeQTree_BoollizzieLet1_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet1_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet1_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet1_1_argbuf_r)
        writeQTree_BoollizzieLet1_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet1_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet1_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet1_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet1_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet1_1_argbuf_rwb_d = (writeQTree_BoollizzieLet1_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet1_1_argbuf_bufchan_buf :
                                                     writeQTree_BoollizzieLet1_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet1_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet1_1_argbuf_rwb_r && writeQTree_BoollizzieLet1_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet1_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet1_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet1_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet1_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet1_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet1_1_argbuf_rwb,Pointer_QTree_Bool) > (lizzieLet13_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet1_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet1_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet1_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet1_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet1_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet1_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet1_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet1_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet1_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet1_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet1_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet1_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet13_1_argbuf_d = (writeQTree_BoollizzieLet1_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet1_1_argbuf_rwb_bufchan_buf :
                                   writeQTree_BoollizzieLet1_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet1_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((lizzieLet13_1_argbuf_r && writeQTree_BoollizzieLet1_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet1_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! lizzieLet13_1_argbuf_r) && (! writeQTree_BoollizzieLet1_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet1_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet1_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet22_1_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet22_1_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet22_1_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet22_1_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet22_1_1_argbuf_r = ((! writeQTree_BoollizzieLet22_1_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet22_1_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet22_1_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet22_1_1_argbuf_r)
        writeQTree_BoollizzieLet22_1_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet22_1_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet22_1_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet22_1_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet22_1_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet22_1_1_argbuf_rwb_d = (writeQTree_BoollizzieLet22_1_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet22_1_1_argbuf_bufchan_buf :
                                                        writeQTree_BoollizzieLet22_1_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet22_1_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet22_1_1_argbuf_rwb_r && writeQTree_BoollizzieLet22_1_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet22_1_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet22_1_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet22_1_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet22_1_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet22_1_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet22_1_1_argbuf_rwb,Pointer_QTree_Bool) > (lizzieLet6_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet22_1_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet22_1_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet22_1_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet22_1_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet22_1_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet22_1_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                              1'd0};
    else
      if (writeQTree_BoollizzieLet22_1_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet22_1_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet22_1_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet22_1_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet22_1_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet22_1_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet6_1_1_argbuf_d = (writeQTree_BoollizzieLet22_1_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet22_1_1_argbuf_rwb_bufchan_buf :
                                    writeQTree_BoollizzieLet22_1_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet22_1_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
    else
      if ((lizzieLet6_1_1_argbuf_r && writeQTree_BoollizzieLet22_1_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet22_1_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                  1'd0};
      else if (((! lizzieLet6_1_1_argbuf_r) && (! writeQTree_BoollizzieLet22_1_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet22_1_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet22_1_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet25_1_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet25_1_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet25_1_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet25_1_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet25_1_1_argbuf_r = ((! writeQTree_BoollizzieLet25_1_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet25_1_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet25_1_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet25_1_1_argbuf_r)
        writeQTree_BoollizzieLet25_1_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet25_1_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet25_1_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet25_1_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet25_1_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet25_1_1_argbuf_rwb_d = (writeQTree_BoollizzieLet25_1_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet25_1_1_argbuf_bufchan_buf :
                                                        writeQTree_BoollizzieLet25_1_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet25_1_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet25_1_1_argbuf_rwb_r && writeQTree_BoollizzieLet25_1_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet25_1_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet25_1_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet25_1_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet25_1_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet25_1_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet25_1_1_argbuf_rwb,Pointer_QTree_Bool) > (lizzieLet7_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet25_1_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet25_1_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet25_1_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet25_1_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet25_1_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet25_1_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                              1'd0};
    else
      if (writeQTree_BoollizzieLet25_1_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet25_1_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet25_1_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet25_1_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet25_1_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet25_1_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet7_1_1_argbuf_d = (writeQTree_BoollizzieLet25_1_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet25_1_1_argbuf_rwb_bufchan_buf :
                                    writeQTree_BoollizzieLet25_1_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet25_1_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
    else
      if ((lizzieLet7_1_1_argbuf_r && writeQTree_BoollizzieLet25_1_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet25_1_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                  1'd0};
      else if (((! lizzieLet7_1_1_argbuf_r) && (! writeQTree_BoollizzieLet25_1_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet25_1_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet25_1_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet26_1_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet26_1_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet26_1_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet26_1_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet26_1_1_argbuf_r = ((! writeQTree_BoollizzieLet26_1_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet26_1_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet26_1_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet26_1_1_argbuf_r)
        writeQTree_BoollizzieLet26_1_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet26_1_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet26_1_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet26_1_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet26_1_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet26_1_1_argbuf_rwb_d = (writeQTree_BoollizzieLet26_1_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet26_1_1_argbuf_bufchan_buf :
                                                        writeQTree_BoollizzieLet26_1_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet26_1_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet26_1_1_argbuf_rwb_r && writeQTree_BoollizzieLet26_1_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet26_1_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet26_1_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet26_1_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet26_1_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet26_1_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet26_1_1_argbuf_rwb,Pointer_QTree_Bool) > (lizzieLet8_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet26_1_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet26_1_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet26_1_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet26_1_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet26_1_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet26_1_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                              1'd0};
    else
      if (writeQTree_BoollizzieLet26_1_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet26_1_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet26_1_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet26_1_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet26_1_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet26_1_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet8_1_argbuf_d = (writeQTree_BoollizzieLet26_1_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet26_1_1_argbuf_rwb_bufchan_buf :
                                  writeQTree_BoollizzieLet26_1_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet26_1_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
    else
      if ((lizzieLet8_1_argbuf_r && writeQTree_BoollizzieLet26_1_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet26_1_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                  1'd0};
      else if (((! lizzieLet8_1_argbuf_r) && (! writeQTree_BoollizzieLet26_1_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet26_1_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet26_1_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet28_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet28_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet28_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet28_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet28_1_argbuf_r = ((! writeQTree_BoollizzieLet28_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet28_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet28_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet28_1_argbuf_r)
        writeQTree_BoollizzieLet28_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet28_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet28_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet28_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet28_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet28_1_argbuf_rwb_d = (writeQTree_BoollizzieLet28_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet28_1_argbuf_bufchan_buf :
                                                      writeQTree_BoollizzieLet28_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet28_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet28_1_argbuf_rwb_r && writeQTree_BoollizzieLet28_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet28_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet28_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet28_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet28_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet28_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet28_1_argbuf_rwb,Pointer_QTree_Bool) > (lizzieLet9_2_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet28_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet28_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet28_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet28_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet28_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet28_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet28_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet28_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet28_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet28_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet28_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet28_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet9_2_1_argbuf_d = (writeQTree_BoollizzieLet28_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet28_1_argbuf_rwb_bufchan_buf :
                                    writeQTree_BoollizzieLet28_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet28_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                              1'd0};
    else
      if ((lizzieLet9_2_1_argbuf_r && writeQTree_BoollizzieLet28_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet28_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
      else if (((! lizzieLet9_2_1_argbuf_r) && (! writeQTree_BoollizzieLet28_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet28_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet28_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet30_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet30_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet30_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet30_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet30_1_argbuf_r = ((! writeQTree_BoollizzieLet30_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet30_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet30_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet30_1_argbuf_r)
        writeQTree_BoollizzieLet30_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet30_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet30_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet30_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet30_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet30_1_argbuf_rwb_d = (writeQTree_BoollizzieLet30_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet30_1_argbuf_bufchan_buf :
                                                      writeQTree_BoollizzieLet30_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet30_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet30_1_argbuf_rwb_r && writeQTree_BoollizzieLet30_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet30_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet30_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet30_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet30_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet30_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet30_1_argbuf_rwb,Pointer_QTree_Bool) > (lizzieLet10_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet30_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet30_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet30_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet30_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet30_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet30_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet30_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet30_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet30_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet30_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet30_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet30_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet10_1_1_argbuf_d = (writeQTree_BoollizzieLet30_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet30_1_argbuf_rwb_bufchan_buf :
                                     writeQTree_BoollizzieLet30_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet30_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                              1'd0};
    else
      if ((lizzieLet10_1_1_argbuf_r && writeQTree_BoollizzieLet30_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet30_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
      else if (((! lizzieLet10_1_1_argbuf_r) && (! writeQTree_BoollizzieLet30_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet30_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet30_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet31_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet31_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet31_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet31_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet31_1_argbuf_r = ((! writeQTree_BoollizzieLet31_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet31_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet31_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet31_1_argbuf_r)
        writeQTree_BoollizzieLet31_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet31_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet31_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet31_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet31_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet31_1_argbuf_rwb_d = (writeQTree_BoollizzieLet31_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet31_1_argbuf_bufchan_buf :
                                                      writeQTree_BoollizzieLet31_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet31_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet31_1_argbuf_rwb_r && writeQTree_BoollizzieLet31_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet31_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet31_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet31_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet31_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet31_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet31_1_argbuf_rwb,Pointer_QTree_Bool) > (lizzieLet11_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet31_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet31_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet31_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet31_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet31_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet31_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet31_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet31_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet31_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet31_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet31_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet31_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet11_1_1_argbuf_d = (writeQTree_BoollizzieLet31_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet31_1_argbuf_rwb_bufchan_buf :
                                     writeQTree_BoollizzieLet31_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet31_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                              1'd0};
    else
      if ((lizzieLet11_1_1_argbuf_r && writeQTree_BoollizzieLet31_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet31_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
      else if (((! lizzieLet11_1_1_argbuf_r) && (! writeQTree_BoollizzieLet31_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet31_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet31_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet33_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet33_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet33_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet33_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet33_1_argbuf_r = ((! writeQTree_BoollizzieLet33_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet33_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet33_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet33_1_argbuf_r)
        writeQTree_BoollizzieLet33_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet33_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet33_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet33_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet33_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet33_1_argbuf_rwb_d = (writeQTree_BoollizzieLet33_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet33_1_argbuf_bufchan_buf :
                                                      writeQTree_BoollizzieLet33_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet33_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet33_1_argbuf_rwb_r && writeQTree_BoollizzieLet33_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet33_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet33_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet33_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet33_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet33_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet33_1_argbuf_rwb,Pointer_QTree_Bool) > (lizzieLet1_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet33_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet33_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet33_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet33_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet33_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet33_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet33_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet33_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet33_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet33_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet33_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet33_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet1_1_1_argbuf_d = (writeQTree_BoollizzieLet33_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet33_1_argbuf_rwb_bufchan_buf :
                                    writeQTree_BoollizzieLet33_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet33_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                              1'd0};
    else
      if ((lizzieLet1_1_1_argbuf_r && writeQTree_BoollizzieLet33_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet33_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
      else if (((! lizzieLet1_1_1_argbuf_r) && (! writeQTree_BoollizzieLet33_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet33_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet33_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet35_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet35_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet35_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet35_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet35_1_argbuf_r = ((! writeQTree_BoollizzieLet35_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet35_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet35_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet35_1_argbuf_r)
        writeQTree_BoollizzieLet35_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet35_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet35_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet35_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet35_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet35_1_argbuf_rwb_d = (writeQTree_BoollizzieLet35_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet35_1_argbuf_bufchan_buf :
                                                      writeQTree_BoollizzieLet35_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet35_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet35_1_argbuf_rwb_r && writeQTree_BoollizzieLet35_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet35_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet35_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet35_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet35_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet35_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet35_1_argbuf_rwb,Pointer_QTree_Bool) > (lizzieLet2_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet35_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet35_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet35_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet35_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet35_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet35_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet35_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet35_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet35_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet35_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet35_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet35_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet2_1_1_argbuf_d = (writeQTree_BoollizzieLet35_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet35_1_argbuf_rwb_bufchan_buf :
                                    writeQTree_BoollizzieLet35_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet35_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                              1'd0};
    else
      if ((lizzieLet2_1_1_argbuf_r && writeQTree_BoollizzieLet35_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet35_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
      else if (((! lizzieLet2_1_1_argbuf_r) && (! writeQTree_BoollizzieLet35_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet35_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet35_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet36_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet36_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet36_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet36_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet36_1_argbuf_r = ((! writeQTree_BoollizzieLet36_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet36_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet36_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet36_1_argbuf_r)
        writeQTree_BoollizzieLet36_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet36_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet36_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet36_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet36_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet36_1_argbuf_rwb_d = (writeQTree_BoollizzieLet36_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet36_1_argbuf_bufchan_buf :
                                                      writeQTree_BoollizzieLet36_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet36_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet36_1_argbuf_rwb_r && writeQTree_BoollizzieLet36_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet36_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet36_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet36_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet36_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet36_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet36_1_argbuf_rwb,Pointer_QTree_Bool) > (lizzieLet3_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet36_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet36_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet36_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet36_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet36_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet36_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet36_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet36_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet36_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet36_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet36_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet36_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet3_1_1_argbuf_d = (writeQTree_BoollizzieLet36_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet36_1_argbuf_rwb_bufchan_buf :
                                    writeQTree_BoollizzieLet36_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet36_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                              1'd0};
    else
      if ((lizzieLet3_1_1_argbuf_r && writeQTree_BoollizzieLet36_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet36_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
      else if (((! lizzieLet3_1_1_argbuf_r) && (! writeQTree_BoollizzieLet36_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet36_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet36_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet38_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet38_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet38_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet38_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet38_1_argbuf_r = ((! writeQTree_BoollizzieLet38_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet38_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet38_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet38_1_argbuf_r)
        writeQTree_BoollizzieLet38_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet38_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet38_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet38_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet38_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet38_1_argbuf_rwb_d = (writeQTree_BoollizzieLet38_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet38_1_argbuf_bufchan_buf :
                                                      writeQTree_BoollizzieLet38_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet38_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet38_1_argbuf_rwb_r && writeQTree_BoollizzieLet38_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet38_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet38_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet38_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet38_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet38_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet38_1_argbuf_rwb,Pointer_QTree_Bool) > (lizzieLet4_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet38_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet38_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet38_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet38_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet38_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet38_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet38_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet38_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet38_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet38_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet38_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet38_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet4_1_1_argbuf_d = (writeQTree_BoollizzieLet38_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet38_1_argbuf_rwb_bufchan_buf :
                                    writeQTree_BoollizzieLet38_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet38_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                              1'd0};
    else
      if ((lizzieLet4_1_1_argbuf_r && writeQTree_BoollizzieLet38_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet38_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
      else if (((! lizzieLet4_1_1_argbuf_r) && (! writeQTree_BoollizzieLet38_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet38_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet38_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet42_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet42_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet42_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet42_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet42_1_argbuf_r = ((! writeQTree_BoollizzieLet42_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet42_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet42_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet42_1_argbuf_r)
        writeQTree_BoollizzieLet42_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet42_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet42_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet42_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet42_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet42_1_argbuf_rwb_d = (writeQTree_BoollizzieLet42_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet42_1_argbuf_bufchan_buf :
                                                      writeQTree_BoollizzieLet42_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet42_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet42_1_argbuf_rwb_r && writeQTree_BoollizzieLet42_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet42_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet42_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet42_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet42_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet42_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet47_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet47_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet47_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet47_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet47_1_argbuf_r = ((! writeQTree_BoollizzieLet47_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet47_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet47_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet47_1_argbuf_r)
        writeQTree_BoollizzieLet47_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet47_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet47_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet47_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet47_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet47_1_argbuf_rwb_d = (writeQTree_BoollizzieLet47_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet47_1_argbuf_bufchan_buf :
                                                      writeQTree_BoollizzieLet47_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet47_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet47_1_argbuf_rwb_r && writeQTree_BoollizzieLet47_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet47_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet47_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet47_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet47_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet47_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet47_1_argbuf_rwb,Pointer_QTree_Bool) > (contRet_0_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet47_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet47_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet47_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet47_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet47_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet47_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet47_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet47_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet47_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet47_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet47_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet47_1_argbuf_rwb_bufchan_buf[0]);
  assign contRet_0_1_argbuf_d = (writeQTree_BoollizzieLet47_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet47_1_argbuf_rwb_bufchan_buf :
                                 writeQTree_BoollizzieLet47_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet47_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                              1'd0};
    else
      if ((contRet_0_1_argbuf_r && writeQTree_BoollizzieLet47_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet47_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
      else if (((! contRet_0_1_argbuf_r) && (! writeQTree_BoollizzieLet47_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet47_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet47_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet4_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet4_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet4_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet4_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet4_1_argbuf_r = ((! writeQTree_BoollizzieLet4_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet4_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet4_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet4_1_argbuf_r)
        writeQTree_BoollizzieLet4_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet4_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet4_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet4_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet4_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet4_1_argbuf_rwb_d = (writeQTree_BoollizzieLet4_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet4_1_argbuf_bufchan_buf :
                                                     writeQTree_BoollizzieLet4_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet4_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet4_1_argbuf_rwb_r && writeQTree_BoollizzieLet4_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet4_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet4_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet4_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet4_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet4_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet4_1_argbuf_rwb,Pointer_QTree_Bool) > (lizzieLet15_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet4_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet4_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet4_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet4_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet4_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet4_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet4_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet4_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet4_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet4_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet4_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet4_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet15_1_argbuf_d = (writeQTree_BoollizzieLet4_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet4_1_argbuf_rwb_bufchan_buf :
                                   writeQTree_BoollizzieLet4_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet4_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((lizzieLet15_1_argbuf_r && writeQTree_BoollizzieLet4_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet4_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! lizzieLet15_1_argbuf_r) && (! writeQTree_BoollizzieLet4_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet4_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet4_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet52_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet52_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet52_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet52_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet52_1_argbuf_r = ((! writeQTree_BoollizzieLet52_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet52_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet52_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet52_1_argbuf_r)
        writeQTree_BoollizzieLet52_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet52_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet52_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet52_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet52_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet52_1_argbuf_rwb_d = (writeQTree_BoollizzieLet52_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet52_1_argbuf_bufchan_buf :
                                                      writeQTree_BoollizzieLet52_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet52_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet52_1_argbuf_rwb_r && writeQTree_BoollizzieLet52_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet52_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet52_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet52_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet52_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet52_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet52_1_argbuf_rwb,Pointer_QTree_Bool) > (contRet_0_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet52_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet52_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet52_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet52_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet52_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet52_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet52_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet52_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet52_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet52_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet52_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet52_1_argbuf_rwb_bufchan_buf[0]);
  assign contRet_0_1_1_argbuf_d = (writeQTree_BoollizzieLet52_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet52_1_argbuf_rwb_bufchan_buf :
                                   writeQTree_BoollizzieLet52_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet52_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                              1'd0};
    else
      if ((contRet_0_1_1_argbuf_r && writeQTree_BoollizzieLet52_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet52_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
      else if (((! contRet_0_1_1_argbuf_r) && (! writeQTree_BoollizzieLet52_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet52_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet52_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet57_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet57_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet57_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet57_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet57_1_argbuf_r = ((! writeQTree_BoollizzieLet57_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet57_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet57_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet57_1_argbuf_r)
        writeQTree_BoollizzieLet57_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet57_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet57_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet57_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet57_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet57_1_argbuf_rwb_d = (writeQTree_BoollizzieLet57_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet57_1_argbuf_bufchan_buf :
                                                      writeQTree_BoollizzieLet57_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet57_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet57_1_argbuf_rwb_r && writeQTree_BoollizzieLet57_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet57_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet57_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet57_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet57_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet57_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet57_1_argbuf_rwb,Pointer_QTree_Bool) > (contRet_0_2_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet57_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet57_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet57_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet57_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet57_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet57_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet57_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet57_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet57_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet57_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet57_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet57_1_argbuf_rwb_bufchan_buf[0]);
  assign contRet_0_2_1_argbuf_d = (writeQTree_BoollizzieLet57_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet57_1_argbuf_rwb_bufchan_buf :
                                   writeQTree_BoollizzieLet57_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet57_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                              1'd0};
    else
      if ((contRet_0_2_1_argbuf_r && writeQTree_BoollizzieLet57_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet57_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
      else if (((! contRet_0_2_1_argbuf_r) && (! writeQTree_BoollizzieLet57_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet57_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet57_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet5_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet5_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet5_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet5_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet5_1_argbuf_r = ((! writeQTree_BoollizzieLet5_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet5_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet5_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet5_1_argbuf_r)
        writeQTree_BoollizzieLet5_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet5_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet5_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet5_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet5_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet5_1_argbuf_rwb_d = (writeQTree_BoollizzieLet5_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet5_1_argbuf_bufchan_buf :
                                                     writeQTree_BoollizzieLet5_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet5_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet5_1_argbuf_rwb_r && writeQTree_BoollizzieLet5_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet5_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet5_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet5_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet5_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet5_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet5_1_argbuf_rwb,Pointer_QTree_Bool) > (lizzieLet16_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet5_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet5_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet5_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet5_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet5_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet5_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet5_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet5_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet5_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet5_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet5_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet5_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet16_1_argbuf_d = (writeQTree_BoollizzieLet5_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet5_1_argbuf_rwb_bufchan_buf :
                                   writeQTree_BoollizzieLet5_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet5_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((lizzieLet16_1_argbuf_r && writeQTree_BoollizzieLet5_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet5_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! lizzieLet16_1_argbuf_r) && (! writeQTree_BoollizzieLet5_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet5_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet5_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet6_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet6_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet6_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet6_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet6_1_argbuf_r = ((! writeQTree_BoollizzieLet6_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet6_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet6_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet6_1_argbuf_r)
        writeQTree_BoollizzieLet6_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet6_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet6_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet6_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet6_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet6_1_argbuf_rwb_d = (writeQTree_BoollizzieLet6_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet6_1_argbuf_bufchan_buf :
                                                     writeQTree_BoollizzieLet6_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet6_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet6_1_argbuf_rwb_r && writeQTree_BoollizzieLet6_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet6_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet6_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet6_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet6_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet6_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet6_1_argbuf_rwb,Pointer_QTree_Bool) > (lizzieLet17_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet6_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet6_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet6_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet6_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet6_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet6_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet6_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet6_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet6_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet6_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet6_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet6_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet17_1_argbuf_d = (writeQTree_BoollizzieLet6_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet6_1_argbuf_rwb_bufchan_buf :
                                   writeQTree_BoollizzieLet6_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet6_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((lizzieLet17_1_argbuf_r && writeQTree_BoollizzieLet6_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet6_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! lizzieLet17_1_argbuf_r) && (! writeQTree_BoollizzieLet6_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet6_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet6_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet7_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet7_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet7_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet7_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet7_1_argbuf_r = ((! writeQTree_BoollizzieLet7_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet7_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet7_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet7_1_argbuf_r)
        writeQTree_BoollizzieLet7_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet7_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet7_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet7_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet7_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet7_1_argbuf_rwb_d = (writeQTree_BoollizzieLet7_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet7_1_argbuf_bufchan_buf :
                                                     writeQTree_BoollizzieLet7_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet7_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet7_1_argbuf_rwb_r && writeQTree_BoollizzieLet7_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet7_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet7_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet7_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet7_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet7_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet7_1_argbuf_rwb,Pointer_QTree_Bool) > (lizzieLet18_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet7_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet7_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet7_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet7_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet7_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet7_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet7_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet7_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet7_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet7_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet7_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet7_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet18_1_argbuf_d = (writeQTree_BoollizzieLet7_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet7_1_argbuf_rwb_bufchan_buf :
                                   writeQTree_BoollizzieLet7_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet7_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((lizzieLet18_1_argbuf_r && writeQTree_BoollizzieLet7_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet7_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! lizzieLet18_1_argbuf_r) && (! writeQTree_BoollizzieLet7_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet7_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet7_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet9_1_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet9_1_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet9_1_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet9_1_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet9_1_1_argbuf_r = ((! writeQTree_BoollizzieLet9_1_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet9_1_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet9_1_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet9_1_1_argbuf_r)
        writeQTree_BoollizzieLet9_1_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet9_1_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet9_1_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet9_1_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet9_1_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet9_1_1_argbuf_rwb_d = (writeQTree_BoollizzieLet9_1_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet9_1_1_argbuf_bufchan_buf :
                                                       writeQTree_BoollizzieLet9_1_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet9_1_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet9_1_1_argbuf_rwb_r && writeQTree_BoollizzieLet9_1_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet9_1_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet9_1_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet9_1_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet9_1_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet9_1_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet9_1_1_argbuf_rwb,Pointer_QTree_Bool) > (lizzieLet19_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet9_1_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet9_1_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet9_1_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet9_1_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet9_1_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet9_1_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                             1'd0};
    else
      if (writeQTree_BoollizzieLet9_1_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet9_1_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet9_1_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet9_1_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet9_1_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet9_1_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet19_1_1_argbuf_d = (writeQTree_BoollizzieLet9_1_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet9_1_1_argbuf_rwb_bufchan_buf :
                                     writeQTree_BoollizzieLet9_1_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet9_1_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
    else
      if ((lizzieLet19_1_1_argbuf_r && writeQTree_BoollizzieLet9_1_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet9_1_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                 1'd0};
      else if (((! lizzieLet19_1_1_argbuf_r) && (! writeQTree_BoollizzieLet9_1_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet9_1_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet9_1_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet9_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet9_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet9_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet9_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet9_1_argbuf_r = ((! writeQTree_BoollizzieLet9_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet9_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet9_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet9_1_argbuf_r)
        writeQTree_BoollizzieLet9_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet9_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet9_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet9_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet9_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet9_1_argbuf_rwb_d = (writeQTree_BoollizzieLet9_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet9_1_argbuf_bufchan_buf :
                                                     writeQTree_BoollizzieLet9_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet9_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet9_1_argbuf_rwb_r && writeQTree_BoollizzieLet9_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet9_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet9_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet9_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet9_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet9_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet9_1_argbuf_rwb,Pointer_QTree_Bool) > (lizzieLet19_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet9_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet9_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet9_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet9_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet9_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet9_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet9_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet9_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet9_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet9_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet9_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet9_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet19_1_argbuf_d = (writeQTree_BoollizzieLet9_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet9_1_argbuf_rwb_bufchan_buf :
                                   writeQTree_BoollizzieLet9_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet9_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((lizzieLet19_1_argbuf_r && writeQTree_BoollizzieLet9_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet9_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! lizzieLet19_1_argbuf_r) && (! writeQTree_BoollizzieLet9_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet9_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet9_1_argbuf_rwb_bufchan_d;
endmodule