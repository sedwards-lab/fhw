`timescale 1ns/1ns
package mAddAdd_package ;
    typedef logic [4:0] \Int4#_t ;
    typedef logic [8:0] \Int8#_t ;
    typedef logic [16:0] \Int16#_t ;
    typedef logic [32:0] \Int#_t ;
    typedef logic [4:0] \Word4#_t ;
    typedef logic [8:0] \Word8#_t ;
    typedef logic [16:0] \Word16#_t ;
    typedef logic [32:0] \Word#_t ;
    typedef logic [1:0] C2_t;
    function C2_t C1_2_dc (logic valid);
      begin
        C1_2_dc = 2'bx;
        C1_2_dc[0:0] = valid;
        C1_2_dc[1:1] = 1'd0;
      end
    endfunction
    function C2_t C2_2_dc (logic valid);
      begin
        C2_2_dc = 2'bx;
        C2_2_dc[0:0] = valid;
        C2_2_dc[1:1] = 1'd1;
      end
    endfunction
    typedef logic [6:0] C35_t;
    function C35_t C1_35_dc (logic valid);
      begin
        C1_35_dc = 7'bx;
        C1_35_dc[0:0] = valid;
        C1_35_dc[6:1] = 6'd0;
      end
    endfunction
    function C35_t C2_35_dc (logic valid);
      begin
        C2_35_dc = 7'bx;
        C2_35_dc[0:0] = valid;
        C2_35_dc[6:1] = 6'd1;
      end
    endfunction
    function C35_t C3_35_dc (logic valid);
      begin
        C3_35_dc = 7'bx;
        C3_35_dc[0:0] = valid;
        C3_35_dc[6:1] = 6'd2;
      end
    endfunction
    function C35_t C4_35_dc (logic valid);
      begin
        C4_35_dc = 7'bx;
        C4_35_dc[0:0] = valid;
        C4_35_dc[6:1] = 6'd3;
      end
    endfunction
    function C35_t C5_35_dc (logic valid);
      begin
        C5_35_dc = 7'bx;
        C5_35_dc[0:0] = valid;
        C5_35_dc[6:1] = 6'd4;
      end
    endfunction
    function C35_t C6_35_dc (logic valid);
      begin
        C6_35_dc = 7'bx;
        C6_35_dc[0:0] = valid;
        C6_35_dc[6:1] = 6'd5;
      end
    endfunction
    function C35_t C7_35_dc (logic valid);
      begin
        C7_35_dc = 7'bx;
        C7_35_dc[0:0] = valid;
        C7_35_dc[6:1] = 6'd6;
      end
    endfunction
    function C35_t C8_35_dc (logic valid);
      begin
        C8_35_dc = 7'bx;
        C8_35_dc[0:0] = valid;
        C8_35_dc[6:1] = 6'd7;
      end
    endfunction
    function C35_t C9_35_dc (logic valid);
      begin
        C9_35_dc = 7'bx;
        C9_35_dc[0:0] = valid;
        C9_35_dc[6:1] = 6'd8;
      end
    endfunction
    function C35_t C10_35_dc (logic valid);
      begin
        C10_35_dc = 7'bx;
        C10_35_dc[0:0] = valid;
        C10_35_dc[6:1] = 6'd9;
      end
    endfunction
    function C35_t C11_35_dc (logic valid);
      begin
        C11_35_dc = 7'bx;
        C11_35_dc[0:0] = valid;
        C11_35_dc[6:1] = 6'd10;
      end
    endfunction
    function C35_t C12_35_dc (logic valid);
      begin
        C12_35_dc = 7'bx;
        C12_35_dc[0:0] = valid;
        C12_35_dc[6:1] = 6'd11;
      end
    endfunction
    function C35_t C13_35_dc (logic valid);
      begin
        C13_35_dc = 7'bx;
        C13_35_dc[0:0] = valid;
        C13_35_dc[6:1] = 6'd12;
      end
    endfunction
    function C35_t C14_35_dc (logic valid);
      begin
        C14_35_dc = 7'bx;
        C14_35_dc[0:0] = valid;
        C14_35_dc[6:1] = 6'd13;
      end
    endfunction
    function C35_t C15_35_dc (logic valid);
      begin
        C15_35_dc = 7'bx;
        C15_35_dc[0:0] = valid;
        C15_35_dc[6:1] = 6'd14;
      end
    endfunction
    function C35_t C16_35_dc (logic valid);
      begin
        C16_35_dc = 7'bx;
        C16_35_dc[0:0] = valid;
        C16_35_dc[6:1] = 6'd15;
      end
    endfunction
    function C35_t C17_35_dc (logic valid);
      begin
        C17_35_dc = 7'bx;
        C17_35_dc[0:0] = valid;
        C17_35_dc[6:1] = 6'd16;
      end
    endfunction
    function C35_t C18_35_dc (logic valid);
      begin
        C18_35_dc = 7'bx;
        C18_35_dc[0:0] = valid;
        C18_35_dc[6:1] = 6'd17;
      end
    endfunction
    function C35_t C19_35_dc (logic valid);
      begin
        C19_35_dc = 7'bx;
        C19_35_dc[0:0] = valid;
        C19_35_dc[6:1] = 6'd18;
      end
    endfunction
    function C35_t C20_35_dc (logic valid);
      begin
        C20_35_dc = 7'bx;
        C20_35_dc[0:0] = valid;
        C20_35_dc[6:1] = 6'd19;
      end
    endfunction
    function C35_t C21_35_dc (logic valid);
      begin
        C21_35_dc = 7'bx;
        C21_35_dc[0:0] = valid;
        C21_35_dc[6:1] = 6'd20;
      end
    endfunction
    function C35_t C22_35_dc (logic valid);
      begin
        C22_35_dc = 7'bx;
        C22_35_dc[0:0] = valid;
        C22_35_dc[6:1] = 6'd21;
      end
    endfunction
    function C35_t C23_35_dc (logic valid);
      begin
        C23_35_dc = 7'bx;
        C23_35_dc[0:0] = valid;
        C23_35_dc[6:1] = 6'd22;
      end
    endfunction
    function C35_t C24_35_dc (logic valid);
      begin
        C24_35_dc = 7'bx;
        C24_35_dc[0:0] = valid;
        C24_35_dc[6:1] = 6'd23;
      end
    endfunction
    function C35_t C25_35_dc (logic valid);
      begin
        C25_35_dc = 7'bx;
        C25_35_dc[0:0] = valid;
        C25_35_dc[6:1] = 6'd24;
      end
    endfunction
    function C35_t C26_35_dc (logic valid);
      begin
        C26_35_dc = 7'bx;
        C26_35_dc[0:0] = valid;
        C26_35_dc[6:1] = 6'd25;
      end
    endfunction
    function C35_t C27_35_dc (logic valid);
      begin
        C27_35_dc = 7'bx;
        C27_35_dc[0:0] = valid;
        C27_35_dc[6:1] = 6'd26;
      end
    endfunction
    function C35_t C28_35_dc (logic valid);
      begin
        C28_35_dc = 7'bx;
        C28_35_dc[0:0] = valid;
        C28_35_dc[6:1] = 6'd27;
      end
    endfunction
    function C35_t C29_35_dc (logic valid);
      begin
        C29_35_dc = 7'bx;
        C29_35_dc[0:0] = valid;
        C29_35_dc[6:1] = 6'd28;
      end
    endfunction
    function C35_t C30_35_dc (logic valid);
      begin
        C30_35_dc = 7'bx;
        C30_35_dc[0:0] = valid;
        C30_35_dc[6:1] = 6'd29;
      end
    endfunction
    function C35_t C31_35_dc (logic valid);
      begin
        C31_35_dc = 7'bx;
        C31_35_dc[0:0] = valid;
        C31_35_dc[6:1] = 6'd30;
      end
    endfunction
    function C35_t C32_35_dc (logic valid);
      begin
        C32_35_dc = 7'bx;
        C32_35_dc[0:0] = valid;
        C32_35_dc[6:1] = 6'd31;
      end
    endfunction
    function C35_t C33_35_dc (logic valid);
      begin
        C33_35_dc = 7'bx;
        C33_35_dc[0:0] = valid;
        C33_35_dc[6:1] = 6'd32;
      end
    endfunction
    function C35_t C34_35_dc (logic valid);
      begin
        C34_35_dc = 7'bx;
        C34_35_dc[0:0] = valid;
        C34_35_dc[6:1] = 6'd33;
      end
    endfunction
    function C35_t C35_35_dc (logic valid);
      begin
        C35_35_dc = 7'bx;
        C35_35_dc[0:0] = valid;
        C35_35_dc[6:1] = 6'd34;
      end
    endfunction
    typedef logic [0:0] Go_t;
    function Go_t Go_dc (logic valid);
      begin
        Go_dc = 1'bx;
        Go_dc[0:0] = valid;
      end
    endfunction
    typedef logic [16:0] Pointer_QTree_Bool_t;
    function Pointer_QTree_Bool_t Pointer_QTree_Bool_dc (logic valid, \Word16#_t  z1);
      begin
        Pointer_QTree_Bool_dc = 17'bx;
        Pointer_QTree_Bool_dc[0:0] = valid;
        Pointer_QTree_Bool_dc[16:1] = z1[16:1];
      end
    endfunction
    typedef logic [1:0] MyBool_t;
    function MyBool_t MyFalse_dc (logic valid, Go_t z1);
      begin
        MyFalse_dc = 2'bx;
        MyFalse_dc[0:0] = valid;
        MyFalse_dc[1:1] = 1'd0;
        ;
      end
    endfunction
    function MyBool_t MyTrue_dc (logic valid, Go_t z1);
      begin
        MyTrue_dc = 2'bx;
        MyTrue_dc[0:0] = valid;
        MyTrue_dc[1:1] = 1'd1;
        ;
      end
    endfunction
    typedef logic [66:0] QTree_Bool_t;
    function QTree_Bool_t QNone_Bool_dc (logic valid, Go_t z1);
      begin
        QNone_Bool_dc = 67'bx;
        QNone_Bool_dc[0:0] = valid;
        QNone_Bool_dc[2:1] = 2'd0;
        ;
      end
    endfunction
    function QTree_Bool_t QVal_Bool_dc (logic valid, MyBool_t z1);
      begin
        QVal_Bool_dc = 67'bx;
        QVal_Bool_dc[0:0] = valid;
        QVal_Bool_dc[2:1] = 2'd1;
        QVal_Bool_dc[3:3] = z1[1:1];
      end
    endfunction
    function QTree_Bool_t QNode_Bool_dc (logic valid, Pointer_QTree_Bool_t z1, Pointer_QTree_Bool_t z2, Pointer_QTree_Bool_t z3, Pointer_QTree_Bool_t z4);
      begin
        QNode_Bool_dc = 67'bx;
        QNode_Bool_dc[0:0] = valid;
        QNode_Bool_dc[2:1] = 2'd2;
        QNode_Bool_dc[18:3] = z1[16:1];
        QNode_Bool_dc[34:19] = z2[16:1];
        QNode_Bool_dc[50:35] = z3[16:1];
        QNode_Bool_dc[66:51] = z4[16:1];
      end
    endfunction
    function QTree_Bool_t QError_Bool_dc (logic valid, Go_t z1);
      begin
        QError_Bool_dc = 67'bx;
        QError_Bool_dc[0:0] = valid;
        QError_Bool_dc[2:1] = 2'd3;
        ;
      end
    endfunction
    typedef logic [83:0] MemIn_QTree_Bool_t;
    function MemIn_QTree_Bool_t ReadIn_QTree_Bool_dc (logic valid, \Word16#_t  z1);
      begin
        ReadIn_QTree_Bool_dc = 84'bx;
        ReadIn_QTree_Bool_dc[0:0] = valid;
        ReadIn_QTree_Bool_dc[1:1] = 1'd0;
        ReadIn_QTree_Bool_dc[17:2] = z1[16:1];
      end
    endfunction
    function MemIn_QTree_Bool_t WriteIn_QTree_Bool_dc (logic valid, \Word16#_t  z1, QTree_Bool_t z2);
      begin
        WriteIn_QTree_Bool_dc = 84'bx;
        WriteIn_QTree_Bool_dc[0:0] = valid;
        WriteIn_QTree_Bool_dc[1:1] = 1'd1;
        WriteIn_QTree_Bool_dc[17:2] = z1[16:1];
        WriteIn_QTree_Bool_dc[83:18] = z2[66:1];
      end
    endfunction
    typedef logic [67:0] MemOut_QTree_Bool_t;
    function MemOut_QTree_Bool_t ReadOut_QTree_Bool_dc (logic valid, QTree_Bool_t z1);
      begin
        ReadOut_QTree_Bool_dc = 68'bx;
        ReadOut_QTree_Bool_dc[0:0] = valid;
        ReadOut_QTree_Bool_dc[1:1] = 1'd0;
        ReadOut_QTree_Bool_dc[67:2] = z1[66:1];
      end
    endfunction
    function MemOut_QTree_Bool_t ACK_QTree_Bool_dc (logic valid);
      begin
        ACK_QTree_Bool_dc = 68'bx;
        ACK_QTree_Bool_dc[0:0] = valid;
        ACK_QTree_Bool_dc[1:1] = 1'd1;
      end
    endfunction
    typedef logic [16:0] Pointer_CTf_t;
    function Pointer_CTf_t Pointer_CTf_dc (logic valid, \Word16#_t  z1);
      begin
        Pointer_CTf_dc = 17'bx;
        Pointer_CTf_dc[0:0] = valid;
        Pointer_CTf_dc[16:1] = z1[16:1];
      end
    endfunction
    typedef logic [163:0] CTf_t;
    function CTf_t Lfsbos_dc (logic valid, Go_t z1);
      begin
        Lfsbos_dc = 164'bx;
        Lfsbos_dc[0:0] = valid;
        Lfsbos_dc[3:1] = 3'd0;
        ;
      end
    endfunction
    function CTf_t Lcall_f3_dc (logic valid, Pointer_CTf_t z1, Pointer_QTree_Bool_t z2, Pointer_QTree_Bool_t z3, Pointer_QTree_Bool_t z4, Pointer_QTree_Bool_t z5, Pointer_QTree_Bool_t z6, Pointer_QTree_Bool_t z7, Pointer_QTree_Bool_t z8, Pointer_QTree_Bool_t z9, Pointer_QTree_Bool_t z10);
      begin
        Lcall_f3_dc = 164'bx;
        Lcall_f3_dc[0:0] = valid;
        Lcall_f3_dc[3:1] = 3'd1;
        Lcall_f3_dc[19:4] = z1[16:1];
        Lcall_f3_dc[35:20] = z2[16:1];
        Lcall_f3_dc[51:36] = z3[16:1];
        Lcall_f3_dc[67:52] = z4[16:1];
        Lcall_f3_dc[83:68] = z5[16:1];
        Lcall_f3_dc[99:84] = z6[16:1];
        Lcall_f3_dc[115:100] = z7[16:1];
        Lcall_f3_dc[131:116] = z8[16:1];
        Lcall_f3_dc[147:132] = z9[16:1];
        Lcall_f3_dc[163:148] = z10[16:1];
      end
    endfunction
    function CTf_t Lcall_f2_dc (logic valid, Pointer_QTree_Bool_t z1, Pointer_CTf_t z2, Pointer_QTree_Bool_t z3, Pointer_QTree_Bool_t z4, Pointer_QTree_Bool_t z5, Pointer_QTree_Bool_t z6, Pointer_QTree_Bool_t z7, Pointer_QTree_Bool_t z8);
      begin
        Lcall_f2_dc = 164'bx;
        Lcall_f2_dc[0:0] = valid;
        Lcall_f2_dc[3:1] = 3'd2;
        Lcall_f2_dc[19:4] = z1[16:1];
        Lcall_f2_dc[35:20] = z2[16:1];
        Lcall_f2_dc[51:36] = z3[16:1];
        Lcall_f2_dc[67:52] = z4[16:1];
        Lcall_f2_dc[83:68] = z5[16:1];
        Lcall_f2_dc[99:84] = z6[16:1];
        Lcall_f2_dc[115:100] = z7[16:1];
        Lcall_f2_dc[131:116] = z8[16:1];
      end
    endfunction
    function CTf_t Lcall_f1_dc (logic valid, Pointer_QTree_Bool_t z1, Pointer_QTree_Bool_t z2, Pointer_CTf_t z3, Pointer_QTree_Bool_t z4, Pointer_QTree_Bool_t z5, Pointer_QTree_Bool_t z6);
      begin
        Lcall_f1_dc = 164'bx;
        Lcall_f1_dc[0:0] = valid;
        Lcall_f1_dc[3:1] = 3'd3;
        Lcall_f1_dc[19:4] = z1[16:1];
        Lcall_f1_dc[35:20] = z2[16:1];
        Lcall_f1_dc[51:36] = z3[16:1];
        Lcall_f1_dc[67:52] = z4[16:1];
        Lcall_f1_dc[83:68] = z5[16:1];
        Lcall_f1_dc[99:84] = z6[16:1];
      end
    endfunction
    function CTf_t Lcall_f0_dc (logic valid, Pointer_QTree_Bool_t z1, Pointer_QTree_Bool_t z2, Pointer_QTree_Bool_t z3, Pointer_CTf_t z4);
      begin
        Lcall_f0_dc = 164'bx;
        Lcall_f0_dc[0:0] = valid;
        Lcall_f0_dc[3:1] = 3'd4;
        Lcall_f0_dc[19:4] = z1[16:1];
        Lcall_f0_dc[35:20] = z2[16:1];
        Lcall_f0_dc[51:36] = z3[16:1];
        Lcall_f0_dc[67:52] = z4[16:1];
      end
    endfunction
    typedef logic [180:0] MemIn_CTf_t;
    function MemIn_CTf_t ReadIn_CTf_dc (logic valid, \Word16#_t  z1);
      begin
        ReadIn_CTf_dc = 181'bx;
        ReadIn_CTf_dc[0:0] = valid;
        ReadIn_CTf_dc[1:1] = 1'd0;
        ReadIn_CTf_dc[17:2] = z1[16:1];
      end
    endfunction
    function MemIn_CTf_t WriteIn_CTf_dc (logic valid, \Word16#_t  z1, CTf_t z2);
      begin
        WriteIn_CTf_dc = 181'bx;
        WriteIn_CTf_dc[0:0] = valid;
        WriteIn_CTf_dc[1:1] = 1'd1;
        WriteIn_CTf_dc[17:2] = z1[16:1];
        WriteIn_CTf_dc[180:18] = z2[163:1];
      end
    endfunction
    typedef logic [164:0] MemOut_CTf_t;
    function MemOut_CTf_t ReadOut_CTf_dc (logic valid, CTf_t z1);
      begin
        ReadOut_CTf_dc = 165'bx;
        ReadOut_CTf_dc[0:0] = valid;
        ReadOut_CTf_dc[1:1] = 1'd0;
        ReadOut_CTf_dc[164:2] = z1[163:1];
      end
    endfunction
    function MemOut_CTf_t ACK_CTf_dc (logic valid);
      begin
        ACK_CTf_dc = 165'bx;
        ACK_CTf_dc[0:0] = valid;
        ACK_CTf_dc[1:1] = 1'd1;
      end
    endfunction
    typedef logic [16:0] \Pointer_CTf''''''''''''_t ;
    function \Pointer_CTf''''''''''''_t  \Pointer_CTf''''''''''''_dc  (logic valid, \Word16#_t  z1);
      begin
        \Pointer_CTf''''''''''''_dc  = 17'bx;
        \Pointer_CTf''''''''''''_dc [0:0] = valid;
        \Pointer_CTf''''''''''''_dc [16:1] = z1[16:1];
      end
    endfunction
    typedef logic [115:0] \CTf''''''''''''_t ;
    function \CTf''''''''''''_t  \Lf''''''''''''sbos_dc  (logic valid, Go_t z1);
      begin
        \Lf''''''''''''sbos_dc  = 116'bx;
        \Lf''''''''''''sbos_dc [0:0] = valid;
        \Lf''''''''''''sbos_dc [3:1] = 3'd0;
        ;
      end
    endfunction
    function \CTf''''''''''''_t  \Lcall_f''''''''''''3_dc  (logic valid, \Pointer_CTf''''''''''''_t  z1, Pointer_QTree_Bool_t z2, Pointer_QTree_Bool_t z3, Pointer_QTree_Bool_t z4, Pointer_QTree_Bool_t z5, Pointer_QTree_Bool_t z6, Pointer_QTree_Bool_t z7);
      begin
        \Lcall_f''''''''''''3_dc  = 116'bx;
        \Lcall_f''''''''''''3_dc [0:0] = valid;
        \Lcall_f''''''''''''3_dc [3:1] = 3'd1;
        \Lcall_f''''''''''''3_dc [19:4] = z1[16:1];
        \Lcall_f''''''''''''3_dc [35:20] = z2[16:1];
        \Lcall_f''''''''''''3_dc [51:36] = z3[16:1];
        \Lcall_f''''''''''''3_dc [67:52] = z4[16:1];
        \Lcall_f''''''''''''3_dc [83:68] = z5[16:1];
        \Lcall_f''''''''''''3_dc [99:84] = z6[16:1];
        \Lcall_f''''''''''''3_dc [115:100] = z7[16:1];
      end
    endfunction
    function \CTf''''''''''''_t  \Lcall_f''''''''''''2_dc  (logic valid, Pointer_QTree_Bool_t z1, \Pointer_CTf''''''''''''_t  z2, Pointer_QTree_Bool_t z3, Pointer_QTree_Bool_t z4, Pointer_QTree_Bool_t z5, Pointer_QTree_Bool_t z6);
      begin
        \Lcall_f''''''''''''2_dc  = 116'bx;
        \Lcall_f''''''''''''2_dc [0:0] = valid;
        \Lcall_f''''''''''''2_dc [3:1] = 3'd2;
        \Lcall_f''''''''''''2_dc [19:4] = z1[16:1];
        \Lcall_f''''''''''''2_dc [35:20] = z2[16:1];
        \Lcall_f''''''''''''2_dc [51:36] = z3[16:1];
        \Lcall_f''''''''''''2_dc [67:52] = z4[16:1];
        \Lcall_f''''''''''''2_dc [83:68] = z5[16:1];
        \Lcall_f''''''''''''2_dc [99:84] = z6[16:1];
      end
    endfunction
    function \CTf''''''''''''_t  \Lcall_f''''''''''''1_dc  (logic valid, Pointer_QTree_Bool_t z1, Pointer_QTree_Bool_t z2, \Pointer_CTf''''''''''''_t  z3, Pointer_QTree_Bool_t z4, Pointer_QTree_Bool_t z5);
      begin
        \Lcall_f''''''''''''1_dc  = 116'bx;
        \Lcall_f''''''''''''1_dc [0:0] = valid;
        \Lcall_f''''''''''''1_dc [3:1] = 3'd3;
        \Lcall_f''''''''''''1_dc [19:4] = z1[16:1];
        \Lcall_f''''''''''''1_dc [35:20] = z2[16:1];
        \Lcall_f''''''''''''1_dc [51:36] = z3[16:1];
        \Lcall_f''''''''''''1_dc [67:52] = z4[16:1];
        \Lcall_f''''''''''''1_dc [83:68] = z5[16:1];
      end
    endfunction
    function \CTf''''''''''''_t  \Lcall_f''''''''''''0_dc  (logic valid, Pointer_QTree_Bool_t z1, Pointer_QTree_Bool_t z2, Pointer_QTree_Bool_t z3, \Pointer_CTf''''''''''''_t  z4);
      begin
        \Lcall_f''''''''''''0_dc  = 116'bx;
        \Lcall_f''''''''''''0_dc [0:0] = valid;
        \Lcall_f''''''''''''0_dc [3:1] = 3'd4;
        \Lcall_f''''''''''''0_dc [19:4] = z1[16:1];
        \Lcall_f''''''''''''0_dc [35:20] = z2[16:1];
        \Lcall_f''''''''''''0_dc [51:36] = z3[16:1];
        \Lcall_f''''''''''''0_dc [67:52] = z4[16:1];
      end
    endfunction
    typedef logic [132:0] \MemIn_CTf''''''''''''_t ;
    function \MemIn_CTf''''''''''''_t  \ReadIn_CTf''''''''''''_dc  (logic valid, \Word16#_t  z1);
      begin
        \ReadIn_CTf''''''''''''_dc  = 133'bx;
        \ReadIn_CTf''''''''''''_dc [0:0] = valid;
        \ReadIn_CTf''''''''''''_dc [1:1] = 1'd0;
        \ReadIn_CTf''''''''''''_dc [17:2] = z1[16:1];
      end
    endfunction
    function \MemIn_CTf''''''''''''_t  \WriteIn_CTf''''''''''''_dc  (logic valid, \Word16#_t  z1, \CTf''''''''''''_t  z2);
      begin
        \WriteIn_CTf''''''''''''_dc  = 133'bx;
        \WriteIn_CTf''''''''''''_dc [0:0] = valid;
        \WriteIn_CTf''''''''''''_dc [1:1] = 1'd1;
        \WriteIn_CTf''''''''''''_dc [17:2] = z1[16:1];
        \WriteIn_CTf''''''''''''_dc [132:18] = z2[115:1];
      end
    endfunction
    typedef logic [116:0] \MemOut_CTf''''''''''''_t ;
    function \MemOut_CTf''''''''''''_t  \ReadOut_CTf''''''''''''_dc  (logic valid, \CTf''''''''''''_t  z1);
      begin
        \ReadOut_CTf''''''''''''_dc  = 117'bx;
        \ReadOut_CTf''''''''''''_dc [0:0] = valid;
        \ReadOut_CTf''''''''''''_dc [1:1] = 1'd0;
        \ReadOut_CTf''''''''''''_dc [116:2] = z1[115:1];
      end
    endfunction
    function \MemOut_CTf''''''''''''_t  \ACK_CTf''''''''''''_dc  (logic valid);
      begin
        \ACK_CTf''''''''''''_dc  = 117'bx;
        \ACK_CTf''''''''''''_dc [0:0] = valid;
        \ACK_CTf''''''''''''_dc [1:1] = 1'd1;
      end
    endfunction
    typedef logic [4:0] C12_t;
    function C12_t C1_12_dc (logic valid);
      begin
        C1_12_dc = 5'bx;
        C1_12_dc[0:0] = valid;
        C1_12_dc[4:1] = 4'd0;
      end
    endfunction
    function C12_t C2_12_dc (logic valid);
      begin
        C2_12_dc = 5'bx;
        C2_12_dc[0:0] = valid;
        C2_12_dc[4:1] = 4'd1;
      end
    endfunction
    function C12_t C3_12_dc (logic valid);
      begin
        C3_12_dc = 5'bx;
        C3_12_dc[0:0] = valid;
        C3_12_dc[4:1] = 4'd2;
      end
    endfunction
    function C12_t C4_12_dc (logic valid);
      begin
        C4_12_dc = 5'bx;
        C4_12_dc[0:0] = valid;
        C4_12_dc[4:1] = 4'd3;
      end
    endfunction
    function C12_t C5_12_dc (logic valid);
      begin
        C5_12_dc = 5'bx;
        C5_12_dc[0:0] = valid;
        C5_12_dc[4:1] = 4'd4;
      end
    endfunction
    function C12_t C6_12_dc (logic valid);
      begin
        C6_12_dc = 5'bx;
        C6_12_dc[0:0] = valid;
        C6_12_dc[4:1] = 4'd5;
      end
    endfunction
    function C12_t C7_12_dc (logic valid);
      begin
        C7_12_dc = 5'bx;
        C7_12_dc[0:0] = valid;
        C7_12_dc[4:1] = 4'd6;
      end
    endfunction
    function C12_t C8_12_dc (logic valid);
      begin
        C8_12_dc = 5'bx;
        C8_12_dc[0:0] = valid;
        C8_12_dc[4:1] = 4'd7;
      end
    endfunction
    function C12_t C9_12_dc (logic valid);
      begin
        C9_12_dc = 5'bx;
        C9_12_dc[0:0] = valid;
        C9_12_dc[4:1] = 4'd8;
      end
    endfunction
    function C12_t C10_12_dc (logic valid);
      begin
        C10_12_dc = 5'bx;
        C10_12_dc[0:0] = valid;
        C10_12_dc[4:1] = 4'd9;
      end
    endfunction
    function C12_t C11_12_dc (logic valid);
      begin
        C11_12_dc = 5'bx;
        C11_12_dc[0:0] = valid;
        C11_12_dc[4:1] = 4'd10;
      end
    endfunction
    function C12_t C12_12_dc (logic valid);
      begin
        C12_12_dc = 5'bx;
        C12_12_dc[0:0] = valid;
        C12_12_dc[4:1] = 4'd11;
      end
    endfunction
    typedef logic [3:0] C5_t;
    function C5_t C1_5_dc (logic valid);
      begin
        C1_5_dc = 4'bx;
        C1_5_dc[0:0] = valid;
        C1_5_dc[3:1] = 3'd0;
      end
    endfunction
    function C5_t C2_5_dc (logic valid);
      begin
        C2_5_dc = 4'bx;
        C2_5_dc[0:0] = valid;
        C2_5_dc[3:1] = 3'd1;
      end
    endfunction
    function C5_t C3_5_dc (logic valid);
      begin
        C3_5_dc = 4'bx;
        C3_5_dc[0:0] = valid;
        C3_5_dc[3:1] = 3'd2;
      end
    endfunction
    function C5_t C4_5_dc (logic valid);
      begin
        C4_5_dc = 4'bx;
        C4_5_dc[0:0] = valid;
        C4_5_dc[3:1] = 3'd3;
      end
    endfunction
    function C5_t C5_5_dc (logic valid);
      begin
        C5_5_dc = 4'bx;
        C5_5_dc[0:0] = valid;
        C5_5_dc[3:1] = 3'd4;
      end
    endfunction
    typedef logic [6:0] C40_t;
    function C40_t C1_40_dc (logic valid);
      begin
        C1_40_dc = 7'bx;
        C1_40_dc[0:0] = valid;
        C1_40_dc[6:1] = 6'd0;
      end
    endfunction
    function C40_t C2_40_dc (logic valid);
      begin
        C2_40_dc = 7'bx;
        C2_40_dc[0:0] = valid;
        C2_40_dc[6:1] = 6'd1;
      end
    endfunction
    function C40_t C3_40_dc (logic valid);
      begin
        C3_40_dc = 7'bx;
        C3_40_dc[0:0] = valid;
        C3_40_dc[6:1] = 6'd2;
      end
    endfunction
    function C40_t C4_40_dc (logic valid);
      begin
        C4_40_dc = 7'bx;
        C4_40_dc[0:0] = valid;
        C4_40_dc[6:1] = 6'd3;
      end
    endfunction
    function C40_t C5_40_dc (logic valid);
      begin
        C5_40_dc = 7'bx;
        C5_40_dc[0:0] = valid;
        C5_40_dc[6:1] = 6'd4;
      end
    endfunction
    function C40_t C6_40_dc (logic valid);
      begin
        C6_40_dc = 7'bx;
        C6_40_dc[0:0] = valid;
        C6_40_dc[6:1] = 6'd5;
      end
    endfunction
    function C40_t C7_40_dc (logic valid);
      begin
        C7_40_dc = 7'bx;
        C7_40_dc[0:0] = valid;
        C7_40_dc[6:1] = 6'd6;
      end
    endfunction
    function C40_t C8_40_dc (logic valid);
      begin
        C8_40_dc = 7'bx;
        C8_40_dc[0:0] = valid;
        C8_40_dc[6:1] = 6'd7;
      end
    endfunction
    function C40_t C9_40_dc (logic valid);
      begin
        C9_40_dc = 7'bx;
        C9_40_dc[0:0] = valid;
        C9_40_dc[6:1] = 6'd8;
      end
    endfunction
    function C40_t C10_40_dc (logic valid);
      begin
        C10_40_dc = 7'bx;
        C10_40_dc[0:0] = valid;
        C10_40_dc[6:1] = 6'd9;
      end
    endfunction
    function C40_t C11_40_dc (logic valid);
      begin
        C11_40_dc = 7'bx;
        C11_40_dc[0:0] = valid;
        C11_40_dc[6:1] = 6'd10;
      end
    endfunction
    function C40_t C12_40_dc (logic valid);
      begin
        C12_40_dc = 7'bx;
        C12_40_dc[0:0] = valid;
        C12_40_dc[6:1] = 6'd11;
      end
    endfunction
    function C40_t C13_40_dc (logic valid);
      begin
        C13_40_dc = 7'bx;
        C13_40_dc[0:0] = valid;
        C13_40_dc[6:1] = 6'd12;
      end
    endfunction
    function C40_t C14_40_dc (logic valid);
      begin
        C14_40_dc = 7'bx;
        C14_40_dc[0:0] = valid;
        C14_40_dc[6:1] = 6'd13;
      end
    endfunction
    function C40_t C15_40_dc (logic valid);
      begin
        C15_40_dc = 7'bx;
        C15_40_dc[0:0] = valid;
        C15_40_dc[6:1] = 6'd14;
      end
    endfunction
    function C40_t C16_40_dc (logic valid);
      begin
        C16_40_dc = 7'bx;
        C16_40_dc[0:0] = valid;
        C16_40_dc[6:1] = 6'd15;
      end
    endfunction
    function C40_t C17_40_dc (logic valid);
      begin
        C17_40_dc = 7'bx;
        C17_40_dc[0:0] = valid;
        C17_40_dc[6:1] = 6'd16;
      end
    endfunction
    function C40_t C18_40_dc (logic valid);
      begin
        C18_40_dc = 7'bx;
        C18_40_dc[0:0] = valid;
        C18_40_dc[6:1] = 6'd17;
      end
    endfunction
    function C40_t C19_40_dc (logic valid);
      begin
        C19_40_dc = 7'bx;
        C19_40_dc[0:0] = valid;
        C19_40_dc[6:1] = 6'd18;
      end
    endfunction
    function C40_t C20_40_dc (logic valid);
      begin
        C20_40_dc = 7'bx;
        C20_40_dc[0:0] = valid;
        C20_40_dc[6:1] = 6'd19;
      end
    endfunction
    function C40_t C21_40_dc (logic valid);
      begin
        C21_40_dc = 7'bx;
        C21_40_dc[0:0] = valid;
        C21_40_dc[6:1] = 6'd20;
      end
    endfunction
    function C40_t C22_40_dc (logic valid);
      begin
        C22_40_dc = 7'bx;
        C22_40_dc[0:0] = valid;
        C22_40_dc[6:1] = 6'd21;
      end
    endfunction
    function C40_t C23_40_dc (logic valid);
      begin
        C23_40_dc = 7'bx;
        C23_40_dc[0:0] = valid;
        C23_40_dc[6:1] = 6'd22;
      end
    endfunction
    function C40_t C24_40_dc (logic valid);
      begin
        C24_40_dc = 7'bx;
        C24_40_dc[0:0] = valid;
        C24_40_dc[6:1] = 6'd23;
      end
    endfunction
    function C40_t C25_40_dc (logic valid);
      begin
        C25_40_dc = 7'bx;
        C25_40_dc[0:0] = valid;
        C25_40_dc[6:1] = 6'd24;
      end
    endfunction
    function C40_t C26_40_dc (logic valid);
      begin
        C26_40_dc = 7'bx;
        C26_40_dc[0:0] = valid;
        C26_40_dc[6:1] = 6'd25;
      end
    endfunction
    function C40_t C27_40_dc (logic valid);
      begin
        C27_40_dc = 7'bx;
        C27_40_dc[0:0] = valid;
        C27_40_dc[6:1] = 6'd26;
      end
    endfunction
    function C40_t C28_40_dc (logic valid);
      begin
        C28_40_dc = 7'bx;
        C28_40_dc[0:0] = valid;
        C28_40_dc[6:1] = 6'd27;
      end
    endfunction
    function C40_t C29_40_dc (logic valid);
      begin
        C29_40_dc = 7'bx;
        C29_40_dc[0:0] = valid;
        C29_40_dc[6:1] = 6'd28;
      end
    endfunction
    function C40_t C30_40_dc (logic valid);
      begin
        C30_40_dc = 7'bx;
        C30_40_dc[0:0] = valid;
        C30_40_dc[6:1] = 6'd29;
      end
    endfunction
    function C40_t C31_40_dc (logic valid);
      begin
        C31_40_dc = 7'bx;
        C31_40_dc[0:0] = valid;
        C31_40_dc[6:1] = 6'd30;
      end
    endfunction
    function C40_t C32_40_dc (logic valid);
      begin
        C32_40_dc = 7'bx;
        C32_40_dc[0:0] = valid;
        C32_40_dc[6:1] = 6'd31;
      end
    endfunction
    function C40_t C33_40_dc (logic valid);
      begin
        C33_40_dc = 7'bx;
        C33_40_dc[0:0] = valid;
        C33_40_dc[6:1] = 6'd32;
      end
    endfunction
    function C40_t C34_40_dc (logic valid);
      begin
        C34_40_dc = 7'bx;
        C34_40_dc[0:0] = valid;
        C34_40_dc[6:1] = 6'd33;
      end
    endfunction
    function C40_t C35_40_dc (logic valid);
      begin
        C35_40_dc = 7'bx;
        C35_40_dc[0:0] = valid;
        C35_40_dc[6:1] = 6'd34;
      end
    endfunction
    function C40_t C36_40_dc (logic valid);
      begin
        C36_40_dc = 7'bx;
        C36_40_dc[0:0] = valid;
        C36_40_dc[6:1] = 6'd35;
      end
    endfunction
    function C40_t C37_40_dc (logic valid);
      begin
        C37_40_dc = 7'bx;
        C37_40_dc[0:0] = valid;
        C37_40_dc[6:1] = 6'd36;
      end
    endfunction
    function C40_t C38_40_dc (logic valid);
      begin
        C38_40_dc = 7'bx;
        C38_40_dc[0:0] = valid;
        C38_40_dc[6:1] = 6'd37;
      end
    endfunction
    function C40_t C39_40_dc (logic valid);
      begin
        C39_40_dc = 7'bx;
        C39_40_dc[0:0] = valid;
        C39_40_dc[6:1] = 6'd38;
      end
    endfunction
    function C40_t C40_40_dc (logic valid);
      begin
        C40_40_dc = 7'bx;
        C40_40_dc[0:0] = valid;
        C40_40_dc[6:1] = 6'd39;
      end
    endfunction
    typedef logic [4:0] C10_t;
    function C10_t C1_10_dc (logic valid);
      begin
        C1_10_dc = 5'bx;
        C1_10_dc[0:0] = valid;
        C1_10_dc[4:1] = 4'd0;
      end
    endfunction
    function C10_t C2_10_dc (logic valid);
      begin
        C2_10_dc = 5'bx;
        C2_10_dc[0:0] = valid;
        C2_10_dc[4:1] = 4'd1;
      end
    endfunction
    function C10_t C3_10_dc (logic valid);
      begin
        C3_10_dc = 5'bx;
        C3_10_dc[0:0] = valid;
        C3_10_dc[4:1] = 4'd2;
      end
    endfunction
    function C10_t C4_10_dc (logic valid);
      begin
        C4_10_dc = 5'bx;
        C4_10_dc[0:0] = valid;
        C4_10_dc[4:1] = 4'd3;
      end
    endfunction
    function C10_t C5_10_dc (logic valid);
      begin
        C5_10_dc = 5'bx;
        C5_10_dc[0:0] = valid;
        C5_10_dc[4:1] = 4'd4;
      end
    endfunction
    function C10_t C6_10_dc (logic valid);
      begin
        C6_10_dc = 5'bx;
        C6_10_dc[0:0] = valid;
        C6_10_dc[4:1] = 4'd5;
      end
    endfunction
    function C10_t C7_10_dc (logic valid);
      begin
        C7_10_dc = 5'bx;
        C7_10_dc[0:0] = valid;
        C7_10_dc[4:1] = 4'd6;
      end
    endfunction
    function C10_t C8_10_dc (logic valid);
      begin
        C8_10_dc = 5'bx;
        C8_10_dc[0:0] = valid;
        C8_10_dc[4:1] = 4'd7;
      end
    endfunction
    function C10_t C9_10_dc (logic valid);
      begin
        C9_10_dc = 5'bx;
        C9_10_dc[0:0] = valid;
        C9_10_dc[4:1] = 4'd8;
      end
    endfunction
    function C10_t C10_10_dc (logic valid);
      begin
        C10_10_dc = 5'bx;
        C10_10_dc[0:0] = valid;
        C10_10_dc[4:1] = 4'd9;
      end
    endfunction
    typedef logic [48:0] \TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf''''''''''''_t ;
    function \TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf''''''''''''_t  \TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf''''''''''''_dc  (logic valid, Go_t z1, Pointer_QTree_Bool_t z2, Pointer_QTree_Bool_t z3, \Pointer_CTf''''''''''''_t  z4);
      begin
        \TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf''''''''''''_dc  = 49'bx;
        \TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf''''''''''''_dc [0:0] = valid;
        ;
        \TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf''''''''''''_dc [16:1] = z2[16:1];
        \TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf''''''''''''_dc [32:17] = z3[16:1];
        \TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf''''''''''''_dc [48:33] = z4[16:1];
      end
    endfunction
    typedef logic [64:0] TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf_t;
    function TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf_t TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf_dc (logic valid, Go_t z1, Pointer_QTree_Bool_t z2, Pointer_QTree_Bool_t z3, Pointer_QTree_Bool_t z4, Pointer_CTf_t z5);
      begin
        TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf_dc = 65'bx;
        TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf_dc[0:0] = valid;
        ;
        TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf_dc[16:1] = z2[16:1];
        TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf_dc[32:17] = z3[16:1];
        TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf_dc[48:33] = z4[16:1];
        TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf_dc[64:49] = z5[16:1];
      end
    endfunction
    typedef logic [32:0] TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_t;
    function TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_t TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_dc (logic valid, Go_t z1, Pointer_QTree_Bool_t z2, Pointer_QTree_Bool_t z3);
      begin
        TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_dc = 33'bx;
        TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_dc[0:0] = valid;
        ;
        TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_dc[16:1] = z2[16:1];
        TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_dc[32:17] = z3[16:1];
      end
    endfunction
    typedef logic [48:0] TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_t;
    function TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_t TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_dc (logic valid, Go_t z1, Pointer_QTree_Bool_t z2, Pointer_QTree_Bool_t z3, Pointer_QTree_Bool_t z4);
      begin
        TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_dc = 49'bx;
        TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_dc[0:0] = valid;
        ;
        TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_dc[16:1] = z2[16:1];
        TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_dc[32:17] = z3[16:1];
        TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_dc[48:33] = z4[16:1];
      end
    endfunction
    typedef logic [0:0] TupGo_t;
    function TupGo_t TupGo_dc (logic valid, Go_t z1);
      begin
        TupGo_dc = 1'bx;
        TupGo_dc[0:0] = valid;
        ;
      end
    endfunction
endpackage